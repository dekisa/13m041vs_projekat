// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ycf535n69tLgcGzoU61/V68pVnn3c5ZeHhmalVLKmFS9zrusfC7Yfx3ix6WZmt2dRK1ijuw0dozv
tmz8I4dBHdX/d29wjGIrUQVsJmyXbsjIt4RK3E0fQ6J2daIw+b3n0K97kyMs0g2lcMxOueS5DjNe
jIAOJGFFu9Qszl+8EZHZfmMtCt8FchKBdXSFXQL5BR6tr10pbyItkvzMandjycbO8u68e7Y+OMwY
LFCc98q+NI8o+esX/ntTrfmtXgA7D4f992oQZ2eu5jEuobMSJJOvU9gCbYVfqMlUSBLNI36bZPDq
8TVHwWtes0OAbuKAMP6WgoS9W4fbHEULPoV1fQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 30448)
YRza+sQcKduKWZaRTUbtKXtdrUipoEuUsUEVfzjFP+ROrW50pQAmHORXbMNMgOKf//Dx2htK2aG3
lS/38jp1TJbvfsqJ95ZNRNpr4KFfaKavIDiWaBDkzv2Pf3kj48xo/O5XOA9JoyqtOyarz//qaTju
iQh+S55p8emX0+S3SOi/z0Wvw/8hG60xzYapKNIy3uIqSaWqEsvXgBBI0xIiz59P8/XHaVS1cpqg
/y9UYkYqn4lCuWQAIw6A52Bgz301RTIUBk1X+igrKUd5cKMwU4NvQ8gvN4uWt0Jxl1WQLi8SkiSl
ZNZIpRqEMOkqqer+Dd5sWkd/RvVl4s3khmt6UxfWwBgsyT80RvjiIbUTiVPBUZ52kX3mxPdCcObq
+aw1V16tpBGSUKwDQBkTtPQfYCM5VyBdfoT03PbZ0PnNfem0Yj/bGJPOWlAgT3qJnGdWkImJGVFJ
uBLSWbfksNzIDIpZuN6svSaNSqJtWl3enfWmjbtAug3eK59cQWVwJ62R7mGZU4B9N+O59SrVThDR
+IbKvxmzo+fDjwpsaBuVjUwmqzk0bOJZs4jIOlJgFPB4K8aXQUqWaosQ33XvtDMqm8c21ZhHAa6Z
gATehMRQ/3I+sP2A+qAIKhhgbgnOr9sF6yQCAQuqH4mO26GBrr4gYu41Qgs89yz4n0imzbzjXAfc
9el3J3PUSFoT4F4HIt2v8a1qLuS2mifJpPuQmxAZZ6KgTsqm6+CU7bA0tXZfchNQqDfA155V/87V
qjIugkn0sVmxNutOmUmFtOJRP7JVJ6E/iWvlXS21/6KOiAUjVKAVTbid7IfJ63z7QYXxdqCNdqc2
PgTvRfGg5kAjeL/kM7+Cq05tcgawnER1gnbK3+oXTUBWo35E8QhpDRSN/ZpTvbyxAl9fNrPEMvCf
JAj0n7ylnwNMXFrgnMNArDP+SoBm7cGOTSk8LwXFFMa7frATyQHhr6fXRyAD2VL0F8UXVCBrPDHL
CNozB/lDawqgnwjU+4spSVXBfMKgaMQmbMnb+GR59+3BGdWJYqRCSWbCijrZL8k8aP3G2VVGO528
WNyUPnCngt8b3ondk83mTZtI8Y18jUoN25e2TeH6quNwT85jzSPheOGQALf4HO0C/6urjOiORY4S
SYMXEvsTOl0XJBt04UqENduAUevcHQyF5bjDXZfhmNj2fxlebO5MjebVFoZ+jYYVaabGqd+4Lrdv
DPiIS76baw5tM1PTsXZKWIDIOWph0e77FNYVlH4fkNeHQh8Y+VNDRgZ5paVRMq6srtKOgdB9TJlX
OdX4i1/F4x0n0JAdl3q1S7kKyaPzitaSfQDfoBXY/QY9pGnKUZh4pj/yLb42CeJ0sTKkXykR0WE6
Gwp2FR9YHNIuXfpbm9o4B9JlzDYyqDZcijslPttsyh/o6XxihRLTTy8RyYB2bdPDGX37RFAKDlTk
RObDm0C+lZnzoMB8Hp1uxWpA93vwMZcOmWZUgLGlo0l8nDC41SSpx/YNNXyXDVmVNLyHUzREFdp3
pZlw1VjF2wLS9kADR1XN6zlh4NBr9A+5+KOqdjxrbWbsAiiEYrUHTfVFq7spRoFk/MT19IZA9mYy
pQxX8CkzQ185HxpdvrtiJlCgfEli0DYe3a8VywpZOrGc9OPEaFqgonc8K+0fQ208Af07dxFdhlJ7
dwq8DqlmKgi/xiQ43L6uMMh/7e+STua0z1FFAaLHy7bPv9XfsSGyiPU6P4KyDh3ZOEfg1CpVtQbC
+LL6DyuV+AXzq3lsy5dfYL17sf8mRo8g6L6Arpcv7sH0txg31xrIvyTAo0XlbROJAIz6HxPeJ06Z
59PoWM63RN1nE/ECVfoJ4YbHOBB9v+jcIQs6m9Rb+/lOW4cj78jZGXtN15HLKyHPjsSlCbxIbWHE
8DQVXu+1z5gBQd/bWdULFDaZxKTALnMWGtQwb0iX9n7GMTW/dVOQN9ToCVTRxPGz1XNQ56fIPXbP
N+UQFg6Lw2smUQDd5tml+XYB47dvKpx07GilVEKo8ay4CeAMVq2Mkl0vQ2/q5pNszdHrJNhwldSN
OyKujSxLG5/KeO7aME09wmGw2jP1Zl/TXS2pZHKoHEpFDDBIijqAZWuu8DY2/5pjUC/3eQ6Ey6cS
9vqSd9RNOU4rn6457jqpsv5dlcVwmbZzXVXBNeBcYN9ETYljaRaPDD9ursVJ+LPzOZq5L9itLwYQ
iSi/g97RAGyAZ5bEeVvUTab6OrYHOj9PyFo04lJIztiUQBU/54S6Jz/GiaPvFiyGegTbaRoXRdxP
rsadi3cSbQiLsVXAMW/UudqEuzZbkHOsXAkRcJUmH/HFpgeQfVlZS5qN8+9XHlmflTy9NCYIrGWm
G1xSH+ZheHaodvfzgm5mJ8zvRHNGCUggb+DAfPOKtdZwqXv0FDoBN5yKtfdq0ZYNQwABqZEUlvCV
BfTkuF6LMRiefqjq7dIWQU6wKZeeOdNweLkcUpLPUKR2J4KnyCeCGMdC79Mmfk95tUYKpB6LL/0j
0JLcbLU9W1f7uqhhjmmf6bOYm6HTONFuN8aySBnSe4h2FyzfGNPvvxe0kgbbbs2nHxufPGLZpgMv
XMKihGHrkmiSQZO0Cz8mZMr8n41LtaRMCVsKQjbh681PxfW7YmFj9rvR7eKpTSxrlK17yabTS6HH
4h2+teQVfHpJh1iReXQo38lGgcihHePSxpRpykjokzrMN7yJhF7vVHoM7TmeYBv11K2tK54yYlBx
1uWgYhXG4feKzpGsskQtLQh55pssFsJzvdbl9o7CW6B5iXQSk/6MBBPat2cXKEGA8D1bBv/D1nQk
d3lhpFdR32+CFcrMTHP1TKQh1+fjY5FpXBNzWsYD1In4rPlrmG8IswCBQKFsOzOWcKhSZY1tAxRq
qN7z9JXpQ+5Egzmpzyzlt8V5eVoeHEGTVmx71d154Yf95QHWCHvhcgeMGdzLBRBLm66qHrum0H9c
ipq2NU6tbRgpv7YXTbMLIprmmiGP/YW70SGG6hP8yrRFsdgRWYQM5vIWeyjrzzafqHEk+rd8kvkQ
aYIIdOV4nEZPYS5XZJddAWPqLntibkNPEGoKXCTylIQwhMkswfsDnA4rRf45uWm9teR7dv9ic4SK
q5H9wCLrio4TbK7UiZXvfO3trdOZdAivRQzqpugHdH8B0iBtUmQsIGoc4Pqb5oz7j+PbPS5SzNC0
LsuwpEIKBzOJzgCPVbAFf94a1X1FyWgbzO8k6UfVGvHPgkhMfqI+2M39AAXTcipRB+6T6KUCpBlS
DpUXP9Lc5cvaNQYT3gh0VpImmbdjI1GqidrwyauWLXboQIt4EVZHUOZoTQr6ruIAlQeU+p+XVAHx
dhzIq4XdfmgZOhtu5G/9S9GYBZ/4v7Z2yfiEWd25xBFPVtNFqVi16qnwMinsCoVcWSfpC7kntVDX
0loj6GYSrvqNd7KfKVhVeJrfG6DajQyD8FkzJTg7nnZO6jE5IxqcdYT5ebEQNAuui5v5SbScVaxu
C1naykOzaBt95BA1Z2jz1lA6KWfuni8FJmD3i+nNeiMyQYJTlc4BWwlZCpeWv93hch4hYE8mv8vQ
w72CrCO8hTmFVDZCGQdMpv9A6LwMk4NuLYnkEm+w7Q0gkVf00rcL2KOcPwgmC08OiqdzfaElvwv5
hGB95WZqGIspwIyNR01TNILn+UfhDiYLmLnWi34CdzjcTJPUKnYkI98uFy1na1XHmCftnb02aPQ1
BsR/XKMm26JlG/L3qLtphgzF0FY8W11AigbVfu64Lo8sPQiuUZzemvs/y3n0VtOSVr25ZqK4Ti/b
HRhnfc/jCQVYk2s4nfAKyScd2nd4CerxC6haEoRBUyPFW8NRTNtvqtoxmrFPIe0FYV4GOrmJ5BF0
BptIbMCuxSLMMiZI0bcEgxgtPpd5O4Su/nxjZMYaHrQs8Eoglv3zTcDbxGqplQE5iFamzrg3pUM0
SJ6Toxc6RcgkPWt9tpfW3H9D20Gej5CvA2Knou9EJBzMHexX36pzyJYbA7ZzPBm6LV83QZX+SKpX
9T3Ip+XhVVz0/Qq6tfqkDmV4yFOIYXOd1qYlTw/suf4IPddO44HoHmj4RMp9JRs9gcuBuqAM5Vvy
1ChFWRTfNyJEreR8tTfmslGrI2+v0btG0TMibeRAyjpgKKwUU7aLVBE/RRJcI2Iq+vqdUcJIID7+
hWo6EnPZ/8bx5NpkacWBx6hBeQjn9hD6YcRYmnCpujN6HK11rwuKYLI4/tt8KYNXAUtBcLLjKU01
4Ajj9Rzn6LPAIGVL6FdxBDdfkz+mFeBCIQKIjQRb8oHCTLdPSOe9QQfcnc1CB262+tgVM5jPsvLT
KEmCeh+atYHVAjefyvsMn05Qpp5nnQaA5yuF0TEnbFBhVAAu2q3avc6pA8kjxq/Em5uVjn/Cscc2
/AFBk4qSZJKwKa/59Ae+U/lCDwgtHNJU0vcW7hf/3CdRmSwuFpmnKiMVgYHpHQqGKzCyGptyvP7D
kp4sHf/m/i56Bk/wI//wb2GscnAmFdkdh++MmG1WJRFDDorGojPYynI/Nrl452qt4Rlj+FFHhCF1
MAaR2MtrehyLdkynLXjeq3eo7HNnLE72J51wTjYgzxEbuM8cSsE/nRMeT0VQuaGBgvPVIZg48UPE
A2fnHg+i3DYIG+ztmWJ5bCeiaX3OSAOs6HFwRh5ehDRK5uK0vufzr5rpvcrIkS7r9a1b+Eus1Lvy
Bss7r6Ea1IGNWj10fuKuPYgUzczjMugyfJZOL2xazZpxnFAsVvy9iQf4phRx3pr07LTBuiZTR2nd
OZ1Y+ih/usD2orMfGu59wpH3itLhzdSB/JkN3wRamN2lMY9SyQrG6CiE2En0nV7KU4MFdzNsFfAF
wYVSUbN3tMn/zrtVZyCT5IQG0axZE/wNGtfK4ZOrXwgbyoXoKhRjwWWO1S5vCRYTac9451t97v63
sM6ofhUMfuR7AP2pns1WfWdy2pJaavgSyHJBG/IfxW9ctqBqKTp075neekQb9FIWG+ffxEDFoDa7
I9zw/w7iLkt2lunPLteIKa3G/jUEubvm5p/AKNZpkRbNVum8ABIOtgynCslxyGHqOR94k2mdXU79
IW4TtuSUXGxta7WGqN8NGfqINDcn6zzBd2zClGGjpZo3uojza4T+lq067uaIS4o9o3ijMz/IMEMw
UEGSsHiiscnmjlU8JN46E+kFgW0xj7ZhW1nSI0BGOOGUGq9EmuUN+XrrP8E77ZxgJF5Npw9Uc0mZ
bRx5KO42AUxlHkDBGb0uAsThJYM8RYmIZ1djKxsVTH1P5p+A7J1lNSJywBDSoXZCypgWjGJVK4zm
uArOYxFFKWLmGaFOyzMx9FVDzvNa4IrxfzLDeWpds2yjF0E9ISfxPSnbp7jnk239mDvNhqFRJ6Le
VOCdoeqFuZtgG5r988P1MlqJHKAmbBNwqR3CnXaNbslnvAtwdGQuNo6Qdh68dp4pdEFOB6b2xvMF
lvgpqVWj0T+BSJIgrhskSopP7uN1pmSSThpdr2cVb6hwx6cRVLnuHoeH8eJGmSstiNK6mjkwhs2Y
BjB3TRJd0E0tGZRaCjt0nkzLnJE2lDnAiGH4VRC+G88+UI5yee1i7fuM5xdmC98ySmw36MraIcYN
tRSqf+CMv4dJ7o9rq6f4exoZF2tcNVFCrnmRNwfid8S8RyVXBQGFRVYLe5w+cSrUnGq+MiwGFG6w
IS9qTRCUji2kYrmjkMpRxHompTX0D71q5rEChTUymDt34Ksv1eUe7/E6/exZtT/d4v3hgSjV0Xut
Hf7+g8PdfaSEVebsuZNSL+RyfowHOBFHtzDB/oDiwV2BlCRJxKiQamlQbq5BFSrH5kfndx+1uEbA
oO3A1gVi9jdgntyWrgO7kFgjy33GxhsNW+G89CyXA2rx3TU77hdkZhZmX9e40RSKhQuZFNl0f7br
+eH1CTycaHyQr5yp+KvNyhX2oZTkHR/PWbHGulJMlzsXHiiTWrlqWWulcT2IPgeqCvAV01XghPEJ
qmy26LowI8PwEc/s9CDCXChARgkiL0XsRjsf1Sir1t+q3WioNfxGMDzHGP1ncoLXtN8xJPq4N/22
5aIs8Hqsh7XP32Wpq1nh8Lv6GIH0JDUE/ujKZ5p5z+GGWmeaQf8rA/gR8WC4vg2M9UCcNxTG9Q4V
Q3bjYfvNGiCgAH+5TCakwo/1PcbAvV+zwer18tmU0fSI+rEilMh4Jk/j2kqVzHRduJCsl50eIRRy
HEc/Bmo8G/b1DQOwKqXSONnlErQe7MF+QagKs43OOG+GX5ecT4Fuowad9RhOQt0C6XMFb6XpS4Mm
6dMl4okjuaagIoMqZG54d6/UQzTeRczHRj1tlKUKnbxO7BZREK2PI3QbZa8yRSa2zqTiF7l2M11x
tZODP5JzCnaBHTtnruYCHXp1itrZAz/5wWJxfnOY5yFeltGmdlPpJFlUDQKWo2kuTqRVp8X/cEiI
luLxmELM2ZC7NAd0rUOlK7PDrxJbvQYmTlVVlcZUBA7yW59CBqc2/Opzw/gt9s0zw+gE8K9bQX7k
a/XmJsq3VMnOomev19/+yumrCY+YYsEwKGzuhfe9pwX3tPF4fuphdIqUqNRbn3f4fVuQwRwuujvC
NDI6nliiflqd6likn2yFOCgj5Yf+gRanFrY3oT8kpDyVN/paOXQy3AP6UIKwCYhBU0yaSMV04I3a
Jsy4C6SFQSWTuof3BiVbzyd/nPoGtlG3TyLtq5x7GIFc0rLeBBY6jRqWUMWqoySZXtpVRnSta30C
+HoKaPKBuHJK6YOPCppfY4VjPJxGcmKthhv6jaIsC/XoddvF6HcohgX8TJ7dS6OPjrOy5zgFn83r
zItJ++0ifhMMqDOsrYu/LKBJE/xgXTF9n7iPoyLQ6nBxKf1KPejmEA9hXjq4W1HzlYANTd+Mzg+S
rBfqOSCDthuuKvVmBaQBOSMtajq03i5u7BK6KLQIimXDRDl9Sm5PUbFJHquTBVc147mshVOTRw54
iw9TISoYVYyczr7libY48iN6CH0p8J6wo+ZHhEesJe7KHmMUvjN/Aob3PWpjOhQ6oh6dl4QDnWmm
hoTUlR9HM5j3SoYKouT/gUhd2XjrXmRtP1W+Xoshwb8EuOghEqqk04FuZ0SA4PRF3FtVcJBgDLkM
YySWr2w33tsrtMnLdTduc6MDTxzvest5HuoEaA1ijEwrrSaGKargoRZWe4YZnGXMB0NylQ1yIw1H
EnlXzE8Kd97cU86ynSAAUanqg0KB/lmn3zSCFlj4GWHv9yiz7BsSHT0gzzxF1c3Ypv1OjJQq5c3M
4HnXnbJS6m44dtRapwBjUTpfYOpwk2guIjVsSFXmWjeuOyCB8l9z/dRFVujp/35TXP7QafICSmVi
uJX4/AGidT71oqMm/Oi7equHZovE1ap47pFnSMlCtOXpDMEcER1rCjEfVTmJlW8hrYYfqsoaQwbH
/2cYolSxM5bV7LbZzx/A3P+Ts+qfTkxwPmT/hhFx6tT5LdPTsPd90sja1WUqVOR7Mq7ZWv5pJP9B
ExFFUUiJR3e70JykxeZTN3cwEWc/S2RiLevaqVFXp/Jjbz4aKhJA66iMhTCW+yvrWsW3DewIgjz9
ZlXbhtTWHlWGLAslPkQCem5YBZXIu9qCu7S9+shUoVLCZTGWBoEuKcaqEfYAk2wa0jO2JU6nWVOG
XR9SSngQ/NijoGLbOzFtqHDANI/rn17l9uUPm1h+yFfgWv7Cc9c9XYAT4pAGLCz64rHoALkZz3e4
Jzy7ZtG+HQiXPb7As6gZszJ5SvAaUoRffqg6X/RgRKzSrkx+HjitahQl57+sm3d/h9Eee7x1tJ/E
MblHBSBBDdXnCfq7MF0G9s5llypRg5O3/ygb6etjYYqEgra8+GqwWsgT/sIa0YZH7s8AlSlfy3np
TOw9Cfbh1TybmPQCyK5PNUn7Ih5pyVciyaMCRG8m+ZJsJlfOevCHEXt2GGzNuxq8JFKEb889TWLW
eApFmiF2logndFBoAbu6gbgKWcaxoo2py8UBwmZ/41WxLJ/cjvABOFCiAk15fcPH6Gc9UQ1xhN41
GMuM2OgdeoEdcVPnlptUresci+DQQN7NaHcTxZoyVi3xkQk1wOFe+985Aql2Kdvk2wLJU7l/1qLI
a5G2mMqJalSV52OkPiLgBC5vEPXWP8FsxstBrIPK9G+k07y0qG8vn/kKwP0psAgS2/VpQW1D9M+7
+/fF7/3SEp+HmkoHJdczoMIzTM1KcctuPI17cFlM9zRZ954Tc+CZfkynVbHyhbJxjneJPXy2f6q5
5K9/iFBb64/XZCmp6mZE+IhhAtTDUNkcsEk/NAwvM2vEHuNePPiOgA3bAV9D2lGEx9fkNWzsk29Z
prN7dH7K0poX68Z7u0cRLHGNpI/otlQffVEBl6BR05sCR2raAtaUKrNTMxZDZlhIYs20khzFMWge
jSbXALoUNMXPRWm50k/G785SbfO41ROYecClyOxV4phKLVukjAVW7JhS9PPT13ObtTeL5ujtA3BM
ur/SGtma7untqJVxReaA3qPBBGZV+01ssUX8pNzD0GHhLIP+eVReVXkULZFuG/fIIgL0CTfqyVN9
mZoExuWSVjFCKeIDAIUIA47lIXRWZHrtDaTpmoh4wHZel9+munU403rmzbxowTPjYVJqBtx0osb7
ybIrkTpGCvyr22w6OYqGorntJcZoZShCaX4rLzUy4PAKRDD6BTHLPbmSCveLwlM+6xbNV6HDT4oP
IE8OlkrG9H75e+WmfO3eNO8iZ93CJnUceSmIXcdwdmO+oDVnx8x9az8LW7UwwThjNn65CqmNVnxq
HiMoSaX8R3lfpQ0yB96xwLuLzIR6PNsE2Rn9PtvuMtLLwcEEsJnsgJkZKqFVJZ+DqUSVYgf2KbpO
cPVM1wS2GAWN2Jtl2ZkuO6dI/ps+QYw4lcLoKrnEIRP8qKj3j7ikGhiul84lHVPBIEnsBbMzy2AA
fU3EIsRMX+U5NmS2w1N42ET9pRsMqDuDRVhg0Kby9wDrdJJaaqhWp05+mbvIGuCTFB1GeEsU9gFj
UOaFR7zmkZrzaAWsiJ39adlNWabSxXVzlI/e0T017kuv031qdxdNs/0Cjm80MEed/V5FTbCl1i6U
LIR6kupfZfKGivB0HIRXrkLxYZBKfH27CIHb3vRnXg0NseazN+m71smOqz5l60sEjS2K8NLbZsWR
nsGfvAS7ocGUb6NzyX9wMomZ1oxDgjdDispR4UiTsi/0InA4Vkvym4VichgMOf+KzA/cdgngQhAo
Iw9nsLm17PO7ECH9TgKmvOkGyNMcJ3osy3pfvB5ujc3jRbbSVh+0yXOhe0S8ozqEwJLtZn7fi/8t
swiM4qtHDu0DtfmO9mtIwJHqe0RW3svTj+mvSTJTUFprCh1cHFVpa2iVi4I1emf5d8WYw0koQpni
PU5Pm2G+UJIR+EC86hU+FCqGkZ939kEqANlmZz0IUf6xP49jdWlpMfETRzPnrPvljw39HLUNlhT6
s3xJqAsD5HaE0QKiim6RBpxXHagbt2tdGLuZLKtrvJMZWO2PWCh/644i2Co9KFOigtBqhRHPy8W4
9x83gAxUnTt8l9ArhB7xGGsklDDwrHNxqeZw+fSKVQb6JQbU378utgRx1WjqhA6/gneY8FcxkP1S
mHyhtk2+mFSCL1I5/8Spq+dX3GkSTrLwkTybqFRgJPmDpnOOcp1RvjWA1x7MSxcGXaoDvcKGFgvF
rCyFkbo0vzJBsPODuuZhn9I+JFJyMjutijoovpt2HsDtW7Ck5aCbqbPTW1V0fGe4CmXDVCxNkLbZ
dzSq56CtlCZDxQa0x5nAYTcFh/3BY9lQ0hzVgF7+JtE0SJ9JqnpNkJasRNmB/515hNHr2+3qSFWd
ERJyVjow39lI7GKoSz09RwL/L1Ooz04fUy8/xEMNVGBAixcrPixXT8M9o8hs49s7XGjD7c7aRwUi
d5ODJG+3uXevmpivjLFn5JpErb8eOfxLCe7meUCtupuyoCJr9chV85OmSf31Zvx3HOxLVZNhHFFB
8l6Lrl9gT6LOyRzx6MrQa2XkZ1NG9sAmpXk3Zw9JK2JTlspJ7muvce8vToUAJMWa6x+OSWmWg7pJ
j8dMXRuLrPEsfvJKiOKFgbRMnRaBukNj8t6Tr46GEr07QROcEs1PJL6sMuAqeR6UhHTIH4qMBhu6
dpLYOD2cNEmSwu2CUmVviDHmf0eMJCZ7DA24CTCn4RSHmE61TmjFBYfiecHC9e/PoIfgyZZIS6XD
tBTgp5tJGzK7sY40IBAkoRaBa4kvF6FWQ+h3jcb5wvijFSPnpw7PUA6J3acXhd+O6bOWBMf9lE7A
cGkjUlG59Ns4hwWuvjxiCqonNf9YWysETe+J6WO89OokMQjx67hIgzM/tb73euC2YGw8lPdt5Jqo
oXhY6wUUlbsu98Qzytu5jF2+nS9B+9O7qJ6zJbSl6oQPpRQy4c82hSAeOCw02uu2qohOgRxnjiHK
tIFPtT9Nnj7psok8fxYvacD1mNv9/h3+8RTcBp8YBFwhKjJu6+gUZ0mWo1gaERLfbWDeJ1XTk9+q
nvwgAoUzRocLdHcGdt2eSHxAsI5zmJ02vWcsE+5e9GsFt9PDpvfOLbvKvQRwZ231U9Pcr04z54E6
JJ2K8TMWiJwJC0AKTM2Vev1DOjYD7ThdwMQA9jJXrgaOakacsvPReGvcG+1sYxPlleTVlPviaVVL
4S8v9s1eBG6rGawLi10AM8kE1gQ2htYv/W8OX9ye1ZKUMAo0jQCnC2yfdqS1HNIi5lKFBBX0ey5G
69T1fCplqoqj+/Md48/GUCRk/53rmy2j1byEJf7/RaolCKkzoW79fZTPpuGlUpu1ktZOyfyz1E01
EjYzNbqEv7TxzrLJRzJr8FV4PsJO15Jrmt0nidIbHATLRS+sgGe3C48aAekeQouLjp6O0mcyRFNM
LFLTlb8wrpxzdPt623aiv8SIaKtRp8i1AKfnWOznaiIeseKt32pFXj4KrhtZGW+FlFV2IgXNSyqt
l4Imu9f9osDnYUP2afGhdLu0tnNASAQhUOQ9W3VoC/0wImVsFYZpuD2HykGGFG5BaWPgeKGVXyRL
bms3wbacY3RnEed8DGasDvgTqmoyUiLTNovq6aXg4jOYrChhlslZlSXf7ymiytxOxnb8ReeO9eNo
By3s2iOrcSQW1q+OHLxtMk482RP81/F6phhgkGIkOBRcp+IRZ3u26hNooOdFXvO0bc2PPa2U8SW2
ftiBursnucNYrsmwMj825sJnbqUZuMooJLmoCTS58n5/Om2JPJy+0TctBbsH9EdE3dK2iQEUWtH8
Ek4DtOY9qsYm7r4bNpLYuCGaf5l8CsdTRqIl0UdN4lB721ghjDPUxSHLWFEsLdAFSdcvk/vn1Ay5
zRpNoNvCGARsdlH+9v3Ya/2o1rT+o9UZi+aTF0oSqUCfbdWZPy7OcCOMv8MEdkTRp6IpbMkRIhjY
DKssjJh1EX75Bf6B5uf6Q9xg0FWMzlTurz06av9pIT5DIfd8OFubaNMuAaeIaMdT2N8wOwnIzu4k
BSBUfEmDQwvhzJyhvHHkXWXB/3qSd8lxTuJqMIQr+nUToMai8qB5zz9I36rgznK92kiOXujJmODs
qeZuMO3jSxdjuYv7n5Bb8bds3rVdSJ5p/kqq/hXNbke0Ek7KhCsZGfIuHXlnzQrm/96W6Q9j+m/k
FO3AMQJc9nkQJ4PQ6ce28H56GrdMk6aPoQobXdjJd34Z6hpc9Smx5e15Eh4B8mVeEjDiIGiD8lqv
ZqKL7esmcUSR+BB4yNh1N1hIq4zRrzh9RF/I5Y8/NiXplQa9fveLxB8GDRIuJ/+b8u4MbKeRLZGb
hGpULWY+OKhOByr3UEBQQTbTqc5NJtM0+eLDMBXOlPBucN/0EL55wtam0OVTJUA3Z8GysV8C5MGO
1qF3su3T/iotf4+7DYBOE3TSZ1oCEBCVDV0TOfxkIXrAlFWezcZGGhHK29DBqeY7sMrBOVsKJKjV
CsUlR+E2kWgePY0Xdk0te1Yje63pjheP/LVDcHsFl3jgxOrycQPt/nHVmU7SgflzhQnggm23tfoR
MVa4jSW0iLDB1jw1nXxkwkUjDevtlG4apJgL9TDz494+wR7ashLmWGdhk9n+cVCK/v2lo/QGzpXg
wlsMB3/icVAjj39n0Sr6n12naTZ+gWO2JS+nO2okAA9nXumy9mFeg/yjP3nF961P1Q5usuH1nCDr
lqYhAHctEg+GhWVOToRa2lcN1ZRiFXTUYu0SG2WtEvpiNStRdAUk9k563nVwBLiX4eosfAejRe6H
1NjzFk74yLGKZivmagA8uOvlSQS30I3F7KMB1vaS5vHRZEFCHS706s7+6vvls0Ko3gxuFqrTFUaY
WinJ/rqrCUvScvMWuLRcKgw2Lffi8hFiepPcLNQyZ5LiAerpfreJqjB/bkcbdFu3qs1ssffuDWvA
VMhikL4KAxP8oUv3UU9qd5gjJ5UNjkGvLRyPY86CKwU8YT3t0P6vFCo4JoZfGYxeJb6GV0AYNsHN
afreXqrpCO1QUQYehRVZNZtPkAWAZtRzW8D19Db0LGt73OOesGDUU6X2Qtj5YCMLli9nRGJdH7Q4
dSgob8CaSPdS8a+3E72YIRlXILjRj55If8LxB3lu6gVMfTrdQo2KY7fEeV43F+C5r61EB6HjegQN
0vDBRO8/JBfPa3GH7NOyUgHjBTBz+THwwh8KWLwyCBc5x0VUzsfcOX+Z4shK4QtlYPzhQOaBWZ2i
JvR9/FaJbTrH8Y4g2qdEFnUggVNa8YhUt86PypaK8ueCav0UBfPOpYCg31lAC57pKZ0JVIwGCZWD
FCjIbpJpTqqmURBma3HZxJo9Bf0irRN33mKPGAVLAkzNh2Ahj7aYLOlBFW8dmPBXdPEH826ZR4Df
sX2ITX7MouLNDY9ID8eHzmGh7+6WTQxYLoDtEY2lwpAgY/XVgvWSMmgO3XFiGMzYsmlaCJihu7dI
ai98Cf4PkiDaH6nD+zKjEBePVNwuKs6lYEfG97qPk5vxZjhqwibfwbqMvBHRw4har24bEXXfSMHy
ls/ZwacEUu6+cAqKo7avFYkjTyF3epWGzQ3DBnYAuZgjBGhuiRtW2uBT6P/IuJFXaEEK4+Z/xkDV
nFvtyU0kUm+l5u3zaGoBTA7ugOkIHNMPPGMiQn/I2s5Rujr5PaGgRfCJ7Ym7qHPmEP5DyVkH1lgi
Q/vFoI+zvgXsZBLPrmIoK7tIzAeodF9S9DSlxkuo+9tw3ZoRyXvPeOzK3HkDyt64xF5bKSD19mhb
bsbUmS1EcrATZ4q1zs7EI8aZp506AHQUdeob2/z+AWe2K6DZuyziKwMvh1mPG5QorwcjrDjQm0RW
e9f45R3arB2rBOljrOtBUVAMqPC4eSj7DFXFgU8cCIXw4I2dG4L8xHFyKjwj41BeO08etlhztcmU
kJ62bLwmiZgeuVWc3+8TqNVJKmU8cA9UfMtwdIwKbDbTgpnzw/8y43YZDjDjose9A9jccZFwqou2
xfDyP+LhvJPNQ2W1DKNvOy08t5l5EY97OAZvDiCRjGQ+G3ehcX+jfdm0mNVASUTAwLlQwNU8ffeC
cgZ1so9T/8EWul+iMUT8Rv4Ywr0gbK2qJTW/AOVRrGiZZNKnktu6EsK0G1v3xuIksLTeo4QnoyNG
Rfed6lNF7fUvg196JDVVMqEc8DuZDiC+HiPqEyvAiiyarrcD6EC5hEW2br5c3IY0g9m6Vgqr0wrK
9W7LQQcYAI3uAwVoeSwj9bXliVlrWOGt9UtxM1Rf2c28sXmdi59XSZnZ7oFisvFNqQE2eq7RnG5k
dRKymL1RYDOhNO0E1SOUeTFuM29yhsOWBdtDsoBE5sYjKbJFib7DdsPvamMp71/2SqkPXp56pjpl
WWeAkJZrJAfKluK670DWEHTcFScC5dOADIKZmqfS6pWZRz/keC2iewUMM1bAqfH3dx/lcT2D9qKJ
65+ejLWHmJnUbJQK+hCiATKB0cK7O4i8hq5dDlTqazDPYQ2bfcFgOHa0qtwS56nRXF8lO+uXVzBC
YVNWZ3SFppd3moRDWA8IGsQprFHN/BJXevLX4XH385Suh89ykxAjT4jZh8U/jPt07wic/yy1dxbf
0miVVHopA9BbJMMrumHfx8KXoXw+ppdHnbc9qnLCi7fMewi64+jM6+zWNHRbaGT8MSxAyM2dcNvT
TeR/+5pWBA8Szua74rDyLXLo37N8hFkqyWc6P168LXgH04SuuY/Z8wuJP4vM+k1BDgClkaHOpwGJ
SQVij9psHRBImSZ2AdX2VjocEHlWcr2H+4AsxjpEd/shjyCYMzeLspDEDK0WA0PeqBI89+B5XykF
bgOOJ33fm55MDDFxS7ksCjN+eE60sHg53NFv+hyp53+KqupBAOpXMwtyXiBAVXQkIpZtb9rLaCF0
7zCAktQ+jhN6Ip1ygOlO5gHTNGV0SXc4FtUjBjZ1n3OtT40T2IsHqSTJTw0RBzAT2b/pRhGPgPcP
uXGCYGgFgfmkSebZQuMOeU682Nq0/tH+KzNNQXBPoIGNA5WUKSZxHnPwuejDiJv85Nwgl/Faks/i
vLU8msRKvQxP2r9/FSHRvMYPPTPj8yQ8FpRKemH3s/hloKW0ZApuGGBv+4LVVggvShcCXcuy7p60
O5Nv+Ntp/8rD6suEkuQY81SDXR1bJnUbDFXFRjIh5IkisVoE74FxZHCezprNjvMWTrnPvUG1fWq0
FLQW+h2GBpkBMeRiVIZrlvocxo4WPVlAfihZZQKjK8B0mpgyFG61pDM5lh9b45C7z3G0YmEPssg9
+1yep4byZPoX/sWLyvRZzaJSfYvmdOvacKXhUtfGSJ4OEleevZt9V6LHmsyzBt1XNrboifdb6UEC
i6ICvVG1LrRE6UuPnB7k+8Xoioqc7Q6nb0oNKe65jslEaxYvaZTd6YNGsoeRsOKgrDA+914UPQrb
2mkETKcixlqSpJdVzYOeZgJpw8cwx8jXLulqJDiJDE9hgcPr0KLm/jzhU5utVhgSeswjbYnjBOSJ
YWw0roUluo0qnGckwB2uGEcyeoFa+1TPPPlF/BqeNfaJ/dJYM3m0FzjPnOcpSbdP/Tw0PtKkbQOP
5YBSH/T81pRX1y4+yusqjrN4S3T5H7oq5mBQDgSuUHaqjVlifuvXv/HrgIdb3pWD57nK5RCKOYtc
xzjTBKW2ytXkt9WLaC1FPO+iLlF16l9SCQ5pk+toAQAZe+U6UdLusdNZISX1EKveWnhcqDiYY5dE
uT7dCI85fg++jwLyxBP54OrXWr3KnWEzpTyb6UDH6xmAcrIXmxzWVoWInge1NH6Yt9pIakgmFJdq
xd4jY01r8JQv5c1P2hKZZdolmIxvffQ1yYnkpZuXP2+CwUOVQXU0wfKhp2i1WoTM4wKNZcuZqQcd
AuSznd5k/G81ajGgLzG9Z7qFDeXH41UbIEoH0fWYab5WtWmDDczRCtxFFVyugzGpam9LbpuISUuK
wU+N211l07m+LOe3gjFlvLazFM30g3WXaUSdXmI1PdX42EU6UM/gs1c+BWYT/ZHwSxIJzU/ApiBH
yN+b7214O8lTEjJFesekumUh/HgdVqNeL+Eo4TQq7GmIBXoZquTTJI1PDidA0fWNLsp0PgEVih8q
74s8MxV5s6EUUNjfwraRLNbeSofP+03sK32TQgX3Um+s7wkAEP19xtTiZ+kfnur/59ldRCOothhE
hL/bS6rfehaR1uodrXFodCMozfrzI88VaTQz22rBh/HMkdJ7HjfalrU0p8pKD2sw77L/VlXZs488
sDbmSdl2IoiKavQeb/7mc0dx2ff/m4Aztg4IVqcYT3Q8OIHdeNO1nuAqHGdFqoMFyQUXevb4Ipn/
Rs8bHSf8rwcFz4okgL3/XmjYSrdcd0o0oIxfEKg0ahq7QOfNUV2DetCh7CADbpRIt17FUwk2s7JE
SHxAkBL49ROV8wtYn1g+IspmHWbmURs3SHRZyLgXqZctBOW1nZAPtvCTRxR4sf7Ho0C1r4BBD0Bg
19l3JTHB7w9I2ToQPR7kM0dEj87gGwoskxZ4rvMKuzUdbTCbfjs/tvOIgjRCWtS3rheutG4EVAzM
OPU9m2CoN1Y3gbLDzyqelio6kjaJgJkdbzXG57fmkR4GTOjfLDRQPoLlwB/1se2ldqF1GSy1eWO6
nD4/D+NMH4s01+XrdPAkj6SNzrwG+3ukrKx0l0MvF+uHd5kBCBbRKznfaIe0AYknDboFZl2ccuyC
b1mIB4dcRfiyCqJgk1UN0UQVTKd5xRwvyjg1ME16cTNcP75fNAeImdwFHru7Csb7pXUWrz06ApJc
scjfVbvbxQgM90JD+tyGpcAuhenOUBwfLwJ/Nfz7LPxiCuocLW5DufHJRXx/1O1G8iC84ecZzwoI
i1TQfPkUMH5MUgMfZWDFf+6W5wlChxiTlK/5u5BJKIm+lj7JEwGFaMSFLhdim37JNVshQreSDFiR
6NPVHrdecnbD+nuku6ltrhraNgw4UzkKKpFUcYqmCoiHMCNhPA2tTq21jssAFA1v5UJvFj6ff+pD
2CZ3j+dddOakz2p4elOboYkSnVZLLuZrYWAs9UKXOD60A8zSyJWYMiDfj4Wy7JhJyH6Qv3aR5Khr
heMknsxlQeeklg1tkbEqbp4h9ZZvmOKNUcRjLzc3iGP2+F53jDU35/6Ih7qVow+kpvsWwwYKNpfc
kZiMnluK+8V0vLBmjVfVRcUfW6JPW7xCAQwD2K1Uk0eb6l19n0K5CMthsFCU8UlohYNRDPAzovpg
isgF6vagBO58YykPrDQZ3ermG2Ha5i2zf/V0N0lIDjyTGUpON6eamNFE2Ny7pYMqekuGkBASYhbJ
X1m6F/Sf7a5sR04dmqZLQWgc8qAJbuwOvvNhuBEWqI0kOPOzG5uRILFFHo3ky2/osoA7zDqakOZ2
VED7xL1XHzkpP7SEWVtsk/54fFjY4SdJYDSfOaDUrcuO9lFMsXnXLZZnCeeXKm4h9Mi7DZn9/txr
godgqKqKjnYyQOqh0dInP8fyFfUyDCgXoqgpd6QaezptobuBaEGYSxYzQn6dstfyIxWie1D+UAVS
OS9xef5bfoCUFEztdtewyujSnE5s/KdrLSPEB0D1nrr1aC7jGYoBK5UbVOPAND/uVeGXgg8wAu2E
BwJHB9u281bt+hfj1YIulhR8GMt+47grfXLVd1lm81XQ5uTVEGqqHGB3MwzQH1AJwzhsM27lJfeC
7cQcvbG44q3EqR0dfWip4Q3zIvG3UXojvR8Q4eEaSuqYMKa63Soevapwh1HFiKXeWeW/i7+0Ql2a
ETnciRr4rmdMobzXuf7bReOkEk9q5igRajX483F7RbgnMlX2AGmjNQwv4Pj5H3RRjqnkPQhSpCvV
2+t2U/1i22OjiWTYzQDy3wtByQKcxnzK1B+PPT/SN3PveBcCROG6IEwogT0iYJSRv9crl6sgEf9E
LtQ5GDP7Gdwna3NiNNlmJcn2De9MvYcua45BAl8jHF6je2KwL/68OaxjFcJEyyr0NmWykopE81+8
26GnmiPT+/CfVFwlQcpUhbYP2pmQrLliEZV7H3Pu2fNZbOuWAtLUWQad+wJiNNWoDD+BAXUcYeDc
32YrtBEYXmLCfZUBHOXfAqvRlj5emuQelYOz8gT/BvtiH/PA4v9zx4AZps9P+L8KNLQluhiRP+Cw
QN3qWY5LuULeSVZkgtkCp/pxUDNQJPkniTrvRj8PIDQxoilXSnL/Qg36tiBGvkI+GSraemDeC2Yv
7wo2wB8zhwp/icepBIg3b/lGee65/CvEA0eN3SDI0oy7T8ycV/l3SYdjQmUOkJJqTmmlfyOnzHCz
Usm3418c22FzoXhFETXSyYEmRuNkx+nlyYBioSRPL9cPll135Q2l/0VJpUJYMGhdqnNz9UZCRn6u
XGnr7nGX0a+C1wRbrAqIcG6x1l0SstDrLQaVVg2TWVyLeupuDjHBonAHbQ6WzsGESSYENom7azub
Fhlkkc7WPiKYdQz70yyut+xBKzpkKiOJyYBD5YQ4H/IjWlSvrJ4qvLUgjh+Swlg7qGEW4bww+bpq
psNU7imSVUJWTHNpqzsOUwAy9aEagryNDWxb1Sc2rxg6kEe49OZ34wRG/6WBgLrCliEb57ES/Faw
OL3yAI7Zs1qCxF7eUCiVzlKHKnHyl6lAyFxUexqbK3AKvnjgl7o7td5/YwWYolcaIXZlU5y4bUmJ
t/8OuTHIFEkPxdoXS1+kHJftTB5I5vfaRWv5EPSCGYnfvubYXqOXzc8PPGjboeB9oWdrdBmo7+1n
1KRQSzmE+o8fwhdaWPaB3XQEZM7CxuvfGPavhy8cvCgyXEmCPK47XMlJEM2LSfKKycnIpABlH2gZ
gVXut+aEthRlxF1QCTIJmMR7/YkUgy5OtDv22JgrY2QgAQtqM7r+jc9H6KqllQA5f7ErWSW+7DCz
XYL9I/rzr5guY1uC1nZ7uEhgp2yCbWtr80ew65eFsHwpbYxIvDW7K0Pf0RxNhTpGg0C/MFd2ij3g
PphxocH2wJ5Hx2HkRBq39Rt3NvqOIxnF6tU4BBBKVpQNFL6SWTtoOLbazuf7DC+uH7YqGFFTf8Uy
Wy5blUalbDgBTnR9naTUDOyXoOmDVyRyMhbVT0fPBwWhL4oFlOUy0O26u/lrmxkJEWA68PMfsSAC
jN17/DAJNOgc14wwkP6VB/g7Q89LhSe9Em0AL3YW+F8dV2TvSwEyOmzXx+He6LaqzdxY9OtGd9a7
7AvZNcoWTWHFcRMExFSN9wryIIQ4WK7XCQO5O8KHVbgtTK6AEX2rLp4E1ce5nwW/76FX2/tqOaBi
MqtcxaST2rq7Qqb0J6IC6su7Jcu6F6iyivHBWdfNQ5Wanqlnlt5fQ2581/Fao1QrnbO+Xb5E3WqF
bA9e94aS54AexMhSG6JQZ1v+n1zXty48WqMYHc4W9MnsrEfj6eHkHjYFjJibClnuacrzX15qdDwE
hCAn11oy7Onpq2qmaIgZ1rA2VTR/JDVZoMhhUrwVkJzAj5lKD1TA66jio5arrE/3//WR2mutX36Q
F5gKkxpZ+iEoGUZnRET1QaXFoyF5ce8XgiVk8XX3NYS9i7PZeS0wYKuODP179sT0Yx+hoJasZWyf
onUCTtYrzW0bFgT3QbeQHT36j0LJUK62wZ+OEupN7+F1Tz/W7+6Vc9KDGoj3P1cW/Tb4CjFE9YpC
+oYPADa60HiQeZBlb2vHMlZeCwJNv4BAfFeVl13vdKgQKzdi36ieAPLmN970S+YCtCMX16aFWguv
TYPlOw1eVv1eeMxX8RbnGvpu8GyZgWatUZUYHcgSulWIG/48aIXIDxS6j6DdxMvmUJRTU96KA5WX
iDX9MYjovJaPXoX7WC5IIOJjWCpwSicTv51AIVaphLhbyi17ViEbAa2lDHsyqTvDheyCNWDrfPSG
PBpF5Xb6E0dcuFxD+BSc3d1DSoxLvCb2nNA3veUKwZgdussnwD4Q68ynJzrcC+IU147Sz4Kpor8x
zqX2OEhFcpiPQ3RWFR0YOJdhxar220SA8+oDm3JdkvowV3bsAKjKoDr5cmryWQoIedvpxJZAozQh
aCKBp8slK2CojqufJLcYiUWQNvlY6aj4weCbCEPejl5ADUQ49D54OCtZ/zTphQ6YidkRA8E0IBf3
9rmVQJrD/UlCHLqc6YFYqZcxfmkBO/+jNVuInD51PvtsXkuT5CbUaoYqqveQvuh387H92my0PXEx
Kq37q3hzgvy52lxn7xoW6nPmpLasb6vfzH70KBmHsJrg4domBCN4bDP6NYjJAuccmJPqz6c8ZIdn
CYAaFtp84ZxfDvsfCgMz64GEVqydzNe+l52PQt6J8vgRB6QeQkzCuExgdBLFlPP5w8Nph9JOeUdL
r6kZoPMvvc5VZHqfmfi/wKOD2OFVVZ36xdlSMRcT8mUMHfrxrmKjAuPzMLCBob3PP1wQGfWz8LKy
7BsQuXPyTYQUjU2CY0IlQL0u0pIxAonuok4o+WY3N49EjXbJUeFsHdSpGM1S/wF/CfNyUDUG7Qbx
3/U3tm9KPx5YqPkb6nxdgjaOX/Xbl0AYeiJMH86HpUgUHMbZgdhPYxr9L1K6QX4UGQWE5oL/5gFA
VcJ0JhEUNHCMDGl3OjvukIL5t3BCeWd6R65eQ0KxIkpaSUwKXMRPw7ZG83fLGZwRKxQu/Cu05nu2
A+4aTRZH3v5vtE4jtIYiee/k8AEYPfyGNDC3wCdClpWhrJNmuuhrgmRygJC8caP1tTdJvZrZfVex
1jvOvCdcUAten7jXh4iMmGpWbQ8rKvl2QW5dAIyaMee59YCj7+j6x5W9h1Fr2T27AhADHB7Rc9FQ
1C/potuNrapDeeSSXytVgdVZAoS6KauPj6YB+NOR24iuxozb4r05sOISCxKiPcGN/WlDMGkx3MYm
asNbEQquqgD9ClYCTdRJPjiJlDI0gCPM2o5msiYsSUE5/p49erWqBy3p/mplYnzRsVjGMz2AKcMa
jjyz8OWDgfcaKVzWYFvtnX7zEuofpAwr5LdJZcb7IPGuMHbjcNdQsouElN+TVs4bdsrrixcuH6oU
wjW3y8Se+R6tLlg4WXzg0m8tWLGtVGM0tv987zCQtbQqxyY+HG4fjN1md6qhXh6iXfJAyous4fJn
ozqugsBx4xX04EIr6YF5DQ33Y02cxJXuAb0rk9UNAOHWmodUIwdZPEKUJdXzoYaHbIAfQAhgd1J6
ggBetr+kz9WWYYNBQXsfW8AyEaMQoT+LpNvfNbjkAJ5Yk5yb1N/ENywKdc5pDkMf0wkFyyKtMKqE
XLLp2aOw7lTrPBgZxdkvvAjBQZY5LsMobYuQXj8AeZXUfxLAZnXRgX3Ulwufp4ZrB5p9hLoqctE6
SD/k/wLwUeU2iKv9vpl6UqWoEaUS4AhaukrbkQnQreuTdvokTDg20DaMO/MgEswLwDUpetHn6pRf
JY5JKh+Nv+GbOdqYv7JOBdKqRlf+m5G2ThCKsdWlQ8qvSBv5K8ejf0PPNhF1nwYIMZI6LPAlNUbJ
MsM1g2ckW3PwbLpQUh5JIczd+5XRW3o8eQNwSPT0hd0ogcYlYVDwmTXhTY5T+CJoEFKDN+gAzcZj
Hu6zgDCG6WH37klv42yYunl4hqgv76Y0y+nb4KZhWrh1ntZnEQTzvSdG0CbKYl7yhGa+ssXNcRej
8IFffX9Dq295l9ymm4zu+3QFJ/JaV6N1U+htJMZ3Wk2dWAoF+k3T1dKtb96tZTjJ2Q25RWiow0mu
dzlNv4vEt46Vr8ZheZvuKpUubWklxHzKhJmORzYdk92TZjkjU/3inNGJQteFCt4ggwNx4Goydszi
9bLiZnlNpkjE2o95tjVquVIz8yS89jgN6qV9q9X45f+h0mEHTube0Qg8yU3oXGGCbICV3N9Ihidg
5wcPEK5DAafgOyXwyBkyNuoJNoAxw/cCLABAB46q5ZrIyXN6FNORYSKTLJgAjdQLQLRzeYJJ1jWU
REZ2o8NqUi7keItb+MTLf+L0aL0eeO5Q8rlIlOAzvY00v0T6E3j/s3BAP+3zk/8ls2Fxy06Aeg2C
P8ZoBtyS7KeqekFhObbSMlUm1BzdTW5i2vz13+WJWvF8/jfSZ1GkP0moadxMM5nNyX+qHNtWTq3h
orObGi/m6J6WLGMLBAxRwwkBY7QscgyqBB3P/8Xhp7XEGzi6UcNwB85K3xbAl7mqZk0H94Udc0gJ
wgsCo2EvAbRW9QDgWP2i1pZAidNoAGjzXXE0kfq1ia400Q+klGI4Hy9kkXuxQo0oIiDFPJbcTzwp
Veq69UcDREQM8velROmb3Waxa4ks3Cxn+c0x9GWD4w37JbiiLyXkMTdxUxsM7jyx7AN1sT/tgrOk
e3d7fQGebPCGtv5XTgTVkfUptLzSefb6bvWLjUUtVMPaUkFMt5AnFSm5dqv+p4Zlnwq9RMZRwoQX
OTXzP9XnWy/0oF+XRuvcEJMjFhL0GeduR1yN1DaoIKguxxrB/1JrsMSPJS8aIBdfV/a4xYxMeLwI
LHhtKNMUQksacVnJD/WuVVEUeNFUQSOsXqvEFSG9h6cMhIIVXMC02fdk6c8D8MDTd5FZakHM9i/1
pphoTgZBUcW0QdFpzRPEmq4Irjs7U+8b9kHYksaPb845DxsSfuhDDkzklbE+vvJbF/VwXLpJ2v9q
g51K5yS8CsTtb3VeSQg3j64qYekQu8lcw/ilI7RpVb+scGSZl6zQVo3Kq5yHzAWm6+Dj+aPFbg08
I9q+a8JCgdEudgFCGEOXgNGq2fxnoc0zmKW9E+A+zzTrAle8+1hz7vCiycLCZC58pXM1CIuHi4iL
ZPPJxktWXUfXKUGvYhvFNrNtRy7BbfwpwXnilXlhbf1vi4D0TLs4vZYOCaWJbY1OU5T3y+0RaATn
cHIQuU0gdzovXe2LXGExyzur9ASifW+UOrHnh7cOHgCvGFH1dYCXK48LouVyYGcDcjBB2MuygdNI
YKr/Lta6HOn4d0Z9o06oUWUx8ASv6xdQUwEEH9Hsxx+azwS/WywKNQjDzT+Pu2Oa/XYDhSPeOge3
xd2ZAcQTfnzPOWbFwL4F5WuTmncLZcXTMUeDrLcmlE/SCxijmvWdAS5Qu75A8kU7P6LNWFPmJRbt
CgQfagVkWk38jg/O6naCmx+CVdIlkhsiGQq5UmEoThIeko73bNDzd81lHV4ZzWeZz8lJUgssohvp
7fg2X5nhbXeXVkYx1oQxg6l5Tp9hC+e12dW0crDWvViLCM/GtRJ7npwbAlMqR6t3akMR7sVHyWf1
KNXxDN3q/dm8EheSQ23mJN3NYdZq3Wty1JM/fpAc8nQ0HORdXTa2UHtK7+1SjcrrJ2+vbJfyqLoP
D5gjxqBXdfm/QVBGuxK04NJku4YC6o3fjb7XDhQY6bu8Muj8pdt0b/Yl95K3diUWaNNgkE0WrEJh
sY0SqjrpXZFobYmQuiRPqyR+QeEdUd3CngLriOjBHJiUKwQt52r/PQL/GgeZQJkPP6NpSpTawu3C
lpvjkUxRJic5GCpfrD0CZxSb93R4tNo0l1pDiqAHIrAzMKzYdwHzF3xmRzYpLkLtgyUemg4/8ZOg
o7SjKn4sz+nNxjXVQhGPc9SRrjH6mxOSxAB2qaIvhJ+c4Fs73NLujkhpif3jQPMAbjynkxkUrPgo
1SWuGFtgaCI2wlvQvMkvYQSDL7IC9epDSdIZyryap/q8Ksr1iVpF7Op59kCRsC4fL0duIZDQcjSW
rU8GXei0Zx6wksysuIB32+pvJvRX+flL+rA7mp7tBdYMp4fBUfl4mHO223F2AxpdxxbqvNszZ9jJ
D8JwMQBJqeSWdjfgYywaqxKKAe6uiA+yFTUy8qYnQ9iwGUCkF+D+wps/e0cSUNq8Ff+xLXCGr0jW
aVa6r8v9qFYW9tOC/JYGiLY8iMQ/WsoKBjqd3Il8YKUxR7o7bCakjA21SlOzaByJsRovQWFigTQr
yRgOBAsc+sEg+WhheXmqWcSzTSwp8Z7FJEWFA0ra78tZ8Z1Jabz1NOKghpDnCbpWlbwMKUydMSE5
0qGeW0LfVrweomg44HQnGoYZeHCPnSGhAgLuuf4SqhyIC56dRTyNri0N2uHlNJzKsI3dvBORBeNW
jLebl36O4TWB/Fn2oeKt0KtIW0aEQ2e9y5B62vYQeWPiEcLLcfgwFAjhK+FiOdhZoXOAWEGaGrbJ
iZI416YCfhs+e6LmlL8Xvk/KTWpA/mRsjCLhg2XD7uIzYJFrzdO3YR8g+XIN59UuzVkSwb7iVGM0
AYZJkSxXfFJb6kxsHGxEn4F2NF0W6UUk4bxZ/IDFu5bN8tNhiRQqF39NFubzhBIHXDb/n7dweSd1
KA7pZlKrwgRDwK46+YF/TxjJWuOuvj3rHFzKztKrt6Rweb0rH8IT+dR/P2YPNaP3977vI7wXeQAp
JGBqNNNqa5yN/PU67Ov2z1O0v7oHnMdj8CnxsPw9yxQrXErPc8oC+7dfcKQSdbXJwjI6sKG+0tjo
jRAi0GkQBwV4viGff/gHcDoG7WynurnvkFE3Odz8egotUZR4297gQEm6UH0yv+ByNYgJ+RSZemEH
jLm3NI+4h3vhvwNXVaI28ij+zsZimhcPiBW9d3Z7z0JAjn5ySnbFUXlzgDjYxDBS3+K9CQA9TMyS
3fRGMyXyA5+p0S3bCMeP2y/Vc22I9S9HGSWVIhuJ4ofgm4AqHlWpEoGxCD2Spz5fG1wVDVQjcNqD
6hhSVsUP3swqlgGK+7O8RuS+Bwo+U4oAQcKlUKYP+kpJ3KoxF4zHuPs+NSlA22NgCL8q2GLEjRLG
YLrmQ1QL/jAv7ttUjqmJWQ1oJWTR0kFP3dDhrkTtGyx+wfhAUwyxoIJRzMedYkVqxAz86elBPytG
bPX6ABF/N+8YH/57plwv/AT8YfKopX2FGQWg3ZvzghQJK+pFIxrOEmXJNpkXhlQ+kChgmVGPmtJd
Pf56qdlc7UAgteo6pipEHsi9LXNW86MLyaM/M+ypM6vwvs2RPbNP9UqHGJ887XyaQLp7mnx0RkhT
yVG8RLHYrelxqQxLheghBnFUA43nb3iIZg6kc1C0+zkC9YpDdQX/3PQH7DAnXZ96Y6w+r3kjmO4W
bI2iVCw9qiE7XvGzYi9SheT2vmQsIggl3IOSk/PawVLqg+DoPF6BYExvjzIwyh/ooUhgXNqKFI3w
Dl+FI6eg7evis4exuLv2GmcFZj0KaTOvW054kSPWixocyPu7okX5K1Rqf2II1sFMte3MQF25nllT
OnfHFTsSpjNyi4z6CXDPClIceore1fSGFAKNaSnH3hAp7Dj7dSl4ZdfcyRT3Y60mg574Pxb5uM76
F/z0Z6iI6to/0dQKHi5tEbqVmFEDy+yriXr8ZGPBxdsq0ZaVBV5gjv2UvzvYNWmLC/zlwefItZx4
K97I45foqUK0yZAu1NDQxxU925nNhN8b8r7oJq+y7AJQ/ZjkH0FO13WWFLXQjC4hYsFPhfjc4DTv
fGUAecQAxTL/8rwRaCbWUV5R6DYNpDVm7rApHjh+L8JOxnw7FSDGpRQrCkluFLz1+j4IbhpZT5wC
Ee9ORpEDgoFi8QjvNqc5L5m+mAx/eHPAvAOyRATBpk4UT3MNoov8qgyyNhrx1y5t6lLZu7eUDrZc
AjJwS5OiJykKPs4eTGrWKT5OCZlK2AWi4nKS4wAwp85WGDJb5po1vvTs6b9YSLgTRM/u0PLFcnyQ
A+RxiNXyCoNQZI2iThIk0vlsEYNMhUXTNZnn0xNTbr5MQHBAjnWuPrel6ItIF6/MXH7XUEO34/U7
oMU853O5+dXkg7fNwgV3KnqFiZym5XzjcVuIJTmJodEyLEfsvxw0rsJ89TwBSqseqYu4f2tgY6FW
G5eYWB/cCYan4xQ3Hk4Wfg1uXmJHXr836loN99yY+yH79axAQD93PAykpu328pyJ5t9bbLUJ63i9
KZQA+maXslfAUi6ftPghbcky2p6smGyJyhqxCk1IZyAgDmmmNuT3AoEiKy9YA+zVjO94eY+U7gdf
Yi5cEnzlX/FUOFBaJTvCZNLXcoxgUVw6t63s1bY3aCg4L5sg4fSL519w8Xk22QcWGb/oW323QufM
Sr+mUI9YQ7LDphZWDvtlaaQEqlQLKf2Ath/bGaCgDPBzJoF0EuPzjALT2TVDs4oeuUFzTRAaor6J
W+yOsiLEZr8BtWjGvso7DoaDsoWySl8qdsIDZNyhiIiDe61SoYg8FG0v/JOe6CPOGjoYHONDz/oT
czLF25mPQhtTFbc7mySd5GAogooyPelpTc+0GFHHfK9H/I44MJ9DItGaoPBL5nI53butYOZ6Zjxt
h0SxBrnyDhyaPiYNhNT7bBSmPz10D5neVXiqLoJbjfI/4W1A3N7Rn/ersewVtOEnttP1uish6a4M
Qn8/f0ZJ2rILMPh2OQURelk4KBFDQQG7gqX83mmYS77HLiVYnskgg//5YXYbNT+EZvNUhkWF3Uw2
9L16uYykXYGGEKxOUsSRHxrG6ttOgGd53Q8cftyqR2AOqDY72bs4OVNGSaFd1KqWjraweUPp+Z7h
GL8KePchSFNP6zeVDYIntjYttEmliU48/T5n0zDdTgsYwZqHIcjlHvG3uVI6jklZ0Cqv8rLLd6d2
sBz9TFDiz6uPLzl+87Ho8cPAcTgtWtInvlGMckVpws7engHtqAB4LydkOnBTrtdwgQNfh40Lievo
RiunZYnKxvWM1PazVUoQ5Z/1J/pMvPkYAhkOInmb8i6ISGOn3i5aGmxh0p0SQZlLRpZ0GR8MAQOl
jSA0/z7OIEwRNns9ivpOimGUgTvC73UlVdw48Bd68eFk1BPwHPuGMBfF58abdjNJ8O9W1nCYph6z
m3KRx6T/URfFU9g7mM1l8pgMOI4C79AD4YclTY2e01r7HwodLLHUBC4DOfekc/gS5lz6lBpKXENe
zc7NKIPNExDnettbRjGlCqedAOy4VypHu/84PWOYEEu73EyvvGy78ALSWDrVYR/AQPqp5aCZLWO9
DXjnlCmS+46oIL0d+kzMe+VwMbEVGEtsLWFy58IjQ3v8++u84AI6xzzWBo0etITTJbTX1ByeiBSW
WBZYMG6/kyGABAy2xosyGQQmpBHtrsidjy6wjZ/bUpFkw091Rh9h4ANTYU7Q6ZH0QQd8Y4bAziXL
mZkOX7Dy40v+obkcKjH70Cd3GAMOMPkbEuvcuPWL1DIN0OSp3IjuG3HWwgR74ioTgo7Bka6OBW/l
Idt4cIbKaB/vHsuaPNkgOmkqP9ykF78bCGFXnjshfLaLkWldf5zBdYFEnAt7oshe2YzWSdE9Rbz3
6a6a7n0M9rO8dvTe8fwJaJga8KfY+Kq+Ze/uts65KuEOYOuLJtsHvv7K3y9drOp7Ess/24vPMSKv
WUZZEWj9f1Rzl3A6LpNYYHbXyo8kINd1zJGk9uMsz5PHcDAh8z7o/Q9K5gapOHBD3pdGw/NFXrQu
WRPBzS4Te1yNky325HYR9c0zXCuJC4JFpFvzv3sgKDkf5JVS1joBrsPuxxWbZz0hUSD+UJ6iStNn
94PfSKejOw2bZ827dXT8bFM7ZcIGrnCDgr5Ojp+/j4d2ILGcRKMVky8CopNUq3aWtVHz5v++0PJq
V/MqOhXmwAOThv678GzML9m+ix1qNlgX30BcerUPWYov8VOxdGEGifmCkedelSV4wdGqQ11pqYxB
kTQPUq2ZxJ1vj/XwSEN2/lH0Cn5gwrBsWPfnjGKHxQOQTpMDMyJYG0EUQdmOCeW94i9NdEfa5wNw
jB644sVrPgKygw/Ng0kEuVzMOl2avPh+4VsHFzPExrYTjhuWRN4VN5n3hnpJ7iH/Lc8pb2P1EQRC
GZOEtUZ8IRuJ4f3XLco8XCxlMwyxNzIpP+5IuuS3CmEUklFSSAGVgb7wDfDpQnOXo+Mmtq9Cfebr
miBwVAoVRh1mlWkJhF4A3q5jEB/oDplB/8JpHiUMo4dksWWIK2zZMzQTFGmOQeTKB1Vg/gZFmnWQ
06T4sGtI+2e6bu8zAg6J7XfcYAf4RDENOyxTvMaBVxKGM+ccMhTEq8FFIVoMVgEIKpQL0d6ox1dr
wpHt2oxoMtAw+H/rMSrqaela6qsYmeQ7tawH/VtA8R76zWJO7Bqj82Una/WoD0bpWTyBIkOueAR4
1K132etLP0EsPGy9CizorJEheSwRl5MIG1QupnZEUzWGsM0ofpDeofadIQ3Ey3OLiulybQqqkUok
Rv9Nv+oAntxx+zTPGoKb0dIzCkfrft1jXwuJYE4n3gPQMRRmkKSAyrabe6fi6NmMt3hoETLyr93E
l/gnVh3YQyMOiiy4tztgGbRhBbFhGHHUDmUfRvf2EsmfmX2qUhxuDB2Anu3rR5k25TtFLt2AW+DV
nzV+AG4oIhUTGkj5kriHY+dvEau4jGBEqHGdjFDQv68+J6P5/peFLVLLVFOC92BxnAc00mNjiAA3
FbiN8+Igfed9R5CIY8fJMHHiVelbe9Ua+1NMgt6wLZt/KAtiZb95SPOqkX2x7oHDYoZjwGfJ+phF
mx9sVmEHLbA111k1jC8oeYx7u9WvzFNc6JBNdfyK1jJawyDRIjtlu82zV9wRnLhxhPVqXO8z10fm
5NwER/YsNle8Wod5JVmbGMllSmBXT0DKpriJLl8FSnbs5PjIij5cFW12m5zsByaCs6ECRydojmrA
10EExaOelfeb1mTbLukeRZSgCWOMKltcrQSjcRfZCnlJvHR5OEh0h/2YsS1zR4GJ/HFjyxAZq2BI
+YFL5zoaPp+AW7tbNygjq8PiOklvO1x524YTqOp5/btC9tNDHzfe8Nk/7JMA8GrGQ9BEtjR7XRv2
uiRa3HYzRQ23tfOhD02QppWYV2oFmWGYPBC05tvuzS/PSVYpL06K33to70z5JP8cGQylr1DxTMDV
X2apKa1rkxSdnrzEW5OusE6L+wqymt74seTGc2FGrJTztHMMSDJtEz453eTjyeH/vyUxD0zxh/Kv
n081dLFeY82C/PRO90a1ENytgRO7nQ6SiVJce4MSsAIW2KTptP0FX3jNkWt/kHwpL3l415snD65E
WR6xRvo3C6llTGq7s/i8ZX8ih87yTGhnPk6E/amPVfSGh77KyC1y+0uwoulUsCmfdXHj4kQxtmjG
wYg07ULhd+i8tpQSMpMy4KHg2QnzcOM5lUQWIaWXLqG3DFaxJIlaBV3a2R5AIiot1BnizhsOpSYM
VYwJHf4g4it219g0uztfaL27HsjP88iB/s7vwTbGCuDOMg6yVIJYae7S/q88GR5QCNguusTf/CDL
iT9U6rwCFm7TuYKA8WBwc0Aj6um26c0V0xyY397Mx/5qpLhplhJr+OEJ3AMRxoWa1MWEtm75botQ
ixgOt0Gj9zjt08ZCoPIWoriaIUxJncroeZyCdwSA28M4vrKlLNpGf1rmoUwCb36dlSmGjnbGGleV
sK/SJ5qdUzFssdFNlr2y0UxhW+7xOCNRUKAv5/QJreTm+2+ltvpLk+uDqK9SfBvWMdxk0gOrDiwE
Ecx+zSl7d8P8gs2BBFRG855HmpHJp4LWejnliZkorPTXMuBdmfFz3GashF3ajNfsmtFvw/ZuCrb1
PL2DzxdaUZYYg/XVr/t08AFatm6WgR4VK2K6IP2BPEfpljpoFZugyCJLLnJe/o5C9vBEDRLEa9IO
4bQJydyQJ8KffqVLEtGykcxtLrRkIHs2WbizjRIbdJ8s++DDx9xwIBT6q8NOLM6or73NTndRzCLT
Fb7kG09DuPgPlp7ivYUPWt0q9iqFb2VmsgeopdvjVEfS3JdsvIxt8VeX/elBvRxDQlnezvacdN9y
ffKStBD83KIH/z8GYYQbFv8x3BTDlwkH7CywImK06RydkqIU4Angpb6Yd26RbQiYQk21yZ2g5bQ9
mOWQKCI4qsfJ8LvMdnFciunJRkuzrx8q8h5At0hnWWbohKlQ3cyv65q25mhpzK12XqQ4+7njk9jO
9C3qE7jx2Wx7ZCnDwXCa6mfRhA+W1833IyXuzxDpzMrhtzybNm/9U42LLngvAJne+1VNXLct69zW
g54vteYnAxNeMDHZrJrmJ2YqG4z6zRd7bno8Syf4mY7CDnJy9wcisk73oQ8/4qRp0+GFOK/mrPAI
aXQXvdIjt2KAwKMWgUGZ8jJzx4qdzDJmj32+ZlHugybtYAVN7nTOOG81N0fwUMAYM2nuVxo93Cfl
n3a02iwjpX2N2ijNklG8+JBueLBdzrPQNXela7s7vPx8R1rGvvxEEtE+BTYApQDfRuX39jmhl9ht
jXcXlhwGinK8wEgEnPIzKMBR4dqybR6cR4WAUc3J1HyW1S4B/2RtmFq4itTiH0n+70V9KNbJFp1p
tk626fShzG7kdCAlpM/La0BS7fpXf1LwTMsMCwV9EqWcuPMtuiGsnsIV6VqLbRJdE0T9SYMqNA8F
926ksomW4Z3pEDkvOIjlW8nCHMim7VfaDEa8v8fzVBHTOi6onCWNSrjSYKYKvm3WfGsvIc4VCE2z
hyHVX3jk1IYikNLBs6vJuveghjVxpAhmnblPvttC2Tk8msRmBw0J7sDrPvNnKnG79vGRKXLY1hFV
Sjouyb7pHUP90Q+F/bMmhjwOrcZ/onY8Tw58Y0QWAlgFXrQEg51f5To4FuPIeUxORf8DBi2gWOrC
wXverbczF7xZdDd9Q4hq5nWC9iIXfLcxcx/C5KZYNfsOZEzy6mzTRN+jeA9KKVVGVeJTRj0KzZd3
FiCYimahcK3jma5WLNmHvnOLZWoFvxzImSDgRlgozB0dibd8N2ru/BjynTFsNs4b1WGa5m1rvrLi
zXrQ+3nxy68JnH6oKOJuNtoJftwUGwrzXIt+Zw/9i5okKvYdb6xuV0O2GiayokHk8GAo7z/3c93J
1PxrnwbnjPFMJ746/PVsy1BOaZYhY1p9H+NTuqwXYAwsirqipTUJXgJhwRkd7HphrWv4rP+gsg3r
FRUiXFslpRMM8Kvx7yZtAgLXK7k3GtQ1ma+V7zmOqcGO5hU9ukrP0ifEvubP+4GcvjK1IC0ZPw9X
FC32gf2I5ir9coeX/AL2semfvMT4WvZ82D00+7A3RYW+t8yGLNYBj67Ljt0MTojMFJFzaEeOmV1n
uciMqr5XszN5JUNxkgQLo1S91I29jSnfL6CRLbBlwmdJzRHwSrK1uVlK7JYYN4mNjfJ856AUIafD
UVyFYqTJX7qzEpalf4j3Ea/flbBBYxO3R9A9aBgtVY97HEDT/diDtvwRKTMv+IxShFDmWPO6yPLC
//1Bwa/6XyPBUD/QmOpfe7szm4PkBdsNTMk9rUHP92VkA7HuYZEmfTJwiFSk58KzPrUGpG+l8Hf9
OcLORpQC30Gi7w8ay/xLqAlwzqRbOjzVREoW1d2QGZPPXac79Rd5YdkiWIqViDjy/4JDMOH9uKOJ
np5Q2k9cUtLnHYV5MDFzLq3DXQXeXTxJaLzNKJes2nkksgJNzH6efdZYm16EWdYn/NO+ILhdyBDw
15Y1HxEkywTAjQyf9Umlb9Bel0H9w0tGcxlv5FnsT8YGb/iJkHJ8/CRL74H/bjoRnbdrojv+4VK+
D4wU+lQnYvps8njXq2WfSsVmNnekKhqlkIs47Edt6S+mVpoinHZu98NpBatxMJfecRcA8NLa1uhi
ij40PrPU9WDzM8gW9Rge1dMWhpnBSSMoE2CznX7WfmYX1rsBhSqk6D7NUl8ROH4E4yMjpokEEA25
0hPuvZyMqOxGR4tT7KYF3CCVi3y4V+xUiMT6lhKSOxpvogE1ap1KS50sWh1Pj4TAV2QHlVFUfjpu
G6ZDecXNm1QBvuEHHHRPdqklBRmckn5tPLo4ZCjv7eK0jVpfXdsoM2+fxe2UYe/82PavCKD/HZoX
XDJ+z8ivcO9uMn+u/i6khEZqgMlfVYC9UlmiNvPRYjKA7lv54dLKtSVdo0CJiYWtSJdxkzUbgr76
tyqSS7msi6QIwWdjnGXreb24noUHrMHPmKgbo8wnnmWMCIqJoWFmmus58fvQNtk9YBs4b+Va+pJn
m742S+19gxkSsqID0kg06vhXD2ljwyuj9QN5xV9ATqmBV/P+rSVGbzOtzzM0yq6114oRjSiW7y17
EdyM9eTBeowYbX1QKSEeY/HhkIOdR+FeE5G6h4zQdvDf1p4hoz71N7Q4Gw8lEh0qqafByex80wrm
W2NqeFl/qetKxmcq52i9F77N7I0KsSDktoRQGby7kD/+VWgfXlIc5j/Y4VKNclMwICSGjmDy0dRv
KyYLKmA3ioPpYQ/zIOeINlvYDMloJLIZh4+zPfxserW/u9xE1FbKCN7x9dW3PRTMI0E5zmE6iKGl
z99VyDie3la9Vbd78KyIXRbmfHSEQr67N/dtsRjxIBlzM3DMkbAn70J4K4MAMDv21KORD5nhDFCh
rJfQtDHbqigw2yX5KGfENcqYE+PqGWmvTi1F/qN0IsexPeFxSLCvFVwNV20hBqIAnsQcP1e0UPyK
Y9B85pB8IyUQuLxjrW3vdykc6XCHeOXD3UdkK4t/H2un5gZHfVh0LdRuN8FuVoLYyl/1TeSTac6I
Z4/7n7kosa3j73g34E6ZczWtmzP4Lq+JR15V8tqTfaLpo3kWIal2hYsR99672aeX+fxbVvJ+cyJ3
locIDvbFG7gZFmDb9c02WsjcLsrg3DHJph2dTHfKBKUEKNJkTxiKOZfpFCpHC2YuNsdxOSLx9fs8
MV+t9Ksu6tz7nzeZa/vtBZecS9nWePDcVQ6XUyA1uEeonQAQCbdBzodZF2qMr+38+up5IdRPbpty
GcHGKb7h1y4vJlaz7OQ/zVqej3FNaLPEmJJVFuRoe4u26CWnn9PmDvSJGBZH3KEBWcL8COLoqGSN
oEh22fvPLu7YmyNBnuc0m8UTqtSsu3qsfBacJVOzuTT1rAeBhmwbAYsSkjBjqhykEKaj7145XbYS
LD0QSVg/r5RyTz+UBfGkQETJcxcfTIShqObcq9q4tKpT4D3kPB3dOhHTwgAln/aN6lSvRnAW+BeV
o5QnUtAtyxBHtrVRiZ9sLy2eSkpRad0Rq31niNLjWFkxQpSssJDFs+ZKTBOIICFAsspQtRsI5IYQ
S49ri0kowWhmay4fzD7XMtQVNF9Y3z0h3YsxRhFZ1yJUUOfC5j4qqx0Fe99vyfnawZi4zgtF/R+a
fUFox79SgaUocZHfY6OyIHu+W1b/xYGBirfT5WZb7MSrKnBgLW6YcOLL6Yo1/oAsaXLa//yDONCm
o+px9ia1lzo3VnF21u7u5WVhSIvbfVpsMvpqYSa2BU+yyliApireUk/7uO7J+4d4CbtuTVA8d/PL
Cj2O8mhkXi9hTQ8qfO75QYNa7AzP7F8sgWk7WlONhBo74i6vnV4DKj5IvywdjlHv9GvN29vRGhr/
//kJ3INuJ8Par6jL+9k0cBBd/nuIIm4ZjtE7ZmMvp0kcKXWQyo/lvgW/brmpTgGmT7rKWd5Zu51R
oHaGVgbjdS+qkr93/0jJ+ZV35Eg4gDxyT8F3l+i4jswkEMEeu4ckcD23fNg6Ulvw4oLaSYbyv3/t
Gcw/QoKiwugMUs/G33k4xEpr/ig7ilhbyGC6GeLQ8UW6Ug97BYUMYDlX0dAYZO2NlPQ2fpdhOL9A
U6Ig283/PpmooL0cuT15aJi2pQElkXu1HkSk+zSmCNC6CbPp6lLJI8oZIYrerg0UJAtUYNEi7BoK
sJeCLcKDLIGfCpoh1cqKD3N/zreJgtt3VEXX5oz2JVLMfAlAjBGphJQAHPk3rk80yy5BLHyM/LDN
LjD4nuGwr+2d1cgs9sewXfvAlpqAJ80QWguy5/Q85/0qYCA1R8OEV7EQFAq/rDirHJfhV4kx7CuQ
MeCWDbLs3GQCoJmPSGgMx0ushhmpE5jJTixQFclISZQHiwTqK45EO8PwU81J2x16M7rPFWLXI2y5
MQkdfERzcgzKet9HF3ncSEpjM6cZQKsgoinA8ZLo1EXlz5AVZc8NN9ycSQLzuUlUJ+bkvQNtMFEL
F9lcbCu3/4NzogjeRJhVO3OKgDtRbyqtwHWXqLbPDh+lMWBKPj9aVPAdvohrZjajJYg1X2nVssk4
IDcnTXgPdVd16fY56NCKkGMfeAiSUssK/hPSTIjJQz1WPRnPE4LqfP0mc7jSQpn/HBSB6iekXYw5
rRpvbjY5FTe3Ll/DjsiFavsSeBi1puoF9J5ypNJcmd6BRK1GqSooWEHB2tCAD9wwu1/QllbMVZIO
3DepkR5mCxZvcqZSbGcH5TgZB12064cIsQhdS1lcggHvGDD6KWnzQRhpLLEHkKLeiK52FcD8dxpU
oj7+lBKBt/yzyX9eHR1wmug7rULGTQd7pFGlRm1q/pKn1jXzoV/WMxEpw4FXDxZuJPphYWq2Eh4Z
GQD8BZnzzEnzNzzWAADv3rxvW2VcTvJO+t2yr41yKsiUuVVyKdo8bqLmk9ARK+ifmPuDkK5yqeJ4
8GV2655lx/64jjQJ4Nj3lHYGCfen7VGTY7xD+otLhQ6kd2KGg71VXRA+tdfQwSvFgFbkL/GfFV4s
aBnwjZqdg3kAm0rj+kKATGL0JMcwPxWm2oJHn9Gy3hVTrYdg7PtnFEYqVOuzTomu1l5qU/8sZIof
YeQQkUWudqbXCtcGW+iJ7uVYe4d1ulia/mPIuZEydTtsg8Oq1u6LpgAtPis2TDvYY5dTdNNiFsp1
xOkCQEcG6/f+nHgn8ZezR578OiKQTmTWOLafSecpzZ0C1ZTSM/Q1Mj49xxfN39HohyWQjGCy8i8M
MmASua0R8ML95PnALIK0qua2aREFpvsgc5zO4A0GdgfDpAjr6bfCmInD2ryWFrNsqA6HDHOXGcMg
ZSapduUibN672/a5ewEoAS5nO6PnMPSLYMZ24LNl4PC4mfh93+cJm6QiyllIGua5Z7Q3TqIiTrZr
864FUuJerVW0pLSadgVN0gYNnmTTS6iPF0iZ72dWPJLjQfIIConvtqHxvjQnLB2jgrGDX+g/6gG4
t44iiESEW4Gs57k9fm4w8dI8Q9q/+loI9Y3kqYMCeUnBBJaGsoc1PwZCHntrVChFxvpNmTDnwJGD
HjcDyc7y57cbzk2fWuFMimzcQttHlkZopGfGvF3CaVq6pRnqsLzMCNswh2PfVqJX7Q2Xqhscv0X5
87oTffX0BzURZdUu4s7w6Ud3GZ41tMAA4L6YRB4vqrAfAQE27SPjRtaRp2jKDRyV0p443wQBGnUg
e4asqMM+SN6Ids3G0ZdG3fG4Ua+CnSbFsg2+Jb1eyR/FTNT7fYb5Raxjw0Ds3DvjM8ewPnelp3+q
PbHF+8zYZMTFLYH+zqUE4Yr4X2+hbqyqd8FOuK0vugf/gKDB2hygCEAwnbYesTJz5VmSGftw5Gh1
QA5eBlEmn2VNsC3vSA1bFcZWgennu9TrWDVyjs7X6kXONAevcUF97ZIU2m/0/VW8lUxQgZauBu40
Y9TKI5VTQ5sUs2J1JKGHVHXKCf0lYGvK5ppMNEii0VZFX8N/70Xp3tHYX0olZjZ/qBiKERCka1Ni
uaGbrhJlJIKgM9CXb9T6w4P5DbKhHPLyG0kC+ny5SxA+eeOJ62yP3WFSJivSy/lMhwSlkDmLYH6d
1olxi8XFMbQumbCSj9r8YGqtE8nq3Stfb4irjoyuE9WnmFf5zMpmVofklhXI9YpR9is3hNi6Az3/
KhXq0RP6zqTAGUgNlgK2x2BBwFa9FEBf3/kBENU5oZ36e5m+ZHmTfMr2SZuIyNIEqbR4VAJFOMnS
U153a14RcLVFZloPiQEzX8l21bt8UOLXxKgzGZ0223ObpxrSAmFk0b2peJC4XLYc21syLwMvdaH1
vqQ80VA9UT7iszQVz04Ld8qJF8cbbVd9MUQAkvQO/pqY4YCvRFeCrbTYaY8HsZpOfW20Ww5MYHev
/UXqtbqr/WRReLZwi0R9JddjWd/uFkKaT/UsN37wvcGzNI7OmOCpg15aXx0djjue7yWJaHFRcveM
4e7VW60suvBIXub/r7AU1K5iSZDTTKwvteSY2q4ngUYHP3pmH9GoFiQY/qcTvOPMLcG1Mgw2Z47P
fiWlY2EfFm4OtA9rbQNR2IuOFVHCNq+kAK539BRcop80Y86aQlAJXfj+T6PmzTyg+TfpUgcetvao
xke//2lU3yxjmCoffg4mziiu7pLQUlGymxilgUZFRBsIWmc82JMau/AP3pFGiHx524C3OrDdhBhZ
kOY6Ki7iREtGfS45d/P4DYp9D8UA4WoET2wrFFMQE2gUGXzf3slIzH18+PSwgwovkVCU3Pxrolgd
mPW5xta5eV7gcUMaHA1E1GfjQDo0VslcPSxQOf3h1FmAfsSPZduI+e4KrJuXuUDt/F6fgr4vhuqX
kxMsnGHVuGTkMODn1dlIVqwh9lnJzpRTzQ7KR3R1vVbBGVDQ+4fJKBv6sLGLy35J29bBappwcl6B
NJmeZJ9lmHKMc7fdDL0tRAgiQQZxesNZi8/jFeLayRRmdsRYM0nr1nw8BWIFrFEm3o+vBpU5noV6
kYHp4lE2585uGunN+x1J32V4EOpaNm7zCx4Kq7amaGCNVkHFVN2ZGDd6ky6hX1P+lCeeOLUA5G0J
Y6NGwBceVpABgoQtb+diLsomB5GS/IjAm3ZPrR06zL+prCN+oul4HrtHB6NRrm3Arx04ihhpbtzq
KREkJv/O/tB4q2DIwiJSmkPsUmShPhW68hNt8P3cqpF8oZW/Nzaj5AOdnVSAr6PE3euXbbNM7nbb
NCTQjN7kKtmxNbRyzeZb0K5Sws6zzt+Hp1/Df6VngZDb9d/ZviVrb2MW5Ia4Uqw4aSkZ4pw8SZW/
HLc26JWNMFHvFBZiPENAc418Ipf0izv3XWdnFMyyozYjiOKooB0C7Gvx4/mb6O1KwOHT7TmD65B+
ha0HLAm5c0kwShTZ7Ng5sdYfZ5UAlppIM6QX05zbu+wZlIa6J/0QaN3JyBHbyCFom4B9IyDBJ3Sq
uenHBDKvAoKf4jRR3GwH3773P1mri+5Njq5n9jUVQdvapu/Zny1PLJeBZ+4bsVbnW/6GGM9FXse4
rrmKlCydhNMday47kWQ2hZ59v+2iLxxZ1HWETnUwDlXPi6EdpGSVJVxMtad4U9WJBagbP33qEB4j
iGw61B7S45fif5HiJjRu0UypWJU5BUX2LVQFrheFFYxbg2wjpDalCcr8i3y8G9OsysO52Ftc9xIu
GGRGVi4Z0/8jU/NC9c77zU5evZTfshkGk8kM/ZjVvISi0Ryjg2soUcXTxUOmZH4rvQ1cEGfzDZzY
Bgul3O4ICbCESB8A7WhpWjUyeUafV9MTYS3xo9ivjwew8jbVccQm4uhV948qddkaoclDFjckHjxo
GyrdvbgSiZe+nUHrEbVYKv+Yq0dRa1fXy3eqosAu3oQZOWgngfmClMbblWVC6855dqi3O66Yy3Ep
VtxmLDmw7C3XZjurC7FrR3Y9fgEqI+wp69QlxAU2wY79mSALUsRQxxruo+xn5X/2WzfObT6nPp0X
MZQK0TJ2zokoOcKnWlQdzAWpd6rOHo8Ymf7Bl0CxUdRqC55CgmtcZg4u0B+9aKr5FUeo+SEOSvpe
3KpB6HaMULaQfEkoWUejcfsCFsWgcKrtXCXW68oRPDs1MSrbzapS+3evs87VmtExRMroElVOMn9Z
IZeWuxBK3ZbALcby9uaQXxEpfTDJailhuptiOaIrHcgz3B0srnO5+hDHpiC7puSZY1NzMdlIZY0G
CUgLGTIZvyzpWueSvPiu8ObCFMMPAyvc41ayUIpxrVJWLMVPkMuF2RsVB95cszmZpx33jqN2LrzE
INMh9PSJJEfvQA52UqWBuQsTMd9XuJkXqfhaoMiiXKZWVeTeq7D5USeWcK8lcxyyuzlP3raOpzhf
2AqeHDp+rCndUb5yUKt307vEzSKJJ7hODK1j8acEt5jiBr29NP/YLBv2UHjR7usqwxF9wFkaVNAT
Xu68/0xX3nScuBYPisDZoarR++wbBO5OBPRaZDed6fvKm3y2n0FuWpwoxVoVLEvgbKmKIjPG96sg
KbeStLLIloPas3K7ZtIfyOs9I1GaS/Q+9MOhgf35RI/u3wcKgOHVCFXr03YEMMEnQjcI5UnlLNxd
BtaMwgYEysmSgfgefOxAdfCIxUCfkNsf6DYcQYMXpSKHE4gunMINOYwMUT8yD+WWsA4/iydDKLqR
TWcTDPCv0wOtgr+nuczPRWrygrU4BKoe5zqLFCRcb6Ony69v+Zo0koI7nr6yRH9kQ+tBdKpoCtCZ
DJdepQx/y4qnkYZZFl5+z8qo8tB4CQbfX1KdGUQO8HuOQWiohHi4Gm8WZlTQ/gntrxirgjf1luLl
MuaYnkESXYSNwZGDlNr9fh7JKe+nfuDnGHduKZFHm4YUqb++5HliAZu/SV+gmSiiRW0i7FpoxdlH
Gw11x8f2V3lh2mD4FKhxoOa956C4WTp7chE2eHqQubaHgD7Ol0WniIjDDMw1LUh+Ma4rQgZaTlec
NAFVv69w/ih4WbSJcnu8NdGKTSg+/cDD/EEo/1OpHgpBOfnFBsYYrfQ+cU2XhlLARcn49k4GZXCD
OGcjJv7rlhOqFA1QWxyFAPmlXS33UvL5A9vvMmEgNzrmdmltD4MIwlZ0oTkLG+o2WPZ+I2wZYXmV
jiGp+eIKktmM7tyrNyOWzNJWlbYT73RQHZW6pEj6HbPi379G9wQhXo6pc8+T3MsjZ8E1o1roMGhZ
Z2MAuZGT5iBtBi6LkrUG0RabzzS4bntdwEYOMO/GgGovqBmoatLwC+6CnPUtQ0v6zDzIs1uYgyK1
cf70QC4pdmdwPzcCYRB5lJKm3fDmd/l1ntgBhb4TjW6f6GPrDiSrtjCeEedWgIUTnjttW28mQZsb
X/ijiSGo493EB6rgOWBEXIiW6JakPEGtqhzX9k1u7N2jgJXcHwxVhhVOhhYnztc4Hoz6wwtspVcS
QUWVQTEqJR5yPvgtc1gwqfCKJYeknSJ0yiVuTHOTdLhmvOAhBdevai9Gq6JU4VAT19Cr/el4JzOn
0qgj5e5BAnlKFvyZoutlVxfT+RJFz4dRuQ8P/hER2BMgyvdpz1T+rKNAenLvIc7DVIxZXedoByvs
foN3tBtvF9Ix57Ype+U0FasbWyrevTAc+0e3nBvmVYeYELrL4P7UUw9GKh7RC7llGlcFVLtUx1qx
7yO64StEsWzNW7PwehNYWA0aTjk9hyM49PS/L16c6luHcI0ZCL2BGBF3EEfv/H2BPDkj7/BYXupD
BKT50xSDn5WTK8FwJbHA7s5xPM+rqhZCQLzKc1AOYQg46YBIvTiYYAvsr5B7D0cu9aIrLd4G5I9R
T6cmBsqaSlDs3wIjRWx1sivNfBVVXxJYeiEfcQBvW6m+35jkUy2WB2yrZ4QbTyDWNOeiurNxWWOb
Fc5ZT5zODBsVuIg8gr56ISNDo7NKnehYgxmffVF6ap8+foR+NyqBL+CJ/DvKqEcK/PfcOHxXNZa3
JUHH1Pwd/ZVAWg6A0JhfudS0KI4I0vmCra+nuDCzKPDrAaWN1xJBOS4HWkR9DurlUXPmM3CZTnR6
Hkt3p7oBO9bmZcTesRcqqalmmh+3RBBqW3AvaNzmQt1IQXV2n1slOv2b8NkyWi1NHmYReXyjY2IA
Tva8fAhweNz/ACuV20iUm4KO7w2QTbx7G5TZ89cDFAZxXV1WtSS7+EYS8B/Xhsfsx7xRF0UFmqBX
ThPQ/7nRhIjh8ONif1gXu2GXwKWmIePeU6eD+HtLh0C8Fdb5I/g5LVykQKx6F8XSrD7s9Vcg5G/3
gzrGYeDPy/5Zdsf5uoMcBgRNf0q8H+J/9PLOmequz+8cTvZ9nj0y0m2GcQYkt8jmJ4m/0MjjBFtU
+jAHAj8YoFPoRJKFiuDpICgx5z7IArgbLfOkLyKI+/qk96z2+yjVdXkWpszw9wvky5/hB0yavvZU
BmoqjHHWo7Q5yiRk9Jsp26ysHK5vnH322Y8jZqfD4uGm73BgR8kvxLUlA3QZAZM64WRrq2GZ0oAQ
9kUcBoHHYx9m0a4HjT2QRpuiwBFz53N7RjqLdWI5nki7j6mFmIGSxLUIxPh4x8qVw+NYTqy6HEWH
DOALHZrwf0F9nW/lWMMM+pl7VBKRKPszT9TX0ie2rb1tY2yXxZh80WaClEa/tgkM5iEX1+jepQJ3
Ul5nYhQWfBwUXYC6MOIs4X0FHtr19iThq4s1q/icwNDdbTVTuVZ/n0djAnt8+T9caGo/JyL99h/w
BcU0q294VL1FFddrWoVfzYiAbL0f9RBl6s3qzYi2kIeffAOyT8OW3kWr5ayqyhd9mCjaRB2y7edF
tDWU8PvOfRWk3ImDo7f2dDymjgDDkp+SfxSm0HvN2T5VgP42OfdcOGcRR7s/8WaKewP4fUgVH7as
A5yfDWhb5vM74b9vChmdcM+3TkIQd8PBIAEU69seMhY4ECIIxVRsQlTsP1Q2XRGKC3ZjWZjatwmX
94e6X2E/cUNnAeqvpTOohcWX8/vM7JkwWQUsVnGT1fRMfEtz5DYycG4XSbMTVnPYwmvbcl/QhZvG
J8pHHGU5QGYSp64V45TrZ/G+uVfbvnFDZt0A3sPBEcAdr3HNbmXrmbq8jZHXx58py44KdVoL/CNX
RriZiHqvo65ZhCU7kss1R6WLulXZhkmS2lndh0l6tzANpaQqPlgEHF2DeDcPmZQiy+MrWgKdHDZK
ucmPDClMa4eYD+QsvNDMqxxNM2PPUX+NGjxBu54Y8wLBMmKEqehlfR1DjN7hE1jWy/ukEdM6Gy6c
TE3xXry8iQFwM+bt2ipxmbpwTRei3DyA9Z7Nc8qlixcaBWo2F0cqjca6VfsuCz1LM7+s9dGhVvXp
zTu8TACw3tp+GnCYerd6JOxqREdVhzlyd9DoQLS4MA4S9cfCA6JGAwcASWA1YJMSbqOGfETOFWW9
SHJXxOyI7VksfnxiEHrBhPSGNBC5YFReGbntDh0moNrmqkiXaMFlKZ+GclIRayTxUfj4Oj32AuIr
SgGWAKOahFDneUfnRGYGiBrbmVhifDuOF3p1g7EAkhcqy193WqRRFqf6APBL5ATmTf56C4S+WDFf
gvivjpijTX7BYQ==
`pragma protect end_protected
