// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
U5PG8yxi0nkc9dEnuqAIR+cn09Pi+dyyeA1YwrmD0pA1BZsYz2eQAzj9Zdkij+4wmVQFMqJ9KuXh
LMqudPOaxdyXelcmFVmgguoWrqb4Iou/zwbOS9+i97JShTyLd2bqKbwou7fwvOHHVPDoOvgNCIf+
7+CZQkAnUaaAmHUNMhVHb+/wr8Xwm4kCcFOqoNpsULM7Bzn70LnZ4VHtJw52h3hIW1wbzdHSIA2d
htjYsXHU0+N+Gsk3o93pWbGWEm13PdqQgjZE9tW3Dwgv1mU/u0swEZVpwuWS/teLa2zpEbKapb1z
Z905WKPy3uOr0far6v37BGbQeb41eTqwlizlWA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 66688)
FCJOBRuyjKRWAZ/LyO6SSFAiQjbcBxrQJzYiGPfzkthZqZMwYbxQM2nVzs25DcU/qVWV7YXCWY5o
I+hVZW7MndO0thtKzRX0PCau7WM+412uB5tZVHhChn+5DZioBWBDVHSdVfcmA5Di2x+rXOiMq4kh
kd5FjuS8tqha/J4aiLWVL4+LsYmVxC8PQ4HrLABGWrB0HIxZyjNFxMI0KyEnbszTEBir+yWScYTk
gR8Xjbi/jlLisPTqwnJBtudPhfNbklNOzTnhDXLVidWQxEJpGQpS39yv4R7qyW4uRtPz4cENQyFn
BPkWpqN9i0xJBX/qRskHxIMQxs5BL/K0fVHrYWNawiss7Uob0EHNbJtmPyktZr72LUTvm+REV1b4
RtHcm72epHW02NPkBZBUGB4fczrZUUMY9/fhl/+Lcb8ODS4ray6DERzpUJ9A9qi8tkrXyu4LQFOq
aDDIN3Do+X+SqMZceNsR7V6S7rcWHJTXJV4IhvyCndw8HL5pnXvdUnuHXv+K9oqwYl7U82merMmL
V/PGmSoY8EF5MWOjS6a49VdroLTn1GLM9mABhA+sxVK67F8golCUwy/MM36Nrk6bQGOzjhxXHCPz
LMeSp/LujcxURw+b0UjqizWLdryydoIJeqKEdVCk9eCRmx/d/sVBIhcouf06+ZHSFuXb27ijypm4
BkaLd2fYCgY8+w0ux3766BLxICQVsOSuAZUrbHgDQL8ILxSQ6/NlaMUMp17mwFDhJJr0fChEuiLT
sPtUFK85Ag4HtKRHzqTy4Z4hnQbs99otfbTwNazN7474P40UReGX1PEMVcGxn6H8YibNJd4WYswH
iBPSXrKmTuGEHmNEBi2fc7M1YiDQ9w7jixhPTz2slqozvAMAFZTvfxX13tmcKlDimk8cnE8xyoGk
ukAWQHaLeqid+/9Oa41m6R9R8rd5Dpx1qtfN4pKf0tmjJwDGutsntPZ1PLrKyiBPPuc4hzQzNxIB
039Z5AGNyUPl8wIq5yzZpVa/5rZvGuDFz7QQ7eME1Zz+arTAhP+H1FWhJPFy1pLulZxHMsMC2w7f
9li9JKZBdiJChNrZWadbd+ZHVy2OzjScRachp35EG10L8Hxbz16kKtt2dCE0eQVesGl5UgFVEbO9
jxTc8vksvhSuJUhbbA5s+YmY7trOVfFkw0sdfLBPonCYq0goqkke9afMDnQMzdTl4dhq5ukydbVo
b7mjXN3UWdVUQ8o4WjGxzMrr3p/CAbFkRqJC2YUy54m6IH31uWYtdHxvk3syyV5D8WuGF8rYVte5
kXqLzMAoILPiz490EH8cQ/TXxAp5ab3jaKfyhWJnfafJjMURLfzWp5O/jqJdw5wtimEelZyyvGmS
XU63sUNitK63oCempg4NLWGvIVMoW8X9/HITmhPpcGR7D1pOj1/OATCeAF0tFcJTo5jxOrqrrGFJ
ihhwTi2bQ/itWzLPsFEj+f8u5Nze8rD0Mr6Geb+QnWu29Fq/rYRno9vnVjY3L4E4Kcrs2g4uU4jp
+QcrovpGdWrQDzl4UwwhAhiSx4g/SM06jAVSVzN2wZmtsd8aI4sTeeQKtTlfkd/UBLLfVhNvrWUM
To0PzNf//UhwDteR+vc+hDbN0b86Gbue0/6rTb4KXOL2QPvjaKO7SX8BZ1fRZBcrXcnE9zTd/Tez
crIimR9tmUaxY9Xa00qjALv1CZv52G51l9WgvoOnjFBSjlP9W4hO4/DgTsuCk82D7lOwg+D8sw+I
/GXc3x9v6WBouMv6SlDELSjutZEKjD44XXnoumYEu70aVZMC0NZAyy69L4p8lz49IIcuFk4RkE5y
NP9hLJTvhujoaImcml8xWx36r2WDzBpXusFyvphPaY8MvjRw63kRZLtpq/oYrzHp/vxEsZ8SOxti
/dEakESj1ux1o+z1XW0UlImqEzX7jqco7SiM4Gq52d3PfjhAisHh6LCsjQHYrNDxR3anwcqe5KR9
uWqfDXnHNRxoY9Dz0r3hEyNqpUoPQvOkJsUIyKwUNj6x3s++1/cabGKufuE4a3VcObQCmWnx/oIX
7Gxy6cc3ZDAR3rLXhERg5XkRa6NUTH4n0LT9qjF2nkun7IyhCc+QhuuEDQ/eW4CIW/uW962wlILc
StV8pgnairTgEIKt7RmyAy/6EvoeYOBO3QJaeVoK05ZUifCh8YcDiNuqXm8hiSwLDzVurDqmzk03
NoRWHs6mNUpwWEZPOSZV1mNKAFwZHc8mw076nLT1Gdvx+E7zHEYoF4AGBmH9HrmteFuoPdnvZWVi
KRSeytK7BH1dNoo/rBSgvfnPS+rXIm7juPvHT1bBZ5SHmIpt7TGU7iqn3MQG/hsViObnu814LnZa
FOm98VTZXjSvXoi6plajGopNlu1aenqn2rZLW0rOuTU+ugDz0DWKTgxbD5ge9U1uH6FHgUA77/Zd
CDULcd6JifxuGQq0tMW8rtNch3aEJ2aqurPoThZGhfJ2af5Trxe2J5ilp1k4qxrxmLP5r5xrVjIB
t2rqbB1TjT8G7v0BYgUYwsEo17/ATbvpSvTwriqCNU+wx/urGBrHawcYq2NScNzUNe0UIE9KZ9kg
nGtS/sCQi9H+hcZn0LX4KQKEklUs3QEQSJ5Mz/1wzy8DgnKq7milhn8fMWPMgJmpQg/WjhWTLWlG
Q0qaWXpOVaXxtUclN9ucBFUg+LdHGyNKquzKTZmPoImh4gYiDoVTej5dQEF7LShMVy6b36NT73I3
LOywD78W4hqqgm9KLJgtknMSrHOYCr7ZXzUqDIEKFOUSxHWVKr/BAtZZHFnCLSBT2UvSt/RX6QSD
xn+gSnZMKGFdd5y2547T9xhpbflHQkLEARFUxfiU3YjzJNty2p5ubw+d3YWFToNYkQfZPEtsQoSJ
wekJK9y+1nur2sET/kaahz2I2ZmVKiSdEJou+mlmDhRtxNgsWY+P8kNvU1L7E16ArN28wbPwHDAR
E4bnD4GJnhT2iarr/ej+qmieHIW6nJX0f0HlgQ1Yy7tatk6oGUX2Wh1Up1Aelcof92t1Zwzhoutm
b2F2j7+9UV7VDtIBY/Koo/JHuDGRdpOBF9Km+r6sTRsjHZ7kdNjddBiXAsxFk9I5LtWr2r4DHbwP
eUN58kOhgHc3RGDwT0HPFsAVzd4wHS/qNxNDR5+EQxbXftiwMku0QWTE6ln6G084RJ3NlE/CkUlY
xZtCZtmzFWuLrlPbnmtXXR7Wm0xG8lZv3LlWhjlpz8ZHb3EfkrePm79muIu/aiiCcx55V5lv/fOO
YzwOv7hcnVsmhhBM9lMJOHrQZR4+TS9E/ooiZS/DJJ6jnLuh0eMcqAs0OO9mZZYPMOml7QR688f5
d5WPXi2gv31aeo/EmmuRPXtTW8w26P2CzZHjERgxRu43F40vSRIz9eOCwPoMcbJBlPIwkOOORAoJ
wiMtWxWMzxfesFOqaRuOesAGecsCw5N4KaAdOUljbv2js8m1QrUTJF1mw6mqjaucM0fz7HfF8ZSD
t30zp3otb3MslvN/8NiqlJKdnw/vKsYTzK4QAZja4JkurrZYtNA8hx9dpnvL8HP+9AAuBcSsGGOC
omVzuLk7TSGsqht+9PfWMT7xNNKmKetPTghwtMonT/3z4dzC1jtV8xLXTdh+Y30yFxqiHm6TFOG2
nPctNuvBjlhBr67PyfEoG39ZCqzEdN/CBQIOI2aNl+2EtkNO1Fs7AkoTWPTCC+oD8lesgJT19lpb
T9shsNEZ68DHbHHYZdqko0QRFmGlFzBQXePyNGF2SY5ZhoOyQFH1vv+BIFiRGjMGFUFhyqijc+zL
GySfw1tgsPXHcUjEBQLXnDqerWCW/tJJjduMO860mV5qskk4LBZDFymFSSqJq1VfehYMzuITmCPI
Sy8i8caCUPR5rUlD77om0rnlD3j9wzpCpMOoVwl4JQXwsLQ/XqVxadDO6zQ0qx5gV2hYhMaOGrWI
/HoIK9mrTfC88TM1xf2pH2b2yfUibyE4O6RaWfr16S5aI1UpODJoWgRK8vgo5jK0qLukDEvkZ40m
HGfzr2wU4J0dtMCLYmrxgctjS1+H//XDV6RMq/CwfwgfmKxcW17cINq8CCnQOo22r/zZ4ksgC9pT
fIbyntnn/pquY6E3l6AMxVSSwBvKgbTUXY0NDxKN/r5F7s/m/Ty8DcZ3+Stp964mSmN55alPlRki
woEWAFNVDHt8x5l+u83c6301LqPRiyLa+IXRqfQfJpeSop0UsCyJifnNpGrKI2z3EoMC006naijt
F4tNVJP/mSVvFLC8RHaT85pTqfsz4X1cntqoxwmMl0lPQqCRxBYnJEKgiWeyvmJPzYGQKBXh4cqa
hDeMXFk6N2i9NKqA3aND049sqmUqhy6yjc90wLU5R/BDZ0zcE2KT4CSoRtZE6nCpiJ6EOGHsyadO
xtlVT71DmeqgnKhAht/r4qY7vhD79nZhfvaA9xTDIJrdNfvDjbJP7sOzwbWzsnWj7RjY5psKpCQa
kITXuYSr5jHQ6QjVXpGqEXBXoUb1Zf1WLQ8aCowOPyghDcfsUYofiWNLFNeFu6Np7qQ3Lro6pNvO
Bxpixq5Ic5mbCVRWObYIgju0L5G6dKFpJbVHvek5jnfuL5HMObH5iV1txPNg8PKb0JBFW3K1ZEJ4
AcQdi4lZ8cJP5d7+5hltXHejtskAJ4f47EukZHekmApctJElVBcCepB2PL+FMno6IL8KCnXION3h
FC2/owNYS1oBkF/BLC6i5iyuceP8/NwRo69n0wKILV9BSO4aLXBrI2CPwLMJC6uIhlk/88KCPrKc
8820Syw11j3NKAmBx7GcoTIxoiMU1qCYopGsY4+lG6npSG5tr5zivlV2LJEhTZta0NuI/mL9r9Jh
KzFRwOTFYbagt9dU1/+i2K8HzsbO1yVDGiRNYeAIxcHwGkRoNt7KqWXYSwwxEWLu8LgwPKgCjw8J
A0268Okf3lbQVTXgA6529mNog4IAvVSIEZRsPVDZfkpy7N0ZL2l1wEkigm5CFZ22Torf5NK3O/vD
EDkTBMZHrHVJRznc+cvWfkQ18j1Su1qoueLEaVZ6KG8VSefGIAx7HtoNyfXVMeNLJer4nwpjmfyW
gOsX7n0+QyKJ/kTaZof60dw2Ju56GhhLuCc839b5000ygX93LXLlubZgSHZ+UZMwyXE0th+atFHh
ymZZ64u6X3VIj3Un83dyQkWfWZP3Pu6vDE5nSGcuN8NYaAClAx6W+zQaezuThMmJfjX8ApeF+DSb
GvCf91XVwuM9DlZvPfJAJR7HE2OwM/mS57Uz0rZgXqUab6DMN/CSDGhyySpEJdW9Ec8T+KP1JdHa
/1EfIkDKQbpTnsBYgMxbwaRLue2jybF8pygmuowyin7JzPf4L1OkMkjO3bd+k/U6rsuGN6M34JiY
frnLf/pySFkAkeRlet3GxOMWg5+wOriyBhNh609fcfYJjueOvdrNZ0EiTYE1RE7NxGF4WKBDqevb
Fh+TAtr9PBWLWLT7JjSZC3VCMdif84VLAfx/DQ8exuRGtAZqAVpOWnFGR1kJV6IyxtCJa3vbpqND
vPebI4DxnWI1i8hHv0K4E5YKnyBj13nr/Ne7UVDeP76Q6n33/1Zlh261gzTL+Dlm1Ob6wzacTc1t
BZv9jocuENbeUns7MxOkW8YZ2Nr6dktPsYcBkOdjtYMZQZ/QeJYSqdbqlNF1DRfbMd9DCCfddNPg
S/mz52nlP1GU8ahQQQNINo0NhSPpk8f0Db/umnrYFpyQMMU9+x2H2mnPIW/LO9Ru2HAwmt6CQUPD
XQVpOLDgolPUQNBP0kivRYbAEQGRKQ08010i8gEtIrowZOuhva3HgyxyJ28LUbZbZSSOa4xEH8CD
nhuCeCI28oT4UpXCju19pud11Md7UN8Rs6mU6FT7CrQxnOdvxNqhjae1ndV9Rc/vWoEZHU99xD/t
n3qYZxK2zkPm/PNUNPXOWX/Ts6oGqUYhf6vsX6oHrfCXLyHVrqU4VI2xUDZR2My0J+flwhKTmi0b
Taofkv1rYp6JmR5DB1G0+sSJmCWtPuWTcW4olBAqAUv50+BQNFHltyPhBn6UYCHh+QQVyUCYTo3K
0LFnHGK3oaYTpcACQGG5wfvARnY4G1ncfG3ezHiPYcJ0H9Rh4+XJcfnZVoBMUj9WZS04u1YDEMdu
K+yidX5Vhkxjmj12WpPuhg1fUy3KcXuzzoFkHJOSW2HTDHzCSM4hjkr5M08PVMDP168o+V/tWLMx
Zz4ge2vnD4zh09OAsgFREecSNBKrToSlKXFQermDPRwarfCFtR8IV+vAC/PkVilEfouDeuzBNAQv
vhT9JJpRVtI5RKOid3RDUpEeiAjbauwI6NV4nP7Q1iF6QGk0dZF/yjHBHzzIEbxNe0OXApSn3V69
ugn7hI5Dn+VuOXu5aVOMoFoCtelrYAK9XbjsZyTudjISPt9dZwim7Wzhmj+b5bJniWFFKbbMDCuF
JyfFGQL2BYGvpHLoYpTi1wmo0qcASabtDd3n4Dvn/GMx78IwulXFS11Lpuj6IXp1KDPEFZdLKizc
rp7qZdmsxtpCivlzi6p5qPDP+IQuJpQ2evj+DvaHq3XAJFMvownla5vl9d+2RTMRRvmEoa/j+Phj
u6W9NmS2pYcNUYLhJnzzAU4/2s+QofrBzwd4xhlotw7nHyhE21ExIhoqvG0BGI/l48Lw8jCb5M0W
eTec+zbeTHIayL/LcH+RDgKf4EiHCXOcoQCB6i2kr6LKVu5GwPXhsn1hgrnkuvE5gvf4Df5nYwf/
VmPFDsjcXC546dTWrsNcyqrgqPZBdtOFbYvpH/lgl4RJRdbPyUt6o9rcwV7OqrNOvcp0R4W7neIg
MFKOuAdqUMffMytO26ndBqDIK6h+lVluQuX5USL8zmkaTQAninK974itN5DW/h199F0FhMeUV5li
H2cV3HEQFfUV7hfDSGX0ECt9QHKQzUqEDIiyQvNcTcpPHw45clu4SLJEj4YTPf/SFEKWBN3w6DBm
yxb5qIcBTaWZRbu57eiriV1V6Mkj0I4kD3rv1FrdDElwvwekHVWg7lH2ltRaHwScWGLoEj2B1Em8
CBjAOV8Zw6Ffdk8MmBwe0QuEqmw6/hoBEzJW9veLBWk2NWdbyhhKg7VXtal9T2ylm+5RUAuo3l4+
rO07vdLMYpXFZWeKbJwy+qbXu5srhBIWx377PV3Bdny0Xm562UkbAgbbtOnlUFhPHU0cSaMfq2xg
VzlZLiLf8aHkUOTh/0Q31SFZecHgewHPXuFkBa4LG6pM0Ijs3z22LUIofrfNg4Se1Kh2sdc9Rz6I
FbggOL3zRrmfIJswsKVZ1m1xtRimG1dlci4jUUj0WxbMBLlwe303DYxNHmJLjf4Pl7mQLXKlYtNo
1YlzTW2BD7CY5f0oKJa3Os/xWN86iCLNu7wz0xY9PlXgRbQko150i6ns1hmsvwJMd+NfR+aD3R1c
fwhpGH7RV+hp9U8hjkrTflKNdkRmF3MTdi0/n9ZKopq/3ufCXK0KSa4MkL/gwZeIRcd0IoygQA3J
PGKflGryAur64l1cHBLEy0d6gYSBvWrJtQlwwemIldgw56JLFtWIq2m1JYgxieryq4gGha/Vy4IS
HfsuP18XxDdJac5cgulzL9uAWtvzvath1FtOh1ugbHlkP07FBFfaOpsdfF0PoWSQEk+YgPlmy/E3
It0KT92Fk5MRXGBNAOO7zU0LYfI5hML9L6aMj90IGk6B8nB49lkK/v92OFFmpV09szI2KiY63AoL
m6yFQlPap+dmpkCa+OD/DVi2VlY77XOOow1pxMdiXfzh3UGT7G4ERP1lah4qcSSp83wxkcGcj1+X
hzh++3KhSXVDfZmcN2OkOpbvAnnjRTS1Wv9ndjRRCGrmff2JJ+dRBxxsugV42/AoHp4SZl10fYsz
14R/EJ1TCgCf1RcbLkxnTvHyO1siiSyTSrHai94H79aCq9qEdQOaFJ346bHyGhbqt4Np+d9Cx0Z4
tliwd2jypxYRYqgVsplEKrfRTvtCPniGYctiJJRXijZcxZqFcKrjS5GECsKEZGB6wlDvYrpjQegZ
DYSm9McXjQepWZT3Nx34FWDrkLzPVpp13XwC9HSKjWgX4hYuPPSHmK8lqRSs7N6dtaVRTRJe6X3S
uJj7kMWspBY8V2cXKP/6qyLSffTszmQdVUiSaizAY/PzXH5G7jh8SS//Ez2z3G2+lXJf4XlZAK+d
y+X0aIOF6buZRMQcfitHd5/Wjg/64xYctyOvHsnYLDrk/XR+XdRxgVbS26FUAGooTlfDtZ/WDTxy
JVKzXGC9eszbPildMNUg4onrtbmZYfdWN1n1kmnOQr8iFG8AUVsJfIlEJHGqbkrIXLDMD+mUt+Va
G9z61g6lYzi2Vsbmh75IXYUh15Dle0hbFsQIHhjoZbO1gKLHUx12UzJteJkQrVIEogQKOqdShgcL
O13N1qoTT3Hp6PBDppey4dPP2uyAzDQaAzR3NZJayN2V7sNCQt1rkzaTnhIj2Y4SX2HA7Cee63td
s7bICiJGp3Laeh9PyZvNKnNkIZ8dgZD1IIdKDdhZ7bQ6DaiFV6NkDmDke0W0SFY0bmtQIgB+RKup
13oKZNvOnamMX24DkRUX6F0PrxNT4a1H5hxp8n2nGFiDx6iQN83fgY3T0PbmClrX+1v2thAQCtmQ
l4DhS4ud0s4D0IKAFgndqfCN0tsBc6c4q0uqEnsRK1jpLxmsfPSYsIrfjFgAg7TkFQcMZVoOS02b
8Dms3jSUlYvUkfCheF9rCkd376MYZ7bX+G8/LTEpsD5qVARzNeQ8kFUZQQ89d3Tu35nqSzVyPGLL
qYohJX3hAiHbrR2wfwnZALxxrTHA5OQw7osau2OhVERrlgT7yzU8K6roPz1XdTVN/Es27Q6sg9/n
VSADnuCszhHm0Fsk9gnoxYwXjxAu2GbgJtPCk1dXmD8HQu9Z/jhsnmrCdD8cRlv3GBJQ24itqgT6
jeQ15+lHm2v8OW9Up6EiJkLnW6HH+KUnvkkKdZEIFJDTVH+wyNxRVpIvw6wbL95aJazXrEsYF4dO
Jvz9j3fjd20gpYPRsfdWcsd0fjYmGznSbiDV8dBolWSxvrrl6CObabJYBiFkR53vQNMRaBRWtbDV
vy400t8EwXI5A6TdkNb3DFlzYTEM8LhuyENb4rRJBpud7jef+6HN5WKJ67HYIyVQJhJYR8G5YmC7
/TU7rAhI02MPGCB/GYXrT1DnlMniPU+88jZPY6DY3N5kd7vdHG3W8k6DWQM/BnErSUA8IxIU0fU5
cSUDVjOyRPJu1gg3t0JjJMjtpJYXZnEFO0FaBGFptTSrta8geBL8zSFUg/BSNK2Lkso2H4QVA4N/
APgwnKFBpy1YrGXu+wEfW/KFoK6zmd1aXf+7jKfppHLeaxaygJLMovnNXC8Yh2EvIi9eXBnYkPHd
Du+TK/WLBsL7xjc3bW1/vu+qTOyBrqzVuMiawJj+PFiGeJB1QKc7hOmDLpCfs4hnqYdAkCvSpV73
/ewHT97tdOHdVhFIsrX6wx0Gv4hILypXJzhLHhCr8a8jqccko6gmG/2mphjsPyyxzOO6sgMWQOEW
111WI+MY63yVOrO82TmvYLh8hN2ncDhFj4GkPgIKcGzHULFDHQ5L1EplHwrcqtFF6iUrOYYpDWR5
zNnK8huy7VGDrzLIPewwkAjMyMftIF2uSfay17lcg4LgDeDGjbq/AK77BuejvilO8rhNFgp79vNi
fPNEdZEMjvk7+AVXAujYYQ2J7DuO+NuwIUG62eLtWnfwKCiQsKLV6Tv9wW/rK+ytiEH6jje3fiPz
rjFCHq64Q3L7jshyshvwK2Xiys6KtJCeYj0bA6gpy5YtZDwA7bI9tPmP19rd26IR4Ph6TxRkkYaX
q4gQq89bnIA7AOEbJy9cwHSpYgDxl/tHPk6JPgGjciKvGGEYoqvbsO56dEf5Z7PfRoJrYmkUve6V
XFiz9KN/ZWa5/XmUR/srTKTZz0SMqkeUyTZjpRTd8zt6qNAOeUyNzeTwQG+xU++BrB78dzkLBMTd
bSMXXtqG+AtP4A6QCBfWEcmuPxEeU0v9wu8rljKV8qoydnmLM/1wgCsKQLgqBU3SrCDyiJZvIYzN
J7rst28TDw//pbHPMmWxAVAKo2pmsivxeMqnYd74zSI8lF/KtGRNzA7GVuvfv1hKvt6U9xxyTxmw
LC+RaGwTSGQGvdWoM9vS3eBXhuGdsknGxoG4wtV4/pmfnbAUuBcuutTA+p6f11vTUyBG+sOBVSkk
PVnoqhcIgM64dAiB3pOwZahZwIeaX4x4ZyMW6aqsrjU15u3frFSdKMoUV+OrbyeusVrAFI0+6FYV
FIa4GgzaqB5aRIQbXagPBh0Hg+TxiyDhjZec/iNaDhcvCaRE+Xe9Ilg51XGP/oh1WIqEV2/jXfh/
nE8ZpgQ3nbtVmmvdO4HBq5kpwdGYl1G/0iIqifo+fX1AXUxuHpYXlv4a0nTDlOc0ERo6DBQm6U0b
bG3Z2Y1I4zSsKd3qOMBd6YCcbVsGClRhvQzkaWNVSURlxG0MTx8KeUblnPjt5HyX4arjp4vjJuk8
V62HuO/+ONUqHZihRHk9NKG5KpGHet0w5XhEkUJ+4sXsZwfgbjKBttBzGiIML/qURjjwyqNHCEaC
E5xnQcbuZeJvRaPkTPtFeiXPyteUQIsuj2ImJhVYJOZflmEXjMqwTRqIfr8rwwNeYNVD80aBhMQa
wp7TcDMZ85jI6/gtzzUAk8SH6MwAR26l+XwS1ES+28p+i+N8HB/dzAQ2oVUQQUAKy1t5D3uyDZyb
zy5qzPDM38hD/56203F5Cqc/ghdKITsFuFgMwGkUWHsrHayFepSnkBzpBLJ/1Ieo7Mohdpv8G6Do
GohLUd2xsYQC3SDPrmNxj2EFTFk950Vn5+iwPcneUmCff7Z3lvzhGF/h1uh+88mMQWNEkraHgqlT
TcOzb1PmdtNq+0doZlVHcQADCboj+mYa1LAaSfT6enE5+XBfE5DuKM4jk0d5S+8S/x8c5k3Fbvw2
pSffbMQ/Xx+x8QhRDkoNEM/afNu8ppLZIEEVtegs6LgmWaMql7UpNREAyf2ChYk9gdXMHp2kC1rU
/6viQwDOQHBYQBSrowmOoBPNmE33M8v/uiRt3VDN64zQUqhtO3S6zAka/yMUEFalz5jlWHtLYmlO
d92cWFCWUU3BxafK2lOnityaJtfjfNzOzCUzuSuMbBKQ2Srz6Dx/2CbjlkVMeZuuKt+/16kVBqXa
z/rYMWswlV3X3iyceGf65tyxmQPSEF60mwKBnv36LIMxzsgm9HabtItA4nBmpgxFkVP5duHevkEn
L69/OeYoPWdPt2qlSAUAHyF21dRwBI60FSF12A1hPUDpaLkwRTG6nEMAc8SF8h8FIjBFazXl2fte
12KWuvMuIB30QdRNEDEQexBDi9ITSvAf4Gbr/iPQW4I56W3/j2YY9cvDagvZQXuWsShT2b4t5PRy
RL/MLGk9JY3nEr4upALdsGo3EKI0GdfyjQjJQ3sUErtXT5rdWYjPwLmsQpJQJyo9YM0bhUdyE/NU
z+QsLI+gxsv8Lwa1Bz24AlfjFM6/90lnzkoChjWNc5ToEwwK+RpnON/jOGtf7X70BlQGtsd+D1/W
3JBSt2maCJUWcOEXSl4vQEm4/F0BN/8tSj2K5FU6Jg34jzKH6kT/Ogg81ka6oJ6bBwLyosJV3meF
kQUhalmb0fWoRdSbMaT70615LpvaO1WCBr+wSSGNKIM59/L0Vg33/Ww7gJzhIeif/l5iPEMrBaU6
H4luHPQ0s4dl15EmvngSY2yJU4EiLNZ/ZBiIhGCVrGHSHaSm36TwX2uOENOlPswTnjwKi1k90z1F
24mRjyxiT8TBCYCUX9u4g3x6XMwYLKSTGkEfpYDXtiS+YVriUIpwNbUlst4Q6iitv2nHSlsbMT+j
5evhVoTQw7uXgQclP38a9frhXG63ikREnH2TYS/KCXeiSFeNZnquq+1y9TUvTQn/VahtgMn1HwME
JdVC9LIU+cUndd0OCAXrL3zkhO5QUelrhyC48HawQLB+UYm8tOTEjK/+N/aLajCcxyJKvehO3c8X
MNdj5ge7sbmZSI4JrUkKvuixrRlz8GLKJsPDpOZQVa4Xc5RX2A5yd30srfa1KJelwHda6pqc10La
Aw8KmYgfwpJnFkXvwDlMu2jZGRV083qj8tuTGdkVnJ+qQFl9eU6pGazOl15XgsWMjxGRAfgP0XEM
T4gSrg6274GEyaiph0nV9thXuCDC06C9/xkzgO4C+YeyNqkzb5IhYn/Iya5ddWydz8Zp6+9bNr6V
4kaZ7JNzcJ+wHqlvNbFT9ZbO4nhklHM17RhuNtOmX8NhPrzoZVaNi+W4L4wXvKLUURjc1taoXZJJ
+5qtT/msZ83IoaPmNbvo5cPLLc5ZrlrTKhtcz56jNf+slrM1gZj5b7BWMn7U+30jx3v+AA4jnjUA
ZG1cm8XUbWGWAgeIzUPOxY6qptgJOJCXGJFmExEGefF+ddGK7QqzYHCexKItECye9K1+ZgxTlk1A
+g9s1JHlN/I43bH72qOH2rrWUj7sAv6KK03exNMWRDxPR+sa03jPlpY0WZ9k+c7FDrA6Yrkn7/fY
djDJ2I20HRjcbkj4HsXL/1cmpCWguYAzzMrmBLkEkl4RFe10jPr6Wf+ZCgrx5k7AJzOFGifQlgWM
sU7+9LhtuV25A7HZ+Nu43kRpxA/W5h94lNX2X0Jt7t1H/YMSqvVBHt7o5p8jJ+huZJhK9AzJAI3M
7rdofL3DO+60N0bIIYiaSG6l4CHdYxOq+6yJFQJubRsfCIpVZVPoG+8GeDrDTp3pX6qJwZLqtgvB
sLdbecUWaggaVo4zz5T3iCfv++Ti+rKQipNjvdA+0YEacXpjhVvxYbR9FDEjByFbVWSkci1jHtYj
9hYOsBcKj2e42rJIIEotS4UaxGvHSF/3lZkRD7WZBMptOO3zMwa5OjYMr/nAlMFyKejbEQuooHdk
HYkteKMggHQ51l4otV0Zo7MyyZo1QXGav6Huuq5jzws0CHQbgjLCU2VzvKnbu14dl2uWZv+GjAVT
l8O41Iw1PHVw8d0e2INhnoB5HRbClesMNl+/yglnOVKbVR2/u4qdHltsvnvVwC1egGkxVk304hxX
eHrnjb9GJn3Y9/HG8wFWuyuxBvqAUjX9GAE5nvvzJ8drjvHgP0Em7191/ocCAJokA1UYrASC3cap
aSRnUeKQBJFITol+zC7OEGPDmVYv7f6H5z/iQs+CcO1iO+0luv7NkVBExg5WDMUtzRvrga/gMr8z
pXIDbX/aU2ooI0XxXsgZo6N/5egxSuAFslK1CMmAuHAs7CveH9whw8lSWd4DwvleXj/8nks8JKdd
IDU4gO/eM9rbiABkmzv1G3mC6l/fRrLsW5RD/PBWenwBcHFFBp0HD1zDoVoqCB4HsrxO0Mls5hFx
Y4KIMvpE7XwvNF8wzjWP1vnX81Qsf0B0CGDzITkAEAQnCcAEuEI2y0XSX6Ramm4I/mHP7H0no8vU
dXNNjBYP2c8vTvnXXeUeSrm/qpvShevwbNF5LMji7zQcmC7AGw6Jp/GqmzkwBhVTOnMj+EZzY5Mo
vUV/S1p6Cahkr4dJBQ00kOdB2nZ2wYslk9LTWOGuTs5B23jJvCXO0rPwUxmp6SG/Ub7pBUHR6pp8
o0D+5QrRYf+1R/uHZpgyQZG4jpy8eTE4awvF+rzn6iQPWNjSKQrJ82erx1LZCm9wejcFmex4WHQa
HJxHr/QzwQVcjB9hw5gnYlBbYb+IZLEn1dOtwaB1I6wEFIUU1zxzGk+RbT+SIP4Boall65+GHvfV
E/SYdF32ROE0+qShI49x+pRTfXuIxUJXR2W+ijzYciqYoS8itKmYSKe3Lp5v2yqZsKMi6lhtXRgT
+YpIezbTdRIhwZJx049hFDwvywnXptBrhdy0dCDqozhhKlXZA0jd1KI+oiXxDzoJ3jNFTPGiUnCD
KrI3+tTk81XaVrx3Z5ocAS7UyeFklThm4H4eg2d5FmMmXmpOZ8FqpRDKfNa4XHBo3Y6Q7NNHOEMj
jN4P/4nc7LTbzLiFN/vIWLWvWTNivWzh1yj2ZiGBoxYE9UXNDFGi/zd/DpUtyAKgrn0ak/SeVR6O
bzqY+RqoQ4xQEa4idAg2QQLvHzt71d+K6Tt5kQZr2+2Oz7plOQMv6YbMdNFwuFmZB+aERZJE4p6p
gveszksNZfLzXnJUExRYFJPyH5NRVujxvmfEpvIuYMuNPwD3jLt7Llgtj0tNmMLxNkPEzqCem71z
BVEdQrUxmV7o/BZCcVchwZa0c55CoEVJ8wQX51n6QQGycWS+dP4efNa/xis4CssnyD4By7cthCZZ
pQYICzHu1bl9X+0Rz4eG5iIjAzNQJFfKmPB3sAlC3SmUFnMuTWCElBUJHUwnB7BQUnuFfWJXutlz
Qz2QziobKbG1b5/TwXz/Kq/RNlaZn7t2febjkcq8OGR/rQccVyVxKi2o4JFEyMI9wcFEEXtBnorh
bBdAlvyP8K8fncN3KaH49W261pDGgpp/lK/FB2/UP2t09M8VPMySdwXVkpzjjziYVnKpOTBZlGU7
NkhLRiXCwuBcPTWPj8iMPV27dJOIC7n54PAb3BdcgAnyLfSh026Dmvvv4bQ/uzVTmPILjWHHQFki
UsqIFI3g989oUly7ElH1SJvUDTBMyQZD02GVRkOKEUW3maveMRULV1Ty0L4nqu3HeAPhy2arGOv1
898wZyxPXMuA9IM/ArMq4d/NrIvq/oWhbAG5OXRy0pypK413PT/mrGLwkchIU9ogsSSkv3wppe7Z
uJ1mYZOmNRUNshia2sB0LAHeTC8KGgEXDfxK+9aEKM/VOIaUGDYUPh78VFqXFlusiKYAZVKScji0
1iE/Ziq21xjHgfj8iAO/a88+ydzn/ABoP92JQfFgicCqVFp36A3F4Oour/FQKQ56jEuKrNYsNDFk
WoBNeyg12oIKYhYqaGX1pBYJbHWGHHCLS/VZbVAOb9BPgY/SURbzYmcuKRswTD3EQ8LSmW9c7edk
F9ESqpS+MPCMzLlVpX8ZDlZ9SnOPrD9w4FGRugUaeXFVZnhZEHjy2QyAmNUmM2xsKA3CJomZ2wHz
WmjWBdIHqdzNc1yj/FVxuT6OHPEpSxl58XpOiSqRjIWq28FX5mDdUvCMY3SklX2if/DoscWFHlvU
dCAquFW5Q/iOF3+9JRXBRiqwnTh4TGStZs8P40cVQXoXRoq2//Nr+HFboqPbBuaWkCkh3mAGGZow
3MqrWrSkg6lYMGBNm5r36ZlnKDk+RovqNrjp3ht73VGlBkgRYPqrCK1najXN1XPNvkVIdkoCKfPq
J8pyhh+yLn/REbE3bGpVD1acom1TPSnCz60R+T7B1CKfBsCL6/2JcWld0GRS9y+Bd2FeNP9YSyaj
HSoAkBufMceffEclvB4lpfO1ELTyzHfJ8AZlDuMlQo1VF+MNdeUqT9RjYm3JHH9DDkLXqg2mqmyO
/gk7ZkmShoisoW3Vw5AaT2bbzrSnSevR119PsQXil1WPKbnXiNYuwk/dywva7O3VvR95vkn10jmq
mezg6lTnLO5MkbNnDT8fYTF3UfiHqWdycn1qomHRvaxUAI0Kqxaaheia5hqlxAkRGzkuz9iT33Ra
CnF7nWGkhLiXCQ9DEC8j+35DwM8PGhOtKQbEg+kEdDktYV2/Geel5FzsVtFJ+RhSUZyxrtidTDa9
Zyb08zXUeFJrADOfF2pTrFncssZxhhpQ/KIh+PkcyjH4H1iME1URTk66i3OtGeWkb/Gk47fbdKLG
79oS6xOTILJ590S8Nnr5e88118J4AiO2fYcrAwvovb0E544KAF3zmAs6KvDTJ+05AW1PRbu5kp2E
MbS+qGuB+h+YZ8OdkGLtoaQBUv9mJLnS0zElY61Dv8e5Qudz7jmPmB/+WqjBS0wZkZxjw0XK9hOC
JYglhqN5o1tpyhB7NWH+1u4LaDIeV+xImyfvfoPTPtAGuNR5/HWaFrHgt6B8bOJNdvCnj2NRYMIY
JMjSb5C6m6fu9xYVkAe1Ywq+dO6uCHLoAZIj9dtITn4/6PnAUqv3ktOUGRqNom7F/iWOwXa3SScp
HC/pXnpVtmop2MJnEbuuXDdNL5sgU03VBTtKkgHPLlrnk09OWge+tjFFr0dP5VufAAb6dPAPv4nh
tsYb3JJwi5CK2zkcVhGm8q75kRTXIiOzBCW2xUgJTC9ZiV9OUKjIYcYMa3tXg8h8wYRGWjwODnly
fQP1Sxr6h2ozurUFe68Ldw4S0J45Dt0wdJW/B+3U73gxlhiM3Z+qyNL0hXBxgyfx7+X9c7+zTaY7
5KKtiN0NWK8Ue+2BNa7YzUsuGJXNbHDfARkxKuQXcJbuvR1WEJ/0XFhaKmm6e6ZGrhA85DAYhMYH
0s30RykIO1IwSs43HHOhsiS72HJqn2BhOrBOsPSCqZN77peJhKDJOIpV+ixcluT8rNVTYRhMRnHD
pa9KK4bfSiGnm+lLncMi4OPRxZd6vZ41BSiXSKVxfZiCP9WQklbrPebvWQIAI0QJiUVRbkNxat2r
DOb33yBKKMhPPKCBW/pAUpmfpPhrxTEWYScCy9QyKtFnYmiHob9SHV5/jh3T/Xti9jnCEhLTYIqP
LIrYO8pm9GZ5dm9Gzu7FmRm6XHf23DfA78CNCO/m0sBzz8W0qstj5v6ggY7FtO6EQkGyDYpja6Cs
88ENf1MIIadi1dNNLOYWi9H/W5EIt/o9VtyGDWqNrCMt5IZyFUiXlfNJoavjrzy5AXuDDFb5nQYu
Fd8ZREEw1z3U0FAiyFhHmKgVSsgnAxtv7XJNf+sqCRYh2R4JQs5aokEPqh7gtTc6W9OO37s1DBzY
NVkzir3Qi8K7lVxjkmdytNrcEboLSkd5drqwYCx6b8sz5uFwULOwWz/smQR2M7oDNBII6acOOlB+
Q7Gh2stLDLBgml77wsiW6duIdcjttyOp7AgbLJngxwSBmM92+v01LdwzRlWlT1rQdc1O3hS5Xd+V
Ap0jBqOcZTy9pBh2pYYD6zJRXffeuxGyCN6ZmRePr9HcPehR4nTcYi9XHraJ0ubed7alJabqcsvg
vpL0zK/KcimoE6ZpxkZCwbs+utZaGZnBlLOFuqyNR6jGmGANNlGwiVeLqsBeNDAULY1cInILmpZ+
n73Yfq8+kGg/Bm5AV7RvGxxO8Rj2uxjX1JEmrHfMsDkzW8MAP0pF9/0zRxKkHCHxxNMZhsvEmobC
JZ/T1v6PbVii1+fWRUSyap3kozxKyZg9ZK9EKsHQcCPbBc0tY3g0mWOi8XwXoJiWFEyMN/oqkQy3
f9sCqAekbC9XMP3M5K/6MBSEVQbjrvOKSCRkKF/GvmBk5pPQFcWtMKA8zkL19A3abbM5cxjP28gM
XZLicvqyOeMjE2kFbwvM+p2wD9kbBuGL5COAD5OLZ8WNZCjIkQHc2HnQR1ph/qBsb018HFlfI9eZ
u9fTibN6xZF+Z2imVcPOvPeezgy2L/SdIVqjGGsv/DJGwAGQMw3OSg1wMyKh5Issc8b5Fknq4dOa
NIDSOpXaNjXzhGDMLJZZ26h9H2fEuFxquH7bkGZOatw03q3hRHPxih7s+rZD7AIg0iplylmmTnNv
12hicLQU4ij8ZDI4w5uvdp4ZTFIrm4YHC0ifc2P+abdDYeDlT1n3ADfaU5gclL/hqaLFX9nRxBS5
KxjwqG7tXUKPUaPpsfhLwbTrQjPNmsL5ymA9rrRKobVwmmyWgyIRARKIt7POMkj1/6GIm6pPmq98
tkykBkp6LBW74K5oSaHIZQxOEEclUjXzMJDFtHo/Po3eY8YbTWoJuU2EprwQkCPZKiULGh3Cf8Wq
IXRYmTUVrSpViqyWRHb5QK1u7gn7gbwkN2B/zambEd1xtCUzvIeD6mtWKg05HHgw9YaRfbVvQOGf
w7EqSyfuPj8vexwcHkq9E4oKgT0+tDyc6xPTkT/gxi6kueQJLCM8tkXI7m10/mbDgWJAJBtLFVIx
o1Yyg507BeJProZfepkMgV/FU8Hb2q3bPfYALnarYAk9/3poYcNeRUi3ocJJOrfHnzT0XdaddvbD
jKidfKphd1HdAhyE45LS2L7EkAwjey4ulDRd2BZZPxsayS5Ra/8MN7P0zJWAwTEFbcLau3VS6DI4
KcyBxe4lA5Icp1ShsLG3ykWe5iuPOAOypVoxTqXIOWJ/oq78KNS3wyqBw606F2wZTohKHeIdKO9J
NMJh1kqIB79p2UtnhJQCjZKrkGDAR4aYLSm7HM2K0fG6sreyiMU6U7LjKZBFm4Kv5JtAjch6a3oD
LNP19GUfXSLUgAmR8JwGqz7eO5h6LviC8/csuK+CU+AufydFLqD/k+72f7KQswPshUIT7oJl/CFS
ZICf59CXfe8ShCwtW6uqfdTWkqDXqgnCX33WyeDPBD4gslTPKHD10nKqjpROYLVN9ukmkxgXWW7W
ThhfrE+AOIYs/hKJMHKRIhL2AxCkqIUGlbN5t9ZVIc9CcGYophPWFPkkzlioAv/Fzd135nNSlsSN
mNVyFP/a8rkV1ljy68/Fx/qUCCTaqzGJlh84xAGLOmsiOjMkJCYl9D5FQRJw5gaBWfL355JX7qrt
+qkfjp3f1WSnDfQy7Rk03CNdv2FAPBFdRuNRsdqc//r/SIUA2lCgR/Pj0XnErX7hsmDvFRoItBeB
hfWt5LFnGBidHebBkYpNNGUgHpE2tdBLjRK4BHSRHlkvudB3B6B8N8SPkWBF8M9YiTGsnVkNsXsQ
eCo5oECHFQJHacQOohNoepH0gQEMsT4s79oSRYFFCVBlRLqBsUlG/Bp7lCNU/M47gHHS79g4JhKx
2328BA9+KIN5zhhmggF4tncxO6JgAJQKFgCdzje0ySD7Veod/ofC1yGRlzKuC64SQBMIa9JNOL2M
AromtzDzOMDpiEdyDrpGQoR3nQ42HgTQiPHjI4pz462TFUKAQKa5wTpT/yy9m3voRiDPjVwE9xwn
kGDsLAB1P+B1n7L88v8KwQrLyHx3cnuJw3vU1WKtRB9JX5iSwVaSYL3+nO2R8C/oPdmhl60Pc2ST
xqYoeicUcCZlFj1kK22QFfzbn34TSQEfoI0scdsoB3T9mmCtXOFOBjprokW7beFBck6V0X1ELhu0
h/NoYLoO1YRJ+AGSga0FDUAY+b9zSlXlZ4/0AoLjWHmSQqGF+0LI+zZ1+ZREoqQaOEtcKbcTTd5l
ZZvhCecVVyP3sj9DETWsqsdNfTSKSHwLoesnKptjgAVcSpkQTODZ9AXiyXOx1X6UXOONkaIzx9F6
BPNbXPNLJ6NzJJ8PRvioCoEiaJdZ8ArKn98nGXGw+LhFKxadsaJs8sjXd2wiIos9uxsxtagVf774
2ZDKC63uNj8QYoyDFxuEQlC/HzfFsKXzg9mggn86dwtnIR99bgr0NP8keKno8XrdHWDmP9gecins
q3p5hhcylKE7AjHw+R7x9RpqOICxOx0lU48B2l5fgW+cZCbUO5TMYUJj6OFbp2c64fFkN3Pu/qzW
ykrsfe7WAk2CWR8UJ7StCSaCWA+E/GQ/L4en+gyTzOmC1CbQHz9hpvSIM3gJmNFyWq5tIxhJAqbw
i374GzkgfrCJAx/b/nyDeRT3QC7ns85cKpVYTJyg8y6NeBBUcTBWopT69BGlFS82HHhmgo96T18+
zWIKykcF2hFLQmcRAbRiS/aAdNm5fWT5t5W2lMnzjo+OdgXoXQFDuwhaGp65dVME25HK3GJ0rwar
JUccIMs/mmHFUUBhwAENOCluph5SqoWsNPRXDSgLrVndedS5zomLiKLe7/BeaK0Yimb5BMfQGBiV
EWxfJZepfJqDzHJBZhSbnAAXsAx+dMc1/AicVRviWbmdydfgTN2EajCHGYzhHhUu3S1xXMbw+yS5
0H8D59cFsI98qAlkCW+9PMbj/Agbszs9lAx94BJ6Q3OCkg4pyjQbkAaSy03sip7mrj8eQg1E2tKa
Gp9quYO4DDOXge+xGlcsLQb16HaAo1RY7tIvY6zpfwraj9Djvrf2lNXY2aOAiFnAfzcFUE984JAz
gE9mcgp08e5MWstSoizbtenTJVVM/jlSNy2b2diNPYQb5ijQ0cqxJvAEjGwOJUVteno3TJP33SZj
rb7hxNRknp1Wc0vM+5zW7v8AJVxYy9VHKVJumE1k4O55yG3/lnT1VV4fMW5sGkQ+2ufXPrdtCZHR
5iw7Nolr2uYkTRJqdSs4TrtaNB06fvtZbycg8c/AQh24Q9k+rU5nHbA5WQgXMmKooAbLg5DjG4l+
YeR3LDOsbYeQGdsXx9nGaYaPphLV7R/G97Ezj5BjyrgnQafNKG27/ePFLKLrHIBEE7tt+z04PExI
H2Lj2AxUG+aG2JOGSL7qz1cQRJDyuSSKReXCMqZtKboiwozCpN9wBC2taiC6ONVY2WVisELLTuIp
j7nQ0nBOrDq9KQ1DAXJosLaa3Aka/9BOHVe5IkYdzavjSMYwJK12Iaqx+20iD2iT8CI0pqW8b+tu
S/LYa+itxju1CrLb4Nt6L1pcGX4LVFZSD78XMQ54jPNFAEnsygRSfdRZ1+IMOYRmFwGpXqXNGpHc
ivIDIoy/bFvjmoonC0IsQsaxwvRt5bRixhJV40S9VNGxzW3PXpu6/IkkxqLvbclEugpTjARHkWRP
RpjUY+9wtW+7escq4hCVVBnyncD3ngZlG/EYucdfW8M/gK2OJOlHJnIlT/Wihv03atteu8BhpU/p
fZ66eryDhvy9XJve21CRkjQzQ7kUek9R3lWApBX4N8q7s6McEJbz1SJdM6FVojbA5/ubqg2wN7nh
788JpoJdPSR0reSbMA4IgnfrKnfVjVeyBLXDT9hdck0YD9Es3VMmVRD+0ExkAATMC1/4Q/KI2EeV
VFydbCBGX2awMOP2n3/Sh5Mf8i5SGTY48UuUr8Wr/h0x35gZ8awOgleauzss/SKLW/oEjAyLvSzY
aUJLv4IGOuI87UMoP2oQZCdGVQ9wpaHRZF8nF2N1OJ3n0zVnxef4T+ddCRC3dtRtKFV7v9K4Cwqj
K5EdW15vV84AbisIsGuyco0Kw+FZQUmBMrBVnjF2/x39PHVoBY2n7rKE5291ORAJvEx+g1y0j1oN
CJKukD8pzM/9tQzXogqKwLwG4sUJsxOgL+wPQRXianlNJatqXZ71uipAPgQ/glgc6JYy2S2F18Qt
WdiwgnoSkiKQJBVHFeB6gcecjiGY8P8g/Kf5S9Y+ofpy94rORtlISTr5gO+Eh2UVAEyQjRJxTt3J
ZNEx5YdNZToj0KB8qlQSI1ze0PeENaTn0mmhJgNVyOWq4J043Sx1ZmkKEFjIjxVEfhFtRlpHqoz8
DN/GzjpSfFJlTiCZPLOuYa/oEnGG3lkwbDJahslqjlNObqyF6aqPsPa/r/dM6xqbcg40S6rt7yk2
NkUmMoebY2QC22OsP3lIavV18cp6OSasSYlVFb6/kV6VhO/dkHlO54grTpWyCD41wwsKpP7h/QNl
7EWMRzNCZiSe6iQ+TZ4Nw4ff1kfsIery4yTxxpW9k1SEz5OnaHOYXWIFwIpwbI/n9T4SlIeq9g46
H+cH3V01tLa+q/NdPnKgSFNktUSIiD5qkDBzJwoL2QTpy+AEdlFqdHSIWMchm+VOIEw4lDiGNXC3
TFZgYmRTTyoMBEg0AemcJkrqNG5/eSnwWjaSkxuopSpHAib/G80uncexrv1hVGbzUgokS4Voig+k
ox1dnjUAIG2jb2wdqZgu2uMZ6i5OlzJI0TJp6FryLOtER67kJPw8bO/JmRxjM6NnTaQhX5DOkvXd
m52PZlIfJA07zWrA6ruV0VYG/UWCcwIM57owSsnvO5VI6HJFf1cjTTQd6oFOgqPYwiRZB4DfUnSt
tWj5W25e/eNB+/2d32bxs6XfpcxQe0sxb9tnLbESqSIDHO+sw0k3qjcRJ3Ry5ntVtYL3KCMEaPIE
ynbGTJlD6DqvDnYqdB9EJNCyWOYioaj0pTllr27r384B6+QeYxi2NmaX94goOPVx4PYm+2NuJ76L
a9OcXD5AKlX87yxpGE7HN+rU0M5s521G/1h6vhfjqb1E0YXc4pKJgsrPkR4dx+xgCJVFuiCw4MMQ
tg/gVjieCQQxYMfaYKhKyhL5T2EUUGby+eUMEglibMx+DCq2GQ3S+Q/fs3AeZjHiHxl+8JViB75/
RaejrTKLeSJo8csK5b1mGpAIej14jxdjciIfWy2PNTLNSG/FSBCcOd/wVvSvJVh0t79oKFL5tZdz
9I/71PLH3+zklpxzghKLWU9dLsr1JW2UViIY+q/Tm/IMVALwg6jwkvfKhP1H6K9czCioTFT0g626
erE9V6EX3yPchcaEGNEW8kcR2fOT5H5UKhdZk4kYEH47UZCtOHClIPHEWCIzkQlxS8EdnA4TFj5t
4kcYUz0HOVw0ct2gPHxA5InTV1tGV+tXa1MzhM+edNhl4Y7zd04toHyatYThcEhgnpDoPtpwKlYt
usdUGOZ5B5TxPVPOzp8fRnpuuYyX2U2rOzUHboX/tplIXazNLf7/NjlMjZIlfJbM0yAhb/QUot3p
z9lPt8GnqpWBolFKhPNWNRT0/3KEhuNcIFubKl+MdXKBKzgda9oC80F07Lcf3bw/5jinNYG6UB5t
vg8RujwjNsR5dHXNG1zbbXLnjcjUhSllE6q6wN9t4QnF4RrrR9nh/R+BQsW7O9M1FiMU9XEyX7Dh
KMHRBQUyOJjFYYx/leKA7psovFOIc0jTudQMKlN4Ut64cDaA+auWLTas8Wv7SmuFx99a9c+EoLKB
iagDc5ET1Wip8f+6yPm310uRC4cw0vu4EW956S5BFXx7Zx0Xh+l5/P0XlbEN1CWB957YMcP905dd
i97mYpcZsptjWI9Ak42GFUVFt1QUHXcQgXfStB1qhoY2tGC9xgpYN7WURQiZD+1UVDbzMGh/dIdL
CUOFEDgvfCy6vsvlYBHnzy6pyqdMoDAj/pnOSweW/XcOlpz2XhQutY0mS9RjkJLG3y0JNjomw6C3
d1seRh5cCRAJ+tA+jsJCGhsAl5VvfVX3fWbQnr7DaeDVrvxu736Vj//Uj3y9ufK4FDuanEeHW1J3
M+x7JWBS4aCKNTtrpthJH2uJMlZt19TcWt5AXWp2Wa7cFSIYdbsXUdx8rFZ+jVVL+SV2Y7XKCkvd
SxZpF/N2IMUAgxxA18avW0bm3EBjs8O0LV/Yhebqc2pbPQKS+7StGUcPT/JdWQrIJynY3lP/T1L4
IQcOVY5RNgku4tJqyRrXYjDaIT1RSnaJujXrACsDKBvy6ghqd/zZTc04wt32yvlmuy+j1IEL7iM3
bFbtM9leUDDfWF+DrIJed/koW6pV5LsNrcCoa4ceel/LnZ++6zjWLfN16hY1eA626Jrbavdw2aa6
s0Zjc0HshiinXTexVBRn1XG7IAhsyRT98u0Ds9vq8TzjL9Ea/S2KSUSS/15surCsiVi1MlNYCegH
KdEl2LN19VAWYJb2983C4Yo0+fkHoxgCurw2ToMfjY1cnZzh/6mk0yann7l8QZJl9cUfpjSnvQJN
IqZ1xdZd8ZBHElN8ODQp3skDmntmDtVs/2jIQq8VblGmuAhtGD937gjrTJzzcJ1ZnK+y6BiDercg
HXos5xQOywOHMvTjzYCinxns3kd7xspQmkqobt4iQp2vUnl4bQKo5QkRVz95R0w/PkuDPiMrPxdg
WsBfDFz9nLOXkfeWKbH5sW0jN/EQK/RGT1/2qRTkiqIupN9i06HNFgv4SDmWm/7bBXvRZ99KWvyh
Jc4vNklWsvv3qq0GRmzEJ1R//91HtHhWZzy3YrvvbrsT6y8z+nYkKoNELag9TXf+XjqryOjsL5xT
Aes7mbjkoafk1g+gxK5EUGa558fivSWYj/FUgRFOM/fjp2zs5dH3Vd+cldTIk3jLyLGJaNeFUwdn
R8ooVulLSSDAVC3LQVbDnW2XTw2tAcPd21yOE0mKYtw9POMRKj9/jLS+f1Ain+S+CTNMprlRDe1K
gNwaqRg5bPcH85EuHFMp+PBT2mLjRXSa67ajPkoZyKJUxlnrZIC5ym02sZLe56pptTxbam73CKON
PkflGVLR2mxZqmc1MhDMHlhcqWve8nCHdayZxSBbKwKm2cUUmMPO5Qrj050v/R1LzRuBpf38RYn+
TrdSi6g6qii6RvfEUuuyhkw5SguFuVu9wkyhxOJnzqNiGv0TKWe3NAWWTGDKj985AfOcQ1GptSst
U9wz9gylhqPsf354ZBmzt9p5fnbPk74LtSNOAUgDgBf2VSJZIt8evOcMvun3Uo55Cr40Rvvz8D00
rljBtE/kkyo9Ib3WtJSPtk4z0cql0ULggwspWoxPXSV0wTvYNqm3dXeXKOCP7sSajH4QWiyS2uwa
DJ7rnB7uKy8+gHCfmrvjC6enckKjHCO+FIF7IS+Dv1bWxKstOmBhQsOApKMr4b9lk0z4QLXFjNal
gE8AU7DVhFqaNzDJGkf8RS6vpWiA2DTc1qz/XPP1W8/ziHv8EoEbRJgUqpkWfDiDyG0FMq+Cjvhc
koEuyJnQDHxXEWGFKxeTFxbw8Zt77L6WYnJffsvyQzU1kbGKbAg5wqRPqpEFcwtLHNF7f0NlMIW1
Rh4WqaObYeywz/w52w65o/ljanbn7XUoEvwLQr7BkRNkpd4KFuj22uQ5kpHZTcm7hb62WMuSpxNC
qwrK9nFP3FyZhKuDDQQwJ4pPyHhqYg8gK2b9NvszFEBLzLSlqgHYmWJ2cWWA5aODLoAc2GySAtpk
lz3x1li2gj2YE8Wdzs1kSgxO7XSAAJbMwdltLVntrhEudZ76U+2D4jB2LVFtwchlS5TY55P9sY59
0kyuQcepH3y7lWWXLOCIzcvSmO5OIxQRx8QTdrLn5PSwcCu8mu1TU7fFFbmvUKhbsubNxInSZFEH
M54ZlhMxBQWkfgtkdfToQy7WBxjhHezAHrH0KDryKcps2/i++I1yUSpNQudo4pHxTfR4L6cj5cz1
ELw1p8eoYqO8VGfc6m27+CLSJ+w+wqYcuI5rRwh+LFfEZu84RI6v2itw252gkTu8eWBsWjzbTRV1
nL2NFY2+zPZ5C3zCfIb3AC8V/RlFo1Lc74HvIK4DBP4pK94dGUtkRooxCaGtCUKpd+hkrV4BNFus
Uh61To/F4r+XT1e2WVOWAPfGxxPyGJLPT0pJVVfcE4g6/P2mkhnDD5gAMo/2Hb1XZlg+iXOlLjT1
3j3Xl2kPZ8A8GmLakzkRiX/m1UTGNon504S2078XLmHmvEVmXwkfh1WtPzNDfFPfCY282kl7JY2E
reSLjPX0XaYORIkOMmeuy4Ix8LQEwAmWc5rswsIM1cTs96+uyAI7LLHAPYo7SuAbIdCpmIS30tT1
xhIolnKNctTueQYqRNsXjkfiJG3ilhSZYfOLS7UXqtTHSwIXLX9kEHbddkPYwJoHSEaZ9ZpqylL2
L+UPYSN36ywBDKBsrfSo4lnASMeALSKJhphIvNPQ8xFkJ8yKGTqI+e4GgP2jIrCpSIBUkKhrg7Qs
yOVLqR/hHLD0YBuigEidIn43REwxAYCoTCvxE52YyA+bzxBecCfqC0lEwzCzLtmlJbPTWe6/CIz/
Udq3khw+XNeLrv1iX9L6mY8IofIiPauRxqbEdH6lhVw8XAsj+S8AZ9d/+B4cTiZm21opixsLO2yW
TQQ8a/mNzaq+54ZeWMrWizExagf8u0u6s7OV+YM10YYYz/ceP+Vn5AUejaiyiZaffbF92qRB5HFv
XIqtbEw1DvQkPSIwbt10qftW9B6OOXkasZKHHW7lZXIrBchxDYesknREsrESeS0AU0t3vOu2/+RU
Yg6ju9N58RSBwFTLYzXHbui9KlLlnSGsDKmw/DJ39ZdualgD0gsVv0UTt5oT+KQaySbgiJvDNWnN
P6e5BJFp41QW86nt0BgNw5FT47XWCfOzzaSJOmUdF9Z29f/MV2/Raomx5zfcboF+LTY2IsMBtJAE
t36BJWp+cLqw4c/tk7xieptE3a/Zsk1hmTf86+d5QSfMnhkGZULLHI9q1ed8FE3XhEF5RI3Z6UU8
S1JH3xyd91Gs8A0eJEIlzBR/+r3YPuAWlrcfR9FAw9AsbNBnukoQPPM2hBShBGUb8mCRuEbOM9DS
1GbmQ9XITAQt038GhdvOb7gMAo3h0MV5iLZZBY8NPdFmNay+Q8ZvSpAQJdeLg8o4ku2fTvJfJD7m
kBJF+QSMgepLaV2SQdcKcSU4VFCWMbYl+Nx+DO5qRiwLUGmxJPK+n7U2jGRmAn28cnLBO3nUbJZN
ACNZx1BzaOqukDAJOuXSKan/BRT4y0g2ZykiAtShmkoZ/6vK3sOBdpDED9QpbQkWKDQr35DPO7bY
2/I7syrhl6w9erZjSRKy1sWUymP5bQhoWd5BjJ2s3QQdYMLDNm23WMf5bnJ7MERP9qz+8jFH+C7a
Ijo2Bae+FHhBiZOsKKkWC09k7wJEzP/zB8YfxBkhZn0ln37BeRnuzZyFi0Kd9SAbqNY+w+qSvrHy
4zK8Tvm5UECeJ/zr0CPo1h0jUz7ZDC0vODVBHrEgRFKYTu69LKsxy+8oPpljXxTsGfhOG/HFxQ9+
EKqPnx01HJ9NiBC5N/Z3RSnvCtiPR0EQ1VA74MyUFPbPxKPMiiWgb+f9WVc+sKjakO9T3z68ihe/
zL5lGpmJAM4l5vPTndWNW4rMsB+JuRMzAYP2lBUzl76NbQL9Ej3o+YHXVxztjp1f4MP0jcpDfEoa
3mkcOcNZmcm+ux/YbjzJTNFDfn1qsS7JAyv2tT026Voba4Ol0VWegDOW7HhlBnGaHRvKEnpE8JPd
60po1vpoLEbc3qoeEjdDmgm/GY95vH9Uv+pMDHv6g6qPJbrf/sfJ4Tbp9+HqVQlM3SygCEOsDN3J
UoL8ce1CqDW2dedqzKCHFXoyei/HC0Z76tjt4Gk0nQi/jrvfD0XUydZ1sto8IwXx7mEdQZZgb64e
OoJj+1hh4hUDQhKISu9ElB7Alh9fk8/Yy0p/C9LLHOQXTvYqIeU6amVZSI0YK1AMRVW/NZTwL5qa
LJOmkEjm2cjnm6+T7F5OtrE24jD/0d6iYd2Pl1ZMsnznGmt1/w50iU06sig15/KX1JDWbQHdtl5e
d413FTYIKsiq+l716I1a0oiSZHETFnzSZ+iOW6RLsUm61UfqPq73ZHTPSzHs9A0txSH96/KSSoHL
vd5WVbcyMpkrTbEpwsvI6rbZa9j/g+r4FdJABsgZkUJji8vsTIIK+JIZrhVBn3zZG4D1iwYhzPmg
ciKZ2mZs1Sl/XIcH5VZmpFLDHdwfRO/3DcmwvsjI7BqQOwQhssvmApRJaIIvug8fC6HT+NwkuUfC
XYnN7kBdLMhInWLhRHYpxbxsca+FY/oG9qz+IjtDy3oU4r4sqLG8u26t1vlprBMQXAVQsR7MqQYI
H6+cF4GSdfhBzt7yhlCmIw0vARil4pUwDbxQsoe/LjgAJUoN1Mu5OmFJHduw0ibyiviW6X6jzKZH
gbSRUb/SxucNUW1twUQk4UuvqgwY9MjrbP4jLfJ9inaiMNlBmVBDKgpXABdm4JBQGkfvnKwfSURK
mNlVH5PgA5fLf0Z9nMOeNJD+mjQybh7FI6DBUSYdT7+MlPvGT5YeX+5tX8BeK2hqCyEMEerp3OCL
I/zd6t1PoByOBuMYyIOvpa2X300f1CszZ4TN7WJe+BnX7trQgwT8CBTtJSAbb8Ij9EXQqJfvXD4d
2o11BF1Lg2fInZ2SZjMK0yUF7sWyxf8USsznYfdJvt2wktd62cf3esVqET3jOL5f3p41z3hMoNjI
UX9Z44BFO9p8/Lky/3gBZzrm8k0TPcbj1uWHKDmYyFIEOGFjMhyC7TH8Eb7g6khdWMbN5RIseiH/
OsrKJoLdwEZZrgHX9cxqxBLBUlJVmDfCBa9ayNgwA7tLT65aQn1uEoHBeFmVZQlkCVJhDOpUWr/t
h41dhCIGbiwGhf1ed4Y8yeYNBHy9KHAavFSgNXKNVFvZPcWta7hfE07iBnDoiMhQqDdQ04PcmAYO
3SVn0UbWw2T0QvrpwOPrZ3whirABn35XFhYn0Z9RfP9eCLkKSgFfZt+jAhHeXpfnjM/kt4dW22HB
raNj3qD6zDqYjYTYgIDpLhhLa5fX0R8w0/W2RHtO9A5NP8tWTQdt7q2QUttN9qOx4ETVv3hkHvdx
omYCpK8tiqHZaLmcChCTfXzxqva+2etVIulXMp5E8TnXs9OjBRHs2f4FXe+rTwIa9dpJFIsVYC0a
UFbNsk9WOX0JfkAxHYHotlmkoHYGNqOnf58RoQ31bYoEmbj2gs5/NMUMO/I+DwWVn1n9Wq0DrxnY
SBB84QuRrMeltZ5Po0Gt6H4CZocrv/HoviSBqeJtouOwcxCgiqPD+srih3gVeWSRv6DByE51shd+
dnaQQjKsJad2AfemIiGE43vinjZI1qybqGxIJhUzL8Ge6fn5IyWW0LgQlQjRw/nnCd8l8W9Dir0R
sC35bXv+ZWFPNIVSSK5/+8/7dFoBM72XrPJut7NNDmXB5zueCtxAflx1OCTdP0Ebm3Em1TeOZMpM
ZLtqPnyinwyQSNLt2D3UKTK8VUEZhhs9Ks5U6VxMR9n59KMahm8ewYnJf5s+xNVVArCJS3++/wiB
mPERDx9uMnURG1a8pr4zgIQ7chslQ0fJ94hNY4tsX+k80Pb/eSGhoFH3h/7K+RrscPcfJicZtrAu
t8MmDvVaMZGpauTIG6VbtM5dKzTkqJdeJlwFyASH/Rib5R5sGuQKf9+PGqNFE8R3n4Hv/zMitUor
qAhbqjklp7Bab8DCZGhfidLwl71lHOMKBNhTeZTZCyqSawUs0kqLToOI6uAvFJbaSyfGgg/fe9wd
WhZ3loMbH/KotcGt3UnxbF7q2H5T/TtmwgxMna0WsQwJaDcEHUjyQgtf+gTDVdKPvoK1wp9PgZu5
BqbtxgXTnK4Tat0FHVyJFUuW743LMVCAQyMrK+OvfVEzj0lHF7uPAaOmNvibUlnU2Zk8UqnhxSqe
k+td4ciFCkjkqSxnRd8HjYuWWKHqa6DYek7UipLu133ufbtpL1h+KrtnmF7jcZw6mwFbNITWWYY1
VUqjc94wGEQUIVJfo2DjeOEEjE+KLJoXbQTSo9AVdcVRK7qFAHxbZk7JMr3roidSal4g+DJiTSU/
wOXp2G7q3ge+MINPWpjAiXnzROo7fmRQL1ypkmqSSaHMBWijWSKouWQNyowI0UKALf4/wawunZGA
hzR/c71Xdg6HzZba788v7BT5qojfopihqbnHh3R8Y96/7JHgLEW+0y6XcjzeKnGBvig6yz3rmViE
zfR0ib00Wmk6gColmeDUxSILqrJHb0xzjyyKvc2fHOHt47+s7nFHady5zicKhliCG3Bjitsxxd2a
f9DWA2VwpyL3V3MNGNtncvSHgLOVZRxXO2s5Pu2mhrbkM2U3HPlmMX6MBGhE5sXQyosWJuX4t9an
A8j/rMbytf3/Kxy78j4fWgK3qfVOZW2DUTijAt9jE8/DXNc7Kaikh8whKKgFgOINt28CXods6PiV
DnuOinmJZmyKMQf3n+zip6AcmboNL59fRB+irVeOdbSZ48awKYzYQlNE5XCA35U14GsfAoNk/R89
I0suedcvWo3rxQSPD0f2qrC7X7o8oG6crH+X1/P875dBV/UYCxyqmDJwCtjzvlGNVGRFUrZbCrks
tCUaZnHr9gVahDrDbdY1CQb7Ylzyh0KdHMj+JTzjJUjmwHPuK0rOcbi9CRE25XPtTF6bsBkkQVQZ
fLy9vtc97751UeFaCyk6ZiqhFx69GrlDFG7qfd6SntTB7Mb7/r3SBN2N2thFEa7kAIXvo6romyX1
IkVVFeADcBhtb3PmsUPEc0mzoUTuw4xNBUWV2VFLZMuTnc7Mt5zPHC/g30dvpV/vhFq8ZJS3SM3X
qHgcJ6K/rLukdpxsUNRo9O7iApaB2/dKxoX6kzV7R5G6MrRfUnIwrRy2pGHKIo/mUvIuIlZ2hzBC
B9o6o6kCO4Gn7QhVMBvhuJYsVq4ZgujXYavaVVIIojzrm6EObfVI7NkEcOSv7mmbICqCphH99Ykh
CMsYtdLSa99yvRphs7LpyNtUqPzmHlLQ2nNUkRn3UxTOtGnb9Ju2ivHVTsI6njDnbQ5NEfeEmqo5
IXwEDcDz6txoyoUlA8FX53JWiTqmRTtB0Z2Wt+7ZgR5qpSqReAuz21H8P/UBfmqjeyPeVp1UOYBp
fFcQM2/7RchCpdjXZcmfumiUGk0ze2f+t51c8qZ94vaQmC1HOt+KOLXctbruO3qN31vsl/Bwizfk
h2zcXXQ1QV4z4rayGKZWz+0lvlfVnxhAbnCopwe7KYwqwemnuuRlfWUdYZYSiDS43w4gl+P6zHP3
OYpn+xIR9rQTZhTbUiHkZWdP3ZnrQ1NxN9cGIRGYb6R6IMhrMY3aDAq4Bvz5Yf8YREihYeyfJfhO
p48GecP+2KStzMKZC848r1o0WgqfatQ0dJR/gC9lCIQUnnaJhoZphP/UaOHnkj+JsFPaKOvJ8tCK
yD78TFk8RJ5kwrCl34llKDvjEWArfKM5Okm2heWzgYwI2lQjWibOuOA8B/bcd8c66CSLbt+73YLo
TAqEO/slcSSHt1uuIkLcMy5MbNeSGMj4kztMK6a5TpOAd/4S3Hoo+j7hiGQ7XcFRGtMIayRChivE
YmdgYRp7UZyEbgQ5SXDAj0Vom3HHn39KaWbvMOBJdvHTzrHkgy2ZUbA+okTQ+JC9vyHCPlLvmmnx
w4heekAQ/YOEgUbcVc55CRzhQzQ2nHSe5qk+kBG4Yjby481c3KJvQ1dhzuMtoj+l9ITmZatDJECW
lQUodNk3a1nAR11XBGfHSGTof/JvGy2uf+eg0byTOYFX6efghAMea9b7SMTnO0IJdPjxn4i0dX38
Qnb0sLGEOL8GHQK/ykHB0VskyoGpTVjXp/p3IspcopQkJR0O5SZEtbjbshONtkD7J3nfgP7LLa74
xZOiis9oBqZQvJFlzGI0s9ROJOqgnWr320lsgINdkWHhiY4f2TnaXnuvmlkPf1/UzRKALDKGZvsD
62Gbioip3aEkuA4UuGc/nAI7/oklHkaEaegDSVfbA0F+zDoasq9urXlEqjLFB9OfgYY+j5ij5drA
cU4g7HU9W0VWWNVjaE3iVXJuMlB52cnsBA6OmiOzFmaFb912o49UYE5UzxyJwPCBVXL8C7tvFDpc
BLNM6Ak9KVwHElpW5f6cFtBxpaU55+9GEOWBUSjdwGK6UiE0Jt5xhO5emDcRzEDCF6i1amgx96Lh
DhFXsoZqZ0sd5xCo2YAI4DqALbMCtXHVTNk1uRiuRihw7ap91nVZreCQ80Txl3XkdHl3FMZIBvMJ
EXyhZwKcUudTsyRce8y/bIheva1JCXr8gjbpGDrw/aoMiro/uofcpbBU03Hs8kHkMa+Q/DYStQ4L
OZfOij0Z609/uV/yfiqbrAdSvJejOK+lUdR5trf+9sQRzQE4AcDhOREj80t3q6aWKc7XQrVK7wy2
G/620JaZBrMinFBjzC4QFRAhZl0JH3ADwzPjkl7y6fGZa1iXl9gcUq5aKL0EM2dFw5Z6WsuqV7r3
NZM/tfyj63w7c5cDeiJs+luPjHw+yZG4EAvQ0qW9MrQvCy4ZwelIrzVSHIJ0U4XQHxn5zCFr/us6
08G5M0L41fxek+EA2Jh6+LuuLTjLTHrPmem7E/O2qpEZef1A1HHg18tVKaoE2ee1Lz0V2lXUT4bX
fEdqIO5yij+oOANEpPTSljgxRT4CXG6k7aBQtN0/8clGgfdvFbXlkE4s6tJm3VhFqFYyxkzFmPaW
qUCP6ysFXMZ6YLCjS3bIqB/N5PpYBU9CzuTu3QaL9DlxV9r8HoEcCrQkNaW20WC+UNt/o27Cth3R
r+JddXmFd5Ug7X0hwLssjgl8Ir0JYFj36lW+mzDjFRcXxGx7AyPXMTNsk7AB2W1tKVsY0Cq8dPvp
CyrDwVrmYTkGtKhQT/r0UupGLlALeGK0jhw+LOpswEoqQQ7au8AFQTqDAxq7ib/qdKUqHAfkBDfv
kNT9FBcP351oSs87omSlFAPdFQxWI0CLOZZvxkvvO9BOdJl1R0BXgbR7m10nh+YC58r58xZ6DOLT
/nQfB4CvG/DChDcQmFk4mpfa+penj82K6ej5SSkIDHpzxwlIz4lWAPn2CpqpP8H1QpSubGFVIObr
YmyUM0NzoX15P17prooEU/qO7cQEut2Jvu63vmNh62vnRWDW+Jl/HfZWOblviza/c+ChTWSDE9lW
QhUlQuAaHwCsgF5mM6h80sqTlbin54laR1s40OYoRT+W+gyfxe19Zy5ket1DOD51NrTASC/ca0P+
aV6j1tBH3BPmE4BoW9zArhfBLRXtVld1l07KFUQb8TbVlg6GHYmV0S/8SnbKTobQ6eye8cH0itEt
+fYp9CeBx7MwjSt/9Oi8uhGD3/KtgsnJesE5j9v3ABYLIZtoPtTM/cCsbX/sZvuHRKs6WXUSJj4u
DK5ud3tcLXJvYpIaPcI8ANPq5SSyleoZZDI8jfnKm4W6wYlIo5CLWpFGi3L9rojAwqe1PrdEUEqQ
qv6jMi7pz/iQa8CGvDpLtqRwPc0wzNsSf35A2wrqm6Mpb6DCug91C90z9+TgdEVGHbeZKR8d3Ax0
XanGTF/JVlxhK29TAJrZRire1dfSeOqxD/GqwpDo8ErdfJ8wNDOCIqqeDdH+DnVEjBnebTGqy1VJ
1x1JEpBduWYKHBcjdhatCQNPuqo+2zRqhFfaK8y/xGa49icuN1QBS0Tzpw01BzYZU/h3SEuLgWdf
p9Agc2yFFs3iKDFjCVHDIzzy+L3dG9IEnk7GMn+ggbJWrxDPZcSxCGUx8CUoZS/MPFxfABhsle+T
FZ7vjle6DBCUW1s5s/OfPskRfe5i3g3bVaxlPmzJdM4vlZ/Un6Wj6eBghI/R53UES0iBcJGwn2+4
zga7LL5rr87vtvSSa0MSK+HsHa9qnoXd44kImhjPPHdOzhuMgDgrZn77tg/85D19nW4XuGjTLsGY
H0YVlq/XUAHNvJH63gJbBV8OeOjCI7FIqR2bEa6V73+Lqcn8J4u9DMHpu+qIVgFrhQu5RHNPfu2f
SRdLUc5BwomXbbVLRp17gziXYcXYCVJbadXLg/8pMNLT6gRdSdpte/FnCkdFjnHOor0DL6Omg7SI
D7bflrfVLEjXubyOJYqoUSIiroJhVocZJ/ox5o2kiEy4xqoOej004Gcpifh5jgEVvnLhJhhXwnKo
487EI9vpX+LMrsqKYn8KQb0kkgzfHmwKwaRRwe+oczHBNaknYV4QlP3u2MUzZpqEpf1zn9eCPVan
Nes1OhxRXOEj0m0VDXXaOy5V06qw0yBWmcKWeSgSvYoNwUA96JKhL9qm5qpoq/LZjFE9MkGbDBgA
97Uj7oJDttSSeuACGjA2PJE1gW0x4cgfd2lZzuBK+c0X0mSFKYIq2lBt54QPzCsyTpTUfq+zPrM2
U0ehtZIQEj5qlrGOtV5+ehBU3YfgeCtPgaxypik4gF2B+l1bzO5Cir5k3JWuNZG/Ss1RnggFRvnt
bKGKXBPZp7DvU9Fmw5OGvg3lW+lqK6GWJQzhXoEDUcIsDXPf7YGtdYnumzVVG9b5kVoPI+rKR1oZ
uCFUkgWI+FySksqDhhZlt9o0ZUMwNlAIfMr+qol6ixzjwQRc45DcpJgeWgmpP5LmxVgqaB/1pjqy
90yUEC72vHXzw9+udnwr07YhqRBtiCdq3mCyqXibil5/sCrjybc+0T4+F3X9ik7xVwN7MeGdVtBS
OFdSeiBmka5vxUCRMVyOTV2tigzr26UGMSY3am/ehXo7lcnZ+YtVoIHseVLD60lriTGjcISMATUq
4AXlx37LIin32OKXbxfTdEypNn5+NEnX6pDdm63UxTSPIx+/uUZu5mHu1PRcFRAXkeS5ktChmkHd
7jkRjl5v6mLLz9Vgw1AmLa3/iGaYgGNB/gsj0icUeWtiuFpWt42226ELMRk6Q0V68dSuv0R/zaav
Uhcm5Kegu8vdKz2c++/TzpTqa72t9otMvdqXXt6n1c5vavihhJTARM/dXff8w1I/PP8QzEe5eQF5
7+q/r3TrCHU+nb4LYw7Upjrqe3aTGdiCi1o30YhORpEmYYw4+kEL2uhUpVmCE9agPsDdM19B0lcM
It86RMwAF1nh6LiXflts2/EIn08xj+CqhRQ506ayur004/vCnFLJU1u2kHyQH0UzmO86rZv8yuGy
xXRFZ6+TdEZvtyFpRF4cvLBU82Tyi00yvZHpp1BS/T38jBiN2PJ5yvWrCYYOqyDS7+157kkorz1a
Z47kJLyuXmZrNomGgzygjnW8mNP19N3sdbzo7ztHDtYAW2pflgzZvMg1S5kxxBdDi5QYT0akmE1u
JIHl/3bZhfjx8+pK3koWxSvf/QqdfFjtw04jfnRAdYu2YFUNepxuDVYBT7qwQMgL3YB1umhSBhfy
bDOr171Y8k849p5yr48X9XtaIg2CIYIxQG2jwJdX3YkT7x+j2Ev1+zMJ0C49mp5+mcafLqdRnc3o
OxxletWWJRKPAn0UpWn1Hr4njjv7jEjP6Q9AwH9VJfVlOIn21vkgjMr0XJz6E1b1iONedQATm+uC
DgWTqdxVCyW4t1E30Js7uM217AxhEOUNH7MDfYclB636517CK+ENpZki0CyMNyjYhY2BQPHdIgOQ
PlxBgMCb21V3lyMFYWNXoiw/zlvdmWgpxQaCjt7tenCooEX1Q3aMlArK/nJRfZBWyWVBgK4kBZ3R
hSc5B1f84vq8MN9OY21Oz3ukmowDUBIyJsJ3BtfGDyOYWiyxtZ2zWUfM7wQTEZy6pPrKXohspV+q
Avjz6wuouyZSlfPKHEFYseQfRbfz8Vl3zFLmk4QJiT0UEscapKxDDKGAXvcnnxY54pIhny1QwBLi
Hgbn18DTSg+MtP/bD+4XeC5mVBM/SZVJq7AJWfSpoRUyr0QITKiiP0yZfAgGYM3AsNhOD3Iy/wXZ
NTa9VPvNH3u28+eE3ih5UkfbtntBXwgou0qqhZaVtcU+rTlxtpqNwBBAlUH55WV97vncHlu0Wloi
JJ5PS9FPOajwKySr9ktV6mnfOGi1bFGPVwbxHuL4NvMKvQjmFz0CGWZBgWWvXotmQHEdYK8BApfT
TUhXohAndvrHptdMSXuB61V+3Mb6BOqUBOYPjM19adcQhUTrkrbvpkzcYhO8wVrIOuZPDM8c5JXw
MUnuOxPtZWkoW6HTFygjeyPG2fPruNaX6EnsfBU0MG7iWxydvy5o4cm2RFy2G+n1WN6uOjWz780W
xXgScZNn8AJTT+cTcIpyYrgh/scyExGpf31E+b56sF6F9ZYGnuVNLEJRijg8sY4dZYYDKcLXWU6q
ws48My7VVVV6LyetK+AqRQKPeVubdD757y9QhaMRrPqMAPyV94h7SwHH/FfS4VR2gJ0bq0eT4miO
waZsmPBzrdMKI0XH4DjLulOVmHSoLMrgkVHhF2tyYInRWUv9ACpSBLm7HGbGJCf0PcyQhHpm53ST
u7pm+fnMb85IrttW7iW6IiJgNLsPZqyYPaNpGYb8sZpCIdUXJeRRrbfU3uxXdhTwdRB56pcWQxi9
TeethTd423bsTSWYrrjiRMN07t9mbr7A6aiDGqaeo3P4fxLc71/O/EyGTJ/1Dug4R4x/YsvOiPFR
eV5qKQO0Fr72eYE+EU82rD2tRO47bPlfNJdJu/m4y/sKEdUNMll12Vx4lCrcC5Y28MQpbTU775Lq
S6NJjcEc+dEooTR/a1kJRaqDhvu+OwMClsXL0I1urYBKwpv3xJfEw5QMi/L6X/OFefz2X9Avl/tG
B8ziypQUOoSZHJXXzO7RbUWxoATq7uxUfL9baTofg3G1XHG+3+TcFWe0eN7vSEQriHWxfoKy9WZH
zU77QCS/3QoYUBcRnCW+8d98509W1IfoZOZl8wI6cJCyR9V/mTvsWXYFsYaMMBIGwJ7F9OS9JFUu
r1V5R1qXgJZ+74laDAX84erxdfaNt4s2KlEhzsKxbF23ipdrWwSWAirhpm2H1HoL3jTctFSNjbbt
sW5J9Uq/khKiMAXIYs/toGqvpHv8DSpY9bjL9QKpojR6R5Kumd1m922aVI70esOj3u9U/J2vAExL
qQBYfLYulMe+rSPgM8I/mb2foZUw8R4FYfU2++aIhmdB2R2hZwEcs2GoRecvbucd+uGztzGSt+1b
ZtxtdzkeUP4S3r2KAulJ3QF6k0YiPePPAQwtqctkRiGMqhgYtpsaqTT6GxthL25gUdM9mLZ55ZAR
RsqYKQwGRgDFv6H8OtmMubwdceuqbocMvluIrrjGvn9xI3t1Ef9EycebSod+eouoMw4ivVk2qUuA
C4dIztsLJkFXAMqWW+gA+3oEWWw7p2hZsH/LxjI+UUkijH+fA8vQlOcernL+jHjrvdacx3uvDW/J
ct5FmLvPM02mEtwf31Xy4sQ+0tI/cxz2w5Flf/ObpfVcebVPBQt/xVXESOS7226nOBwfcGq1feSf
mGX9LLXW99Mz56/RplPGCMVRrNX5pD1fbFpJsP7hwYKqF22r+Xa6MORWYlqPB1pycxoiNW+Kr1a/
xFOuHnzvpiUns7h/OwSQ5H6iUFsyWeMXuajdHOA9Bv2jHpVjbMcPhI/DHwQkD4Q0zY/xYyLSZCC5
4ipvm9oyyYuuO+R292xEVj+WpMu/7K+kKhLWEVFj6Zk+yHzIQBYoTlu701ZLCiYUcrP903BOuU1H
327yy4DDQ/ufeG083fujJ7UChIxKmBHGqUOtMyiFbmVt9/1XJf0ElRMqxOwJDH7F/wTnzosAf9aT
9ACQKpBXO+9rSCHnBq5Xareiff3FG69YyJN8Ekc3WidDlDBFYZl0GAr4MMKD3N4QAqIxDmn5ROa/
XB5TQysGXBURpGOYvpVTl5PPMo0Us8Zjh4ypwdb17mMmNzeB7kQEGGX7JOOKO8QRB4qIi71mzJS0
UnWGmCGcmtZiBSOWM/KKjH6rKuxPD6Q0kbxj6SciKNg1tvP1TnSMt2fpw3kIBeBTFuYf0QaBcL++
AIM67xdDXQp6433f3SXExLtlUlzCSWyHO+YhJiuWGhrE464xReComTdWdNZao0Qc3hp1Ek+WGBn+
SBqgb8FytNkQ+4PYfCwF8NCP8sYNFzaXvgbBPB+CQbFPWgZTD0GxAGWrwOXNG/e/FbqRPdCSt/Vo
yM+ivjwC9m8+i2BbP5KLNIHqKcAGZdJVFlHSDc6aNA3zyfdxOKX/4TG+sHlNxVN8ErRFbaN1gHnJ
Q8LRWIilpFog1mnIFE/pXSA0lK4cZVUg/wDq8NYe6VJ8YwdBCcmpV4EHCqDw6g9y/DopmoevHVfb
+bOWD3e6E4WdI/e+Xmx8dafzzwPYzHvwBlEVq27GqMtigbGFWFatH1NffEXQCQCFxuV4fdT0II2z
RZRLNkI15PuO3JfE/DisurjfU6gtiVZjxb6GnZm9fswiPAEPfspwtsXcNwlkJrJuW/V0Ig9uBbl7
mnS3Adxg9nTVXxxRxKyRvDWCWVdxB2U0VMix3U6NzMbi+Ei2Q+M4mKqnxzh3wu4mQEs1YN1KdXS9
UWZmYcPXkfpApFyQ6ftS8Q1+EzUxsi4BvlFtfrf/15BBMHGd3oninUuZ4CWCfDmonLiBBJckF97d
NaBmEi3NE30+5LEtIAC4H6a9L0T0h1jyQAJpe1F5R15hh4mFyRP9onBs3K/cZE5v0rBNwbj/12Vm
LbVVPLiOJoeV0D/Q/cN/HK0HqWzbgyMVSewmdVY/hMY6wnG1mNrE6R8vf1bo4wQG/cdBES7xvMN0
UBjeC8wGaAy8GOYWJiaNbgUPzt5pVPXPOAf4E39ATIvFJ2hfZhLup59ESt2oVdncsP5JIrIhXZ3v
ht5BeQIe1bqu4744R+DyDhMBAPES7Gc69wcDP2P0JLG2CGO6iijnm8bRWZEo2OXDbuVZuFjASIfk
Bli5ljHoT7yvfkKNxdtP+LfJWlMsy6YFpbsjxEI2Q0gCQ1tKU3gQR0wapUB3GZQlyEfiexmUeooS
i59Vj47jmK/H18vsQmi0aIyrBh5fhMNU5FTIju5KeWV3RGqsqT0jVs91DfjSf1Z3hZDXz9eszcbd
YJjrFheM8avUzGgJbwVNQYlVh0f/i6rSBmJ5wt9UEQrmgkXGJcMecptKnJNPuN7D4mbd1A4ZpUFG
aHqwspZezZT5LYDTRs1CyHcJM/ukn488mTiC3ijfM1+Fxj+fXkbWzoXg1Ghhj0847kUtVSQDI+4r
IpcRO93/bozhcBQ3O3JrLNYNZnK2wQuN5qfuvKgrbXiwskPH4qFz/NPm7Vk04dFK5/pLikkpQ7a2
+wOGcYqgFJIiBshuFAWXpG6YyJsIZUZkM9yWrLFhnUP8fHcNgdgJhVnZttM0KCUD0VedbZhPgG2l
K7viDUGQdOHbnUH6/x8wj83hiwnxGzYdFWO46HITooYF8OIORuZQLh0vKt2Nll49VWs5pWXKDaM3
reDVaE/4IInTR/TPZ9aRpdUJ7b6vb96VtYcWPLh93Q+FVIALAeFvg0OjBfKdS4X+IilL+qj0NTL5
owrYcqnMnLVR//bxdkQ9WpLdlF4e0u/p5Z6J0nxLXWzdZ8VXq82YKvrReCy78chTkJ2FDXvhcMf1
LraE3PQqH7Y2FIcWAZbv3lS3ahJFJ/LU0cTHOEX7p21X9Up7KMB4DogYO2R1WTkf587hgnRA4aze
VvFw5LB6ugZwcB18Nmxd4rZEHtKnEl/2I/ovA9wyqejDRiidM5yO9psaGsHj6DP7xltXJOJ8gKtZ
WRVwYQwWcOWvq94rBUqo0X0xup8kLVdNyTWId4mswAH7N8iIixcYJwfLXo0l1358ZR4tebAJpklJ
ZKWTuD2BgqfhOTRf/IsJ5eTzOeUrFEZ+eT7DdnsEBxyObmbtrchpadRVGDrVh7fnP9HcMu2LwLI1
LG9OeNHDKuyLG8VuiAY4584wCYcnAQTt2qSyI+X5yLs8gYyiAcHleD3gLMFZWPrih6KOLpWqmxnj
lbr/+zjui0ozVKxcRZN5A1KsjyKw0GGv4DtAQ7KrpUZTtG1QOY7CVngyfGu9f994b8nf8g0GL2IQ
D1wle6BNHVzPhy5ArieIJqOwUciYMhJ//QAZA1Y9iGEiu328ugWSB44Y7xYrDcoeVnRTPEPTZJFM
2dJ7f+5WJa12rbS/oYMwpgaK7G7vXTsz3VHgjfB3DN4vRpwCLNmYmBUPqn+T8L5FQ0S896ah75ur
td1BhVqy2fC88DTbNX6yhA2H+VU/XNlwtcKRwl0yHBuEKsc7hVFeuZyKJj8YwbCscPW/+diN0u75
f5AGBSsi4mE0AeF4sagp8piSc+AEN3Wu9M79IARxQn8R4lEpeeP7Z1kHrzza3ZC73+cli7iV07KR
OywlwM5IlETA3/2299TkBF1T/HIhZ5fYfHg9ETuPWWuZh0L77E2m/nekM3dEsKDqnD/FCaSH6Hrx
6AEQ762Us52RrvamsSwp2/QLd0MGPo7jQ6k4An57iwX6AHIhiR6hFjW8UKXvVQ2kiLHTDVq8Q8dq
oyNbf5LeprDsIut3WNqUxCX6RyNS2ZpSWQTyNCw79THcoic8nALKCjfTCE03rCAXempiZF8Qykg1
9DwAMwjdfzkzvwgCl1O5MXKtQlPX78vZ3mj51+BB3KbOJhLw9ydcfL956oMiHhKbZTxPwO/smoGR
Wq4GGxJzKEgjRyzvzXDRA/RLUUsw0vXugKMwhSEDXQnSKS7s7cgNf+KOvlizAlXDNIxqPnSOvZLd
6cJE+Yulsri4jZcJgAwoXxsbdExdMOgrWlVBFwH1sBznvl708cZLdHF4CZJ7+ilE2vduHxZL/mcD
68agpasoGgSz418jqOyO/hZownaQTmju/DHxGT97y4ZZ2CiPePUvNMNqFA6AfdJ7jqWvade/BUdS
/uPPTzfbYI696OKbXEK493WUR8wUJL7r69QAILIW/nN8KcdR0Bb5dSII3FAbYzbEB80LDVyHnGM8
N1/sAmwdhT2Hxdc4tMlKm7eRfmIJREZ508lUm2CoKmotU91DCD+hSy5s0xhlcim7p5BkxxZO+mvl
x0AyRMIKwsL0nxx9PQUYrowgQwg7KymBKLFCfjG38gKUsLcyibnCfeGIwzSY8UaAqELtfcm7LsUA
ddHOIGPkV7hahwD61NFbhr1yQDq4s7AnZD9vPNlMbR0T5WR8NdsanqJ7MLyxevZQdJ8rwti+6pP2
f7oHEeOhHaBEpP8jh8Dk3wv3LXq81ZbFcizlYVtaCJ8RzjozSW/omFp/PY8mT9Jwj1GiMr7OUFRd
2VeI6+XJEkYTori71I7Thhrzg/AHJYNtkHIMARSbqYLkDybB8AcE37hW8ioXq7QnmA9H17Awr7tc
mu3f+3aZvu0N3HS0/yZ21uQvJwQMBhSmX15bPFLctofkYvA8HN635vHR6opahBhndTsiLkvxGHvk
gQXHuHFoBNa2Y0lMEj1ZbhnnCn3YwBB6keY5kOE/tChErEM39xslcawsNscFWqEm4SRl8esgA9qD
Ph0v2x2TTcEHs/jtJ1dNZsyDt5ereLqpAyP0l3fz76C9mBjx3s/c0g0Ei4yz5DNa9aV4H3BRXfOO
YjVIWSjO/zO6HItp2uGORmOaLbYmexzQiBzx69ENhypGAkr/eFR+cLWzVnpFn13LomiTgLRdtlIT
LOtm1aVzAswLgG+uTGBElcrFETF9jJ9X5P0q+ttMK4SFeZu7X7tx5NPQqyyIKgF0eS/i7Fg2QNxf
qenanrlBnAhdt6iRKKvXKMZ9MScPGITi7LWg3WJbVpbxtybBAaqY2OQ6LlKUQDj65AfdLyq7td+a
78/s67rXDE7hGBlCT1f/X1ml+fIeT108HTnHuSO3O1SjOdgBkFfiHe74UDhpUtV0QKJE9I7DPLTI
jApF98Lqd4xUxig8o0KENZ+YTN3/OiDgAY9igaivE49THW/ZuxVfBaVeqPPp2qhaEpZGDoGG9w9I
WBlhKgQEJirOYlTBogtleTHVeeBXkdI5xEbGpOiFnrH5AmniVeF3SgXaBlA/9nY3yNeMutqlkndf
EH0pRx/1tcW8AUdjtXg1KsL5D6HHwEu5UFTzj7pLu3s9AIIk16F1+Sst3WM6r2KhN/okPhgCezIY
pn122SIujJQ3kshjVG4sRoU2v2Hh+Ifmn6xzmZFwyNJF4RD0zrhEzJk1VJci2sgrXDOnMD+8lkMQ
6tqKirfs0J/9JWDsN3un2CDy0IAmkAyx+VFTPXFhUGyDXSGxKP4HFISp+8UQfV8uRZPun7VrLxxk
ujnmiuXTNK/OT5izA1Qg13oN0MJXoatfW7VzM4lBOAqqcj3ADMrPQJhhkvVSlWnw61IMZ+IrVvZI
ji/F9KfOeXT9NejKAYWSTQo/a5pkSSlM4bly0L6H1zsSUbQDil7msM5RgGPAIbN2GdlzlvE/QTNS
A9vXXUaBK1H83lHd52JDoYR1YFeC+c2Y9V1buy9kH2BgW1g4iYqxnj2NvSD7z9QBIvbjYbT27yqo
WnKC88IRii4QEEHdpUgiR9fpp9io+OjUziDzAvtmxLlt8A1hCELyp0vId9c0+NTvsb6ocK+34DH/
VR2WlBeZJOHDUD/muZa5TaNf/knqHUVNSp/dlh47yFCv7qpkIrJW9VBkGP9U9FeSeL4432CgFU3a
X5L8ivS+s5k04CW66CB8UqhOTpFGIY/UqMjsuniTDZBI/EoiU6WwA3+jm33SmhM9DScatQeQqRxc
cauWkmxUgijZnGmLr23GYvTm0kmjWlyja9e2rAk4zBLEG+2Bw4qfiqtkSWkyqTFMMXqZ9YYWK+EU
NhRuqInPYvCuv3kY6/t2URVlPOqZfI/9c9yXWeP+NAQcR65wa5/K9ni1A6YN7nxYk9bJ71DqNL/f
D5r1SeaRnzxTEPVqM2QLIarlqePKoccwBydY3Ivk6FZE0b5Jx+LUAAWRr1Y693TQKdDq+2xReXXJ
blmuYzqS4LF6bTSQH7+3SDHq/w9lK+lIh9kw1erQpQG9jNTv/Ofi2HwnVqOlQPFuli9DlXEsFHNy
1YOzXt8gCUWwj/g2nAKYvumuz2ONJGZyuAhoJPRNoFJ+6V6eWzk/ZwzTClTRhAwzglFPCaXjYdju
80J+PQdZCHJ/zhH3KhAjOgJwsnHf/1JqV0H9YrivVHYOzPUPCgxgx8CFRySyS2yKeHPmDgC62wA9
HA4aDs4Xci6Z4I6obTXEvqbXMOdkLrz/lVZTeOsGEalKzViIWvJHjmdKCvjGSOWDDLKQ098Jh+3x
JdwZTnsNzlRZ6I5OFeQSOIFbprM10X1irtYWAfV17xNiCaceJX6azNXR94Rc5HNAaAY7WUTCx+g6
dDMyEmB5ZUfy1iQ32m4HAFoFjubW67QSNXOaISxrGzyJ00iUteVmSvC0JHYK+Qe9ARLHtkCpzhi7
2o4HjHkGWg/FCEccVMfVYvBLY9oYfsfWgBSgErwoYS8VXn66mMbj2885abZjv9tUl8Sa+A+ffzBw
6oL3tgXCE6AB87wqu90pE+pzZ9QFXDQBCJbk9kyxgIp+XUfUnu7VdyZNZTwihlry8qL7M2YILgk8
CAhChso+I5QkgQUAI86cv4xnPa3cTzIPjMcl2ws1e/pnMMXRghHWkxfEcjodlb4FvmMr+kvrKLWg
mEOTk5MlymIwHq3NktBPCsI9D72sCLi9J0hb6uBtrZ1tZzBd9yByqxqhtDUDgw1S4Q8zkJm/WYdx
fpyT8O3R8ONVHFnWYZldbqLdO0bl4t50h32uYWB+HqxLyyFHSnhoJLK3rCLbrGrunBhDc9Cq9ucb
NCi8HTucjwpfycqxh/AqVh+v9zWP/o/kBbeZIpapoXz+P38prXLdPB8QNhL32KHT4IGf0fRdRt10
7zC9Qz2InIxjFPxE3hf42a+VLCs/hfkAo/Q6iuAqzNWU1FSqsH6sPK23u+NCIL6wVyx2ytVzk7c5
FBvfLi8Vut6AwMTR1ng6oUVrZj2M7od/lM2rLcHJwBpWYPb//A4DSAbRLFn5DdTTRqbdTAQy5RuN
eUuFtRgjmFzWCq9Dzj4KVLW6SwYfFSY2jafErt+Xjg6feMzgYByzj11h9nC0pkxGSTayIL589VVw
OwYTXBVyjrh2KtgDzE0PWQWyOpjLD0tNBs9m0N6drRBPKtLrH+kSnyTqUVnjRCWRYtCwP6/Y3TBj
aiyq8GqYfkZtxx/x3rGoDfSmMBvC7+rdCB6Wi8NZ6i1EvAGJ8/3VyGsTiKTUDcTyydJ9G4WCP2gs
gb5LoGEJ4an9m45bq7YhvKx9KiBoOsCwKbEm4c/ua5bg3pOPVCObxXNwNzzboSY84hviq/KPrp3Y
ge/lX3a6sWJMb8QeY1uUHRdRg80kL6ct+BZPemxGgGQmjs41lvwLNX2RiDS+CbEFvTO3OgyYPgZG
vVtOcs9Su6CQJ6kvsIjcZ113QkGPiesjmEV8tWA377/g1iGyKRsMwoYflN0EKZFuNlCs2Mn8FUwf
UgkGfmKTDI0Y46UOXVR2HZmQEEFBlY9Jg1bltBFmXOhgJMmSbE8n/JBVpB6RdVG10jSENAyFYtv8
+Bo+1QwCKtDQXNcq9W8cLvPbPNEsc3jk8TKfsSw0p+sNqvPY8dtu4I0uiIlqFJ9r6wXNqmA3rvCx
PBQBxYEGidjIyMv2hyeFGXOTSvsPu53VOwb+sa4wRHShIe8MwiljU+pHWGdndUI+824HcqzHU1gm
k9iUi1jvr8aCzvlzvgzWpgVVZZUlcMAiAlpJ4QH+jwERUu1T6YjCHZwSqItOk7PBf/7vlcaVSKKI
FoAlI41pJ4d5ChkPDqAChwfeoTV15yShsWtDnM+aGTUerwzio7WDTYu2/Lb8QXECdh4QlfO1natF
jDSmpq2FE3ifwplKiSASPsSyiXSxWqLiLIrU6gFeGCB9zNKWr7O5jQFIRNmiYgA3vR4/lIRU/KVV
Jbgb3XDYvZrgBQBpyF6AGUW94TzDsLbTIXbZAc+roAd80d0GSTV8FoyIpPt1sOUjb2gyyy7QQnCd
R8fzUsP5auSa7PhgLsuDldWTk7MHb9VNu+bd3FeO28XebiGAkD57xLc39kyfC19e+BIrCdWESI1I
oH79u9AVIiYHs6K6pgBLWcAkxktyCncYRvnu15ZMCYzCm2UkzK2KAS8926rp/VMKhrjI1+pRw/T1
KMSpujI7rNJLMWldmBWW1I1ceTDIKCtd4TBHCl3H9kny+kkHqm+SFMwQvo2hTUzCM45TqaG/gChn
UsA52xgBwqbNc6+fULiFBueIrADGs+jtS5X0PE9XztVCy/7NVRq+PoLhEjGJsumjxNjR4NN8co4W
TB0vX3XA9xyBQlBP/LnZn386brZU2Sj++GyRjQ1cuD1WcjM3BIRIPjaVK6RRyXS8upC0X4jNFLVn
dccSjZ13/kNJ1Aj7Ms6bLg1LXXXPkE2xsCq7jWxVu/j2dcIj6po2u6e6dM41FbMeBJdwopNazCAJ
JtZuGcRqpOsRBqTpRLVKkBorPK+oB8xbzUg+Ubzz3D+jCCXCYP6m0mnMD3CRgql+Dw8vZGQCWUOc
ObRKHfzJgqRRAjyPprzBlgrMM0p8vw9VZsq3IrNLY5teHUUXmbkhRHQVG9kuUnq6J74DgsRUECbB
pmomf4ORlnsls8coIAMAmTbTPdx36N5qqblLWPqK602JaHhr9coZ0K9xdymKbHFBWyjf1uC5CZva
8nDetmIx+yt7SY4oq//QdtutblKDQ7jg0ezJlRto5it4obtzt6DPA6ZqrrKkeSVdaISoKu0hk+Oi
xxTjLmzNu79WUmfYeMWkLP7ULqpaYfeO85hK9wyp62n4b/9Pe/yCtlqKaDv0U3V2S/rsKYf7xTeX
s2pSrtKRF2IJLadXxPfGHHvNnGzrOgYo3lGyiVLkWeoCrF3xzhmCP5pS+iObqxeNJtH2nCZ8AtJM
ax5iN5DVXfT53qf2SOUXZeOl/e8qD5Ftaw57q1u3fBVI4h3e4EPQIW5kIQ66RtCW9RmP5YbxLXyf
sJIK5mq89r2mH6GWoDFNbpUqf6wfTAVBwNTGWdSHPIoXr4WAkULWwlO3pZl+BOSd3QNxLTkfIfMO
JNTSPVkh+1eUzb1+9vcge0+gYF8exGumnAvirAGA28N90G72W1EjKx3tvUZ8BPwP5Nik6HB8Rm2K
gZOwhmEUwjRR9Z3tNZ5wl5Ya1yxh85fPy49K/DBexxgbRr7qSlqaceqD0UqySQSfmqZ88k47HKEp
R4PCHmPHolh7M0LeWGq++8PitKV3yflthukP7+iDxhONCr/+uA75d69sCzgcyx2Kp/s8tpU7DFVt
Vtv1q44K1HFa0qv5r7dYUjLeEbBk97B5e+x5D4Je9DoW8d4BN59Icxo8QT5jcrCtSqTAaIee0siD
Z/7bJvtJ9YuaR9ofEfP9rCXt3UzdTlBFvRVjXTF/X0VQIPKN2APibjPXKMghFij+y+tiLwtccOu7
jyCbc5pmBiXMqnRSUMBzxk0rIWICOqtsq3GzoAVewadtZrfomD0E0iLxTD88U13yfW4TayiXb/SQ
jvstP3TdEttPLEDMtDS0Rq9IOWxLh8P/GodVr1+V1/akU/7To3ytKJLh0skyUWptYZFc+Pu6/sUf
ZOUFQBe3ofhdT8eaPbUGWdUtuhqVIoWC8M+b3Re816qCcxb5awWS/QzwhuhpIpG/cW0epphcit7P
peROdyTsqUB5uE2aSH/r6h2T2IadW8N9WIUCeEhUgeaq8rZm7COeKQpEFbYbBwWvWGlvx8PwzCoT
V72ppuoWf8DiIKTTccyNfL93VGoQ4q65z4DdqMmHTqkc8ICH0siWp/aJtwa4qiCikXpGx0epQi/g
WMrhQkTxICl7KNtICnFpKCvmX8IAtWWHefceNxmvBPbnESf3X9Btv/uQTdb6uP6z3XAsQ7V+mhRO
pKUh21i01w/B7Yxa1G7aiXijM6obvqUXkSaHndXDUNDhpVT32b68RUrlWlApNsPpfMXv9CX85Oyz
9eOeJwLSnQjMOIW0MtqyNenH/NC46yHq9bF3mIKOZpp61JDsfyLBep8tw9qDA9uI360UYu183JpO
uIkS1Unnhb3gxdfAsmt1+pCcmq/tU/tHybYy/e+DgWNHHtjWNfEj7H/8EJaTxyvpjSjLOvGBwp/i
hE6+Q7c6nuXFsMpRWr+dvBsJjbYD1BvyP0JWn7W9e3idrEZtbPyd/u1Xc7EbQmdD4DDXcdmviY5a
Mqk59EcfDjdqwsnzh4sIRQ067P6vQE1aLGceN76KnK1vyxQpDRDLaVSSpDPq+TkZjDDhg3lItUlg
py7G/+GE/iDULnOMOidVcLsbH6FY52604CjzjpoVrBCzsSHBmfOJaLVZrdi2OTqfJJ9JgzqQtB2l
UmRLmHspI0Zn5Xe+fnkNyF11amktqE5SXRDbHFBl4bTzKfEUB7qGdJqJ4LubFnw+sbBmeWeFY+Ji
jZX6KvDKCEW/tLdzqEfqzi6sVoFO/meu3yP9UixWQhzGaPLlO5QOGc/CIkq/NK/dVU49XtvcJAg3
W6Y4XFfiHMRqZtvGZT0BUS8oFgggT27LLR6omJp4Y5eIUpWUTKtkTxKRdMjvXcBrJXrNmnLy3wLm
4dJ4KSmWCJM6BdFuLsHd0m6ZqjCPYZLVpntlOIU8iXb8/HTWfnZG+L6lFOvLaVvbQKMcRMq55Hu+
Evtrjp35rrxtmAZjbdqvEbaXwXIQT6Zx9bNLl11/xSfTJeWe3tscKOyDaBz9lftLy8jKah3QGVpH
qXzJj3Yw4PPF3JRc5vpDuk6/BHcf80IyVAdLE8mxEFCDzXwamSzFsRdoiWoHxHr46ySyl09TPBHf
Ztj2KDnPn3iesVmVSjliIzOG5094xIMZm+UNCmiC/ZZMnScuSFW4nznWC376qbfsbRGP5jDWujlB
Zg8iqt08W5AFtvf4k9E7J4G38IOrffsX/VEnsXoOoXsqXM38A6oRObPdlMJ9naICEQh0R1qWk9wK
rGpyYHz9sGAmwDXcNIkHmCc6g2/MVXKqIPIVcsq4cd3yfMcRrKy2Lx2NRXCjD0knzNp7p/ikfc7R
V0w/RstVa9egtUCCl1KbAs5BUMxgWsJISbg+tBIyjj/LqckIv81sNGsQrMi696OddHGVmwPXePec
utZK/lTB1oP39esXi+fsdUbwewPqied+4beD8Q6D+rzc9a5G568W8Insvw74hm+7xgYAdVmZ8mTm
gK7eNH+fwk2ZmIr2gZ7eKur2Ysbt3ZPlJGcI2RjMwgd8jIeJfQz9aQKqgt0oB2/6tS/xHrSQy9+u
UYvJF5VV2A6OPnXgYNP2DXVsgUaTByF1qBwTOSoPUBnrUBNbH2P5Hgbgx+JK7lVRGy1GBK/dPPUa
UMqi9gryWSyFKLonFi/kfba6eE/tdPLaLQB9m9MMYwqvmKK3CEb7O0hegWeF6tUpjAdYHnDxOhnL
FsjEJuxm1nQ9KDPw8l5Xj7ezS4LBazEic/PDpd+M/IdS0esefXe8fWIUNWbDw31hkkJyPbBEtqyq
4OzPM2+YxGBaxezZ7lbFpHdebIfnz0Y+mZe3haKlcG75aHaWy6aQBuO940WxikJe664ejeoIRNbY
OsgCaU5/vGFrOv6cK+M7t9E3A8GJ3ts0qgHsooK9R9cjuSLBHFTJf2kPKCrwzQG+MhRO7q5YqSOS
fHP3UV9K+/pC/t0F4SfeXm2l0qSc3o/FSwuh6+az2KAQpsK/Y5E0YpTM/FxA2/wIqxHnVtWV56qM
UfWk7lotKaJpSfvVHkTxuOOJmNsDKbFIGbfzItGQNBTNyI9F8BRIzw1GM/MtAPPj/uq14eMeZ7UQ
RiITRNVSK7hhMJ5L8Pd6kDKLWM2JQ8CQ2owS8kjakeNCpY3c00KQNX1kY6kidNRtPxXq3IXLmtmL
z8KS0A+M+uFFFtzbIz0jysB1KzgEKT+Y3M1YkKDK0olD2hQu7QXi6nJb/NNeBLVt7TOgZwjpzax6
G7fQpNwqlZTJkapm3QB87c2P6FyTfohjjDamti/cFGUKqtX+/2wQqk9O6qxUib3/i9uOn09V4Ty9
Eqwo4J3iJJN06ujFztRiNsgDoomXNX03VFoMdcmWKlgry8yKxfJ/f6yKlAsM6DhqjdB607nznpIp
U/Rf4wE9sJTb9y/9rfSaJrwGoEEBix4BzmSUssduHg3yjA6LvZr6Q6EVe91615CaWwMgJEMWVL0J
gbpYBl8ZdDYNtPN7+loG1KmYVq9DG1K+shAJWC+eSr0/yf26l/Ga+OB7qWgblg+HlhxCJpANgN5K
fKjO1OC+PCc3UD7Bj81h3nXNsuDFgQxTQbaYoOH2znvfkCrzIGvyR6eLe3fN4QlPnMgvHgFd4A9R
y6JmIYhOYV2UVfgX70qkPxlonkNJb6o4l9ffJcpxWGtbpF3Xm2FF0oSeS9qAHGj2ykvkbhgcTmvm
ne0S2gu4SORuTtGF2sxVAhCteDCweqE2yKxesOdCMHVBETmUPrGG2yL2A2gr/8ZiYXDV+D60h7Ze
/6A9+GMWE4s6BCxIsStXUy5NB7+HjJSp1ztdM4ee78VaD2zl51wD8XgIvNBE353o2RYP9G4UGp7S
aYcljljTg8wzPA2ISVvFHagR1hMajBF/kE0vaqmNsjgc8Xtw75M6aX6WvTG6Ae7xm8eCvVDe0hMM
/aR8zGGROmkzU6iL5aG0Qgjhp5iK1qiTO0N4BX3V7BRyC1B4sZtNOW09TaGMKQbjGGkgzA1qYGVo
laCeTL8tKll2ZK/QaBoNNE/qbsqlRkcSlSb85mnvnT69TpRlBKSwjYaWjYItpYT74nHGkyJH8zQe
E/heMSGGg/CSqdMT6JOVak9OyCo0MrIzVxNc7/oUsFci97Vv2pG7sv3RD9/wLwnaGz5cQXWuw3Fy
sBEoAlRt9QJomCKiOrij1EQ9HcnWqhS02E3FprVwvREST1nyYxJFp5agvuqGhfTCi7/wuOkGvvdZ
qWtJhbZPoDAWXheOg6MonZeIsejIwJF6nM1TmA7XZ2tuEaZQTh+ziN/NiZg/nRVt+VHGGJu/LsNv
GbwQCpEwlM1BvR+EiRFDzkwYn524D8I3tuFPDIzoyMEWvYIPc7yayyXjXYIVmVB7L1UDgYGidNqI
MhELS+FJh6pR++gz29SFvRDgLGG+nQdvES0riIG8IEwXpNknVUFzT5wFQhbKFJuA0wmwvfocgF6C
rUx9N/fOdwyzj1/sGV8NNm0KFpJaI+zrnOFFORIv+xWLPCPoFAlMYiK0vrZLNOzFV+ZXWKTYjNf7
Y6iGsmOl9swAX8roPdh/VzlXN78pm7/UIQsB8+KPAhpOQGr6KZ7ST/X1i4suM7yxPXt0c0K8hLVH
StX4Lef3ecyrP/ESGT0lYDuEX8hDKGKhnKRXXTjrhmdsRGQXVnmLKEgzQZW6l5izPMoJnUgFXL3l
wAFQFXECym0+urM4bRaq+YAP7Se2ISnEkO9uF6aHG9oRyG2VKUTY64SuMxolxkOteZ6gd4w3lH/d
zKCRopaTfnqKm2RCdwPQIJpB8UlvOPwfivXPO6xKnuz7hszFc6zjhpQInQRXyUStJp0HVlTQpnCX
rPCHSdkFEi65+uPzmJkFBDBLNbajpC3gafu9jly5XEKhYw41LenDxWXRYEMBGckg+zQ8tEEo+Mia
52BcG6Ty2kWJXAabpKvX6o74cKu49wOPOaIHbBjJEBMr7ZE+UZZKMx+4+9/pwWNzeZESWeOeIyqb
tRxP2OzHGAVUlNVud6T6G0epgitQ3qwxufGnSs5OIER3v5XSarZQb/Ypqhlvnyo3oO/Z3FSbX8K3
v1BQCW1SEW2V+3EWJv0v38kv0Gw0fAlERXPC32R8JWpCWLEgTPC0znRCBq5v8xaD1WGBzRHeS9T8
gu7U5Q0Yzxa1nTRYVA2eCB5HeLIQjDvdChCqvGAZizCWYbTstNIecMUN9gIx4+8geC4eHL5l15Lk
yriOWGN79qDbb4nIFuGi5cV0SIewDa0C9aOFyE4/WUjpaq48czfeqxKglFGEJTnHI4CGrIsFex6v
XDElklAro04aVgd1N52vhtRfl5LnymIIWr9Bgl8ilNwa7DjSmHVaUO2QLf+XnQw2UFkf+i/kdKkV
ba0SxA4Jms5iM7+vJVj9up9vxdH/J4I9lUSEYG5CUh7T7snthsb5222woA0kJzgGG4A/jmB5IUh2
van4k2EEV+vB3yYVpzRJqARkX5zczFUfBXYhTNg2XdmpkP9BIAS4U39AbBVubqcPi4nWO3cFLru0
T1MhwFCGX0yMQ2WjydmJeRA1QKPiIsDRvW7tY8CWK+cX945n27iNU/UG1LTIsBlhyjxWs2vrXgAm
ZaksFAn/V3YT8SiOhVdzqZ3Ao+uioFoUesyU7itlGJNUI0QChTIeMdnptflxZtyukjLRyK5Bswez
d2h6weMxDyaNOfiVsac9f3VQdyciWStn39u6Qzk8P6sASynD3UsPfF8LM2vjJ2B8lu4EINorLk8S
CYXJIh52dcNhAOuV4m8F0xJVqFDeS2b/kk+UchiLtw/vRHdkAvE6DYM7bqLI0DXBjIShp0c1lMjS
Si7/bUX+vhs8ZpZGURlPBnzSQ4GnqRVX5lRX9Bcu3xgVrLVhfjVRL2HSbl04y0jIs9K7VHQnmHE/
G+gpA5Izx5caNdfyFTI5Pdyked3WV5Rqc1igzx45G5iUCgoZ69qmHeFXGlhiA390Yp6yUBl4ydfl
d1uyB5usArHJhWE88Z6V/g7B8Zxlva/idMyWGmPS+DiFSPD53HgxOtVsPoywGKqMJ7IqSx0oZu2k
Naa1sD7vdvr0jGiqHb2dfoKGphLWLpR9TcxvA+T7nLqXs/SoysdkD66xt+WkVxgbCA1DNxPkCeK2
0Tjb806ZPOug4gOVp9Tq/GigEyuk7IbRWOcRTz5UAjtejoJIuO4lzZju907VhreoOhsR1PwIaKES
BWjZN3Q6vpCNQAp5jp/q0Qrtr7RHTAvjzgx75kLwZtl48TYBc6YjZKfu3dVRJ2njZb5oDGfMLHd+
12y4xSm6Ty+kmRot/qeGb4zBtKtsugkg71hChtDx1Qs4z1oYZmseM0gmmw42Q8gtb6aGMHBlCeO2
92jcie8MMVWCFJRcveGzH9TQ6c+GJydw2/PIUWpDrPzYiBPoV92qdmep39cvCeZHHYx7TYs3XnNY
FX0/IOLjDDPTfwa8wOy7RmcyuszBgDqN71pwSraB754m0/JiCpenXeq4pfPmmFXh8fzH8RPs6PxS
W8KdyO/c0FBzLcUCVhkOUE6tRuDGHKg978PIjSp/xutLYMY6BMdVIgPF1og9yP++UhvTD2wFZPQy
xlrlAyvFi9VONoXsgIt3cK9RDRV6pjtLRR8wV/KaOWhEVoO+qhquBooHbUmI1kcqUOxiVc5TN/ci
kMUwoKYMNflX5cXoDsALbi3E6WAixC/wfjmUdF81rzpjJ1w1Grx/TVxdyXF4TuGwDVfcfh+WYyWR
uqXuqFZvxlGH0N90U6EZpLM2oHyAwSCOkyhbFPKcWgeT9GTtzmye70OgvHNqi9w1bfAM7tJYsGbu
jlzWwYgzZqKjGrwXd7apKuv5XgwANSruEMkCYt0fet/ShlVgxPN7brWA50TCBUq8iqmUdP6CsWV6
+BAqfn9BACdGcVgSBOakWlN6wRwZfJe3kJOSE0dYUN73X6wZhkIBkbMDEsCUwHebsv2qo+HJkFgO
KgpuYGR8iemuj/Xf8UFHXIPiPOWBdh0qdbdfcYUNYu3g4QJp8GNq/3yBH6lZbYuYY59drOwsci0k
6idhsF5EAxSVHEiQtoTTd28sN61qaRGo7Vgu8LnkKD7AL49NX9mAapGOIeHwfAKumKwQ3X706bpQ
SGpJNvkAKRXHD2INsjcXE8RVSjBw2Aenu81OEfzrFBKHrfpFXPFuPnRkOCAolC69hxlJrsMu+WRQ
1MK41QYr1wyE6TZAeh/wYK0HVJb78NYuKu5DdD2mgocl8x5ssQjH95t8TAUZ4tg+9XDt9E7ADMPv
70mdpVY+kvXTsFC4ICOCjbswzrHLev3qkqNIyJHFxa0m1w3WUnLQdV+fdv/DxdqdxunVXNc/1sG1
zD/6ohB18OVtRF6N2TAhnrPbgEt4ZxtHUXkwUE9nLvVvcr8LlPvnB56Hd9wsCktCfMCLG396yMuO
OBzUfA1CchSGdUJb/fGoIoxuU39iuW92gGB+VFPqSworEfHS7kzPOTRmfH/7Px7FKGC/pahrV/GF
8d4Lu3IKAfkMpk2UdHTG15UYEc0oq2Z1+4hLJCfCxHSn1ujCUTC5G+LIuFAx9M/3qFCtBibB8/H4
kZPSgIauEVdDNLfVEYzb5SdfSYN/Z6AsmZzP11pOOzHPKEOGxULcLWWZylL5Alr1QQa9BNK9dCma
YlzwKANUievtZ1AAhZ4iYC1rLFilWS4JAK2gX5lQzFdWfzDSg9ZfTYEaVuzjy+6deUIhAvYBXPnh
Ry2X5CswkJWxUrFP58/8B4Cnex5Qkt3/vgfMsuWtKzFQyMYK6PaTMEFE8xCFmZtualcMMtEOVljo
Ma/QuDcsbbwJlLtm5MaKolzj3VslD6nJSpquhdxos7TVEzR8iHjup5kM+ohz6m7HnVsm6aHisJgr
YY5j+zQOSLk6OFBU+ychyt0G5zK9GHQszZ828c/VELUQxE6PiaDnJtgE5pnxf3V7fCNztekewZe9
Y1h1K45y3T01ncUMqhP6806Fozrw+uVyPVsn1bCsZK10Cm48m24/tqgTOHFrAb17GQpugjwqr0eI
fXijB7yoaR5m2okwXWqdXkUaE01vobWjOMBsb9YGQx5A60/tgexp6j5XWeMHj/2+wzd/K+eEFoRq
doMKMznC76FKqX9ZtLDXAmgC2rLEGrNAY/SIfI8i+8yfIDlGS3//ia9dIw6Xs3GvNZB7kg80bThB
ryHd0ylN7p6VLw1/OQMqPoyMWSoESYDJ0qVNnnmwP+mxi3JtoMXmPpkT04NtilFCBVuvQ/MH0YZx
iY0pIu5VuLD1AQvAi11y9vnlxz/5lwTlVgsiVytpq0u3+3JH+yvTknT1M/f/tqGvffCcBjELQbk6
lbqW9mqQqgeTvjd0ru+LzyMwp+hvnSbpkkX+Sk22M6aPzKUCUkX409CGnkE4eqOt4/f313iCIyfo
5/PERYDF01HoyX/F23Esyv4anpiKRzxhazEmfCNxuLHhOpImm538jcqLivjV33pQoRJRIXo2ZXdw
9O7nOPm2a4J6aTu+29Ny8amdRbzbxtD7vC7vpGDBOii4403wFDjcFjZZwEVs8Xzebm2in+igcwoL
77k4xK0Whk8tlyXBV8d4sgQdbz5Vy75Wl2NeZrwpxxqcOiHddHt9ZjNRhEbfwlUKZULGr9ncBaka
vRyhBfxkk2efeYYIbh8DL4DzBqYlntw6JtENJW5MPJ/UsqdMX03ENq9YGA24s8pbnM+kt2gajtbo
GdWHqPK87DcnPFk7xRREfax1S0BPm1VvnicydT0VpAnAOtbt1H1umA+lssI5Dcu+oUIF+8mm6PFr
hSJWeW46LTSooKmwlOUTHJDFjelAi2W3he+x3SGBoPtDjasomlByA+m+LJQ+uo6Ziw1LqG0X3b9k
LXyx8+XMe0r8h5OhOWfs4tN07PLUjlQSXqdW2PAd1Fyo/JJps/zW81B9uOxay2oV6nbWrOCCypJQ
XV42fDRjrrKGUv97Vbqvtpl7g6Bw50NKKsVGF+JB6vax5jxuAyvFELmy7AIeJQP8gAVQRblm+jtj
DxcqvrBzyD+H1MwNq6mRvrIwUDjD5xPqBPHX51rnpy/4k7sYrarXGiyfQKdJlFCHQovrM3mcDmMt
C7/udwJmjq+++HBFTOmbnSlhSokn4Iof2IYjyKKUSnlHem7mOObPpc8rKOjcaZRlpU8BNkak8Xba
BCdD6H2vTcC5Q5uXne88KwY147GgzI3n2LNKhskZQsd+l+ZwqT22I9M2gXBLRLtmm1GoaKPF6Khy
sChEKS4gbNqMucKIsnfM+8XZYHFEdYElfMyJNh4DPzoj6mKuzzmEbuzWqoCG/mfugDx3GgUkH0uK
c6swk+PmU0i4zP6k0bUoKwBhCiOqnsRs7gb4FJqga5iUvGexoVyj1X2exC+f8Cb2j2G8F1obMAp4
eJWFBKQ5juVITXDNY9LoRDorXapWbdK560ywSyf5+JE96yJ7n5BKOwPnYJsxYfxn05Kf6WlOz5uP
mtPtLRdRYr/tyx3DtvUM5Djx856xsFo6f+bHJGnQSOw8IQVNfGpSC42T9lDPft1B+YNIti657u2m
rvCvxr1z4oIUPnxKikQXdRQXB+NoCfJW+ZzE3HuyUipSTJT06whiBDSTpTaq6Z2AcOJriW7b3Wdb
aTgz9Zuu9bh4GdKIg6IoZMAn2YeL6VLYy+2rRoiBwnxJMBPNUlEmaTcrmp2iyuVCamxzgmv0kz/I
R8UYrUxYPfwlds1gxlo3vnr64/i7lxCdI3/IMZZSKnJTbtGfuIUhvRsEjRFQW+UXbk1lBD509dgd
kCF5pra5MvP9gOaNOpI0RidoF8EjhumWcDncdIU5OZU9IL21fQYMewyLlbPSimtvqtmeMdbzL/Nb
sgkMYE/dfGGZtT2IBCNH4dYwphZJAY+1nC8zEnhtFWCqmqyafEoJ5iJ8a8lq+NHikeyUEOK3MGWR
MrEQS4i9vE0R9zRXBOvm8fS88VcoZfgUZhvmoIeTqBwZZU06pNrHQoHIYu94hNkI2qe+AnNnBRD3
OtFZHpSXz0/jhfBsC0t9TGVwJ6ehVtv+dpZ1/5OquCKkxuTrTWpEL+eP2J96WwgZ5RQ1lnAp60H1
8TyxmPEPy2OgNRdM3BSQJ7j/DO24aD7CFoKVRoc/aq135YD7kGxg8tzxUxTd5/SKPx4KmCJjnTnB
r4VSp4A8ni+hxTi+V5lvNnN+i69zZbnbicqUB78lR/Xg01sPNeO2yLlgM5afl+vbD1LBOoMaPNuC
YwX7+qdb3qOWJyH8byzzhXPPTOyptyIJctZRqJbKVS7LfWRyQ/m6TGGqcYy3Fo12pGYairejpvDq
A/vgd5x9SviqAecR/CGVHDBTlAJz/+Gs4U7Wi1g1jgOs97ZDQSDqnpHY4dxulFE14rT7NstjaoeT
gVTkqDmINoUVqXLpKPW1lLAk8LLobVd64hBtBRzxTUkg7fwboWwI9Rx4PO7MbQVhnbGlX++MlmF7
nJQ7it+YkQ5r6BDgd0+EO6BJAgmAH/l4QZPaNv1LtZuasdzFO7Y7rRXqVToN9jWR8GPEefkFg4Jc
2/neKGUenSWWAiDpTdKZWR/HIl9dIMKU8GPGtMp+u72BUsk6jJDQU1dzU9+jyAi24v89hyX9qY3m
Mu00wre3nhe0AetwpKCxuQ0WMV6AyxGbmmE3+29xhvBWQd1I2qmvpqacM1I+B4dGJUWepVYfK31x
gsyTcxl2IUMMERSTo0cecyLQJQYJVpfYZMZokQsjLbKZXKKFkrCGz90LAx4O0GZWa3c4kT7JrHhX
HZ3hfdNmyFxHuiqI+iug81B4U8A9ObSqb9D6CJFMOe3ZxsRvGUUdoIXsFUF3NH80iW5umbZfHlBU
FDtE/2LUZWv2UPIbjjWZqqfq3AiDeaM4PnGO8Z9U8XFMxNTnMu3j/kzT8zgbiDTrMAdxuNU8Pgtu
x048G3lpOHL23m8Qgp6Uei27U1FjnLIkMvGnazMoZDaMmRdJO9ch+RoUXo3iz+R9bVHM9ycmYKkf
YxbOb1psrLI5aa6IUDqpA+iXM95dN4bjyzPEAqePYwGcrDqWuNAvp9xFXXeLMW9BwEoL931MOigp
NS/IBZUOlv4taFOYk7OfM5jyfP+TDLfW6wi13k0+0l2Zszr3BoUYBNcvxesnaF/6cVNWyK9j/ufK
d/m2ouD7AVpqrHMbE+m3uWPw0nZdAWp6/wjs7B5b4OoZSzNGeXqW6f5jdDzX2fDTec5MZPiPXbb5
FWNjxG5scAgsaDV2fONt8iyLZpNpMe6TcmYwtiFknZTF+TH0jl8G5Dd/Z/toAep++a/rH9Oxgjkd
onI1K0wQ3BgnsJ9mo0/wZyHpmx8BE7N4KFqIGToxY888cV7KvQMVmegMUfVZCEEoi5PZ0P6rCzKw
viCbJBhODMIE0GzNb9aSu7V0OI8IaNDaDdMwYUUNz5jDPRJcNIkGsEL/83IsDrqyIPljLqaFOnlg
qulru2sFXB/tr18piVdxDdUMZ3KAXFii4Mb9lsWlOq9Wh1vWxpe6FiH1xO/UgoyTMaMbRut25z7r
5uEDuG+vA/bK4DtfRklwBBLVCoxqydwH2mHPMUw8uYzRoijVaQYGUg+iAwfjfI9EWkxAUg4co5t0
4yFhoHJ+mC6rK/gUvz1weadgTNlKgU1SaQUffsfbnk+4meplqW0klHDjqK56zwWW843mfdXf6iFK
IvC0AeicTGtlatmODZIbsQ445Z6zGOUvjuxpfWoxcwHqxv3+UPA0KB5c8UAhaXr49EIKU+AWKIIq
b7Q/ZFsXU2X6nSKXiLf7UvXrsys97IHI+rw4xqH2FJ9iZ8aOPZn5p8Ivd1tTxGLjJtpAaFP9J7QY
wk+mLSXB8Y9+o7RV4Jv34dZqrboOzDO76oHEUNthzda9DSs6wALZ2QoZqkPge1AUlS7tp/aFxMpP
KlMquHyp5mdsumrSri3/mK32GVqRh/VwD/4jymAbjvV5v06H2ndLiXHSsYa6JjfOdkyQfHpJsx4J
kfOVC0GPZxZfVv9+9jLznX3fI8LHEW3Ctr0PAyTZwArEW1wLD0mIKC1R3gp9P/l/b0mwBWBG1UcW
kaGTPypcZzrkg3c6SPpFlr91XB6JhRjjm5pUFDDbfRkuD4EOvm6uFd8EDISk6pRQ+6oiQLXzraXB
7BkmOoS1UrWlBwvHACGxcHWMBeJ+9axyLoWcd3dNXTeQOhhk8RKr9S3LDvoXKIdfSjFmj5VlJH3Y
ihWKyYshVmPeDoH/THnI9eGxQMOZZ/WMaZPWbDG6h1+ZvfzaKrqE/0mfHMyO+AboEWiCWVBoS2vR
VqLRgtsLxBgDvLjfguQsin7PfUL7B4HYzIg2z1PXdVrKtq3CjWLpv+OzKaKbMQpj0W0R3iVN1g1c
XG0ppSmQRIaBqF25VLUIjjoXNnlWi/zwIXKtHUbq9lD/Ok4COuolr4YWUOVwzJqBMrxiB/PAMANA
ROFEyoH9HwKOaC8jLvJOuYXno2HUpJZUzWuFGYceZUK+gFQqlZSdrvHv2SrowvOorIQG0FHhaG8M
BdVbsWxTNgpw8mV9pPQnwNcE1a7lS0wF23wshjShPLPJskURwvGUkfwH3qiSY7kwLBHpDknCLQ7W
Mo0qCYohNNLEJmnOOCycOf3u57w03Npo1Yyu1WC9iPmF1im0ShxzT1MzV9iy5dNW34HaX4697nPZ
h8QZmlSy5INSuatlm3/Ca1V+wL2R5O+hBFA4DzFlrPtuBDMklKDpM78HsUN1h4CKxL5WFgtmk66d
EQoykzwAYwEa+TIj7w9QYhG9uEX2AzxYQcBi8shB096W2xmsw5ojEV9b5mC55lCOJ15NUlvLX64m
yCd73eJdRLgWwTnPrraEU3UwB/qdOYteEWUi4CzTxcxI1HbgAxuBLVYoiAseo3j02Xb5So3SiC1K
R25GxE37XxDTouuI/KEVeNmpMQuoWoliIWja162YnL5Hl8raIhxrOQzNIYi1qJQcbfadChQ3O/M4
jLSMVJZd/7NQsF/8CEaX/Ziuchqp+tSujVxUMvQri0XRJv+CZQPBzzLmtvep7aZAKZnsXOW0bPxm
T6ukrZZ9IoDeHWnaUX1Bb2syQIZik/Ip/QrZlNnZg2xBId/UG3sevfcVASE4IzwFvF7aKa3ZgBr2
McKuyaRxTsi1KjiKTFjdhbVA9is76EP9xfjAMYHEiAu/AUoc3T2UPlhyg7Vo+KVev/suk8l8FINn
iF/oASHURxTzMl99MNYc8Hh2Qj2B7gN3cOjqDtuwlbkrcM4eveQDK24lKwAQbqIUJzZOwEuCMJ+L
Vq6IxyZiLMfzplxkmojPEk/+zwlq1dP5FVTTxzZwa05hAmD9M06WNul/asO3wsq7CiNZlNgHqD39
P2EBoSXyrEosEtCRpBkOGPhPIorHOOtHx321mQFV+u+vlseZksnKoNjjRgCjzmjsVBX5fVuVhTwL
T/LmgSDs69bX7tEcMJqNknSH0lmegmU8oEnaArTSZaxv/pMgd/34qVdUWP+KmstpooEzRcqoLBI1
W/Zq7cUpHVe6dq1yt7PNJno29q3ORDJZsex5DeXNjrR4qurA5qWxBfvelT9Ro8AouNWrbU2g/AGW
t9XVH6uVxmIvmYUyIqVJoq7y7DEmROvi4rmzM8Kkt9p538JVqnIHHBP9zM1kewGG0Tgi1zV0vuIr
vLt0pd+VwMdPVbH+cJA0exjXUNZxBOeTcKK8wUt/8/jGQ+x4rszcsHw9A4VjvTEVPwRsT/rHD0Tu
Vk9KGKweD78aYCTVgbxivHr/sfHczZjOVG4aeDkiBH/5jvPgXx4qd62DkUSScApJZoVuMyL0M9gV
y7jl9ow2iYMrO8lNg+2chsTDsiNQJOinmRleGvJHD+MU8fA9o/cP6LaNmoPbM9+/c9FRyIQY3GSF
RfnYO/tCBaZAoYJcJg2E9xE52tqnx1vxmsU8/ybPtolfzgrrEm5+/TAcuOlQM1zRuT4FF4YN/QBQ
doYwj1Uupei/eOlM6eScU+FR3ILOKNm5fTdkD/hWXBWxIOEssky5AQcABPqjeYWGFx61G20hOrc7
ALtlY2A5gfmedp8nuuSADHzPZt8MXjk9PJuwDQvL6CZv+p7xXLdzu/oZHjBBelFro5V5BC/5Tkpy
Tm16UxCyVd4Uup2U8iTF1u+PJCDOgbPcm+gI2e1ruiPARikfg7uyt/MAapo60TK0syy+tctWbwZk
0GpaCewTzC1jVRLk7nOVUhD9XqyDnBI7u6LohEqSxMeFREiZIwL6mM1vkdbd+eJs4BLZ/6cLscDu
IrXlypjYPRPrnf0sjYY6OjgBjzFUQHl9pyDcl8iX9cJTQn4yxdy6BtwZSOg7HgExQGElJec1SSXR
o1PMdW15yx/47sBODs30216mMpPo4EtqMYsirKTLGbTKP/EMvQCfKqYlH2A/UgSACK4W405LuO1o
8hr2jQGsaC77zV1fl4146S7dmYi0hr5WzuKBhdiojj1nJ/yGJrLrkX4rNawAWrXFL58/WlPDm/zq
yFzWyF2Bv2M5c1EzXWMBTNtiBWNbglSzBoJZOcYfljeoxxL3wgymqVBdU5AaNKlNcT7rP9RJHnLR
uSITLoWCRkIb9xozLxm6CwAFS47eHfyIsH7xuF0woDtznObeJRBqJH3ACk4RLBKweBnJKz8E6ZRn
rhWV80tKOeXkdHqS8DK3WJEYHOKy0B1NTR/KU8+Rt1FP67p59Nv0ht+4gyUh25ZF58Kv6Qs+4l8m
9fxdUwXopAW1k77koyOYMn0UcxNSt/GdQWfqef6p3guwF40A6qe4CJnzSoa6+6Au0rd9FQVO0fhn
1IryL4Sbw1uOWBkf3gLAxib1ocDHi/fBW5WiTb03WZnvkD2xi7Q1WYHoYcmVr44Okjfkjqp4OUCX
zVM/O7mWG7dp1zz4AZFTl7Rul1Q+w2r84UoIXwF2hyr297RfaPWvByXkAKIGFfWNP5dNJpHz9kM1
OS7iEJN6cER9nSm7vye4fsx1yOde6z53oXWNtrA9w2RPh0tyMDK24m6QCmrYUqt9dmSWKpODYTjk
97eS/e7Ykk7x67YfFvSERJmaFYuOd4qJQI+5RZJdzG/K9l+oinMCKsUf3hO02daQiYjKvkNRrzf6
zqAhmnp2K4Vwcntzidf4y1Z/ROliz9km/I3n+rhu0VHH9p8kX02bLxQExEj3PVw0pBJ1lod+t7aq
kocxqAnwjQTggdeDwJnetginP95GWe+L8oE2AooC1rdyO+RaOBpRzZJxZPVnL/BzaU7dokOhBZv1
1F+xe9eZ89Ri9CA1X8OSdfFz9/0G6TcrJ4xsusYr8VFFnHY6Q3T0bthC3wi+rdiKDtoN7W/E0Oyh
U8pL5tBxHF88u8afog5h/JqBfqAynnBh82csszLeKfcOU//TNxa3Obea1n4j4rt7iQ0UfPvhV5k4
XJiFx/iqSlLrdpN1vXAxvN7S+CFY3U+CX2+rEhNRdErxbShQuy7zBBC5HMupQk1qmMp9ySmFBoJc
bpEFk2l/zFQKNrZhkN42oILjJYKRqA4drxdiEr+4qAS1FKD15tQX6Lat9wX2sl1EeHrrziEMNsXS
GksIiRD79eWNfKcyIp8QIJkZEqBAmPKmT49b4NzUyxkNE9vlJ+TOkZtdO5cnEFlSLThG+TctY+2s
PdnQdqoaiW68vLkX6cvLXgtK6rSuZ8tUm+bSV4izXiPmMgsefaAV5HmESHVer6/0QuKySTI8A0bV
5U/SekOGarGthaFm+jSbyeDZ/1VBGh2j6eUbGONVeotp1/QAsjSn97yGXbk5fXV8SMMeQ+PMWelV
wHkO46cUci1pO87mexhZFQBcstpqz15yGCL+ztkvmy5U1H9I7KwrTwiw+FAGPWGzCTG+V49EwR2a
v3mXDIHdjQVxTr7B5BispqOLwzumbSAiHfR9pLksrNfr+6/4Ur4BPxmoA1itXI6I9rXDi/3EIFzf
ZZWba6BDvJ15RvA5UnkdUqxkynSIJFBT+X9K31739HfOAFMQ2X5dYjw26dObcEQzubW/CpSCnz2h
KuDkkTql/iuhuNvX+e8B9StBh4HqSXdRtisFgoG+3psdcK6YY6m9y7021ykbcnVbOXO4trMF24r0
iz1QbncBCCr+jcIa2KzvE8gzOF3TWz6KLeyFBLhncKzjrvfYgJgEUVhPYo+XTp/TpxkkioX9E0gI
AXCQq5t5AYSg1h4Wuf/oif4DNsQCArLRA4z58N3Ohq3b0PqV/Pb1xoifxenaA3oqfMSFMTerPvvL
CAKrlOcQ53APlbGlszhSqNhyPwfOSc04z9dcf2ItfObKXeGFzUpLHqOoGqf9F2xVrVRwfsPZvy/2
vQIrWmGBatjeLHNW8FEMeaabLoj3iSWVbjlUglRNvdQPeT2cVniOEZwQcRmS0/fh7r3scPiWz3hY
sad1MvE0qhqHqLLK7sgRq7evxKlcGvbSXEDkr7e3uW3B1azpj+Ezzd6Rm+MKOexfcgwjYawVGDsb
NM9aaK+k5feUlMwCC/D3H5HsHcN9m89Du1DuTLMOPRmdNQ5dfro/aVBSbS8k3aob1jOUdlwKRGk0
rQTb8IE/G5ShgvzoKHYTF6FlZs8qWsYlwV9ADcLtJAY0IBVjiDjUUZuRnxCgUjNq22Syi8Me46D7
x9glAfVQhb9LKJtr7lwy75Dgt9kHX+VqWduPQnMBKlqkA9VOqYcdx9Y7IQDvjA69vQUKys5USF+r
HG0UquiYpR9uWYhkPOkOzBbEanGfys6A/Iv4wvc6cwWgLKMasfN1zQS1y5gRd8+/v3w1CR+vp9XM
a6WheRgbP6EIRBPC9ss24nrtyXRWjF7mqpGYcuW1NxC6SJQg7emmMDe4CGkAjz57e5M7M38AGb6o
eEV/k8DvISQlKE1g3PIpNvpRe6fOoqeFt4pGWxqpUA0KwwH2koVvjbu45rZduPX3BowGrc4FUdRl
djWhHpJM4HaW5/EwTw7DkMlO2laNQFh1NkRgnr9xIGzh+ZVOcD+5hbzib/6eJvVc1NLUZW48ueeq
fArwZiBgpOP8/TN9xk3oZabtPgGAHCswXOx3WDZkNY6BohpojjJ0AfxixMuQ+AlgeaYCWx/1B2eD
OJp1QFZYCY81Nd7thxEMuaDuokvPgWuIJ1cQP4YnoOi4izC+CVF1OSIzL/qsyvj0E9mmOXn5FxKi
9n2Lvhjz8OK/u4TwvsWdsO3UkOb/9EuMUJ4r1AeccgMzf2uLGPpoRss6hnexmQAV7O7rJ0Tqdk/R
hwmTqW9kPCedHdvuujR6Fv2Z4v5jyHLM6EifI4khQ2M6WOOvZdklIpestQgUwMc/x4o+ijGXFZ4j
qsMWYQdmJLc2VK/xiNtpk/2oqtx4Cuf9hkJlhkVkjxjSZndoF0JyT3Rb3r9AkVS623rxFzlkWWem
Kxd6E7v6hmbkCmlwsMK2YE4N7KmGbAByaM2vJCDh5OgOl6X3oAqmht8iAinyWi5TL0BC2TBf5QCW
wrtgypWVWOKWC36vkfQmQCtgptscWw39wBpXl+yZOzBm7DJI3anE+d3gx8xCrHyw5AWEBEPIjFni
E44BNxYG+4haY0SY7JI9ivCs1sfbKsQ9uGn/UjjVf3q1KeMNiNRG94czItztRkSdMATNbDoZrzg0
30BVdwmoCqGIKnS5Vqa8nqrieKxe6kQ1lOgyFVVtMrRwZpGhDo5QTodnmp2PR5bffn2uwcb5yRK0
PLuIwoZjcWv/80wFBIrLtOvTST5lmTkdj7WnM8Op0esKeySMR7ZHmAZ6MGTkjGld7wtnQ/5W4tSm
Ak9YJNyCDQQWzjZU4fEs+QFZHsJm3OmOudesTj6P1ZkPLHNUZbks+IdR8nIhfDf1xd6uO2J765vE
vWD+8aVTRzbBCoQwgMZKzHhPy5N1ApuzkhRT2mugXIVnvZ2ZW1hUs1pg1rrC1XRTzbG8T3sOY9bN
SH+pIZ0Ryekn074t7zdmv1sYbB8anqmGFUouzm8Fkfm9f19PZErf+ThdCaqMO3XeDg8qCMrvoSxR
VifyLOWBiznsB4d4G8PDkUULnl+8V5kv0glu6ilW17/0e1iVTRT7yf7Oi81eIzQkqbyZI7EoBtUE
Pz9vh8Az6BEwG/A23RVNMdWIq1iMcJuvZeOmKFjrCQPPx5D8kIzRTG30K0gJUTd7nja9QP9ktmcm
HdraxxFEONHIGEg3IY7DCWtQSrvrsaj3B7rIAeiuUjjkM+iORY/4Y2Q8g1V3lSJUkH9GfCH7QzcE
JH6XGnenwBcHcC06djFFWo5lg+8O42TmoYu96dvc3LCLXGDarmi1rfBVWjO+r9bh7MqX3jSYSV7M
+tzYeDgbOX1F58s7ma/FKQnl+lKfbFPoRkjkNbuUw+XcdBrvI0g8CJzK267aI23JAotdRge+L3n9
weFrJY1NV6Rd5KMffneoVVc35cijiIi4fYhqo45Slj2O042MIuw/xMctJA0ZPk4Noub8igOyGNm9
D6i1gpubX8NRx/ckrgDS42CGyGbggCMy+XWwLe4YwRJ1ZrJwAIv+mXtQcfTT2xlMj3hwzjm4a1dx
c7PFL6ZojvYMkj1NIilOO4Po+KinKDJBYf8v5mrpdlHChTejxXzSMZSAg2aUfY5opEG547SCCFIP
aTAWzPCG5W4wH+SJeIjaOi88LOJIj7VFRIEv8ymHoFKNXTHgNa0Z1gufegFWpvnoi0f3zETxoJK/
l1dnGfXRTBKd+Z9YbO6NwVtSsTZXdcJ18ffm4AHLfPMuVkM2wzlo8VAOwEEAJq/U1cLPCLIQ3CVb
iJGX+Kl8BrLSmt+T+njXOU1PsU3r2AFsQhN8unsTIrblsKjwos+rpEZQ0dPbnlvb4XSq+CDMFLVc
vA2sXqLBiCK5xPMtemUHBPX0N8im11Hz+vLRftW7i0sCX5YyNSbRxsPtVo3XzpCC0jLZCkmia+iu
Sz6pkNMYoxtD0a/P25fS7MP+O4UQRuHIZ6wzWXwFfrm77Pk7vo+x+J3Vm3uoE2SLPvVYivfmqdr7
s7/t9g3HOEZ8KQOag3AEvyRihFWNsgHvUs0ZFvafY208fYCIXWh0D49P0SFADIZ0ujGlkKByoZfb
UFozE5sGQpPrXE+TFCS2eZPPbdx9VhPn6OnJMkMBMHvBUCEjN3zFnqn5IqDwIknCS13yhW0XBfr7
6YM/Hkr2tlEqlYV7MPl9BCf2oTvdcwjaaJbBus/5RXSAcmY+sX+LmFLVuMN2b9RpXEkA9LEGk8LX
TqbDbVMYoPhjOrnzIsUQajYmNT4s0FztyiEb7ZnYjs+KUyTrBbgTS6wand633xtuQjBdeYPKwhiG
CTorHUIZyDeAMwjhImlWeqNbrCeUgoH+WUtMMT8g6fBGfFv1rI31migN9RhEJyuziCciX8b2O0tX
MhkTWDHEeROZmCQC8Eiwg8iOdvJG8RfVZjXqV8fekNnkiZZiotx9RmZmp78/J6eSJGJIeyHjrRmm
j/vvu/AWeLfEO/7p5KVhSSrY0g2woMhs/5dCOP1ueL7cm73nLsZwFn8Bx0pnI9g+FsB5cruGuFxv
r3SRlxjlcXug+9PcmB083fbugbMSXZiwVVSfe5Mf0wIWaj/C67ZYBqr80nqdZfKhEvaAgZr+x4ij
FiLHQgXLncl7HKHV1hnjV3HuG35Hnzz98BPBdjLzCpn3lD5VZ2XHBsT/cq6AVL6wZbGF9qfNezkb
nt6/Ec8qUn/42xyq56dHeg5dJINRPblvqNM2HdQIBpN3WFew1p7si1hrLnvvnA6yivN75UfW+vht
pxVfIG/oesR+OS28KQ77W3i5wHep3z9s66XN9TKzNulrMpu9t7XgN+WJd80705MsE/KMFpEIhs07
tvnh/B9gFiKcFhw5mmvX8oPUMpzryaAJsqfCzQDd3boEeQ5ruMT7DVSgsravFyTNd7qXXiM8JpGV
q2p/rOYKlEQ+7rAt3DdlLLEEWOxzARFyqa0QHmshERHjPRWv0t1e9jb0ahRrVXlayU/GaEhLUyTE
UcZmZP10RwZkhtCfyDjYFPymW2O8hJFwRTbHjoDvwVvYGY647MNyXILYR94oLUAk6npQh/A9wmCs
0+pRC61+RY11wmBhjP38YIoX57BNytyGeE7k7faOkMSuRa0IX98iNZcI6Gn4+gi1KIom2+45mYGK
iJn/W8MqZeMZU5gi2PhhAmjEW5w8oKaFUJvod6A4ar4jZkbfFOP6jhNMeZU8bvpJP5AdF+X1pLjx
67zBDtMlvhr8c7ELGn6wkaA21RLwX4wU3pWw3bfg0Y25L/7hi/C4+MDpzzdFoMvapwdJuvSN4kcB
bbjUI9kY5VU63++xULEpaya9AAqJCInA+pItUAEuFgXA5UW8DWRETW3ZVpngRJvAjKVdZ9ROova2
FJGocfherpQ0xbS+Wq0yYebekf7zGzB5mwmnotfrRv9/f2pdcNxCRXlTs9UbeNMGHn/ypN5M1U8O
Bxzi0dRcZQUvW1hiU1Uhjl5q5GGHAJNWJ6hWea4nP2lsNSI1zo6ainXkvEL50bnUD0R9spjNVG24
ST+Ne0e563PEYx/UoJi1aA4bXiDNt43d6zNPyBzUXGkg5+ydcXlvBJQK3K+7sRkXtdmTaIqE5wg4
xK7ZXPRQjuz1m2jwbEU1bxitXJRzgFPxJIBXsAubBXneymKXAZ+cmGoH6AspDRRB/EFyetyxhkBq
BTtApUZM27QOWud65VNxQqHueoy2TxOS99s9ba+CXqS3SZCeGHsmuRxEi/NeTNql9pBi46VCY4cv
4ty1Xqu14TUIGcMMGg/J8Tftv3YKFRFzgj2CzJ8nn6MjDO+QQ7T2z1lEKfULYZ8G7oz5xm4Ne5GZ
TEC9070rjM3S+RwF0PkL1RYIg5xVipB+xXDwqccIzZUoJrmsDYIpSUr8EWhsDA3sw61kVLvwhsmi
D0tWLqJh5PGY9BGvf/6thLB7rk3M2xiIoSjueP1e14HbZNnk5CX+9NFQXERlnri9Q6dlS3ZTTfu1
CQA1eqks523AweJyDDxOnN17DiMPeQy6xLjykE8iOVEyzgh9z5ngQmkjEDuF2KllLmXvXNNEPKx/
StYj5qQToxqbvYrDrbu3S3mFg5xp+ku/OO7soApQjdO9znsDATY3YiO0QSNClbcKIWlxVTx/idFv
C41pK1kAar7nRtB2fsBAZUH7zNnmMvNjAAyJOznNcOmFfS3Q8q38VJMjS86vT//fVFQNGSQeiC+e
df/sbmza6jB58Wtst9El83phQz8TYqQP7zblLQYJkmwPI4tHaiFrZEkdFrGd5l8NBXLtzKRCWhrK
qyyB6ul5mdn6J48ug7vMg+vqgPaqCl/im9Ya8MQodJ95SKkLxefeCfUliFIHIl5zR783oQ3eJq9I
yTiC5J07OLP02t/r0bxXKOnxjm0DdbmqIuDTCnUwiZAc2K9XPi4+4hTN6pm9WC2mB6YRzTOK5VS/
bFd8lAKtwwAKBlt7VsuCaY5U8Fd6n5v6S43cV4aUDsI3899msLceBXeU2IAkoTwo7OEkqNJDY37D
5ztGWvwVQjQ3PF5RviJ5VDRuQsuCqnZVditqy84KzM/2m3aJHolAQ+O6J26b4V0mCJCcdeMzlh+O
MjndiPbWQFihlTjRu7ltfNDk6pDeRTTgzNVKsFMyAJArGIBsv4UrvZD4xLgctpudFRKu2MsKAB42
I6ekf7fkcutLWWXE/bBhGvRdLcRVepXqIZmFqvYb05gS5vX5EHpKMLkPXNe0HYhvYndE2bcrAvGy
vgvXGCYu3oH2coLn4D2igEfZihrjGxZ5TrkaM8VX72uA/ZvXXbMriGAlCEzjw28HcUOBTmhI6PLl
YYHsNoRAQwrYbu+dXr0WpmZ+qATFfiKMj4/C2kRbPBsD1TJez+fZh93m+lRRXUG+AKT/L4QEnwag
OWsAYEtXvI+uuLbBlQnNZGOKHbwZkH+EHgJzOMK/zDEVVgu+R7JjrHwdTu3yzQFF6xcwU5mUoqqF
HuDYJqn9m33bOCRv/pFiXiRlrNOnIQB3znf0YZeV8VCicCjanPgvFBiS724fqZackLz76jK1FMxN
syosWAghb4p+UedkXS3va8bbXmzg3DG04oRzwD7l8+WWRQRg/Ee124Q9sDRPfSzL3i3ogd30ZN/Z
AWH8lNI5F1/WAKlgQA42frY7NMRSiXu5yOToNFNUylLVax26SobzeV0PNn6uNAqC0DuDlD1joBXO
vumGTG7nFKVYquPZNWfAXWVz5yGTmDgkLhBjGlgxmRCnrnC+aGodrj2U9TANbMdOzpBlM+eadkyw
wURs6sJqhj1ohE1K5we3v8OsU30z7maqyitebgFTQD5k8Kz5mhzjpwok9d1mnGO+JSa71H8OsK94
SIp/SsZKzDjIYyT8I3JKrgKbzgQZbMVPnmdKlqz5bwg8IY0Hx6dqtNe7ZTfEVqD3h3xBFYZydh+X
UQJp/L74p4UWqa3+BCf1lcw4MeKhBnu245A6HP6mn5A1QIrvJs0qfvwK/Flced4ZY+oq0G1eRjMN
uYwNqIacm8H5cdXxZUq2leICE4I0JkiBEDOSF5aWWgHIyDvDldHzpYUGORT2jR/YbiN7mUtN9Tfa
oiN7zlicUOPTI+UzRmsaXOmVF44dQPzUEcP2rAR9abVcneqmCX5Qo8paiotu6unFZMckcrrCctBm
Ud1p5PxYLNud/38mwG3borD/4G2/rtRoXG61xyOAzZ/tcggwp1sCJ3XGi/WxP78N0oYUaoDkwvLn
svBRayFvUIcFdO8SOCLFDHJaBp3PFOupj4ZamXPs3l/J9eBwQWDWTW87Mi5e+/AxPJay3MzWI9C7
7IWQ0GkvIrle6TiWf9xcWsjdZd+ADJ2qd5QuhO2YqUWq/8t5+dYcMU19/QrbbOLzsn/sk4N8/lyZ
aiwT/sfhqWOAYpHOcSBCjtsxNlTpJV6u9aIaFAa3dK13k3hd8iYj5A/hCFtJXinZdqqoG/T1APKk
O4Kq71HPSoA/lBlxHvceCaH72jhTYcPzz2yWcNetQKP87k6eYvybiMsE2ROr89iCebvwG9lH0C1d
5D9osd/qpgTtFdD8WM/OSPgsghvDwM4o5cOAN1/5a/DNWJgAvm16uFdhbyI2tlpnPXs9KkxE4p9k
Knw+aRWsqZA3shvFLrYb3EXj6KnnJUitPLr8M3nFrwUgtqr0qF6jr2VDCMTER5sNsXf/j4UYsiw/
rQrBnbjp3oUkNFz83CG4WSYo1bo36bGWyV8pOW3L8FNFzbjuM5N0oYM3YcYZYHLE4qaWLYhG5Z8y
OrBEC22F4S5ZzxegAIKD3yHvsyyyRJa+zEluywJEzj5RwhVGH+1ekrM1PKViMC7p0oNRJJKfMG/X
fLTIuoZZtDfYqINO7MnMcx6c0htqHu1nQcQzXuu/1T4k+GV/aq4oMEsod2uJytVlmEO0fSLFn1y1
6HCYVWC17NZqKbkoFnGTffin6PE4wtbKZQcA9bSCsNRqpDswlujRKhs7AKi4dyCPspDWdtFI9viO
x+6ez5Y9n6lRPxoj9NBMPWBayw5LHsKdXqxEs+QweEjA1mBig5ebIBiHcnPaUGLBB5Nu9oCE41Yy
dOAkBM22PU+M+YMq24oArMQvLrhYVmEapNmi4Hs6urhF1gpRF6Y6BluBMZ3IBRjysW2r+tcnokE4
31hKexCE8UMi5nKWj5TkRdrvLRvc0542wtrz8C8/ullellqKtC+yUO/DKB4xl7gMJc+/yQa8CqoJ
lyIxnKHLs0qZ+7pYGxvXU5Q+JVt5LbLhsJzC1o5ci18q7ghruOaeeFUxGDJrlGIor47aLG127OBm
q0C6UkuyWxkTYNrxkcf01Ybg17Rn+Lap1c8VtFRXG7oKWC7/NesNH6RNNW6Ti0KIV/5Bhq+t/5gF
SCn2mlhO32aULzhiL4w1eF4tEK5xNVf7Usz13MLofs10g+1lQLp4dPxBMkxpHR2AkTGhHvkO2lQS
cPIjT9Wra9+jHAho8Mz5XthOOoN7ZZ6eqexMw2ac/bBX62kL+jOq7T0j0ba9+E1Tzpg9gBRjDlp3
HaXD1XLQewVBC9yjZSVcEiQwu4Tup6lmOdg+XT6QkUU49Jp429DHdEqzuEPKQjBmVQQqbGmZ5aqC
fdtT72jXSKKyO2p09N/lO4zqG3GT/s9LafTZQ/Ty5iE8uTgPmP9fEt5oZQMKWawtJFMSgNy+QMRC
krU+pkM2UZUyu02faJ4EGyfdJvFHCa6lO3u/OPpM7RiiZVmDCbVKe43ZmqEiHlbU6SM0xTBCtj8N
OJTSX82zSbs++bYHF6ABq5sirGi170diWVcJOyX7pNufQV/V5JzkGEV+MyNp5UlBZabQvPjPU5EB
PeYOjQ1vh4uavaxwpUhiRT8bBwt6guyFsLVxqx90qaBD6QI/WAtkzeFvUkZV5QFAP7YtMraVK4+S
BguQgAsj3ykTppDLc6nUOxNEJVxQziPMw1q8+yz6eNUevFjT9i6BqBE+iQyAm1keTxglb6E7DvX4
fqgzVPYc4pOAuQ4uiAzsX0zKac02YmjjTRv/3QlVbBE0n0RwZZnzbQBDMEum1VOw0En8Zfs8u+G/
vidCdN9LEpNlq7BmIHhuUwlxgn4pKIZf3EYvugCNRoC3gjcJurz6iakSWmGjSTWxGEC0fIvc+5Lx
M/RcbYWJmMUElXwgcn+EpFagnOtYkFz2QBoDOhXDgvPYQ3gG2Bc3bksvrNRJnra3gowyAkQz/SlH
et/OZCE86ozCvUjBwZFFMTwoUU2xEt0kWX/lz9bbSudr7RcRQ3WkLgAuxU+lZjx7GEkhfA6RO2nG
mQQ9W89gLnmMkBVgweqJRk8o8Nyere+cz2t2tlIbR+IyRTgg68h8PW5AdU0yOo4vWhf4rJf48uOY
FiZo/c3zrOas4OVkHIred79xgnQE2UkMhvgstvWgfpQiZA9mUkdAyNWjewas+97nEnnqw3iyThXR
CUsZPIOFu7MALQDdPpg4EwNbw4Fq/95J+iFLA9fyWzmg9WDi+mb5/FM1Z5njWHPLI0ps7PIZU7rx
nqMBU4FNP+NyLbuyFzml0DfPcKT3vfR+xa9OtnD3pYtiS9H2RI7iD8jvIqwDbg7QUMq7tPKJVAdY
29jrMP8O+5esy1Mh2pvjtMJ9F+/yr5C5dH7ljeitKiX4FZzF8vQ/NNdzW/xsaYfPqLZARDPV1loX
GLlqHYknuVWCe/EQqNejghF74lnJDFEKVdko+yJsFhxfxReZF4sD0R/HyOlJJjpP4ZR02KqrKKX1
2zl/P6zv2pqQ6tzundrWO6g+jN57l4Owcv6kjq1j3tJLjnvMh9ktw4G/wviEG2WsFXqu7ZGUvpdi
sxElC/+DsYqq8BQp6wQQUSwhG63656mxbWhJxu+j9+s2M/JOXYUFi6sOj96gsW/ipTeAtIWxkQiW
eiBhg9zI62hGt0Qo2/q7IW3/sWx8IrO6TZd8CNGMulfhoH/Ltoqk6dzTvxleWzeTEPRy4ikAQSkt
HahkaCvH8AwnZAHG7HIDWHHFIRJY2EEDCdIg3IyrnOwIH9ILQUBbuvWsFcmHQK2urFggTAQn0OX2
2h9mLb0lGG709Vm4m9cqs43oWQ7C74BZaqawFDFy7CCZql2dAtRP0GQx6PWwdej1a8rvzcPxJ82R
BhaBq37SqvZDnpGe0l0ktm55/hCH0qJswm7QRHUI0jjaePxJGmg8YkpH/l/IlsLLCZ3QM7Lcxesm
wkGkfMGuTYTWEpIR+He5l9vgW1ojsVE+LeFVO3YaBD4yLMa44V5GTPGPRAZAcx9QKi3tKN76uweq
+886Mjax+47NidLxrdmiM1Jml60eK40q+Nc6Ui4ndVLKpXrLwyWAgoqprvmNN3E4xwyQo8sKyBor
Y9JDxkwE0DrLBZc/n68R/y1bCZrCD4+icFAEeySHEn0Zl+vOT+cBKWtjbtezDHslVOHOgZjJAzEL
vw4dIrpPrf6Um54maeSUnt7R28r0n+/Ja6wTZHX0W+w2OuIfgReL5vt+qVexKHexNiCVbJOHk7Ut
2fqub4UQbci4HOs+F3VYqISNZIJE/8XASyVnRFCsT0UPi5QFghmT+2FjNwN5vdzlkZKBIemFqhEI
gCLJ2GXuIXBq0WxpguzmbjtqM+5DZWEsLfHVOSaoUcr2gtv9uKEebg/fn+FSPWfttjmhmOIvQAAO
mD3aUBSndJ7EvqI9jbSXYPnNHH/XZGbD7F+N93yR6KiDTuNCrmpM0ihM31n47sloSi5UnnOZTWAZ
RVVqeEW3Kk66zr9JkCYhiEImMrCD7+xBYw/eQ8598ZZnVYZSZUC4f/87kw1T4N3rAlAwB8P6EnPY
jHiKR42OpfP3l7T5mmfBJ4QjJh+82BwrqTGHbhV8OPGeueIctF30NlYcn5IGPdqToFkz2OpPguK6
LSiQJXz1X2GByPMmuS5VqGmGWlnBZYjEUGDj+bGdNfMwqpsjxp4d+eDOh1+BgPTS6kJltfzTjPEx
x6p7/T+lCcl1pBbzW4CXVOgY8uTNMEbudagK+/MW1+Bc4MoKPCmlRag5yzFl+7Dm6t1XaDXuzuTc
zfaTXMO6Y7Gp8DOFq9VBXB2DcZZ9KDZYeGZorOSu+2CnIfCB60TNcNQTAB+becxb2hAgxk4bZ6TQ
kUeApVAOTjUstm7lkQLaMqDqBTQBFAWyKdjeMWRzjjiOHl9CQJpDaVWJZ/bxxe8jUeBGfEWl6FMv
zykKIHQX16zfC98sAapx6j2NswpR0D/ghm58NbvYxOq44dF4j+rrSE0rAOqhVhn7G8aHXtCLlLrJ
BUVXvTEPZpP/5DvqWG8ONYw8MBjpcEXwFPjA2hFVvU2HLTcbA/HEgBMVKPx4YHT1yqKRMeuS+wIG
/qCb2u4QEM6vjAe+Z+f5FnCuj3852598ouKEJnXyTUfPX8gIhhbjy5fJYE68+6QErVO8utjtK/eu
C0FqdN9k0kldfUVoDLzLoXmIPVjjMxF2rE8zv2CoCZlWIcPXpPuv6InYdJPQTMjlrNfXpIb8vgRT
41DwY7YCJl+NhY9NxopCuGulF4fnYAXxZ4TEBE0Z7jXIGj74PFl1g0MtAw5t3c3mzQ19LjX16lh6
fhlUBJoCGebbfFm0G0qIlztQ62OAnwS/1mcsSRe933KHCruCQlZPagAjnmXMqlFim7BZ7AJFTtBG
jXHSzFxyWEbeS5/IC1jAfH5bXlnXNaMm9nPKUGU9o69+zA/26JCC2o+zRGIbduImK7i2WrQD3xU0
PNbproFNG377HO7U5tXB3r1V4Xkb5aALSbYii5LBB2lt56xLLrdFNBF/jV8XNsuehAHCB+W1rKgL
HQuDJ629e0j+SIgiG0VaxeXenolN5p2j/aJTg67d6IUvyPaI3hlEd5brVH31qccXAD/K9IB9anLl
EtQgs/FXoXK/OmoHT3pxXKT1A2BW3Yievn9MajcaWGtjT76DWgHz+AD9G6pUIeBlj+fFdUvnfGRb
KamXLKunk8b1nu7/lJBZUWv+i4NXCo/CzLAF6EB5fNYHHc4H2Qn1KzbvoYfA5H1xS1SIwaO68Gxf
GLO7Vh1eln/QNTDczWwvwCjYURNkNqFyPRU0WeQlz3sEkgfbteoYQfXZAxrhzl9UjJBRCfJqO0I7
TDtqEeRdm3Wj/DL+wXmHZ4uE0LdwddpV9wFyGkF+Ju2bMW6K7FDKSDxv+BslSMMYeaSgTCsayp9B
78/gxM047ldCBcnRXQErg5YOx0nbpobIm93SZRRblWvdsNv89bbtYJRv07i401+7GX9wBmfoKjgi
nbw/lAaP5OAsfV1ACL4Y9N2qgppOAD79F7OlMa5WR/Wlrq/2cryFscALtow7FOuULdGoFf+yqw9e
kg4itN9cBFzZVklg/fdLIdWaP3/EdcqVpKWPR+7CXEJmq1Xl9lFb91y58nNPgY61JX0DH+0xvXb1
tV3tYcUQafIZ1OfjP4UY2rjYJnxsTYJxNEB0PBZq8nRGPFUlnrnm/935+SBQdT2n9VmGd0M2fCxX
B75pEVwBn0RKTwaZwZUScLcTzcqNMDcuLiBjQiPvBnUGiPvbCiwQ+CNjckuP7+3dsvFAXjJtoTJu
i1icZC/laArzsOPvMBH8ENqEaGkVNH29thc1GKTHK7Ce1unAy2bBPEJtB5uFP3G1XA5YS5tdNs0j
nVKCQ05JouDRqkXmgHQZ2vS7alPYv6FFerHLCfa/w/SxyMRdOwaDFH/dddxbQUS/HiCbb52ul11P
aHLrLT5i1Vkj3ZTs1yK/hIJekfLRFe1levgPlGO/GH1sBgsSCiTe0KkzmjcLGZO4b4v5+gaViEs2
B2oPMEdw5GGZIwK//IoQ6XFoudVDi4eIafwJfA4zYURgB3gPuPhsWtpvm8SPLV/HWSxjI1ZSuBFA
6XMf5y4CZaLTPLx60arFeQR43IhKGnCUS0y/fTdFIuGOzNGAL/OD43L0rATR39tjgwHIrdiBTDdV
qEPwTCY9RafaWkHIyNHYwFDuvWSZV1hUEgB1J+hBRhgmHICv7m07qvA+L4cT2Ja1JCxU9gVESE2S
JLxjn+u9Q2yvpKvcfrOk2wpuDK9QaMLKdxG6BWjti6+Cw94UqCAXTyOBlTacViksY0kVQowBUJMq
JBwFK4sMmO805V9o/2iN+GiOzcUo8ePcpc1Uo089P5x3FCK835ZVXFRnwKAR5zJjgMe5xXHj0t55
NE5f+7k8TW6wjrPpe9W3hYS4PWKJ+PbJgXRNztJ5OApdyjOBNnbFu/LUlRSLcmCnfniMJfQaogd/
yrR1fOMxrnhJUDf32xEBYtwVIIZ1kC6Cg8pHWp/TejTF5HeDx5aLM3SNaZp7fSZsKd3Nrd6u2zCy
okO9Fsj+YK5f/HEqMZ4b3jTyhSMDMEymteB6Wb23ua3GNar14ZJqse1dsaf669bBDqlK8YwvJzVC
UPRrUzfLpH+KAF3a2CTWkD72i7Ce9YM3oqcuOtfLbORzOuLlTTjBoKB6gOmr2PeXsX3AjZ6arqk3
WyuJ6i8rwUY+tmjfhiE196ikCSEgLKWlVVQhG9/H8XjeenNasiWwr31ekwaj3MM0ywqR97JAU/+U
e0gBTQWfqNsQzp4iU8ltfWhA9+bd513AmnUIotvRhoCwVeUYGNNGsg9fUQCh03xa1Ve378Z1/lTl
TAypxKyj1nn6l+4GX30ZsII78leBaVDz/eArdhvxaPvSwdROr5k+n9BaLgz+nK8CS2BxjPMdrK3t
Jf6gsB6rD87xC0kUJPJd2htXHHNNab/sf+VEzP1re3wRPj+tED4IL/OK3awtQU8PQRaNHMpLXRNa
1TF6aiKV9151VGPtA2EJsUJJJ9TtqymnxQnCxb6zyqzkpFm+kpWdG2x05+1Uxan8WCu0dI/9VmDL
QZ6neW/FYoA8k7zhTCq7DF1isXTqhkz5i64o2nbO2+Ybm8d3YtTFIe/OUInEdRkcVxAlphCgiaEK
1OxXJekwvJI03iXyMlP7x8WVWSBcJY/QSgnyjEGPBNfmAzCwLkX7GG2huuDb1JXgQqZGw5I/5apD
t+SqW+FRNxE+YzCnTeaCK1Nk36wanORoPsUa18tC3Vn/uMt5ns3KuQn6VsCZaJ314r/IOrQEmtcL
2b4JNTpJ79skTULEFahtYHlhbIQb1n2JGKQHvYwAEfbf2iEyTBiEbMAPBYQ+Tkn8QH9npGw99aSi
x5vZiPwhV/9K+AdCDYZxj/CKGoFwYiRy/pkpDezoCztvquL+QA3tBYXGJ5cuCzx9YRkg87QPyL2G
7XhY6XtyWkmv9xmcAIWAzpV7YtKstwbamiA2uWBIBqFYZsPh3WiMILkWXJAjloLLZxuAPcW2Bm8A
6/54qYIL/Pq5YK+RrhrLdHPSdzz7MuFSXDYplwo/5PHpgvlhA4Ngx3SgnnjFocM4FGF4YaEs2ljx
ZBaD0CQNM0sUVZasX5cJjT9kxFZlgpdT+nMhioNjjz3hOhaxTSMAxmpM6bU9fNT4bvVrvkzhwV0N
FdF5A/ZHnbgk/1tN/iQd0cQWUTctRVQLez111GVITguZ1RnSflCF63S3F4q6qxEf7AA5q64Hi9Cx
dUM22X8aaPkjk8FoUaXY2M5+QBU6dg5SfSGXWeqEZs1lB3PMGnC4QXBbgZGLC8eKmNBlIdr9bOIn
zQFPO1QeVVXFaHryLOnNrBFKF3EMaAc3HGkHhYm8kQg0k55k9hdj7+byqAog3yVA1+EgTYG4Esqu
7lIWMGAWdlpFkMYLc+ldBKSZxr5bO5jLx2jkchlupbH5Hb9VR6e3i0blzeVBBKASCDVs3X1Wdrwn
dM0yjl4luwenJ+n8fGEQqWtupbbKW6vE5YwivovjhiXGfhA1L1YcUF0Dfx1qb/+DB+a8KXEs26Vq
vNO8JiZ9ZMLO9E/OT7fIb0AVtO2y04TYetaj/9NgzrbjiQJMB9TECvyeXgK4L+cpfLRC+o8SVusJ
bZ+onSxaNUKYPWCuKfd3St4oAGrcQoOb8r1j6bBUOjhyZZzwDtc8Yw0h4OxLQtwel2liKHlzpUew
8t+e3Xra/rBYQvrzwWa7yBIseLAkqf7BjWYWPf0MSbZxkiAgtOVLMWPBON65Z3hiUqaZcYKFPdch
FRbCJ5Fmsh2FBglLWuJ2BvhLOeVpZ9XZX9n0KyIV9MxfQxIqUnAUfVmDBJWGv+P1iCFvksThAQD/
ZdAPQfDdnsYkXwAPgLJacW9oUJmKkVPc1RshsWjmMnZX7WNwcS/8ETE4sOoI+r4/OEHTppmJsH3x
CS4b3Y4CbELjb/Hys3acl7byouqmT+ka69oiQ4YbRvV2BpY5twV4UqlBX6o7h+cE2weOE5BZzqXD
IHf403AwcZjmgj3QShBoJ2ur6tqJ/5+rb1Rv23mthKBJznaHiWW3Tmmcief5MhdJNd5PUa0DN9Q4
m+Uk0936hAdrxeGTsDR+SyVFr1Bvjn2BsDogKZaHx9DnW3xhgg0ZyhswSFv/AoC+CY4clGOtFutX
aufJiadByvy5PXQiy2/l4MPyLuA5KayzsvnztS5Ef0hPOxBXjcQIc7VTCXUTgUAjJk3Rz8ywM0nD
k3GQ1gC6uk47FDlk7oC4xYH99PEb3reficVjuYre+5a5j9dSC3wDgLZpdry0pz7ejh+dWP15stjZ
eLq3WQ0KuK1SkWb8+P1pANQBTt38bRxwHA5MfY91SPT7MSOmWms2WCVqptEy3x4mpq0xzdX+97ol
X6LQJuWTxiSNzdfdzhV7RjKjRvT4wqvlR6zb66eLnms4Th9qesHj1JcksGL5lqZLhD48Y/WtDkML
x4NwqKz5Lwpbj22vZG7Xn32ZnZ12OE3ycVAVk7hhEJKX7oY0q9R4Bas80dyJC8+V4+Tb7TePmBrA
ojtxTx9Hz0oqQFocxi5+9tW3ZGY/Qw1B6QXq27Ik2ZXvG69OmpxjcjB8vdqxvzb6gUHyBh3V65fO
RagAp6/EPn8MvFc9UCJB9o5BD7MNv8WUx2o2DSjWOCyV5Dd/uB9UYURhHJ+q29pyHYqubDTum96T
KOOmQOqbMRSc2cfC1hrCf2EdzuvN/fzE5X6m24ulqK0r2xzY/bYHoQn2+P0CB3lWE7nP/yw8zfFq
jC0M+BJJKk7kIosgQULOmcEOXKsPQq11biCnR7zIQNzQlFoXbZs0Y5mRDM/GS5CLBoP3WcOSQOed
KoteA31GwBpz9G10JPTNbf49zvC6S1wZk/vnMjT8Gg1wDtCUVUr4+xeIlktTg5Ij1hGqiH6NiauK
K2aSKPjgS1vaAv0BBS917ClKlqFcHGtlkiuuE5kHNSlKf/BOaJLlQ//aBu57FErHxWIU/x7o1WOP
tZloM5Yfc0c7yJQ0xYCR+Jo6Se1XKfQBno0U7wBoiYR31gMH0MeRBq6AISuvIUIZjbjkuzbIg293
qkYCMW4qEGAvYLU8hLJFqp0ojPIP3sHIOxfne4pX8uRyTSlqz4OdqEno6ZdlEzbj7IC3Mhf8E/t2
ufwzUF5FPiR8tiinU1IrVicPpGZii6BBgCFkO3ZxXz3/Irgrm1JaCPBGU3HaivzQLpJ2STj1+rIE
Ml2noZD3E7ptuV8dnzMo0NKlnIs2er/M0mA/vnYgyPOTvuaX+85fgdlS9O8f+d6s8BDMoGbOiWXg
I5kQ/uREry3dSsxcGBhM+11sC+k+qlUS8H2qsrbZ8TG41p0ZoSlDWdY+/wTyom+EJBpnwh9kN3vK
Kq1zVvy/ZO2iZm8ORRENYqt1htGQpMf7/yJAhHiLQLOp7SXlR1wujfR4xpz76QZGH/XUIhHnY9qS
5YCOegL9SzULTM7z07iAIR80t+AJV6oyFZssJ/B32T7TYhmRp1mRhtbF0jcJLwUKhqHxAHX50MAh
5ItGBGKAt6YOe2RPRHfoFRd9j+dr+JBlQSGUAAbmPTORcs0boUtfFbUjGI6Nj2gx39jmwEBSTRTF
W98lSQKZZMsRzz/I6XoEhRKhbfV2Qp0JT6OHin//pqzrrW0Lrm0qSYMVJ4n6VPdnNtL3A7/6Q0hc
RmpaaoakFnqKbtU+UVWW5pHggU3dxhnXo/nkiakn8gHJ+LM/5ar2Uie/v+a/6hPvpb1lX1u43KEj
m1kRv9bPJPVzb08kX2PRjZ3u1xn2VpzAu1H7TB/nnHWlU3/oSiNJMRSPndyPVXXA3GRFfyXxwWI1
QCxHFq4UqvJfsjYy3ME+vQ2c1cvxgmvA1D4ma2UGPJXTkC6SEWq7FjWkyf3B+w/t/0BX2pna6yWt
+SXj0yyaa6kMgQl1U7dHTxJZG3GtO26UePikRsZG9hyS4bkhBE7yDHbNnRXixUNLlJULhsmZSF9k
moYJ4J3cgF3RTQKbJ0/5HRi0hHCoM+cazGhX8gCepvoDLeBrJe98lF2NE57sQCMKOheUnGnDyOeY
/H0UWjvQf5lK9gLIyFr7LC/5Rdcv1i2peG3zfhBaDPEZ0nT4+dLe+XMcv2iRjhr8L9A2PThM51V5
z5LEXv3U7fAHrpyH4HtwPeQLnHjGgCvn2qmgPb4ANBGVxCS+X5uAgtqU/mWuba8QGNei7wkq3fdE
Y77f4Gyo9HovITfzTmfqDS2ipEnbs8ntblmCPYCheFYhH2N6iphWZsvFQvnOwEmciVxW1YvSjgTC
zYAnATmP6T7I6js/TzkKFU8Yb0WFRQw/MFAhZQPq/B7lisb2rMjk6+XNVdUsZymDXlHs8bwVnf5F
q+CKEu/4LIqj+xzJrKz+P05CK/XNhoC8JqqKxO5BPrqL4oGtSz24ZGPLYGMpzABVHzTnJmO5eDL0
5ealVdDaONC2kIqGHgz1PrqGYVi2dJhrw9rOZ720/9iLKbpQwBnq+2H8y7ZqQxDk8pMS4M8D7+N1
JsjD/mGa8RS5O+JNG9PisPmBhKrziX6Wjf2vB/iWpi4QD9fXb9RIUUufJTSZE+eIMM9SRDMfCnOg
af92dYbCOaxnQQnYOolU1pVTJ03fBFBkSECAsCEtCoI8UCvl/zda8gOj8TdDGUeYxw/+0rIoCkZy
qHJca63TSyOhGmVR6AdZXfuFwy84DoTAmctH3WB6EZ5mee9dKdRjNmlhWj+VOFwcIAmXVbCVfREf
0hMvnw9jjRJQKgUYN6DCGWOBxTZGY/ERVdNvYsAleN6VVUu0qv+EEYkkrpgQzAsZqoIO/CYtWzta
IJMSbxoiwpW7vNst1WvAsehgLl417xeXK4zsB99uRLliNMpvG5UgjJ62v+bgDsjHelNwKTznUckw
9TfhdEPRcfHThOsET69JBudFysJCdlnLu45bOSL2pHAweGKztlE/DpEO6xcRKLTC2BN/f/26B23y
wLwijnjIqN/E+mUipGuXMmX+lyUMAFSnqp36EdGdvG3ABvZ1l5YdxLhRviruJTUcBux40XBYZT4m
Qos68IiR2DiwZEaut6wTzS4yf3w5mlhixEBIxbBAMEfv4XAsXCZ5aP/GNGImNRSj7utbLNgPqr+w
jxa/1eYMhrTNoD0asX3qQ1Zs+gfLRaHs+paBPKC2lfyEXTGQXr2lNLfdhJKUf2mfdBf4JJz08f4s
17RDPhPBnn+jY/Bl10VGzedRs+GF9EbzEyA44qcng4TYG1XAVvYD3UyUV2+zkP2YrnMR0Xozia2W
gu8U1wvu13An4q8N9OkEJ8H2tBxlGlFs9HE/KqVIgsOrWvIlrn3B5lwbsPhbMLroEQDZEMYUd6ba
rz0EgG/DThf3JxRDphKjaH/qcLYgwaipWqtizNDmOLxcR/p0/bw+Bk+feofkak79PBvtp6XvN1zQ
4KBMmwSdAyXB/9xCvncHb3YuqS6IVsM62User2NB9mVEbSNJLLNhb3DxEezvGN26+ZXbo+5C6WvH
m6/cNhskKQ1X4b3LtDw8lSYhq0ZsIolRMEkoOP/bqrKQO39vAK57DJFu/mZOlVTuKBvbYyBPeSib
MWrCs+BHl5KxT+cN1/8pL9cMhfi2Pk+2o+91mqmCbbqnlg/Gu9eug9edD3BP6t7QcVYPQ/+CaYC+
JZ4SIRe2rJiTBK0lHu+z4xJQkQFvMKVETwc31DMzPD1BsQcNm0t/NgEu38j+1MAlic46gTQwV4t6
5B0p4awHkxM6oGhzbCzto31CIYVqQ5NozkUlRHux8bz/miK8ahcD0wc7HZ+/jCVfK3OgnSrD5uG+
meuPivmpH5JMXgFa0bpB0UCevYeds2UO+5tqKuZLd3DC4KdAV72fljcZKciRoMus+4wdMlgcj//Y
K3haFPQj8x9zfeUWtR6zgoeFQRbkj0VKo7+ogR/oMA1hghQ2GYSQSvIQu75VSI8ks7MHWUqAw1MQ
XyiiywxZROxqdHwCBUS9EHzBrrrATrDWkMuLxgX66TIuy1jhD7wtJt8iKPpiAtmlgXw8SE3nazvF
3HY2+nu2KGpuByPmFIsIKHmCQDRQZVoONdfiyOkXeLnxnAgzHlCxBI0o+Y1cgAieAS0n0R4M8ge1
ggJNOJM4boG7Mh8vJ4tJmaNN01zuXVR5JQrq/becA4qdI6Ooe+B+0UxVxRTBSmCagzEYNx1MhbkM
cT3THRjkr/WYt4mvHOUtdhgJN1D2BItfHKo+uENmX5ACeW/UQ8S/WFLalJDeQ9hEDbkI/OhEHJt7
zXmEWJXo1/1SN1878N1aps3CGYWUhJDsQzUEYctiU3X/f6Dfu4YRxtc4tDMcrfBlQIKM72xoMbM8
9IjklncG+vZuOFdH7nTswZu4X3T8KLo37vsoPw3ZtbXwgRS4InryKKqWbiutdq2gXqwmM+xPN+mz
rzzY0/6hr+VU1YJk9HJxD4nL+OJwR8sc0bPWk2HogccP2aRCzIQh8zi/7LfcMSf4WjMpcVzPv8e/
bTdKjKqkAj0PoTdgMfKwhai0UPtmk9JkdmXs+JTshNI7HktwOFcwg5EEfcIbIw82VndWwvJolpKD
3AC6Yi6Xi80ah0QGQvbwophCB+RfRcEiVw5awpneRndmWj401/uMSZzBWRrMwufgCZmFoUSX9iQ3
wFT/zJm/+lWw+yj7/TvCZGU/SvKrowIKhRXTtkGkgrJ9oPMV/HXDbXD6+g5/rZ7/3MzGURYXvC2h
+IedOUVOvIXsQcE0ETzRJSvYHTcNfi/puM9yfC0onQvSkv3lozIypwignuQcLvyX+Kox/6enz171
MODl9KQnTxLOz/agNYdA2JeJVF1XEw3WfRNSdYT6k0vncD18pccMfH0KXal7mvoxZFrYPfLCDcxR
pXWSYGNRPWQKZ/BREAHZQXjr7MeuBw/LQUpGJ2Phv1fyupN/Ph7tR7u6JE3Iqr60DEQTAPfW2LAe
Hf3v0ogjo4WGvtzWB5r8SKeB0OwccQg15G8zrH61J/KN4PmQEl6JHzl9ptLkCE+CSTKT0+jwkqMZ
ppuGAjZOMiBLAjyY3A/yqnQbJMgqok6Kr6wFk0k7SobGhJXHDUBOfVRqcee/0EUuaOsZU0S2mA74
N8LYA8p/cdm78tPOiS3iMM1lwI6YzoujtuytzqylIVeOJOQ5ikPNbb16yBE7hot1rLCTX2U8ASF2
vh07P+95Dn+eae3Moyb0bzFXk+OIEC8pkKDoUpbMNOlam/fzFjJQdg4V+hmkm2geFY0/qZSKiBDe
nC/wcB4bSNE1gAzLkLjTZ9mPl3olbUrmoTxVPTcckHYE0eDR/mgzsIOIwYtoH6zwe6qx5yrTdX1F
3mnYMuT+BKmekj9ZQ4lD3fLk58d+CLCyVN6yyab6ESt18e1hssIUrakk5Ea7QIUw4IbiDON+Zmz1
yR98CNNamJfSsB1X84qfu98C5Emn2rgU3tsV/x0B9uL3PAPJH9ALRvBOI4kSCqACy6QAg6I6lLRo
h2n6xBTNTUNLUBfM0XcvjqN3CI/pCz15Kc8T5tAKRjmWk/rZ/xx76Rwu+OQkkV7FXhqwm04M9lUk
KpQA1kKXn99n+fNzX4R1lpxHS7WOsNnsjNrwPTlC6Z5MWGQchlz88JIPy5wbDbbEwf7a7wIi2uIq
qjRtueMd4bN8GcaWmSX8qS34xyJb/oJF9uQr0dMcU2zaFrS1zOPk/C887wdI1vjSYJN1uMumKaTN
R5DBstDFWeOv3pJ1ObT5MEf28VtPob8OPhQ9I+W6vF7D+EH1aDTC1BNNBuk+CBqlfsP26VCG8SU8
ueVDC6TCbYAf1cmSQJAHlddgiEODrN+cH9J1XrDwhWt2luwjMJpHAuvXwrGLqFQnqe0V39XyvH18
wc+eIzKOblLbkM2/M+OuB3VXaV7XLwheJV4jJTDf8Ji9iiMeEEZumPQfhhDWiOXF5QfEqDBZHC3D
P7DaqOv5VnZhDPBeVzyVhQcb3LfxlXZfP6wsp4auPMR/mNOYs9Ois3GNFuzGu0tgz058Yyb8aajA
UTLxNv2zdNk8gDJOTfA/d+3jx0r9BzYE8O4QYRdZU2AmgJUwFSLJk/rmw/H1jF05EUOHzxNrIoBl
eJhWXJcPifS1Lkd4hLnMmOd2KV6D9R2dk6pVYG1Uwpa0O2lw6Kn55i1XLkAAYdqOg1NB/9SmxUtB
o0kyJVU4RqPnpsBjazyD+VujYC6ql2/4nJxc/hcsLg3e+KvgvRo3QrlVf8plj9CnEcWHyFbzGzXs
Rz/RhuV6S0pLmXTGrsQ2ndWlb+NR3a71YI3DN+6kb+1DyeK2nyg15Mirbq/l+NgFtYUfzKeLXWZ7
4eqx4v9vS/fJxaQShA1h2uRsYliNF0TSiFXradSFxfLR7pPiUO7Lpl8YJgoqnIww0Vi0YR73V5+A
xgvlClmLXrtETDjezR59Vb6U37KgNG1zYWpbWD8mTWCiIxhBVhfTgNMEosGQqigJoeBZ9KFEyrAB
LcNsNhZ+vr3F3wQTEHXxtCHYgMDeAnWD4DnyrYaBCMxyLCeylcYCXAZAVCnJDGYwN4zsGtOKuudp
cthnReLaeJmJmE7/62ze//VuFnRIX1UDTlei9BBBemoajRfvfIR7Ihk9RAwdQ2E88GUw90xkK91s
NiGyjj6nz5rz+xvYsfYeUqKa+z8QQaCt1VH2EmUkVjVlebyqnmiEovSEXm03I94v3LT2zGIjgglt
MGBGjNFl39p8u7h5mnz99fS+UBkOb5ECkvRvXtUuWc/qnya0IltzUt6cIjtx7OjYT4usZnAcrrhp
10obg6wSeIRCt2HzsLpHTc+xdpwIRSHFUHlNewmjZYoq7BC/AVUKnXuphKulP7z7TEB81XY83Z04
HBNZMbD4ZdE+vNxR0rnOqLPWr46ldqMu8Gq2VzP3iWV9IlHxFPFKCo+uGfyS5woeRJpbkB+GDgj0
c5CjaMWwDP/lyq2CaPUO2bpUufl1u/t4hqvuvtL7gIntw0Z7K3U0eGzSMV70r5FjHjdBjT6TXITf
eZCaWMg9sQgWeAQrkjvI9FttLNabjUBCnKGvvBwZcF7MsdTIotVwvSE4fv50X68d/CERDWVu+vs1
3P2uPqCyNbFRodoyZUDTNfi9XC/uXJvkPqgpwNhEAPix254rehpu8nNsEjg53rNyKa8LozKSA0Hw
VboUALzdEONo8WGmpuhsU9UCWyJpWMup31Lk9Rl2UTtUH4Z4XcfUnVRn+VoXc+Rq+fjrM59Sqfi7
z3GoxPGxoGimSEfZel2mo75XTKwnPzDgsXcGt72TzbFZtFahuPbA2B30oQQVlpnqLSPiId8nqINg
f66p5O8QmAtXy39Ma4vLDWz/2UIHMITfu9tqlqPH7+Y9wMdEpzqc87AF+kQsPIofSEgLTmmWzBty
3U75UG5yMIB021UC4pQOfbrs+yxlXGuSI47U8rsfyZwaa+uQNapkD5xWsUibQPgH3PUpf76LMuBO
P08ix3EJkUlV8UuG16JkYg2+W6RerA+QglZmbi3knKUP4hawdC26NBRtp5L/V2Ue8Wj7hHe8/OzO
3BQSI0S84k5jfkELz7mPt03rB9LCXaPz+3s/wpVsfs0fDbbou0WmVDzdiw3e+YRfbmItNXWJGNSQ
nURa2m3NoDGUAJigWV+Drp0jpVBTayX2wW1Xu63AfSle5YJIHnJuMWCrWcEdqsn1zg+NOUMt3VsV
hP88mgPH2kUdnjzHIHQmmvt/SZoU3zV8CnjyTUlS9CLz6V+xqNKJSuI/NNNmxHNYa3kJ0CASlOHU
ZWKlB03myT2osJiHKEvDQhVWKCIrnW9Lkz9FBTiF5dKRF4PKDlclgNEU2hywzmcz/tUZLsxAm4R5
LRJEEZ3TPspM9ggBFjTIVHBX/QSqwD+gehPLZdGmFLUu+Fdwit9XSdq6FTWzVVt89dgad8cqlYRx
WmRE4dr6lQtGsGwWDK8ZOmFfL75nyKCTVxwL0eHmv4q+SghpchRlGligUMgExpIj1XfBPjDvxGl+
pIFgN7V6DmUqzxE5fgP9WuxRjRDTPtEwQvHZNue/CWmsc8IxR72Sqroki78rw7pBW6fJ8t6vXlxm
tGpR454Io3KAD6eJriz/lorVDsu51KQmDULV6bo4GDgGk6RAHW6pMfq2N5gwr4ZTwowTDtAVkV78
xfyFQ7JuNB8aeCtbYIQ2gKHd6S+UZiNtIMk3ZUk177BVSYVdcpW434UVEaiaBPO7cSe4GtC3g1+L
ebQm9U9u6QKb2MvUIFbznalzZ2dQCDJfnBdECn8pbjR+4BoNyxVIyL0OnKA+wRO11bzOzYmldXrG
myNk86k0TMBk0BJOFAKhAI//igY/nVqN4yyyl9XIlPjjCeYakyveHBEbkw+DohVrirTSddT1iCbO
UQHydJ4s8jlAkiCE81BUYcxqOE4sC5mYXnUG684EuJeF+xcFvvT5WLKgIcMtJYJGyH56NRj447Bw
cdRwS+GeUHJLQcAB3gcOJDnkBjyVk9XeXomrvghOtagjHkzvdZHfLssZ2ElXvPrpJexCYVqLwEAn
vUu3SDS1pGlHMIVx60bRyxo2MYQaEE7O4S4wi1slCBwJjxQiGMztxPt1R4EDDY2HB5g2vU0/os3f
oIqzW8el6swrSxbSie+rrLP6BrGKrhdqvYgUmqANPuKZNYgx/x2EXKzB+Bcj6wPgakh/dnbfRSU9
87hjmvSDEC8SR7nPo1ywQYUGO0JD/pbYaGrL/8F/9lwROk9r3FNYesnRg+0zJ98Dmm0Qih+pMCNB
mfUGKVHc8CjUCtMrycqBTjV48LjsFCsB5E+nysEIoYbDdRbqphO7+ElC20ihk1lCfSVrIv5kemjH
fjRZ7AbiC7IbwrwEJ0sukXg6eHi4DT9U8ooslO2jp3oiyRCPeTaoEQukSnKz471SY6rMoCjs2ro/
2iKRqpI/+DAUoqUE1L20vkJhCQW//UprPVaow8OTxffdZjNZZ/vcS5brZzahnLhwerKebWbuXRZ4
XXHv7dSF+ADc9eg0qMwQiVtRxXf+dvwuamwmYPLlGEbmM+ViZeM03vL/t0JmEAqpOqvypdio+3v7
GWBeUJYuXs/BiehGvT3TYapGqg5BKWvr96LcZKa69LnnA0gv/8V6vJwdic7+xYl7yHQpKAxlZQEo
EXz4tdPScw2WfUniiqww86x2zu0qKow+oGgZM8tZDJfd9NIvWERBjAzRDelkFxSwnegcQNo2t7n8
IdfXb2WdDoFpASQpM7w0/z7Kts/Ier/CAYxNxKEuBH2RJ5BKL8qjUwReLF7+jXHGAX3y3GANqlfp
NKIKNoFFBOff+HLP4BMIGi0DEcjz1etoNGrzRtoeDnAkxjFK3tKM5xS2V4NzELHAyNDzFY9KCkay
RpK+bmakurBF5ZwDR+NlAtzJxliiE4nliF++v7EkNg7xqq8363Eojn6ukxXz5NpyryU2RpF2acsg
nWoj427d5NPNiVOdmxZlXou/Yipf6zo0+w5cjAfm9lPUyDdUDyhLDOtJHd9tf8p08gsCcArl0Z4h
DrOdjjIo7DrnfDJfCdYnDooQg7rWh0uS1PDSjpf9vQGYLbWsUByCOSNnPRtviy3u+1PuxEpaDRk7
TnsM5ucjgVion/AYefRaOSoc9+C64ZQeFiCcBqom5frd1uwYrDtMSBFLRGfb7dnVeSi3SKq588gu
3rl9g4zj/olc2MWjKH7c+IFk2u3yvDPyfqP5YdtPCi6oOzWwK/m7k268kG5Ks79CA6l7cLBLzz9J
vWA/kIk7KOvbX3TvOn3ZyDST+Pn1CqFChkV/sVmmsKgjs5vMAS2GUFx03KtlLNFb7oyQ4woGhvQn
J91ibl9VrPicsJlIsQb5OYADdjyrj6c0rRnJLbYxEAKTiixwxg5k5ToLKHty6IK3IraJzb96mLl5
xrjjO56wPJSzUZTW0nNzU7Y+9OmE5quYU2bF3L22IwxKRSUmsDxkcCm9qT/kFTeZ3lmithzmEPrX
WLK36bRQX+D5jOhXJjcHFkt2VtySVvCXMql8uoWS8WDTh+eN17CFCkZu00fb6w2pEKcvjx0vXOuT
XnJjVeKOfSAhfo/X/06ZYfbU3DkiGVLmoNoK/3HqfUcXGI2b4X3LM74Rzm+OUnsIDYF+RoEEd3mF
eJfmn7pJ6rG76k4KApgGbnO7G4Wn7G97QzRAdZi9NveFs/a4v/IGzjVICLWhUQxkZlE6QevfTI2w
J9ZgSgzTwNzen63D3QmgSaItCE75xq+XWUgCraH/Aev/+03TyZTuRJrCSjRfvuCTbdFyjPnyUXsL
1rUNeAeb4aJRtitCa8YfKAQYZ9FQutWAddmqAqtIQPqL8/r1tkW2x5V2+U7Xo/LplOU2d28RU9Mf
K8WdFsbJ1KjCv3y1bQ1VW1PBIN+nkK2uHFT6hskCHbC+OqtF13aHI6mTVzkMJfvDQkmFyjKfQjkI
b9aoKoktYCV6NgQk08mIqm1nZH3DoF51v9TJXoNhe9j+4O4uJxpZEYFuVeyaZqKrCIGAYMRMQLQJ
IPdn/iEdOhJW1kU/fiXRkDxaWmDzE5pEaoPWyhT6vjt+gQg2MDlPJuuYBg2a24GeuCS2ZV8jW5pb
jrsTzUAWhpjTPNAOnjLKdJFfdq80my/WWjqUNkFWve7XD8wrFSWaZmqUYUrMq1OycuJSKpFVekFq
QvXiH0p+2GaK3n57EY6e51iIFu19nd7/0T0+6pvYPbu2+xMqPOF21rmxX0L6gaApJu5mgebnNZYk
3N1J/BXQPZwW0c92fgAz74H75dmxzq02TZHhZntDN7nd6YUROosEo4d4GJwhd4VxVP/7bCKIdrhG
e5vpbXfG8TE3jmmxH8KlfrenkuJ1FsU7046NqUBpX5VLGIEbz0/2FHjq3+fyPZTxG5+EZwiP+ZY9
Mi++j4AoKQjbC/+y+wcK9XpTKonGVltRMxPcadKu0kfxGijWWuIayS2P2B1edfHtwcT3pUYqnpUA
Qny27yhLFFa8bS5er67JbqxnAg7EhxsGWeHARFwecr6xl+mVRpoj76GcUQ728458bqQkL6pvbvDf
60w2oGcmWcN+u7aOo7RvcZ2OzcMJ+2amV/E1UuuMTFJJ7Tqrn2g7EnTSWJFhOxlV/+Rciv/XvdLB
ZidpfVLUJQQ3sjSDby6UZ32Y6meAQrzI+WfUqiKYerD2XmHqUnZ0QXQZZRIkMbZND91bkDcG9xYo
H6jPNjw2/nl51oQdIi97KFjvFPyar7buwgsVM8zOhefWXc1TULPg82lsqCqXMjzhWqdr6c1Asxmv
3lN1cMSO2zcnpisSV0cztP33doz9aUiW0CA8nwe3bJppDBVQkuoZUWPktkq40dOR8vwGAdlizovg
/AKEDFW0WLj5lLTBLBhCYfnL5K87yEzHdXLYJ1zlFcdR37fzeAU293LSs/GV7mxSPD9jJsHRWF6I
X+LEU2yk/2cl+Xe/fqSI1vp2oLzj6amOrYpKihZ3Su3SfYNnlDGZvy0yq1FTtf6adctBA/INkBa+
4vXd44paebkGQIdrMN7W2+R0WiPjwQUW3xaKfJckfFbnrlat1JiLiWJYjsg0LWdfZWBaJrXDwM57
O5ZcjSP5P23zySQ0oIxCZ6Wtw+PLDUlMTBzE4xI1JquA/WYNSfhOGxkqmJrqOhUQ6ReLfyUTlUqU
ZzrELwM4H3ncZgfWboLSVuBK8T7dSJBB6+v7fdg0FYid39EPEszZaokW1OjGObpiRhqZKFiQdUsu
rrBFS7xVxDdWoS+qc/4EdLESUVFcPIFqM1Uqj0Fzr+cWARIpIWZuHW63y/wR9c9BmBG0fmNg4eWf
UtWx5cEX5aTrdCDgofhYNZgC6QPaJMdEXIyKFnRFK5QiI8aCPlWj4sJLloNvFd7wopHqG5rG9+nC
w6/aaNsr8XCEz/a7AwPDvbjyOgb+iQUnRuXf4N7yTjEqaOQUgElFYY2x6N0peJgmtSCMdzMI6Kn5
AOqB60o/0XmeGY/7916MiSKv086W1IdW1yJTHErSb5qK35BdkO0rbCUhv0KhdPPpxFw04Pq7a6aU
cezvsceWDMX2qiVDK4UaUZxBHHvCy6zP7vSx2mnnz/22TrT8wBvbhfIgZ+0ON39373YyiVJapYqh
tvHAbqrEtstpO3XZopSDzW97G1LSYeviPx+o5gCx3NWmBVCLBknZo8wJDl/2U4s3ZmV7xPvy2AFm
XwiluXb7OfjIC61hzeAgkzuxf5flwyuYAfz7m5EPfMJQ9+hKgiCwdP5oRCVoVeTcsnJqG3AXn2bT
u+4QuojW4HvBsRU+XmJE0GEAP+pIsm/qVM+BQVFotB3qmunYjieub0PZLx41AIr78eU4GGRfNOi/
VrpgMcerb7iktEGuBzgxZe/OKbPg56Nwk7w7wHwYFA6o9C5Yww0pDW5wlIcX2K6aPoiCIHiv5w3L
/BxM9WGanr0K3eZfsGB9XO3iWMBCj/pCa3vc/bAVK7LQNLYR81rgJ2DnrOuE24mhbLHTAZf7f8hf
qN5CzrixlEk/CBv1DXLBQvKq1QQmO/sSZQtV+jbbUCpEo7wVOvVQYMlMSscRXMzkW8Tv3gdwo9Mh
jJfssBziDmYDFO6F/NgYXpRUHliWlL1ClsKZHIk8wwIJ8NlZj7lF04abFSa8SxP0ob5kH5oAoa15
+D5LvpapkFR7dbgCR9U2q9nyne3hx+YgMm47+FAfl4+hp3Z7f57tbW7IUj41SUwEdOufwqwRgHO3
97wk8z+7TAsSPFRgr4qPSYAv0WHL6EZZ9WBCouz7acU7FkYMfiKyKYPiAhkKWbNeCdOlhFpaiC53
GfPWSDUrqJXv3dW/y2uEnpDknPmLS9my3E18zieh1pcH8J0d0nUe4mbgO9YvCrYNKRAZS43M+a4y
Ykdk7UGWZ/emn/oqdUehsDGtDF7NDxFZbcsa5agOCOyyPDGn9yvj49fd3aElLz3VYPHFh5y41rn2
iTjZPSQ4XdZT6aBSz7AuUf5zkPsH3vI4guczFdI69C2fnCSQknBVcDiuRHekUUW+XYHNTgIXXqui
NSyxSzk9LoTtfuLCxpf6NfnaI4dzw4dq1khcg1kBmQaIcu0aH9ugxyEQ/LYKiWPqb8t0jHpl5VwG
j8Se701nzq31VSssas72IdEQUOcOeKkEdmem55zprxL+EZU5hUEtVWhTHljzqSdv0/vItHIpj+DO
Vhi+pLfl92Q+SysY05mllRHiGaZj26CLnakhU+s2xh9EWwifh4ebHfXcRvaaZULkcTYd/Q3+FFzn
O4WiOAphxwvmfmaWfO0BZKP+ZR4NayWbWmYssFVfRcAKqEXGomFnkXllVHUb5X20FaJP2bDRYFQK
adfWYtK3ElpKul/JGvtq7mEkWijyrNVPqX75RNKumUKz0VOTlGgVuz8C8vk2n4d1ajnaK+uPlg==
`pragma protect end_protected
