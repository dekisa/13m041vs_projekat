��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�@�w�4s%�mH䖹��F��Զ��~����Te���@��m���i��VP���_:��	H'��hjgm��\��E��52s�!��%&B
^�q(���|����X��5J���F�tصU�ǣ=!�-������TXXo)w���DF����~xv��vF!pB3�>�6^娖B������BO����<z�g�	��ܤ́A��P��E��E�"�V;�%W�֑}܀F�����xx�� ���}j:A,��k���!{T��J`'		-�)ˡ,��<\�,�d�_J��#�#)�Ҿ��18��ɑ�NS�5����^�p�!����7[�R�����)x X�LN^'/$�9l��]�!Wa�}�8d'ٍ���I�N������ȏ8���~M�Ŋ+"BZ��kd����~�w�P߀Լ7�"�3&&;��9uz}��N&��y�,�5_��}�8Z�Y�a�9Ru.�+�~�62Q��XV�{}6$��ؠN��s)G 7C��x�Z��+�z��zD	>n.��뤫��٥�ؓ/1"C�i)�~~<�3i3a�Xw
�	�-���[QS��j��#�b��ar�Om��U ɭ����S2]k���nm���(�r����cN{�v2���[E��6]K���4��$uչ*�"W�R���~�b����L��Z"�=�i��d�L����ni�-u�:�bG0XU��=�r\n�	
��.�+/VFT��r�R�w������w�l�R7�(N闯�bBwk�]`w.�����V�$�ݎ�F�{i�N�:Y��H��v�����q8r��x|r>2(V#�\�kY���?u��؟��Ս��8��^��0���E�~��Q`,�1|��"
�!.As��\ty7n�wW�j��0�eIV;��i	a��7�M/���S���?EC�?�vf+W�|c�BM<L���=i�Rt���<�A�J�y�`��3�%��┴RG6�Y���&���'�&��ь�]L*�3A3wj
ؿ�?Q�g&.J��%�-�����@ �k��m(O��6M���2޺��f�Ml4�oպ0 U�h8�������R9#�C����a�@�����Y�7�%QK�C���/�
�3`�����B/�����#�jy�:��%��XKW�uwn��g枘`��%�ؔ	�J��%g��#�!�.rҐnq�1o�y�Z@ �*9ߟ,�dϩd3}��H���-yr�43��A�wC��$�Tz%⌞���g��b�L�&���Sa�F9��Tr\���=S��z1$,��r�&D�,� ���!!
���5�KE� �&.ozV�k5J\��-"�Nj�@lސ�.���L!��=�+u��O0�yBq"�*/�.�'����vE	�}$~���l�����D��C�^�ϝ�**��T���/��?�}!�bm��{���-���b�(�Ӗjq"���4�0�z^N���;�+k&$�h�+�B+%��I���`X��_,��(!��p�V�QW�s�9���)u/�vf(9���	A14�U�	À�Ԛ���?�fs�ߨ�1�Q%-x� Uۨڠ@u��qoh�}/��y�%�W�ڂ4}�wZ�;ٝj����3g3�r���y^��#r���Hr�����b�1�hy�"��$#&�y`�<���K#P��Я�kja�1�^+샼�И���*bN���	m�+~-�������ET��Rnf��傉�-��}�9ӳ�����UTU]o��%�=�7�y�q�q��07a�'������
���������!��Sr3Gl/H(Z$N���2oǎ܉���V��g�� ��H��W�"'��=�c��yn�\��%غ3��\I�tƞ����ؖ~5�F�Y��Y�#�d\k��X�n6}`DO�1��h\y.v<���<��L���7����SA9���� ��?��z(���yS�Rq�Ή���;�YZޜQ��Z��y�=::�xt��f(%dN��q�xF[d�I���@M�/���{��hu2�/���+�6���yM��ر\>B���ٰoѧ�?��H�1�+�p$D����Z�]zӴ�Xk��@�qL���g+O9�La��r]M�|0��x}�tʞ���A�0��F�sA����%��*/���E4�և�1Z�'��-g���i�ˮXW��pm���`��c�M���i45�f3���q��j��S���@#c�	[����w�����������sɻ�J�qPG�������^�<�$��Qp}�_y�~vL����iĈoZPbJ���M��o#���o
�ٖ��������G�o�L�������y^|��q'�������]c�E؁.I]r��q�ϝq7���Gܹ
I�r� �8���]�փ�=������;���*=Tr*�]s���SK V�(�$���c��Ll%i܏O��R�N����������m7��}sm�ٷ�6�����p�Hp�^�b�$������t'ۯ��ӓ�7�ۨϺE����;>X���]�P��d�$�MY|2�(���C��8�C3	_��L�v�K�Y�$k�n��?ٶn�E2��DR*5�b�3��:oZ43g�ѽ�14NH�o����1���qc��1[p��\��ؗ��y)GU�Lz�����@�MW~֑=q��2449���63�H��dL��Xʒ	��/KYA�'�"���X�Y}�8V�:v����s�|�b��15"��
�R���xuAr�Hx'$��/*>R
������}��}����Ɔj��2�/�B��,٩"t-tQ7ͳ�ܻ-$���#���=���/���K%�&��u���8�eJW�v�=�]��K��nw"����|ex�!�$H(%�s�휇 �ۮ���/���yE ��K���lc�����"���*ӺL�������{��[@��)\ۜ�s��/����u��y��£��B�݆;���`�谊��b4����ZS�=}��h�IS���m�S߹ʭ�Aȝm�<φt�GM�A*�Bq��g����j��I�;�;R��o�4�T��b[�"~�$�1p�	e�v�.a�X0Q�~��{b7_�<ۑ+�.O)3=T6�7Γ��vp���@?��-jn�����֦���h}᱄b	����N�C�ZqҌ��G�Kw潺�-%��Hg-Ub���}�os��� j�u����VJf0�&���{��W��pz>�k$�KcT	����g��܍�+�q���)���Zm8��� 9��g|?��ѻ�B�)a����D��ز�5p�kJp���l�6���:lXy4:��p���Fs]���3�n�PS1��']BY�˂?���F<5&���L�D���������{�c~�ʫ.x�AC��Y6�Q��crK��o���k���g�D�&t��ٯs�] �����(4��+/-��(?�"�H��Θ�/�6�=�,��8xyg6�@��N�f���4�>�1�B�Et�e=���V�9��O�4����pG�ndZ�1�߄�;�#C+8K����Lv���h�-&ԧ���"}݌y��e!VPHCM1� +����Fμ*�Uॹ����c!'�k�h�YUA&��B�<�Qf
�����s|��͌C]3�yC�Q�	�����O�UM�^aʱ߭dp!��?�乢=�U�lEa���*�@B�6�;���񄹹FK�t-�sv%�W<}�m��þvqyZ	�\}�qX@�v�������[�3�;���o�E�c���D�`͝��n�uf&������beG��ic��r0E��Jw���:g\�M���G@���s�ù�t`#X���Z�ۙ1��#��p/�ۋ,�u&n)�d�l}�H�Ѻ�<����XG��K���F�ǃM����r��G������ �Jl@��2p��l?��l��{�M��� �	�6L+j�kb��S�[(�[�&w33�����m���jXZ���;}�<�PK��V)"n����[9��8�$��VY��kp�'�,�2JA%Ρ?�h���E�7N�c�e��ϙ>�i�#�T����p�m�F��ߔ�a�Ս�2ҏzO<��&'���Jk��B����}�;a}�6�z��Jg�
�>���h�O�0���:�-P�q{.�[�	�g!f�!�ዖ4n��?A����}�I��J������\�����Z�v���h��$�����W��]��z���5&.��|���
V��� ��¢{Y�޺p���}�+�Ŗ>�f�o� 
A��JX�,�4�N���Ӳ�;?R��8d��X���B71Xn%e�0c��$���S#�L��W�uy�*�XTٝ�1��!����̅:�u��9D�O�����V@��u��GR)��x��v^fqu�4�zǞ7;���ˎJ_O0i�}���fd�������?}[W}-�Qw���|��&I����(E�ˀ)f�����3~�W�kqK$hQ
��"����X�.��|c,��y?Qz�׺���o�8yG�����YS5�ݍq�JM�c�~�T��~�h��\�B���׾��c�٬�S���խ ��A�-W"{\n �^&B��I�rT�@nBM�2@�#���7��U���!h��z*}�fT��K����ໞ��k$^��x�xs�2Jԃ��-���	y~��F�Cl�?C5���zj�܋K��Q~�C�FڵN|�� �~�]u	u�4xg�>��K�'�:������a��,e�m2�lwV�=�ya����x����澲�f���s�-d`�j&!<f�����zN����P��)�Q�����o���������	�o�s�f$,��$YO�>j�bk���Lhh�h����ʳ�{PL�%���l
�txU�3�/����չ���p6�Q\	�wSl3�����+y�K���~�&�?�L�^�*є�L2+	I�!�`��k�h^N�5v=j��pdk,&���.��������W��:'+�TI����2�H�J`n;_U�;�P7UPv:BY)�J�+����*9��sy8�	��m���hV�jO$�:�/R�d���^����:z�ø�=��Mc�4� M\�z�5D�
��W��}��
@�x�FƓ���w�p�,
��F`�m�.iy�>�6����`N8p2WLMW{��c�v �r^;������O@|��(�dK"��qj?�J��sd���Lt�,7OV�Wr��ˑ��l��@'�q%��b
�7�n}�1տ���7HjD�5f5�� cV~8i	9����J�?�:�PrT�����$j�jHb��--�n�Q8ɮ����M�ҧ�$R��ke'���ȼ�C?1�~n�3�5ݔ�йX�Z7�)mp�� X�9���9[���KV���>(��J:�Ҧ�wJ��c�1��p�Csv��.����/����V���W�-~zG��Bk/O���bH�<x�'�fP�a�ZX��&y(=Տ�z�T̶����<���X0��N��N �l�W�;0	?��KO2��ь�օ�>�d$�"����!�s�����,/Ok�j�Wՙ���xD�ss�y���(�qH��ٳU�r���[P��6���ˍJ$��L�.�;2���IZ�
��(��x�ϲ|��BCYeu��`(����F+�~`�F_ku0��8pU&�Ϟ�!$� ���D�`|~�-��ׄ�R��B��-�v�x�9!�ef�i`�V,�'�#�c�E��:�D�f�nXj�e���\�%mk6��7����f��F<U�k�j�-f�N�1�#Z2�Fj�e��>�#a�S��:il�Z�E$���验X�ɹ!{�vFD5�}/�>ض ��Zn���Z���3�[݋!z7o�4�5,�5�?�_��t�䘁U�♬lz�ҡ%�K�"$���&��oUdC���h��p�a�̍��� Nl�ʇ�:`�)?�1L�S�����%t�`1����'�};J��k����j�/�!)����}�������k��Yj,m���h�h�^��'4�O̩M@?[fE�Up���ΦB9's��'���^�ev�K���d�Cs�|D�N:�@�C|�i5cQ=S!��n~�|Q�H�/��8�jT��44�%Aݣ۳��UQ���m�'��ڈm�s��d��Չ�s�Cd>$?1:2GDq�b�ߕ�����=���P~*���i�qJ0����ZfU�.<��/s5t1$��C�Z�ݫ;�s�=WM�S��^��KsX�z�ղo1��'����{g�m�tͤ���&Owz�1�`�`ҵh≤�~��2=0#��~��n� =�����^�	8���e��$uMo�%P��"^�R�TW���%��������̆s�q^���ϳJ���6$ε���n�S��W�(�#E��'@L.��߼V�T���M'=�;��htr��`yo�{6ӺᰏCtؑ?�j�Kj�P,L��O��x��/����� ���"C#��[�Ї!dp�x�w��V��Z���(����bsT��̾pM�!�eH��bn���8��]5��r��.ģ�$Ne�Y`F�"f����M���\+Z�4Iծ�cP�c��n�I��4�/��X����iR|A��j5���'�L@�r��N�=ńv/��L�����������~�6�>#��^�y�u���6�oG�����P�q��J`�cR:��{�B/��pg��&�O�~S����f�&2�~-ͺ�ty�Ծ�ݟ����m��:; ���<�?R������s�����1��ן�� Ce�CH�S���~�{�W�&��({V"�M(�I�8&hb-Z��?�54_�X�c��l��M�*������ٔց��X"ɐ,�����fΦ�1�l7Zw<Ab��bdڽ0]���m���������F<�@A��"��]2��G��{e�+qL� �E����i�J*~�4Ƚ�㺟�ɴ�C��|P-)���)��>,|9#|�Q�e��P}d`d��$���dmƅM��E��T:�������yhONT�w5�DwP�Oē\&��ɛ����	�uo�;n�ܖ;f�q��W�.^�����7�!�R�^$b_�����9�*�>9>�̿��_�*8W���8b!ñ��2��p��yI?�x�	�����j��RM�J���H��{���I�AY�	B��v#����v|�v�A�wڏ�3k"�����&�@�.��? ��H=��&��D������B��h�&n��q�!S�ǧim�+Y�3���TԴq���h�i_|�rq����*:S?8��t�^���&��>%؇�闬/�j�sw��z
\+W�J1_G:N��#K��Z���"�^;f���3z(N�˞W�*5�x�y�F�{��Q���g3�O����/���ӑ�n)?��=�1�bʏ���hsq����s��mo�5J�}b��~2KY�J�!B�s�ne���8�@B�q��c����:����`�`�=VョЮ�J��\R;b�2�3,�q�6��^R�`���v ��Q����+�C|W���az�K�b_��0LЕ&����<q����0����Dt�H��`��~t}$)�]\2�K�ڦOh~:zQ���p�͍:�.�lsU'O6]�F%*<,D�i���*o+Ek@��cMi��b�ex��Ԫ�u�J����<�d,�S�>�}@�n@nW���- ��?A	���@���r6��Z�!U�Hz��!����혹�!���b�ǰ�Ҝj�O�n��{㫶�KF�y��e9 #��Թ+��^����ܷ�X�����
�+a`���Ф�p?_���W�XG���?C�d)L������!��{�ݹ#KOy���Ah��S��1lAg�6�p�7ɜ���f�跷L{Җ�2����6"v87@x����0��8~��1����0s���qd�-+��5��4�I��I)��'�⨐�:#�w[�h��.�j�Rb�%�~�����g��Ղ	���ϐ���9TXHw?�GƯ!7����bk���'�@���J�+�5i��Ζձ\��}�օ�!�S4X��Vʄ c�w��eNS�,>o�@yFK,�R��$�I|S���"8�����;8`���Ud���ѻ#.�,#!A0E��JƇ���sy�Hn��5@��ʼ/%�Σ��V��d3�OR�<�QA���F�]����?�^�#E̶EvC�Nh3��rs ����-yxd�=P��y\,#���z���75G���4x�Zl�+�tK��/��S��7���a<>��O�EH�>�s8=;���ԯ`p/KY�'n���t��!�|\��+��w�n���r��j��%(�u��s������a�*K[^R=	xp�xJ;�z$�x�i˗��n�	��L}
<"�]�b��W �Y���n�M�Ĭ�E��bm�7�"I?�I>�z�!���'%�4�'�cdz����<9FӬ�k{QS[��(�Z���y�%Q����%�����,;]�21$(��Y��
�Q�/`��(p5��+�>g�CHT�w&1ad7��9��L��}�dwԃ=C��-yEy2$��P���~��L��mվ6�9ȸZ,X�v�B7��㏜Oyْ��v�o�����?[�k�M���l�\����vEٿ���{��C[����|���9xv�Q���������ƻ���G�捠|�-�$�kN|�{�A��׬K
?���ޗ�U��vY��X�ˋG�=IZf�u�e�5�����ҺE}'�`�F�K�N�@�>a�/XO�6��t��v\����7W��`�r�c����Z7Wsf�b��#|��_|�c� b}>��el��R�E~%�l�d��H������,x��Q�7��{>FSL#���*KBƋ�D�&U�t�w{4���~Dl�v� �yd)�@'����#�˪AhYM�*B�J��}04^��0l�,�����j���_{9���;����ع���W?�� �SX�~␼��%Y�rycqptt}E|���oBt���h:O�%(u�ac�{���_��=��
�)��U�~	"}��.�ѬW5�+���"8��8��C0��3��	@��-W����gi����6�"w���H�ݱ'�Ia�`O:.}�/������H@W�5Z�Dm#����զ' \بr�����i<}ϡ?�*��|�l�X�c5g��K�\U Ki�	O5,�n\A`a�%L��lJq�jQ���Pxɉ�Ϥ����]�.8�s,�u����x|�b���V	GQ��2Ɏ�OL��ڍ�E�/�D7� �ۉM=�	�kQ�u]}^p�Gp����x(�mw*�D3q��H	w��7�gwd��	?��p�K�!�B�ķx�d�uz�����*�e��]��Jb�Brl�� �N���V�&k1�	6��d���Tg��h�b��!t�T2�΢/)��?Si�Q)��<�
��ۆy���n7K�j}�xZ��?�����n�,P����H�\������@=��:@�pzYh��!����6�?����6߿*E�g��26v|�ܧ�E�E��B��q���R������q(|V�����8�"����)a[�U���//w�]GX���b`Y�hAl�?�F.�960�����&-��*+�_lr]!5��)��i�2�����+�����Ǉ�3��E�K8�c*1*���nY���������O��6��Ӏ�;����帇���q�����-�t�h�c�X+��<��� u���(Id�o�9cy��|�-��eQ�����*�Z
���Dp�~z(>F��r(FyI�(���oh�¦v�C����tO-[�G��_@rbc��y�v})��n��$u���TFt4�W��&�g<Gs���#���Q�oO?����&��Q<8�񱦫����N�W��O>�#N�=��(��@2sUR!��/q�3I�0y��7�bz��
�S�pQo�O��,��n�e\g���Ca�!0(Sh�Z�ԭM��%���_�i�_C}��:����Y��K���T�۩)���(�f
�M�݃��'�{<��}$5R"@q�s��6g��X��[���}T��[C�T��ֱ�k���ُ$�|�΍����5a;����{%���N(ޗ����&D'V*�x��#�E��$e�B3�n�Wc�1�;qo{�Ѐ�nGv{�?�DΕ+� �:�j1c�F���'+b	#��Q�4��B|4cX (��@n��f�������%�� K{f��<���p���ll(������>�^�~i��7�K�n�!!�7-(Al����!��Y�D����+%S��e�@(�U�A���|��d
��Q�`}�b�'�^fpi�xsw�.�#M��{�ah����a��IG�ٽ�-���n.Sb���_�4�X����~�1�-����txd���=�>WmFq��(��z�����H����I>5\���U Y*=��68�t�z�;��εۂﭠ�8[�Q90�~��C=��G��oxVzM�7#4��B�e�nT��	J���+T��ӌ�ύR��t�)*3m&cvǓ����&._��O��ɼ�qV)�!���[C8s<)�<D�,-���{�=�'2	AR,S_�h�'�Vb���~ﴪD>�D 2o�j;]��C��/�)�~�YW�|L|��A��'"���PA�M�PVFp؈�u�!5�= �Y�CtҵE�yr� ��V�V�t�K�T�}L9(H�g-�%G�w�~�&����L��eI
>�-����_4�]�F�w����#i�Pn�(+���f�Go�+H�)ѓ����l82/��?�1�-W�&֥~{��BI�L��})	���3|���o��v
������,��Q����;��̝'q'\�B�V��L��	A�2�l�ezf�Ox�4����M??�<��Xp�6�5d���㋹��>�K��ܮ^��-}h��C6��޲Ǩ��G4zfUwX�Z\}�}����h+iǤ1��!���x�8Wgc4wH�"(�l�.D���)~ �������c�U-V�I��2r(Mڳ�8],ûH��V��a�eY��q���v��Ž�G����i��M��O��� �/f�����D�ﭾ�IX%���;�%��oV%��3an�'�r�lO�� �TL�%"�M�]��
���L9����R�.v���[U.��/R��+�s�}�.���8�E9���ni�F2e�зѺ�F(�ṷ�J|w�kKOEUG˶#��rl'Ea�ly �X	aH� ���œ%���M1)ܼ@�E@�2�֥W�,5k�V�!X)!<�b&�����V�
*>��e��H�2��x�����L�����/5b��XS�0��tv(�1�I�S�){9&�a���m���:el7Uʮ]�91S1*�������O!��������[F������F@�W8��0�"]5��q���|H޾fY�0�[Cec��b�THi�է�O���޾I�� ���`��k����P��;�|�@�~�Ϥ�cs���L(��'����Al�-���#(TR��M�ǅ/]+���l��@=�F�^��3 PEu��x�D�o��ݽ������� ������d�Oէo�}��Yűd���4q6�