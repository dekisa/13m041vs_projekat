// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
evGBov2uC2OJOABlJMxGAG5mvouhpS0KaMEydI5EomHsOxvo49dtOBbSR+GL36bJ
JPcLG0TZZU5ovmQJQSdV6gTXcVIKFTPhHwPKGY0wWbByGC8P67Ed/sRy8uyuvjNX
YV9QsV0kurOtplOwmjv8zgA7E9vPsMXXLsSUAUDqWs0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11952)
7A33ANOAKLQ5XGxbDNcA2Q+n8TcgjYhkjUUXtzspR9KXzRWtK5rLhviyz+gqN8Yo
0dB/zxChetwxe2MpMnANn5NDV5uObuCDm7ZJlGwn2YDCb8BrwSevGLi4FYbpdDlE
sc7gfQ+Dv9qhph4s7sHpdNQ6cJ8NvF02djDnDOd+A81DIzMaRwoP14D0fmlYBu24
4YrylsECPq7w3YTCZpbi+2lmKsGhgJm4PA6AKSFkT+STSWQVxDkdJMphEWElBrPU
6a29K67bnIixCACd/9zCJok1nyRCrzDcFbnacXkHn5Cv8MQXVssVzJZ4Q2WMmFnZ
26PFJ2jdO2GDHlkdCCApw1ucm/jlsqfVCDuOuxb3CVRSK7m+5pjZ3NlqOET6UQeW
7bw+ztS/YjtJuGF9oNfjFc+LjPYBintqAWYNzNaeMw85wBo/ChU9bZoh4fg0ycl9
et73TFrXapd8xDQ5PCt0gaMUWp+ZjyeD16Y90b+y/1FZ1TgWEUduR7gFTlTKlTI1
VzIHLbJ4dhkZm/DZ5057rBTJZ2heTqWgxcpy69ZF0EvXkRaOVVKgJ+fcsdMy94WD
+PqLTNPqEMRurubdXSGvyQNwKNCAG3ayvAV9tSU+MJtUP6Lnjv2hhYZB/eK/47nW
w7SFW7IINh4MjYsCRde0T/axpCD/s5YudrihSEBphFL7gtE2qOU66IxlZN+Y7KZJ
NEZQ383wNrGnULK4ATy3DKSXDNmkQ5eFDPyMyRZb4Epl//GDj0vCVMOQwgwTRd5R
PQ0zf1zZYtKiWDyE/cWG0mDFd5XHI8jveVa1AUjUOurEbYK14PxKHflocI7AHYrY
G1XyT8RYU3Z4UGEPdauGQ7+0mvd+QK0fPJij4lsIZW28G6LMMcbWP3YNb5f/lfbX
D6iZqJiZ4TjDm3nPEA1pQ87y08HH1ZnVEfGrLJvOq08afR2u4Kh3EBz145n3YXX8
FknTz6XhbY9d8sage0ABsopCPkOhebYNDtQWMz85IOEiK1QQnyJbMCtON1nZGAWO
ZWHsyDe233bxDoInlulOeDzB7F8Gwga/PMM+EfmGkF2KNDt8PIRNeZzarRG9ECfF
3uWHy+GKe0doqhM0Ug9KRnMPX54xa5n2Hyg913KskT5ZznkGIRV0+cBMEU6FOgWW
/2niIsGuguiyjYf/Qs3y3aLNgFeJVpCFJZOGTfziT7qNZYMoGyO5UCz6NnmNfZgH
Y9+v9U0PrNHAkHWWW1qVC8EO3YOnzfrUVc9RW7f1Q2Ww0se1ZH6VCJ1Gg8t8Dxf7
nC0stqkKKLpin0x2tRE026re7pvd38iEBbM7rX/gdqRnyVnb7DLAcGaip53Di0er
eFTDpoZWcoqCaX2TilikvGr+W5qZSZIRvOkto9GtR10dO/3Q6aSM9ouhlBYX1/ie
WqgkGDNIFyRa+NImThopNPCEE4fmBDfxYF40NP2LhsmH4grI0XqB+Spi6VXgieXo
oAqc7k9qVslzQlmNm2aOK4ss8et6MwpthTi6QcGN/zOKYGDqMxEMXwVXCibfknCg
kz4M2ZHPNlaKO+8/dLru+O8cNQ6I3kCetgOkuNov8k6YOAFT9Q/Yeae+QFX78lTP
9QNyNUUfAsfJJ1DBWX3L1vLHfpVech0u3pSTTDSv9WmDeSUrakFIqI9muAaqgs53
kK1lwlGuMheFshcMm0xVt+tXLlX7E0sknAcwAGqRWGVCvoHkJez9asNid19/Mv8u
9u85tgAvOuGSitW9OnmoWGj7iRVkdqmOzPmw4gM3RwoDoW1xh6KcgK7N2OC8/Pz+
MxKBWqT5bSLlJsY4ZMSd8KCfoVH8iM4nKpjIKtSH/VBRW1QdD6nrvT3ZAOSTmwKW
jq/oBWUDYSgyV7ZmJdwu4o/sG7JBaMTHc2bV0ixNmoz8v0PD/LRf8bUK8+3+uuox
zn/zf3zizU6cDNqRGYz1aCs2RLH2f+EYI+WLVsI/Zc3uRaS3Qfi3PumqAM2fwT4T
apBiw7zuW0gP+mhwfbGQAYBe/6utxVu3WPmvPXsvPAtEzxCQzDQUgMwXYaSq6L+/
RlmTmk5MB7hjcpvjQTNUXAcakInTQ9L7RIx1AaXpCq6l8GsILJ8FuS4EBqWGtBPL
wR4HUXkUIque185y3pf1PEs3INIZalPDRBvAVAnQ0vmxNKIAqdwVrZGqSG9SUn2O
XFiqV9ElR1GN2MwS0xgCLNiS2LfDOc/LwaiCLqjvVwdGm1RP2IudzenzaywyDDHD
s8t5AbKt3243upD43a3IniVxs3HUFc16Xg4PMhzbqKD5tQ4YjWNC61t0bRR3RMHn
e0wpUVybQcEC/tHlRp/A9H7UCD6TxIx9d6yxdYliDC/JLqh0Pi9FCG69fDjuOkIl
NQa9u1gsm723LwK0zYcnK5hRicH2PHxkj8p6NdguoGEEBKHg2cVs+GmaTZIf26Um
BFcrvcFyN6KSvssgVkJgxQPFiNa0ku4o8yVWE/Xd+vNnD0IfPvx8b5rDwXQ0rGGU
Nzms+NwmZGTAuakeqKETFxM03UKcgwTSY4lt4xCM03r7m/PvKcb8HwKFSR/g2P4J
qCOwKCZRJYNKxhXYOqaiY3RPH9PgMYWvigLbf5EnqdJQDOU0uEZQl4jdeKsVjNiC
lR2VGItes6EuSY3TcPNrMUzLmVwITT3ESs678Nwwn1yB0QfQkPEp8EqNS/lqExvU
HhhFIU1SI5vVEpUa6xayPKWP4nmcXQ44UgF2jzHDDgvfrvqy93gnQLygfwnkDoVK
BnnD4XWnisXSSc2Sq5/LmhsIPhk9Dt2/Ru944Oc42jsifDBuO5WxRRHyOcDoA6cN
2U/6n/UDcu0tLlfkXaxOubf52wmeb1Ojm9/fK8jclActPQuMOdToc6lYG/Q0G+tk
nNYSp3L3UlLGfuxi5lZX2mp6GYBlsNhbObqk7J1Vm/gEycuCHxh6CinvcCeKImif
beF7aQuDESK1wAJXf6Lm/OuiUFf3oJu50jiFiDOTFH9jBH4Wk222T2NOD/UYBh5z
eQ6+vriGoNsEKGUhMBCmtneBvWbwuxY+62n6Qwz6EaT7amas/Mhe5kxrMiIeXJk4
oG9/1zRnJ9UzBvuOB/FA3NnVys4jESDOs3cHdAU04prYeBbzwob0j1IPdrs/o6KC
k91qv/BhZ5wmmmbOqlWoNzlSmHwHsGEhxLZWIxhnRvrF9+ePRFp40zUJS1ylGWJt
oeOGj7CdgxwJ9eJUvpJtHz/x5kMxGYvTYm1zjCdNX4EdZmI9xdfdKi7sAnlWd+DL
DBLpda6l+GNHeolPSgOxOWvPfqMdv+t2UbD3f7iLMVD6g71EnA3YqYG6eZoHYUr3
4z6qv9dUsR7UKN/L2VD5rK6ycXSZA1thLVUi5TBhQ3IUUhzhv0Y7RfB0LT1jdFdx
WNrgttEL+SxZgbzoR5hzmnvqiE4Rfk41FXzD9wx8i12qqzTULI2Vf8ygnTG7Fwop
AFgLveLHaU9s5abyziIdD1vNNUnzxAF6WVJl2F1Z9soQC18wdSh1kF2hgfVIsH31
OWx9A5Du43YgSpSSFXDCm2QQncp+RH/0fivN2s/cBPWpFStIerK5EcHbwUbiz3lt
FECgWrRD0Tmx+QDPjaxj89b5QVEQd1R0dOcwqByezp6n7ZsSkWCbqAq/Wol2w1d5
7+49FCeiO1bLt7yakubkvkWBtqTLTDd1DiRwvGE9i4cWa+ezjjl9t9pYiXHv+TkB
xDo0hnULEWibDQlOQH6we/njMQh9W3DJvlXBL2B7kHayZPJCtmuAIITlCWDwNsSN
PkYfOkJuVZsGpH41tlqg3rn4GbihCoR4u0IXApJXW3oFGEYDc/Ot7vawOC+YzepW
PO9zjo07gpbS1W5tKZoGfHBuaOulevSTdiJDyyByPAJZx1QwLbZHicvsFPjqDOTw
ELOKJU3mACByZ/U81t/2e8hlvH7PE1VP1Z0R8hVzsw1SxhPE87s27OjSEqqnFnPl
7C69zQeRNAfKujJ6lt4NGCWHQ2LaB9rVRjreoKc+39nxqWCk5yao93yS67/Fx2C/
fRil91Eayc9QFn/Z6EEKy3wXOps814EXoJGC2PVsr3FNxzYiSwpBJfpOc+eczc1r
N6Y88br60igxRmI/fp8c7TOI8+kNLEFSYGlDGvihNREHlVqx0N+d9wZxxXJ70dQg
So083knyR9GE2ZX4HfRhiePNhzXLuYjGvyTU3kPikqg590cykJD8mmA5iI2paC/T
AkVsk8E/r6iwtxFfw5gdgzQnTbilJzcrI9WnRV2/9SAzCY6JVIv+wdFUZRHxkGpj
Aq7UjozVlX0/aHdfW6XWT8pbVafIRloYeK+MSNPvK7F2mXfvIDtG11NbezCCRbB9
/xhIzLSy0exIom6ty4Grlo8za6Kl7oxotqCQSu1/eZC009uIxljh8E+W092PKpcv
Zou3wI7vxgqHLU/PYGeBTtKY2dgTAz9bAPxaSJ+ppWRUUIJTpE8v5McVK6dvSqlz
324d65ZPUIsXIWEJ8YE9zsxNkTqNkZkDmJ3mRH1BTq7te8iSsl92WIqtAGV+Y6aM
LK9b0BLen8fBhOPgQ7doNKpV9bIHRePhKcws8LyYABWR+SIjLfESncqEJLqsEs8D
Hh+zQ509QP8ppC3auH/BpKTStmk0c+MxmPHNsruKRXmPvW3DCM+HJVnfUSxkyIHC
k6yY5z8lyluQZSmUL76rztjq/4A03mZwFvVEhKCeU/FeknEIGfVmj35tHTeXKyXT
IWKJqf9N6Xtio75qVI7DzjNU8CHAk2R3nrs/czSCtohMmzCOlNpRabAZ4lkBvUc0
N14w46PKeX/2Wt+l09aFfzlzAgU5a0JZufMGm2pEkMKguX3E4PW6geU7hMU0UdaQ
kaSvi2vQvU9FfL1xvlpHTAIYvhxzm50pE3BRtpKYOGXK+eliJKuKW65RlYSpDW3e
7xgrCYGHy07Qyc+QxIB7vm2vmrWjb9X2KtTgmfcHGJG3LViu+/elwZ0+4dDafWXV
3WPSsmHqnIOyZ1F9DlfuJNX9ZELuu6PiJ6sO5bhadspfNCUGLhqu8pccgLMGzpyu
jBnCvD2odNW1Af6q6YlI20jk7LtnMRWCr6SxMF6JYasPgJvcoT8vl3e3sSvZcCg4
0FBYcR302xl1bQCoAFu822fedzYrRfmXvLHaSEpq+VbW/Xnuh76hpNpR0LwIeznP
0T3LQGTbb/XvHoj5V1s0rLNGYIb60K/edFx/sipNZ0CJkHaEELd+IIJyN5D56Itg
761rFTTc295eXrIh79wv3T/liW+n8A0opmTS/x4Wxu11P2WY5pVcqY55DvSJixVt
QwxJtI+K3vhzK/cfaSSw4xp9kdl5O+mXow6IoawAUfsi0XA5F2atcsNN4qsuZpRm
f6d056/0WQG7jDUg4tYYAOMWNIOiiAhI3wmXT2lTv71QecHv//tNb015URus4KlJ
VU6TztSAxrA/bWat55eGsaaLc7LWBS2ML7h20MORdw0hbyH5IqChpRQRoirDUJoK
m//wBWd7d38j7YCJGNf47HlEgDMb7jba7SE3YIA46kWe35gh1JXjGUwVtEBzDslV
BdID/X/JGy2w9eb+luCgQoJ+zZ6jqNhAxHcIT0GuH0pfAyazCgMMgFi3i5bJwmKN
cz+mmf0UxgcYCNCY4uxRNhSkc7SyPMN0sfsgtlZ6p2q2c0E5r8Rdezcj6A5737rX
1w6FLKv0T7CBtr2FYcuknXqCkOowj+j9fzGPR9ZrlFF6qlCXbhA+v26pZmVJezkN
d6j7f0xma817pKPRLwdKuawTtyR056MhQlysgOgxQy22w4sGWrF6Id4pIgge9Tkr
2bM9efL4Qws8/QLhnVdQfS+CCiFXiRKycyFxV/WykwebH/bwrToNL4t8WckhLRD7
1ZZjr1V7LaX1YoUK8l15DZ8zXNf0cmXnJCtupLaQ5EtqbKtJufToj244nfAqN2z5
Jc86d+CTqIly5Cit5BbozNp4fxCuHuplxXYyzEnaTlKTTp+/lODIwRd7SafAWg5z
0gh+NjnCTmWheud8SdIiIs1tTOwzrPg4cwQ4ZThM9ZOJlRUhBuGUBuqqVah1Hte8
85anoUpuhtPvi5l750DZHljQ+U+8qT+eDuTByNP8trkUHXVTAnqO4CRRYIVZNCCy
sWVqTKmDN1BK1fWuaNvZUEHVcTbJkH0jTEbP7Ax6BE2GlVvDD16Zoyjt3JltApsE
0tqG3mex4dCPbJmQcym8OnaekYZM35X01irhDEdnWNxDn0vVgl5js34fVmM7zEQp
7uywYwcm6Cxt9lm7shxYdTfRjtMQ5KyMP8tglfZUmlGsFTUnwRgFSTy1heOSFQ9d
5/v6N43OI5B/R5XBz3qTwaD6almGAk7MCm/uqZfp0KZNrWugczlC6dRLPM4HaX4m
yd0zS1ji/o2BscgU4c1Up2rDno57Nc4JsdW6aoy569n69AXfX076YMtIeVNp5y+5
LglWJkZswWkI2w8yxZRab/AF3k/bOMTdSI06qtA0HVeFNSkhbz3U7wPbk0nSBNDv
biF3G09svYH0HW0lxYPrsGJbgtkhcl8yG1/Xq3fL0jSC1Dkrtg7F1Nal1drXpgEc
UXd6T1Z6953FzSL+osk8zU0cvb7XN4n1GhUV6HQNNXAom6ypv4hlOGDswu9+5Bji
vZwdQJ9LyoNiPUzeYNBz0wqHK1AXuPs4zzdmraakxyhYk6K6P44c0/w2trj+Y6E/
bTmPCdstNd5R0DLK0leo2o7+sXkYzLZDvpR9KVOq0X80EtoA51gCwWZDNpEiUw0D
qchH2UY0IMqAKLdoDJLRtD9VaSTXI2KhNZAfPaLtIy3Bwu/jBmGEwDOYzCz5KOVX
M70/y4uq00GuDXXa5Jr7HrjdmCvTcNIt9CvHJncwPUu3oMFhVYuM47TSCrsGMCFi
EXtTn9AbOMhzrAwpyNAnSgewlJOzD6viTFRPJ0ze2OuoIYBYpBG0+MPka5WJrKRi
tfCx8HLBQDbWRVRYpcXaFIRqplpBeYGe+w0p20fpOcNf1YuslwsPI8zjvB/5q3z7
69zJxTsnxKZVB244Jqvl+GYn+n+/qtmsry/KlsLuSpHEsu6q/Kxl7+ob9uWGCqT9
b5J8fJwnIpNqDiaI6arhEXwsSL1OV0fdrwen2gifpEM5qTsDihM8Uy+OPnflFbH4
0g2hJOGgv+2Xf635LDuzL+gian8BIoTmyi7E16LCQ+XfN511gZnAmOe2j891ILi8
ZeWXz7oP27vrNKXhN03ELDXhBtU5TwaI28H3RxK2V8PjqPxW+7f/jEVzWIdYycCK
Ppb4Cxp0zxtTMt8CGdxoQ8wtZDd+8Xv2wmK5U5/oKMYEK4IuPC+UDIGuWnGhdyC5
8ekjmHci/CjxElw1SvDliUs9kGQ8hflPe75UkX/5jymz4SI0rOZ3znykiXJzTVpo
3uwB1lK8r7BL48T2mb7u+aWTHt6ziHn8730yibZbvvT9ZesK96aUozYZ91r/FJjx
3+Z0LLWX/B7j0y1cWBJocJpsltOQvCDtS/e/Mn+HlNq1oMdRQAF5EZop+xr0unbJ
XTXMIflZSM0Y8OuWlSxZPAcmeDDji1Zm5Sz4IYGssIJ/KTFDi1bwLK4LGs6qQQod
y8xW7f7RfL+CUKR1omz+z+VzI9uEkHJRLXwZjNAaJYdTtxi2EqikISt6LaYZH8TM
Jm0XPTp00VKIyq8rs7Ar4h9GIsk6zmM2AlV4UhVC1fzz7olwfI3mhs5SKnlRFv/D
AeyKGVEDYY4t//p99d2lYljqC4v4cNWssfkDexdW8siLjsvD0r0TNDMGbR+qhFbf
iiQJx3bZQ+dhXXw5sdwARIzB02eR3ic6iz6RzbGnqcCWMGZkbN83jDQInaFzN/xn
43PAW/q6SZA9POkefKRx+AquIk73QWwTGDvSlCz/7sJaTy6xrbrV8L4id4XTNCan
IwnETlXBTtRmdP8q7ZNP1WLXUGV7ztsWHdwNKe3IhwYJLs1tSzm59ZRKZ9ZzSq2N
DvEPKl7dswG0MvspCByzeUhf1kxSqMruvQe14uA92RBVDL4c5GbBzWKyy1rKD6Xs
exGM4yNm1TkIDBHsIUcTFu1yGH67Rg+D/9wDFFBkSHbHS+Q7knZcucOcuuc30bGH
pBB53yzYxN53fHdrwPOU89sJA+dx2gE6hFSk4MgF6i9MV2PY6mle05fWdzhmwY95
7tsVZKYoNbiiSO//ZzzwEkV68Z4qlBwFEiFq1E6TLaCmzp4xfmgmgpLoFafg65GM
SZW9yhm+wMTVcLw+tyvlhSdQ9ibxxIyfC10q19ohYU//N8SpqCYOxW1I6VfKspD2
KNUBOqHRrNu4gMmbjfiyBDryXkYPS6hHP4TV+sH6HKHjcDBVk47me7iAyGuvj+EY
IWG+fP1aJx9ZOea6H3lKF6KaLQUtsA64jOFux5exMXlWyRYrTGs9iPL3WplBxOn0
sae8PeiSi4kOMElvsFAogDaYVIQewQK9hdOwNZbKDyy/u4zAMF32g6kEqOIz7M3S
3KFQ7tudbVWsHhz+q0j/7zuWr3u/E/ahOpQdgeF1XrvDe+cfqexbdSINs4BiRTqZ
62xHJqOfwaE8Q/iYmF00SvMt5qBS4pzTE0Hz/ehaSICrh0c64bZ5f7tlyAJKR+M8
f62Dlxduz3WJrPi/Vz2claT274u/vEQGtZnrYr+weGOVfKXHuVybeJbFYTx5JOTy
XLE4mYK4neOwzqKN3o3MX8snsiVK2QKSufOCljEgy9hbN0GHmxT7jlRDyflZaJhL
Lfbi8hRdkjp4Xk4I4JwgKauao+VTcxidfVtRIKTAZZWstcl9ev2pqLdUXb8AN//W
qWfXzc3KOzGJUmGirEhSppzXKrmj3MG8/RDtDx5JCf4VwacBdn+6oKmRRRKpK5I8
eJRru2jFObPz40UlzG9/jcmCaTDuMRACK/uO6o5SY+NRNxKNozgFilXSGtX3Mm9i
Lxll0h2LKf47oGtHxOglApOZ3cswtomFkQh044jjfDJN7NbUsVSNKwzIHUC6BvU0
U6YbUfXDbfkZdOrxZBbtBfCEklvgM8nCdxwnjjFyuyyhUbDkIMGuZUUyDIjwXJY2
iZcZiUeeKlmh9UPWT8TgtmT3QwvVIpJNAR2ZFrHfOupvEDx4AerMN/60y54cpBKw
3BxGb+49VYpcE5259kpE/SOxoikGl1Gm8BpB6hHfWhiLw/GxkxA4haVE4AYLKvWh
tCj8SR27AzdwoK/XRDw0Afx+Yz26rnuYSXc2v6Czu3x24WtA3NV1OngIs1YO/660
5hPMTnpFeXzh7wGV56qiyEulMZtMjQwyTSp/ACiwcyVLg5wabs8qj8OZyUQ374eB
wObysINpKFPJuBJSs4S8r3lIWlXrMsrf3nhwxGJnF8ZWxa27X3NejvYD56hrpqeh
sGRyOfZsRbBDPfEeuRe06McVRixxPNDT07P4Ki9elf2ns1b39t4ntYCACBKt61zW
Od2xxvwwpcHl9TWTSRiC9bF7zytj2DIb9hAA4BHfbr9JI58UETojKmSwhHLvOSnC
WYqFlYV4jPXa7OoaAueMcKGpMKe5nszO6fy6DpoM3FkeQRY/b3/h3Fc+zkpAPRrq
9qUaSN3fWtqPubOWy1uJuTcG/Vl7fR4q/1a0t7P7N1TLbZFtNFPkA14oEP0jyNRl
/0fD3V/8pabLeDWhHBqytCy59Hn63KhhxMNibttFZHEfd9TNDfPWgaF+V6b3l7bz
mRfaagU8+qppFSV+hEVUEHOKKWKv+ihqZKBwMCGQlTzG4qAvhfLjWaEcBcl9olOw
tI9LeumTlufxo22+8iV2WDoP7R/B1Niz5ooaAY+CmKRQ/pgecnPEIItyfHoh0sGZ
VcscGWKE8u/p/DWHaNFpfGAs8uiKwmwGF/yidGVXiVwuB2A/fqLoIH4K19/h5cNu
wEIqhPuzvmxU5IJiw8ws6/Luaw6SQ8Z4s4YsQfhbj+bJBGOE4GR5OwWnzc1xamX8
hrxMqCX31FUTJjmD8NMD2mdtdpKyR+T/ocZQloq5c4JKklWRAT0fi8h+QsE7fERG
0NXwyekxUcLvSc0IkTd+fq31ng5Ossc2nwNZlNvNY14K5RdkWMP97iTaZhbyfub8
OewooLaEujm0pJQ7VFhKUYJPDMZRe0PVWA+kY06dr9gco7S2OApj4mfr5PME1DHk
Kr8jW7EgiB8Qu3rQUq3n7y/JYZ/zeaENQimn7YQXzgArfUrF0q2k3zzisgV04Lo5
0Nc48/9ARwQAvGffdQdQWaq8lxz9kjQxBHwNvzE5kgTQffndYOt9ZZh3l7zXERGL
/atEI7ChbN9JOUu0sOQODwU0ZEXeO+U+H98BQlLbg38muEbwviylx+j2CuZMzyM8
arfZVZaZoeHFDR0kyRh9+zqFJubGJe3IFHk0aayyDkYCiDmqz4WGU2qf54+6m4VI
72G0TVFazFTwG9kmTJjX6hEbKptqn7Q4gDUsKaxHPC4SFQTq1T+u1JjCVHeka7cb
zZ+xledHgxmRdz1iuYS9tRFw8B3V5gMASTW/rg4R0pa8A/25AC4ygQvaxIZUthY9
qGl6K0XotUEwLZu0qPULKW40bRaEQcPF+AlYHeLGPxLayDHt8Ka0791Hs8S18RaM
r7JnGedOHK/2bOiLC+NmAETblx+Zd3O9+kmS0pfjNGDp/RKgCqqS8nFznbsKlmK0
9pJsKU9eDi1dbMnuK5omAAjH3oC/XRT8uwygNbS74gKmGLAIOaPCroTwDJiVcllg
g26hg+CuY39bobi8eaYdOxsjqWabCkwUqqmusnVtGMCBdbTio2SqCk8/27nv4y3F
pO7b48I0ewnPz6R/WkCzznXl3j4lQ1PiDOmbnXwV2C0QLK2XJSPWhktoF7C5qHQN
Um0ZL21PjWVMuDX1zlGSNx+6Bz6tftugV1/EzY0B8uLygTVMxJ230NQGHVPf4zIT
MFquCFsTMXZwiIOwiX285oasHpDB5sNeKGfkCVW7VoXsE9YtQqKJYQpCqIrPs4tE
xRWD1bT3b7iMfOjpg6+QXQBK/t2hStbQVOdoLtB4R5Zr331Nr4CJWjfszW9MI3H7
qPyFZDRcCKGc588SvlATfmt2TvohD6NoTNhUphE/vXNIt4q4JRTS0kUN6DnT9Gqr
DKd4brF4dqt22RB5nW4EBQx9Gtj2OBK/WtSX2ogB3hKNOL2rUwLGcEQd5iCz3+3I
KI/+wq7He4D+xKkeEifDVLBRJ2w+9v33mUo4KWkKOPtANal73+en76VryNztTMD8
6aOWwk86TE2C2C+XkKyPVhUyGFS6iz/IWlUVpnxLWQSbKcnRnc9JporqjHN/L/hi
L8X9xasg8lDmtgmKC8Gh6cPVhEUBsnhaf1Sxh9QlK0bm5lwpVIzeQmYqnQq5JS1q
gUxDhuiGaP5PB1YigDg3Jk/7gsp2JI9z6nb/JLLPR4fS/CQOiLjSW3KxZVWwrzvd
THf4x5BFhVFEDQRgxCeMFCI3yKqwvpM/TrepczheS1YffS+vOPmE908mvMFhDZAk
Zrc5qSqToUJSBGSKUSwPOVHaVNWUrMM2aN0WrSa5MBtNwkCXVktkFyM6YjROshyy
+3rJPwNJHssAx84RpNX15c+LLriy6+srBm8yUbi7r2s72EW3/6/lzYdubDVZKS+H
kO6GByxIZwsK20zAhU3/3JMXohQT3Tp0igMQemXI6XZ0+Ok8TyVqyivXAiEDAX07
4ldfk66LOqOhNGE4lL4RDXvKlCZbfEjmjBNsvc73N3rIipNz4u6kuqIeQ104u3sQ
tb8MPZmD2NZ9SQkeNm7eGfk04M1m3Sfh0DU4Kmf4Sd5eW0J5Fge1q2d4iV8G0SN0
gcF9g8347cEjPIUbaTX7KbU+DMOW2VHlFdSiSr1Fb2zsg5ctEgGpksgJtPrhZq/X
rA28rzj0RwshlM/H0Lux7zzQwYI1jA/cEg+odDL1v91zLUciWKVbz+7mKblEH1AN
sTn0x3fBZmCw7oI9cEusHXMFDKFZElsruiMITpArAsDpxSjbhzyycBXkYVtHIxsZ
yDlkbkXI9ipGElt/h7T2qwFs/ogJG+XsosEY4CxbDTOrh2pEwMkCQSQUueGi/nyv
1hUGAm7Gx4CVCjv6vR8VCFiTJ+ww6ps3FIfZC3AeqK/4praA+WazlwJ1AJSzbYHc
G1sH5a3/WXDmW7A98UbvYTYFdwnhHZ3EanWBe6AA5GnL4j6x1gD/90FwAZVAKiZy
1Q4KAzUA0ZaEaoi6GUOuKkeYYuvd6ILVMK5LCU/NV9rrw4vPVX38Batk8ZEYDpAy
DTp/OY8fbqghMF0NyFXFpiz7JogUsK7TcdlU6AJRkk4VZm4CEXnRu8u1ilY2GIiY
cmNhUnVwm2XXFA7e6sFrKjHxKBL1XrT5mNWs5O9virEFjMFTvvO2J4MNOQ+Mh4MO
YgRzhIpyPsD+fSgDRtm0O80RcqNsVQnIEXSxTs6TiAuU+NSs0yNPF+qwGsSVDzBQ
6oJjcpGQYkB0Gr3B8pb4P5Ym3Q3ia2TBHLTLQH4TRADZLbxPotk+y4f+S3I7CXIQ
ZpbPI4YX5dJQqWne2lgk4WSFcJzUWCmIYWsw8ujUBdnCYCdFCmqGOlBrVCSQtWpL
Gh1QQMWONBuZi/5bRSgqTTD2BZseVXIXCLtPsYnEqxLpGPjDEP6kRbtbJYlW6q9P
rywuqWdP10XuGs4sasA6Wo/FlfctJVl9mSo6LhjW406c/QIkOlYaKHnjoJr32GQV
MhCLJs5iyJR9w0WsVju5uqbU7/MSPkLbHpAEaOn922ag52mmj6rYMruZW23KErDD
EuDvKznEwpdRHxFylGnZlOneLUVSMdxJtRi1ZN8qcKS1YeXUeNmUOdgIeK4xqZGw
oI7gSVnZXoPZqYki5SQjgSbHMGEMwaV3QYrAh+lG37o9JSA2v+6pQTmwx+8xXheX
osN6JPKyJp5lDHSdvrfj23jl51RlGVYsbm0l8TaMXBYuqmSPDvv6M7KAQBvgEDKu
duK/LWcbGGT85WNnLgggXBKHVlFtYUUhzndtjVu5YakaLMyYLxyzSXO8T91lIg1H
WBwjJx4pUtn0Gmih7HcxDUMqLNQmWs48va3J0jLfOfq9meK52KNxIJ+P8pBmm40l
yxjm5gXB5lT36xhvL8T7HicDWPVLYRuf9nlhhC9ssTQuMdqeMltMwS3LbdD85Yjb
AjDr7e/u7bNZj/41Awdb8kEZu8vXoKJfnAbXkUiyRiUOz1bqw4gVaq4u1y2qFMJH
+fBetfFKLWFZEnUgtGIBAzLbSYNOFsBj2E5hNcaov1ta4r2zK3Odt2uTa4aX+sV1
rLS19cQfLyZVgOqNONFupGNTcf8Je5nwIux76Fexz9wvqYb+znTx8eiJEvmsI0yq
+HZILopCLfnvGsXeZJLg+sv2kTp6fRAdAPjUe1tJGbdy5j5Jwz3ZobMj0wfvQrcW
oQVC6VS4g2c8cz7QF0gPy9J3GsZzqGHKCPiw6pZcj2Q+2pa2iVSbI9op1HNdKLCe
vWcRdnTb/YWnC49dndJwbrKkJHoAeXS9HoZfIRwH7GPndVzOoIoomDGm24yGH3iT
D3XICpg1l0CINYfpVp3OtM0GaQq3U0fNfzmGIrVmu5obKUk7hzFM4nbyLpMIUMkh
ZpsgSKvCkq+5ftS177UpDsoa0YhBFcrqPk/n8kiFVNeU+6QtZ+CcutOolvc6FiCK
AqgWR9T2I9ScVe4z5/PHD31z81KyzPM+FPNida/DqsKhoLAaC74KkzRlsq4HsHQN
PF8HRUM3+jwRBKzQTa0/BUts+wRCtH4Dqk9e/r+pvPaQhNuPxr5fOrJo9ZbueOKO
N5na5nkkQchvR+WN1ukXQnxd7/4ZWzHwbocPFfuO5AF5qIlhNLHSH8vobl5poQ6p
LdIiX3nhstsVk9K+8Tlpeer+mRZ7/3rWnXzAg7JAb/IIsPG/ZPuwlKhR7OPLdQfh
TAr08vn2vu0vUqu3KOUtcxTbupRHp0ZzmXSHemMGpabX6Ue+uQHTaqy5yL7yMEq0
2g2zi5iqVVN3/TpI05SVlG5M6ZNDjDutj9UdyTwje5mapPJVn5tGDtPgwXvYSL76
OaM5LmtaDO/+uANDgIKWdrZ9ETvGA8OWCNupZlW/a+VOIwDu+F7Ld7CqsDSevXHA
eB9AZhQslH3Y96TpFCVEQMVUUGh9tk/brkhdKVk/IWGg18zwv27Ia939001CGfA1
jgtmHaSmedfbQBOaEzHliWxBA7sEqa+rGA8WoGoBvKzxpPWNK9Oz26oYH3AOVQcW
Qu90oWEt8SP4wuEYNWp+ntYNMfzuX2NEMqZ+WVoPAoB9G68Oueht3ITv5sS/HD/B
D1N3qNJO1jzfgsTZWSGm1TIHRtogRiACIieClCnLySwzlk334AlI/sQekWtJyppD
+85IlqqHUPn/n4KoMVOwupcOYSpdjh2geC3VqR3TwsCgkMCHwir3Uq31zD7P3zG2
L2DFqJfchJyElOFQYBfv3DSVquT/axrsPlrl/vErMFcTnrnAY8LjtagFrY+5Lwpx
JOk00SOojx9XfMJVOZTfpejKtp9FJCAlHDDwMuuokquFP/Mbl0kpIcj2TcXPNS+k
nt/dICbeq8AlWhohGDFnsFT8rHwSOO7YkRlhkahWTtBC1CPHACX2ADHEFBszP2ey
T34DLpe51kzCL/3IZZkGDl1plcz8x1q1p/cC0mdvSqbeqlySJPe2vfjwVIDmazPY
KTgKVmYgh5vCDLXSsnYlTM+aR3xyhV4tRIKTJMyBGjkgHEZ3Cio0+pkNR2lxJ0OZ
X67bBTq8hPHvchbAx0KwEl/djVlWvOhwzvuyo8zCVevIZkUPahh/9emtK7wBXmkK
wnsZ95Uhk0fg8HcpiESLKDe+TLPTv1gj/e95e2pi/MhWihD7Mxii/z2tX0+5YOTq
iZWuuatqGncT0RofKHulKbXcvfw5uY6BFqe83taeZomF6v7eb0pnwKBJAzXI0UhH
Y7UTfVAjt195LXH9nPAT336c94YGmuXfUUfBY4ZO7E9JK0QGs37VatjnXNSasB7F
Fhn3kwDvy1s4fYxsdXpMfcfEEdOvZK9U7LS35G9uFfIIuqjBXQdul5RspwodWbJQ
uN5L5pBpcPvbJsLHGhspPyTUGbxhWvWDmbWrH0w3QOFsJxKqtAjBb7JajgI8tFiD
P6v28Z2e8gPvghJF3MHb5YQ6pswzLcLMMomkp8/+7K12uNz0iioGKeQyRXtBLaBu
RDPy6FAFD4Te2qsfu+LrkvNmlnoL0W/kqlCStR7L/dp+JfUu5ADElMhHb8KoeI2B
dMB6ehyFFcCCf1AmSK8piSSN/Z32eLu301dkVFDbtnEOMYl5Y7SxwHejWgX08Xyi
tsXcvONRxSXD93hjOegzpbGh71KbwhrUlX7h3F6lj9yVo6EDia2jYU12zMVx3dwU
Ud5mbpvphoxTJwpaPZkI4dg3qIEgiIB768ZJr4/ZnxioYg5b/aSs7Jvbis78zSvw
fW36LvHvPbCe9CpfBtvCVc5rFYsyjCdQuXiuI2YVSz0+JxfU4mYXtg0NxzUpIf+T
p+65D3WDK7CkUPoT+QtN2Y7BW0ZpY8Y1ed1kUEeJayXKb40wq3rCL2gt5EPCA5Az
vboSn0VhPf3K6eAJR+ct+Kcr0hGqHYRlvf30lmbQ4W77fi/vHq/o77MEr7OBHciV
E3gxJDgL+lsdKJBlRbwJLG0BOoD0bl7n/S3MVDRqPK6WsYuQa4fT0iQUT/Ylo+kY
R34A0wOoyDw3Sm8Tx2Xk2fB6+ng3+TiZquSCnvb/MMA7Jxfh5HZM1Arz4LYW8WrQ
STQ1dw911j1cnlAm+fZ6ilLZMNfjg4zYVYYMGnLU2tWriIlyrW9QkfPQGyzbYD3J
MNiNWKQb49KyP1oUgHVT55NTAM09jrRL1dVQ5wvFV++Efq7zZRguPf4tpG6VXCVl
`pragma protect end_protected
