// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:19 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MR8l+wX0TU5PCMHpydyAWfKEO40EqP6vh0Wsrsm1CmMa1hT7u+ax+J2G/4XOcPZ7
BXeI2ofDwNZLS0p8fHDl7W0FslGOh0gFNdCU6SNCKbpVp6i1EAmoY3Y0hkv8kXCg
2rC+fI94brMUmKrBArZ2d4fspePDpM2bj0Yvu2OawKw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 44064)
suwPMSbMGUqK8w+TeEcQrQdLyDSfNkp2eDch0T1VwA6FqwwH3/E7sBESkxRbAFt9
YhGz+gei046lXFBV0IEvwW4XdDaIBliAGcb8GRPhIOaRdT1uBRz2IHwYQvv+CmQx
Y8WOMqsjUpHCj4cYvqVZx+WzPdR36UvmtEYVnLGHzuC2S7YlBtCbHACEqaqsP9Pb
0j9KVwEj9aLrjpOQK1bN4ru2/AWy4+5ibsYI0tVp3u1c1GmVo0sSdGb7wJ5ZTnYC
h0Tr0BN1D2LGyoR3GyDl8lVAgyYuNuE9r2RBOyADF3IOjkCOrDbAlDEGpQg3allX
gL7pGiK0oFN45R7XV3FGB1l1aG1QX9pTBieIhz4FlciWmQrKZIBVB/R6+3HilNq2
x08q2Vt7ydMBOMCsea0Zv06JHfbp/nB6qaVKu7YSsscz6W9ikfC14c6/RdRbKhSx
i69vWahJDRLq1M8KLitpcVTDtDxbpzKfpQecnKGXJXJni859Knk1V75B7L2McIHS
Aaa/XOcG2beQEEukqMlkqdSPU82oRPXISoYbqOwubHogrUfZGMoP7w18oMxiqaPv
e/r5Vwu9Auerl/PCsfVB2AgyhX6890UXtyfn9biUV3fcznNLCGylmEJy5pgy9mEm
O4ptThPErl9LtPfqrFkO64hrl23LDKNOXZb6U1kUdLeohrEI7WFC5FbHkOuK5DML
vGP4/Ef0DDT5mVJXZbMy796+sngPBFNMcFOTeJWgmzyuht9g9lR+YjEjx2oPdMjv
K7b8WohdnthkQrprzQSQ4b8HNDQaHQoKr9gnWjlVlka2zHlrRAkxmkkCFJFFtBb9
8MPZAzRAo9JujY2p9ds4k0nTlTw72X7tQ9mV1+HFx+/RF3FG8Vrp/1mllhx10gtz
WPtPZBN6mrP2pEqVx+9nBYAPJUnTrbkeI8BxaTdGKnP8BN3vcbUAbzgWdR+b8nlv
fmarOO4hNa40S1xNvSCy0Toyag5ko5fdMCHXGcX8mBcM0rZEdB+GYFq8p+GYDEjs
3toLLJ0rId/YLxpJxreFeNR5pIVU1fFe47MnEd8Wao9msc1VBRdgQaK1XK2FwRSN
1tCPFuQ4y0U+A9XKp3PnI2/MCslnFdLjJbo04J4m1BiulqQZqJaZmFiuK58LvQZe
bks3guEq3dKyUd9c4z9SDXPft6UucYtgN6hZ7b89DD2ieX3odoUVxYqJYAREbQjn
cG5bvnYbIoscgBCbLIWH5Oz4NxReD9Q/xV508Py6dy7fW4ffUAhWZpC424KqWpcN
8SED3bSRoySgtR2qPolUXxCHh+Hgyj1suOIqqGPyTPqxU0zBQqefeErMWif7r4tP
rAyvmjKPXxj5gfFkbjTNLCB81KmqeMSEZNaP81qJ6GfG+6KWF4zwysyBq8v+sNwP
ei1LUulHjnZp/A8eib0z1D0SBgIjF3mAOP/mENdrRQzVpCroZqSsE6TiDv0DqUSo
2aIx/FtGi5qLpW+ZNz7zjkkL5NPIJjdzuiOOKrH5p55zp1K1Lr1hT3mDEL618M04
bUxI8IXxxv6f91JqKaD/SJty83doZ3Frp6Po75kT+dtgmpWywA/TBC+9MKh+RqWi
hpykzliLPkmOKyAjeYJOqNj6o5NrzOcHRtzq0it6QFhk8h/J3AHtudDx8FK7lqgl
UJe7L6sKQKHJPT4JEQysGNecCuHJU5DiehLro2dHUyhREVKF3aNEr06l0Ozhxh1Y
t8LRDhToD+8OSjwswlHWDncCRnW7fALMyPcmX9Rrl3h7vnllT4grpwKxwpTofPhh
vLitxsL9gOWTKqqfFUtEeg9bd3j8LQMYljpN96h59Y5DwfCfIoeA8DShaamjAJq8
/Dngxd/sdruyM+Y4JQpmw5QCJSYm9MOEW6qtHxZbtCV0fPjHpeP6wczIbm3466q1
Al0QxHeGVkPnJG7te0OOyn9+AFSgLTB0JJXBwo7nnWKashkFewq49BTEC3riGEj6
auFcT/DbxcYwv8j2GZ2Wn/efi1XdAI0z72F7X5LYJND4IDMb4lUquaeS8CRN7Cbu
ewA+VCpQA5AFOZxJMvnUYwbW9ike8Yu/krpXFBZeazCXxPrUJuI3riziSK5DG6gg
qMFh9G/OrnrWUGHFf1ZEobAeoQGTM7sdzQVCa4Vf7bK6abKQ2Aey0wMKhDp/i7J+
6JdyrRcuYfZjiAkxhhRITl6cFs/a5Mi/21yOy0lEt8E56naZw9y4rRfS0Sy9+DW5
MoGY+AvvscgkwU4lzDMCocli+sh3DxWgvTyzAug2Qqb+IoIEKq8wPO9JiZmDr6io
557IQ17AdM4HHtLhhkmRFjZJd7uZyddsEqWVRflu+1WEUqqNR4wlSNCEMLranDNT
GG3/tgQ1yamJuPda11ByWqFPgYBymb/9APHxnhST6nUg3v1NPDv7OwBy/Q3yJ5xd
2AB8CfNH/wv0otR/BVfEdS5LPeb+bT83RRiVgsPLxqeDRSqnztXld6t20HkqbGbM
FLwL334nfAgjMiY99fmOkNbtZGHrxaD26N5mfxZQ8UbydCUCZly/VXgup2/ETmHd
qL7beR8Z5qnRSRrXKlbsN8sHm/N2nolA+xVFTE5bTadFY+8B566HQdEMzRxID2In
+QFot9Pf8lbxGnMPuWhpUYS8rPo/VMuKYdyThMgobxbLx/mIp1asXwZxtbw5ddr5
eAfUAcK6JEeSXk02Hd6XKs6y7hLF0ldWPc2K+biOxV28+vufluOmRlezuXE88iO8
ifDE5NyuJKWATVX+2AOrcibhU0zVD9TB+S8EEP9O1FfjZuSGNa5sdOD+zJ/oT8qs
wQwRL3/8KoAP2GpgBGoWn8SD2pqAuYooejjS3Na0yrgap+iFB8EvUbD2rkqJHcdJ
zvxcrVql0yV03tNwSzA4NAPCQdslaQ5cuVij3y9AUjA8oyZKVZFaIKK5DbrfHoKA
XlAGjoQRFHTMjFWX2GPt0L4gJQE0mlUIAJDYPnqhJmGftTD3AAOf153X2D0DF3vN
lB95bZubId4SjMaLqNJaQr0brcuoYoXrE3yGnLRtBJA4DtKpvfWTJdSGB+a4jn4i
M2J+XUzfkKzlbygW7194KIZ+Ryv6TI2EXqZC7ytg2JB7k0cC3A51gu6p4ZsGf81+
n6N8WPrjgS5ilT/Sz0o7YHwhO0S41+108cX6QAcgg0oyvxL7g7OmJY2zqMGv75E7
eMQlxUZS0DaN7gVDP9Ypvh5a6n6KW7a+Zj18wdIiV44z+78ETF6xpjCq6AqUcf20
gSbvsIDRc/PFuuRQ+QgKbZGjolku7ryTApZ+AdPa+BFnt1nV1uYHcLmkLtb9Pogq
gYih5oPY70Edd5M3m026Q+JV+Ou0Uet5Gq984WGGFR56XvKDx+S21RyORYu+wakf
MwRmQf2aTgYSQwo9JxOaoHLkWYGubxDgCTtdXyDjaVMDfWvcXVJdrzfx2k6K19eO
eO61TRGDR+7jBwIDyYnzpjrysxhAmYb0TgmcuKbKHpLpIi0xFQj7+KFBxEKQDzJ+
nm01bZ6aaraMKDEBP4mjqPPIQH/5ZqAIBpEGrla1ENgb3xc9rv8xBMhiQQ0xIVGe
l4t3Af50NzyCbC7xk0tHbw/6nZmNpzxHI5X9wm02uB9zBr2VeuPadcEf1hr5ks+b
EAZsAzkFb9Q6FvIYjmrXQWhgT29rv0zP4F7eGi/XIBwv12nQ+yGKW5Bt3mYbvM6i
+2cW/pF/XEmnNQcrsDX4Bt75hw1/37/t9cQl3SfyWNX0q07gy9vAfd+d6XAqYHL4
hhngCZ42Sh8n70HTxknwNq+I1tcInryqXMJ/yvAdm9ORVMTUGiKbEZOYc8o4fBsU
PkyFXeX7CzL1KHzJbI6UfBabJGxtZrRrymA2e/Rl+NXhW9zP9Y7WPlqbBABjsJDK
HrruJ7lDwESlfdKgAVy4QIlpPPPUDFF/a773ZOSdmZ5TCcZvfQRbNqO0MeHXCLAe
SmVwY67IgVhhp8PZrQhaqfVhq8qfQmqvZsOqTruRoHHrSeqcU/rn+TllgZXWwps3
p/+uiy2f6s1oZiHoSWuCNRVmQ4Op3yBeBmEtOWuRIHnawR+UsBDqIz8IU/I8F/sv
SC8++iIXqXrnhaa7i+4pRHALK0EavBn09DsvL8OMKkKbXcFzMQMZHHwd0dKn68Wo
Y5ipa3X0EPlFQ4QgG2X6ScyNF57zkDKQf971uxZqrGSNbAjMdD5jg7n8aayXMkBx
rprKiikAXW0dfaDNSgPuirKSvPlgph3BlUSrvmrYxuitLnzFmnj6zxSY1S4UWi97
dhdczllho0TblLsxeUi441I0sQm9LrBJdsjfDI0epHcfrwKVXAJyC05GW2qu/hRI
81p5IHcerNyWqK9X+C712yF4EVnq1gUpp+A4KKhuet8fx4ihgxSAAsq/eAgY6t6s
zQlsthgT46S4WikXsu8x0fwerhM/3EXACFzbf0c6H7/rRoRw9pdFGsip37ZVBG/E
XoYdJGa6/HGGXxZT9ms5Li/+K1S8H44HohUnrtXjXfQQo6FmGqVkL+1OuMbOef12
ZzISQFfWSdRwzGGwViOW87iya54+vSAUCaz0h6wIIl9pbxqHdQhU9hvgj2cUrMQs
D/g9T70qNa2p5ZyGF7p7XxFqroS3liYKDS4rybJ9uqNJTo3lYpo39G8BvKtgL26I
OCOI0lSvqial87KXewfqtNNtz49P7RvYEgxzoDsV5kYJpbAtU5lTB8P3XLWDaIeK
1Ae7UFo9fHlCBlSjsF2qoDFyjoLubVK+2TB+E2OyPO2jlLn3d3wDxsBYl3QCKz19
3WHCJj7GYxw60Blg9Z6S01i7F0DX+IkvsV5y32cSE/P+VnndJRXYvogqVV0TIKUO
l1IYbDuw/43XhXeeuLPnd/5tO7x8UFLwPn5Z77hDGaIS9K4CbLHSwBZWhOfj8d9J
6zi763EuP/2Su4JdYx8rk1heRJTj2SabdZQ5lkp3YgzP2hALzYomdw6Y32qTJdfn
Xe+KIYKJgtFOelFFOmi8jwlFfXALj4wI3TkYz1YWByQmnHfZ56PVPQnazj/wxasA
2jAhjrRwhNyhSZBBoToRL0EvZsbTpExuLcLXJHQqgeu+a80JqGf93b3MvXFfYuqj
xOXRmNkDytuxVY65QfjOzM+79n4P0O1QkgIPIgh8SJ8OLPAGh6q6+BNsIjRxr91b
q+AZOLBB/cslNzQHpHWKwPA1+PiYLpUgYrL87btuS1aovaWJnYw1p2BwiuY0f7Yi
eTZMsZYD0ip5V+bROT3DJbrwHQkTeCow2LonGIQMFo4VeB8+tlzLkZMEX4dZqHAd
cLO3e7GWeIGEDOojWWZPm4cekxcXmpFV1+3gXoircG/Ou0p6gHe41Cvi9Z+aSjIR
fbYYjehyKGoqvwwUQeB6HMtTkq/59yp9Kkrpuqd5QynXKnRUtiR+bEErQ+wolAtY
ypfnQ9OZIk/almBVZMDGwvywoo84TCgpzm7nRHKVFiWZ8JJ6/SR55Jn7o6+6BnoS
57kem+G/Ukk6cW0/XaNreIH0vdPF2G6no7PGgZMS34dkkjpjhKnoNQbgs6gZW7Ax
ZlUxc7f8IRgPdA1aihUfr2kBsP71ObWpej1D7h8wZMjLKi6x0f+sUyWF+2rlrvjl
OyUrVmEn46HBgtf5heGL7Ed0dMJIAC32Uq4a13gl9ErtvXtJaFT5yIi1o+xGX8HT
wEaGZwkrbTIZg0njKG+6L6v6uAJyxrjch4Rg17iLEstgubYWNarZO5Hzb4npVcsm
VMAT7B4By+hpj4HaXPQh6oppyIpHuB/yC1K6VVa5J4+5L8LBmj/TFiadFyZKvbhv
+4BVya/aggKKIswjtnFcjRgoJHRTESypWQCrEN+PpbBIP65awxXUgI5uJgw3FDPf
ZdPfNE3r7HQroNlKilcRs2bze0O2QRTSfOX+mXiilKM7XzCjG5+ZHakoGQ8wsSHi
0LDFQnygFujzd5mGqrZSkqgeTOybysd0+w+dbBeYfRwX+KTzcC0xDe6CRjhgLNvd
yok5belFuxCE42Ne8BZXLoPQt4daXD9qM1qNZbrdtHCtJGvttv+XDGGOQlkDlZG6
SbEhFCIG7OVCFndyMwN7f7wNgMtZ7LyuZYX9JI8j5Whv1afpZ+PIv/WBQvONwtbq
9JdqId/U4RTCfj8k5IHne22YLL46AX9BJuB2qJnS4CsTcO7PqmQ6MewlSbN7az0s
Ii52N7I+m5LhXVv2WenXgK+jMjQnrmCDk5ImN9//L1RTUwos/Ju0G/U85+fMU+fE
nMBK4xMlh4KrNuzoI/s0UQwvTkfRynESQDfUz04NUAzcTUcNMZPeMke4bZMZ9Bmh
CcEvPkDkXmCHFWuy1+SZ6UGW13IMlb//AIEq3kA+c9Fps+VpnV4vcVNtA0dqzhRZ
1OhYuDt4SCdWHJLFQ+xnGcMFgsPaTopBWur55kH3iakdJIY4vs/D/jpCj0qXiSn3
6zvD7M071ci7JkyJ3t6T3hWCseWV6zBNw8BURKjozA91ZAf4bXQkjvbHHaAYvt4O
gS0mN+4+NXNhwFjhLYicT8UjgXDbCqpvbWRMEg9mqgSiVakMcRhnWsUIzx2mwG5/
aRzFsbMY8As/PnCezFZQuZsQ2yoxOU49motTTupF9/AK1dZWO4pWbgRf1YpjFMcG
8jxSg9bkm4MSI7bdph2gxPRB5x6Jfu8GqAz5znCJS/O9MN3Dvdb2pgROyzU/7tdE
Bzdn7qLxn64M4+Yq5Tdh17G6WLfLGHtk0+JWrtchXMF4xz8E96mEmq3huxdr3twe
ZUZnPhueRD3cCjhDcEvDOz1wTcq1w9zKhPVQc0japuy/qXkGGLNrdMtDg2lIyqWq
en3CaIt7EYsvDnLJVoyIHZsitfpjiqVlIt/HRZaojXn4EjWmo5hxIcWcUYW8Y+Yv
hij39Qtiar0za3WoWnwGwgxEomQ96vA3qo3Tdj0FlAbSzSZGnf59OiBgoVRq3pPN
cjkQIOo0z+3Mom0jR4F+3AJRth7EWNuyAiMIpKljBXPTiVEJ+uo4lf+5iL4qQPzU
XcWzlPcAqUUIIJBqNouSiQi1kctsjIgNZ6665GKiMVKkmvPfyJKSfYzmdm2Gp/Q5
GY/rBR/w2bGXBu/V4xsabDrr5bq++JEYMU97/nUYwNl3hBYcg8UGd6nTXnI6ayXC
5Q5wJ4dxv5Fe2z7PB2BGWYRfYYZmy7IsNPs8ETLIHDLIJthg/PpPjtZxX42sSoRP
nSP5UOdCN334d0DhcQCVnW04V+UThD+W4LpwR3rbOvRmsZJYtkBRB5a+aeRaC0j9
IjV8SetWWbnGjugcsvinmCjXzx+il2xWT2beZi1XD2hKq/KeEZIg/ZaMEzMgzvnI
Ddr1mhuVUI3TM+xV/JiW9icAnoT+1qb7fyXbCO/brpH3cLQTthmNDLO3dfegpUcI
qYeViy6k4GNjx0DBAhjtVVa+N9JmIm4KPw24+Vf0vueVS6BL9bk0d6V4P56IT1tA
tHYWyziX23Ei47IqZcMNXH3naCmO5uWtq36C1tWTI0ODFY7aqHOkoBq0UcDFPgIA
xzJ4dPOl1N697nUPPbE2hdbMP5TRdHz4AuR/A0leP+CrmUcXrdT5Tf+gsKZ6gXNz
roZ8YgepyaCrhhP7S74FtksoxljBwpVohIR3ch790H3LT9Zk8hhq38kVHYfICP6Q
hIQ9SEpZZVm0XrnNxVS5iYohZB8abJe6+6Wl3yDCjBP6l51bFVquKZyqw6CrZEXr
WCXfz2Y3V1NT1uL5gK+8lFkrEn2KWT2UIiYX7Ztth0iewcB72tGMhh9cJmnjg2n/
9he4YCOnGIGDjJ8QLxT1S8MlVE5qbnQr4hwij4jpEb5oq49Bol8f29yLlt3yS6oQ
xuiVqs4bnoRJ9jUbkVhdV19YiT8c8Ql/FLcCAmV7/7CXJnBJePa1lOivU/j9g057
NJ0A8NfmVExGHWz4Di8Z9Nktrcs60Y9+jZDdQq1OBq+ii+JGf1nvnI6RfloZZEoJ
taxavns4lUm3oSXMmPb4GhyFAwqcUvrUORAol/IXqjWHScYZv4Fwqg0ltwnW44Ey
/9f/qWyCBsX4ZAV8YxSFbjAvu02dwBr/ZHIIFMEfMeJdKwCWjhHueHvJXvUgukLS
kzl71pOdQMcJATxnfCPmYBd/m3KDEgMlHYxaz23zRYAEre+0pw9qqDA+CfrRQ+Wt
3XSk7QcVBMvaC021pVseHS3er5n/d6IO8zhpAP8CKEPCA14MuqNj5wlsGEJeHAQT
lyPRcOm8Ov/iU3PbtfvyRx7oxjPbxXkORX8FA4eTH79ADLjL7owckzmj18VdQ/9I
wb9+3nIa/wbmItPHwBq0Fab6LYgBhG2OtFAW0vfj9/nFEcQBENPidQYKjolva2iI
FKqRsbcnG3CcXbVF210/lWuSvyEJTZdHmRS1sDeen/fwUIR3liJVVPsRn4/SBa6V
vP9/v+U1iMtr6pxc3Bl0Pa5Wm8eMzPoUJ1/Nar64dhra232bGUxItb6UaWytVXas
3SfYy5511PcaUHJ+bX/VjobO1Kd/ZejwqfVhdkN+1Qb0/H5pI5MO8m844bZML3pk
agBUKbAIfuebvsSmrD7WlMqsw+aruW1VawvF0v/6HpRlDmKv1MF+dZPjZY4LFIUU
Dp3+d9wykkHwrw2jlkvuOzrqdfpWZPVJm6KZ9iElHdtqf6w9DRJGOdKboSRM6n1L
nlL1STpXMxntrbz4LpTizepwk7sTofvJnHCuIzeIrmHfh4If2cjeVDW+aP6Psu3g
ttb/VtVTMoidGhp5e1V1mve6eqSP4DCINao5D5b9+x0MX37AItzZSrWcoClqi8hC
ZB8458XRS7fSvs4QGoK0Cqoo8ENc1JRv+ZeY7UIjKNLEz0ImJi4yeOk22rsxwSnu
W+crwIrNqmMuYbWHmsYWPOs+mPKoo5O1a3jRwv6pruljrKESQnMbma03jLH8/hci
AuDTpnt+HBKEzTl4TzOBnU6jsUl2IgmqYVbTDKXrs03pNb8ETC2VVHGGRmp5m96g
BGpeVEkHKc9sY2J2hjbUU9pBO47GBZPSVHuhOsxTsVTpZCUuJbIE9pTbf1l+91KM
OqavAcpBKg+cD0WMvbo3wI1LRGbVSXdRGo09Vo2MeBinWd92q2clnFQNgVk46+z3
BGFTDeH+gLhb1TlS8FgT+olzRl3/fb7lg06HTIdEnQaFoJGSbUnFG70YBoVHPIWP
htgwf3TTOqPrWYS9sT7wNAar53w4d2uc5+13a2XB6fhvpvBT6OygyT5p7b3YVmnO
iJTLtw2IKP1dwFqzrZ+rYbYNow1tAQ8JjM3wX6Kpl5UdhaWDsTl1IgEQgk+A42BC
9wnpQ6dqoFiQAGGvR+enotlK6w3iAioJaySc+eWNtyjg5wZfZKoAjON1/GXoLfxl
3HoDPmPZsAA9LHQvFuLUc4JVk/dH7GfpvHv32r7ziN4FM209I48BH2Al4rjJWc5J
8pjsfEKjpprz2kVp5MvGOn8GHocF0bGXRSYe3FRmnCwUYKU3gVI/Vf7gNF6mffGl
ke4RafEKFQmQuEjF1rSRStv0ZIQBsRmcy6aKr9HI8bKlOKvJ2UlgxN2J8ce6cfQi
ZCJlyvGvS4MZKv8bgYx/eTF8W1Zuw9LTOEdieWOd5GDYoqnx9f2/9/40HUUtTdoX
ihOrKrv8iR97CnLiOoxWMDp/FBvWyqXIVss5cJX5pRf4/pzTzkMDDn2Ys8l1S2aj
Nen5S+HobBfU03nNMz4zpYR/GpiOl+8KjnQRiKZwmvuBt+dPNA46EUQL3hDT1nYe
Nlcf0EZqen6F+3gS/6erYVIi4rKF+q2SoMV/igQtjP/6TeukvRpJ5ecEVQPq//XN
jMIjGbBz5goAYlKrCOHKjFygiRwJHavW5sIiVmamyOPEBYpRmg3JGnyu9eMfJjVL
QXrkWtMYqm+XOzKNQZPfOeeONgvqOYnUXggoXVeBSRZbHza1WytFSaMIOpGVkTC8
bV5LzGYTpmmxc/0wsJopZtnMtyNIINAEX6dQIRMwHCzIt9e8/CH7U/sQi+0AMzHp
sfD3AJxAnghznQ7NAq0dbHsdCursk7DnhCD8Ayap9DvAK+eAPVPVG9bpOhwy5dFc
xo5xQL1NNcdV0rCXjv4TJvATA15YMyGMJq00ulVwyW/kMIqqcyZia3A8abmmXHHg
ZQtZPIZ4Kk4iFWEa1iDcf7HEA0AgnYZvS4vUHfeLipADIFEFfAF8djdt0Q0FO0wq
yed24FE02eDv07gDWWj3LjRRDRCL5wD5DsNypf7KHvp7pmZWZYcHgj2EXk/NPnPY
dB1KSyNQkCHK4XrR/SA6rFluo172UaLe4l8AgXxx+5+uuWjAIK6oQhSzwmcyfPja
oR/mCREfcIutBIoxTyTgRb7LalHlYxXLhMdblylzInE7VWGMwK1FfDTcKsY637ki
rUkFyAkMKotho+1RqRqFwz9V9zlCg3ufCu0uXNil0jDIWMQw5Bx7xgbGedWVOC8Q
NPnSQy3BiA2N+ye9DkPTQs4bHmQZxtJ57zHpMHINCERRGMIEmIKaipT7opXOHKVH
dMGHhem3L/mrq4JfqxfN97Yq7qqWqKbnN/4RRd5JR86ZuGZU3v0gC7DDz7uCLaL+
OrkmEUTkOIQFG5sS2aLhQJRWYJzm6fYbK47lA/A5H5/hGKVX8n5C8lFMsqEwzFXu
6IyigOBqOnoPI3pu7CgtdYsJthIt3eMHEpcdnLxz0a3cWVTG3h5/6g8WMUsmH/kK
mzhjMzpiRofILVKXCScYk0BsL8dWD+377nNRS6/USBQWISwD3VNmrytTaRduJFMc
PyjhFM1PSuhZlNx7TXhHuyn5zgnfjXXmrP1CcUo7Px9nZMn4+rmXfncFHnQwsAti
coJ3Z9/md6BFR+xY3QviZC+ljaRndtJSgXIGSfqcXfUOZOzWkdPYcqbYdNaMA06v
1vpL0RcEYKsRbnqWZTGXz+bSsRi4Oo3otAztvo0HWO2K4l17/+lqXLOzAAsDCAD+
DucIYN+rUFzeXfuO4SJgH7YTHk4N4xx8SXsLmF8wqEkW2iKmp1ZcT7SpCehEd+N6
lXsKTctYUWYgGlxoCqOEq0+aS7cVPMhWY82eFuyHWii/ukux3m73vu5athAAu5o3
Fc+xZJKYtfUeY6flhF9lJLJ2RRyDX0rBQA0V4uxC2bxYg4dWPc7HJvWrS/X1GKPE
HaFe0OgumxA5DDUPmizF/q3q/B0XALUVGFlDFnDAtZqIABzWcSg/IsqWSyDpo37o
ar8lAQ1FW3tj8tE1yDcrJ1egQvPTDfPca9irlVgakH4IK9Gt2WBAA1bPFX+9TXtg
Mv7PNXAKoflA3SVE3AsKpPh26U0uBG2/lmzbQ5NPBb2+OPcYsrD8eb5pRjQgcic+
qR7wSJ7HOgHaiAege/Dt5cFkIrTq9P5qaczQssy0q7xySszO13HCMrarJQVj7tkq
oeCbZSw3c1XjZZuk1bkHs8Z7J1NL4omDmBUNW5kK7fGF/04ofKTIceCMmAEAlMsa
QzcCpQMCCnPw7z6iLfdxCuzj5n0acgZW2X8amz7NXzQKymrC6HhQzEIk1W+J/Eg7
ZwOQELzJaWo7ZnrMjTHAKHZK9BxLEvrf4z0rT9p97DXyL1z7T0f60eMzO8M6ljrm
sq9s31b59C2mNQAauwrCNXD9a2gAOrDalYoIwkQ1RMAywK9Atw7huDvQWLrVz1+X
HvlDbAOowaZU5cwbUd3LwhrvCast7srG+tc6PB6o6ij3cKvIz3iKgj3UJH4zapOa
rTH64ooY4S6PRvHWymnpJpXWpPlWylc9ZbeqdG/9Emk1laFtqeWYMLa590ilt8A5
Ewk0nGd8m+O+3X7YGa39zyQJwFluRpNe6Q0ZfNC9QMk6vTohdki1/hQaOLqqmyuQ
PM0qlXp0zJEE+ppbicKIZKL9zSK7rqbMs/pDxVkqwQqZj3UIPGChUTz4tV8D1D7g
+8M5VEJjb+52MTrkywaSFF+vkYCudfVCNa5E6Me3ZBWzeFgS9WCP4yGZtTKDHRTa
YRIJbCCbl3ojlIDDIi+BlmomCRDTm+6A7XF+TM3uviEcYy/2juHJrk/1natvevz9
BVmjpwEriQB9ibZHHSE/EVgZyVlhnCvwfqkjW3545e+t5f9ZeKLiEB5qLE5jGCUv
WRyA1dzdICsY2EqSqvCfVgNWR2BbJtofNbq4o6MDwjeslM4PdLg3ZWSRCrZkGASN
UWwPiCSZB156vVEB91x3H1g+2pWzNxgBjHwH3Q0+wxlMetmdg6j1hkfsD77ggsOG
/wLUyCvFwdThrFAfOO4fhbRtZEK0PACz0t/aluGbCWaQQp/vJMmc2/v92uA6nSev
Cf576B1KHlB9shJ8CGNcH0k8gyGbSUQ8EFnKbMbRBgwJ3nIZY8fxRzG4OS1RznyX
c56zDbJHSWvt+Q6d/8EX2A8bnpIBLV4kF7ZDl1KHM7tkRMvePap8gaYjpOauWrIV
Xvkkka7V3v3kZmmExdlbBzRJYix6dMZ8GHcD7lDHD7eDjB/3s/oh6hEBmkeCC3CY
XayAkut596J9/sP84yEoFMYLqcTQx+j8Gm67YVAaQn1qxWCJjUTc60EgwnYxSXqO
u7klI1Jf3lgWC+mp2SXKooqInZgaB2FeLOaUytwGC9Qf6Jaea9HWtoIrQG014nEr
xGt1F5cIVGsMNyQUB71CNpXM8STbeNf5NqaOc8mHBrKVLiyy3ypP9OFSyHEiZzo5
zCId/ebDDgh6mXe9eM6Hh2O216Zy1AXYqGwKWhkNS/acct9zdArYj+TKD22YecE1
aU0bxrwGaFzCiF6RWNpsbwuPQyZjHpNIpqVxxfvwqf65Vx+qC7Y6N70HvXisvDTk
G0IPNoHNj+6LMLF4mVekszAUJi8XQTjzjuMw5jTpB8LgM6wFHQSfE+eGeU1WhpBA
8QlivEK1fhwleX0dfdpV48IK2Mh6C/Z8Q1Dysz8q4iNw4wUII25PaaXkzjFCmV+i
1uFzV1TGlyQkYeG5iXERVOt2RXugSWt7N6NHA2TWE5CMdDHTqwBNbvCM1IP9uAIR
/TDPLwG5ziHWakmGGQsDRQQWaBLbhpIG7/AYDBH+wuG0T0NLcFgFGZ3HPPa4ZQiz
jHI8soSAhOExE/4ZP5e6wPn7FGHHuamgnCKqGc5pOp/3R6nP6Y5nBSLrGVcXxe/W
ZIda/XHQcnQvbgqjGqN5yD8wfBB19O3plQz9WOocp45j8vXXJIL73Ip5u68McAqg
bxoJCdtPZ/bUGxreBM4J8bU0OMYP+bkhTYvh5DJGIvZqrhzbJxck6ohJlkOMVeHF
/rhTfdsjL6G9P2c0NfNs3QkzhoFYRMZbhsXyWYN5Bocsn9caZkWXafXK75yGYlEf
w+qFswYFSWOSfgWLlpFdbv5y89NKe+VbiwWRXzVLNGsAuqOE24A2AZuiViICn9xx
RKsjMw5D/c5hJw/08yYBZDR9zKFHzEbB34hBTvwY4bb+HLHCM1axEK9e7eVD5rPz
fHyChawAk15AfcJQOYia+ZDjYpsuAd1GwWf1mS3HOYigwZ/y8hjEf+5cuahBcID8
f/kNUydhvBmnV1FxLvo4NpXWRQptIr8cAUPOnqxu5P/NT54isBAEOs+4voYj3KLz
CdTisgCBmhtXAazI5wlGjgjnfJqXFxTeXgqwekAhuXAJDurMxNuT/RASM4VtvCZ7
uj83/lM60Lq+/tx3oyOQcm9hQv4hLwPZMr+6gTtVQmR4oUCpyOOqdOe62/A2LKkR
Dfs8HYjZ00RhbF0hT0Ef724/xmDssSwZO6qZC7pm0hPNT9QeBelwuDKR89dOz7/H
ylTZmHTJacMTrL9rMpvvYrmwDaW94uWdjal4HtHNIbZdZGc4RLsv98HhFsjotew5
/U7qPTU1i/T5b0tgHSxVWQbmZd0ou0tgtzRusFZkbb0zb3oIQ/iIXa8y+IHEGWRw
1hZPB44nSJAWkAApVIY4Q6UOQiJfQJgAk8hKj5+wUM+GdQ5oa4v/iAc2CkVoBjH6
dQb7ZYOAh+IIa1oVoxHBKezOxrGUniQbw3sY6Lh/K0IE2v7iYoQLx+zkWBohdB4s
KGloBmbiYMm7U8fiVeb/lVek7YjYJ0lel6lqPmGXFco34ijYn9XJffDnSyb5vU3a
LNJADRoKq9E5kamcrk1Rrk6OUbB+RJL3kSc4dA/62mGnJmx/0O79+E6FC1z3U0nX
2iLjnhEQUbHymn4myJqCrxpfWdR6ZrUuKhh5cuaf2dbEFseRM7r+0m+G6IJlkse0
SQey0DpNlyirxRLC3Jz5YbksFz4ckfmhEaYvjG/YPPxR+8uaugL65i9Co0ttz563
R72KZ30N4tNdT7jb6X40NEML6xrsXrxhCJrrS4SYt23/jUFrNf+4a9w8QkK4U3yi
7Ja6+Bwbow7v25NGIJR68jvRhFT2Omh9Rk81tE5VwV0jsDvgZgAl3nNCZDGXSfS2
d96rHyMYtDucSkUig3jCZ0Ct3N4S+OHRUbVnqFKVZtHvrmWWj3ROFPHpX5tphZ28
CjBrkCNS5ePncIW5g/EbNOKYHv8qzaovUZEt6bgM/pHEfaoj87dXA8qoUapjVtCI
CClX3d5L2dYkNdmnhcYhl/hJVIQ4eo0y06ZK95mfYNl5W08ye48/nLUxiAEo7c86
RpVEyQXVwefrDZ9RQky1EGrUZl4CPOm1BO111us8XU/zb3Fhr6WMLB4Bf4uOgtqT
+CJgHutbzL2GkS6KtT4tgFqStU/ke9SBQawcRBTsRKMBm4Q/T8oU8Q8e1zfks1bI
QJPlwpBwc23QkDiA4+F2SOPOvu89iXdSMSithpoe+iAd8P3TAwD7So9Nb4wSXAHm
P3fr9Q5b3a5FfauYG9prI7ouSqjBtDo9xDzGvyERwlFT8ocO30ZCG+2keAm/URU0
w6yQUsbG12CUoOLgaO8FH+7MuzX77ok2GRbrNVQOzIvKgrbzXALfUf2HvoRt4DJU
GQvgG1xs9PrCL52QgLwpRXmYUNEntggNy/S4aL+u56JYOmhW59FUqMI5vn/2xZGM
Gi9DOd1e5Nz4KwZXO1lrnpn9lrC5Fa8Br+mDsSjRe/WItMB7wEIxYYWi1CWhHpGQ
IySDYG4GpDvg9Emz57iZlr2/nlUvZSONvM3TPSp3Oxey6s1KeGEbIDsw/jSc/vCJ
5yGFl0uv4ZttuNLeckaw9u4WccYrnvaJoFFbmXBePJB5gyXDVC7uM8eekQblv5jn
PMtCX+M+p1TLML5z94eStr8c8Dl/E07X+9ZiVTIrcuB1sC9YUoP0Kou9VETdAdfS
3pxpqlOkAMOy/bP7JRn5QfZ9UdQrDmG48QnaOFtcYJOA9rnpuUo8EfRMby+VkWdd
N5blBRPp/J/fZU8tk/zzw/MyqC4wmOF8dwJay94tNHi5mvWNOVcowiwmaaBf6lV0
APmy7xi01bvI8uiff0WvXvcHESaiqxdN2F4GuAbOJcW6VmA2piNyGtsKX0VwLXY4
Fr7QGHRpvxEyObay6kCB2Tqnrrx41+Lm/peN8SZWGsU5mzy1yZLbnpwafBUaoIhW
bWhm9ltH6E7GvhK3DYyRldsP6pemG4Z+CClkwcQF1+rBGg5KkGtxVWyZj4xdJ3Yo
6Mwsv7Z5LuuAngx5OLxvhkdgeYtLTzGmK6uqxARPoiMF4HEY01LrSUvzYZf0rkE4
q4W4drqyyxRwyt2MAy932NSujc9xvj/ScMPz9ZaDy16lAQwFI/NBJ49wQMuDNbeY
6qCMbLo5LC1u+EQiFWNXBb6jbrE01+NyDn/kfg0/HgmDzLlXDZaGHxC4ql8dmfDs
UCv893n0FIhrivF9IR0kgzNPf4YVyFBJUYkrK7agRPMY4GPIRpMhwh/JHrCZN/Mi
3fb9+rFYxipyC3+kYevkHveEQlpW165Z6VBO6uhdoNGNdIJI/CDA66tSj3JjJfCj
a5bgW7+RsiCRhpd6vRovFGJ/lZj1HX/e1jUQ0C9wyzLSYhCDljNhFCTdLLxWybfm
2UEw6Glr1oYJ6X5XND+bUWsHox9nqZ1CZ49xaSmbixiZGUfCy0uq5bnRAA4z4NQg
t7zQ1sIZF74LluMOhe8K4u362HF1R3QDlxBkm2KNOssQ47rPUKa0Zga5Sneq5MxW
3wuQq5sZ/mb8pDPvBqi47Q2n5rhMjg8HyU1HUdmbXmdSDNnZxFbLTMKY2baB7g1w
fu9i1JSEBesGHgg8p/JkxbpXQvS2ohP0ul4L/0wQig2/sVjNT+9f78/JUnkWin1l
pe8u/M0tx6nXUJPXwg1Jkp/ymaq7vVCejAh3xyQ1qgsQIYvmfI6xEJyTiAsNZ8+d
WoPKnGhl9FSt4lCnCm1wREFCADhMNaPraC+IxRgK0+nibbrQ0szuviuXer87G+1n
azhm+CdlIJZSUiLCg48TmuLG5ujNHVm5G5K//9/va7jsZjSzk7+obpI3zlhC9HGz
ocR1haerobLrJRGAceaLW4c9BDzp9lcZN569FCdh44MN2+8NR/c/ww4DSRBhytcu
FiJki7bhTJEpNeVR2Thfg57lWaWrq/Vh1HVBgVyPj5gVjtgVQP8QrR7vMWcftRM9
bjq7ZjPCqJ5mYiLdYdNYxiyGNSRJJ9YNEOQTCZbXJn53EehHV08T6iJoRy3aDQCp
YD7Pk79rIl7RX4erpfSJKH0nPKYwXemSEhaIc23ArLsSwig88mNR9RFgxGhVs4j0
r/95I/p+mzVPA7/Xc+fOfVzgGZfq17708mkjAEYU4ZCk/Li4WN7hnhyGTXY3qKmd
cPTVbagtjtj+5Io2hVKd59HAzLx0xsZvJBXDL9Gyia3OxFImJ5lB+XceUVP9UA33
wUag+Zx10TeF0n6UjRTD8gRtc+eQ4YJlDnXMSyEKR2x/Xu9MB4LDyFxzlsZhSD0l
SUJyAlA1mEs7tol7zFm6cPgcWEYtwWEgbRlgDmyNvo8RK3IXcNSMHY67rTFDQqs4
8qSxpIQQk6L04oXUKGuOGtDvl4EL0jbb1BBf0du92d2r7/UZRXlAhNur71/Ft0QM
Py4Zxi3pDP3UclVvAfY0d9/QpxItJxQZK4ElOg3FJxRYOnJRvVwdV/ZOr1MnhGbf
W5yxN/Oc70xXmTfVD05H+IeN94+xp60mto27gEg0G/FZW1DHqH2H/r74orjXQa1C
O/7auTDoXWCTLv707sQVdMMlAzGLhL2pb+KCG6eJUQffQhvzqyS/7jD2XJN6vJS7
uvSuLltWhbX/KGBrtvxVITn8cxk4gPSkM+YEYpmvHgjARmjA/yxF3d6DjMZqGRTN
Fkzbt6cYaQp6eNRvnllgSOrgNXtPVMGCzo6djSsJJOusG9gh48nkLb5yTBVZfYyz
tBdxCcCGi0nddx1MMDzRevd6cMfR3Yc448E6EeGo1HCetHcFakQaEnp/u41Kk64a
XFwNpgOtTMjTRk98OOdq9tS4rjC6HVZkxkwA+9VVXoAOg0GkoFXBEMnnz7xljYGB
K8E7nBn4mDzjRgDjOz9HwFxk5IUfBR+VfoD13rupN77/7WoA6AXAU9vJBZMtBfAj
A0gLptwr05WZFavXvcgvZwEN7U6J89keOaBB9FYadShTEIQHdyvJJPUsrMF7YN3w
4ntHHARDyO3oniZHD9D+k0u2arnpnAL2JCg+VgpgQ2t0KT94FRcIxK9oLSBf9xtL
ZVsh8wCsly+7Q2iw2hbQB57JhN9/H3P0a1LgIwk1r9ajzhwGSt+h8EgK4fyww6lA
iYxehZ9d4J3roXxVNwvHs67WLHvHdKanZ3Ymp06UKFHvZ/G42wTIs20vv5eNSdU+
40yAyNv4Z7B9HVNlvEOP53Eo5qHIKoDuaSq64lledn6GRnsxs4R+dzNGBWX5RQs1
LnzU1HenLGHgkBXtm+RAiT0wGbZMlmInxwyNahD51MaqUsgE78qgCCdlYsZwyjWc
dV6htt3p2H0JXbaqMZvFJSOxj4GU7aFn3zuoi64LaEOVpRcJ0q8gMHB3yRfXECLc
WMIF1eNZyfMlTAKG3vUn2C6h2VDTFI/PicFHf5934AhS2AJcsFId2sy4ZNELdXl5
PaLSVqPqIWdYLiK3gXjibsSs581Kw4DNPEYrrdTm5lFl1jcStnJgM+rT3D9BX1LP
Hz0rXpzPDGxvp5EYHa4c3ompp5SPZMMX0ImlDpCokXDLVnBNU591ArsPrlbYErjB
ba2z8nGC7fbs8W83wdm1HM7sS5mJReZ0GEtfay4dVWXYfyMsWErIOgD3dmLn+VtH
uf04ZwAbrj5RrCBUKdMPq6yXgxBSotNVeMDZMKoUL6+Vi/p15ke5ERoiWXIWvKCa
N6n6r+8cIPCWPEb2M0qMk9NF72RLy3fc/nhy2GriUCFZcNCFAoO30257DGj641zX
kbgAY40WObx6wQD98SR3hjt6zHZpk71myK3l3sUVXqNKTI2WSboHr8rddTob790P
P11iIe5zHMJm5xC703QzI5qVaoNGzweW769H8uNNc6qejK27RHjZ8GXU5wQPORmo
2qBeDNiyRIBSkIxRJq+AltUsiwgO5Iz0GPakp6FhFxaH3y5acoc4zjp9oG5J45xl
JZU+QtGz1bhe0lUfwMRu9QId0bf7VTvBTS1rEggXhDxh66NhAPhSs0bWbVoS9O8F
+VQul6XVxGhn1IWem9eRepHZH1oXgR9mwzl/Dj5UDZsvyZaMWMiTJsA1/0RklHx1
OkImAGh9UEBTEpLN4lbnBpR2EaqcT4MNcodTrD/1qempOX9Ah760sLosS/S1gogz
cUNprKO30CRN+hooAgNPd/0P7UDd4pX1gaRK8AbNOUIirHEy+KZapbsDo0W0zHz4
mrKUH3Q0y0hmZnQFYbQgjqlQrKbJBzqhSLQdHYZAye0FpbL8SaqC6T4wE36MVEBC
Qe38lasyBsFvi09nd0wnmWEW8DJTJ6oDZoOa1L7FxP65mVulaUjP14jeX4cNP3XU
umuGxI6pjTW3OO6UweFpAcym/EeaFNCewVeFurjKh1F53o332l2NK1X8aEWnO2Ew
tDeKhGShkozFQ1gz7t4u/BnCAIh0f7wkd7rpocXTLh3MuXRJGU2t71LQ+gA4UJgD
TEOY0voW/r2HwR5ZrxHra0p/9xUOslULm3rn4NKwKMXr2THQuFYkHDwPSwf3FyFP
R83uZYYxqiQzrUQ03335HvZbUVZv21kDV3Q+5wAdkV8mm5fuK0gfD5stuiBuQqwZ
Upqx/taYZdt7qTB7/RwB/a8jUy0tVQMrBt/kS2I5gf71Jy+DNwTUI4ycw3lTgOhG
oXPtON7qgMWdy89hQr7BdbVa+F0mNCFUAcNoZBiq1JK3TBfAkPLPJeW7++8psjNH
rXBRBASmP8s2u8GB2l11fYtL0VFGBXQrZBpybIhBljrxnAA8qW2wIWcdH39cqJem
w3TK9rVfUMuK1yWDwmpGSOd1SUDdLSs98naHo24H2gXOuoqzdq73Rr7Fu/EIkvAW
/vqYKu1onE2+MEimFSg5f5TBkNQECCAq7fJYOlVVF6EwcCt9ZvQmVfoZRazq40PE
S/sz+vBeyPDYnsdhW4xcGWkB/JG7dW2JQADZGsMFe5iDX3sqYmsSgjYsgeF+TT0G
bDUQRVbD4QcJ6gUB1/uzNBPKJ3rplXY03s7zK3H62ejB7AsKOddZIS79vEHT1rkT
0NuYK7wlXz3q4dwHAV4apKByAINDjDd2E+99dSYP9CSGtzVU7oRvELp6clIIpp11
i02JtafDl1HjCTK6sjWrCoHfqfu5A5p4C/SEVEk/6YkxrxPq18zUHohcIZH1SBvo
dbGGAyLJOQ9iJ0XQc656JRT6Jvdc3lzqB0pmQefD1tJTBYG2jFQkxCL+65KAArQ4
K8z8LQ9BfUSg1QoitronIV1yHyeQ74h6CxAUAGk+f9HS3XvnRbaMUzxOy2gDJT1r
mVdqlc0svmr9omuaBluyibXvuLRikhx938cpoawaqsNz3+vFI1n4TFLF8LrJEHqn
5diN27AOVBn6upHftGye31726qTBB+GjHo4QNS7tcoa7Pc4z/JpWGNkGxvAvxrTo
YRpkaXUnX2CUb77YccVxd48QbTV5pzqOWrMKDm5Wy+WT+KTSfX6AQYyGCOGKIgkU
pTkns2cdCH0ri3lhjrZdY/DJmz4bX79NSNiyXIT7EDZTfVZTIrxqM1TbyjiVYOD5
TKWAQkqTKSD/nh8FNOMOLrZ50g+i/SE1E/bfWn/1ih+zxce0BBcPtUMYYWngI5gr
D3Ky4r8cT8m2/+OpYhcwmGOdhNz0lboCJ6qw9FwXR9ZeTCIhso2bnqaBMndsBfS+
ctMtXch17euW2wOXdkDaumXGBhyB9MNjlveXK/rlpOQg1Ghq6/1qE3RMG7jx7Kyn
rLU3CmSl5J6ZXDXcCIXTkwHHUAJqNeFM42Sj1rPfpEYJZ/DesXX0g//pmRguO5PI
kJh0POeBdLbSjxRPzQX862uUCalYe0e9AenMQbSNUJtSgFUX5JJekCgWd46gqYiD
lR4QFCsDPN7vnyIgs+fOfIgb3NDDatpIJTSJtXcrKAWNOk4qVMRpja01Pd73d0tb
sOeYESyLk7hmZwsne/H/GsluthBVvJT9HtmtjAJeBviCdlj8FThHfyqmNSdr9ECg
Hr+ldV85DzAsSzYNz8TCCmrKHrzsKreEV8sn5ReAsirvL5yPt+0ppg0QWqtEbWfW
qC+o2jcESPPLrmQsSXb+C9zwmfAB8r2CmT66u2wFGoB+0sEY5HI6Y6yd6QepNkRc
na5nLLrH3Af7TX87A/2cfWK9E11v3Dhd1qKIn4GskFHULNdZ8oga+SVe68kh9VrF
TiJCXcFKnFuoqSm4hnDIAjsb+QPqLGchHfYY5Z3q7Yg6tJ8smKhlpL0CKlbnKpaz
85UzojE7lGlzeOEc7g+xYcpMiHT9Agia0m9ttThQHv0A8RSyvMsuZQNu6AFF92yd
oZqKYw4JfoOw5AdbjcEmQURxqzBK+c7kT6Bs/U6a4cgsRVUv2fKrrIfbywkTVDED
Qsxhox+Xe3bmAr7iLIbhyODyl1nOcNdKz2Q0mBMYSk6MYdjLR711mg2qlZ0D01e+
7VanRj0nPsJ80e52aImIk0x+ryPnlQwIe0DmiytDFgh82Dj13LXimqxxNwe2RkJB
Irox92vi4Q4ejiJl0miBHn0kEKQUUZ9pxphmJcrMvijVVduBPppx/v4q4STwgti/
n73Tlt7U0gN1W7+YouQUicyUZ47aSIiRP7MBEKELhO/mfIH7GmKEnUJN6UhOsEyw
QTGr6pH6HcBi/1YDVNThsIn1DAnZbvSAFphGAVuyWR4PTfT8MJotYkpHn8+uVNct
fs6/xlV1J9iJX9Xoz/isH/rDvfNtK1LalUsLqbB4+X5858TeBRbRztQDxkM9yUoo
wQ3VS2zg3nIpBbh1KVfwwG61EHO4zTaf4Km0hIs6AFYXHw25/bK/s5dPm/cTBayb
9P4Q9HFiq/RYepyNH7esrHknregV/SKyXXmLLyv3yP2MQFMNAkaErg1duLkOSZQt
HXp3gwaCWq5QjqNwGF1zpebRPB+FoUhY4ZNEdI7SzhPvP22BUliUoy3EhmZmYHDJ
DdbSZ/Ip+ivE1vq6J9++pEkmB96MbO/u4QlWYXcOib4+Utlu42OOREyohv0jxaJ0
ulZkMzaMgu4yaqZSmllPJdQQ1qmBcWfGLLg46j0+UbdjU2RKpW8YjpGPigDcwxfY
YDcnPpIhRb4/nwGA7LeiTWAvt8V0NLkIGskW1lwHb7G/2Ytf3y/0KTY/tO9nOeNA
UXZGodUGmTFK3v7z4bPyIE4RZFytHYMm0Bf/p4tXxSJQBOYUXBml6WorF4Uah1D8
82TIlzjSNv4XIqAc2WP8lJxNt7MFp1FfVCRnUqhM6CQeJt1S49RWByjtnXl0R9gp
qArmiUu7VN6zzojjGdeQaCS9/4U2G4ld3F96VqZxsFu9r1HYESvW2mH7JCFgFyUr
fgBv0CnIvoumochD6rS3okeYl1fbNNEVFefbQm2reeMmkvbo2oYSgJVx5Pr59uk+
cdNvmPo2gkW5HvF+39lteWwx4ZLEEYb8D74V0m0X7SzdMCfptsWwAFiQ10H2mMLl
f+envbLq9Y9NJ7DxcrOEzKuNVWdxxw06fh8oRMV8cReDxxLKuxSXIWiJNpU7OcZ6
dyD76qVYGMp+mMkrKcNhvtEGM1WwhAeOtlLwq+9CPpKI7ccOv+KZegB/F/VpJdgr
n1/Hh8zpfwF5Wt3AQAsv72bvhyPuWfskOGOzIfTHYO941EPRnmqUujU6KNEz6AOc
MVLU/OuVfsy+6ugzAfzMhVR/nYkbKx9uh6ZJay2vXViGxd1rivMwOw5INzb8DpKN
IDXKDU9UiYiBr2AoCHWjY4Cdexu1q921ms8L+6bXksaF0AYZ+7nkDIfUivtnkzqa
Qke5gN/gPhvGwDDpwQJsXIseuyVeGNGwu3trPbCyGi+PPhb3G1PBVgNjN5O7C4o3
PJKsXQ3uoSaDW9wcP85JC3pCGaiHfoL03OmPHjqAz5tJALaW2OzjATnLJbngqdYE
rVqxwmSFxBrAFFOJLuPGeGUjZ3YGDJbttW993lHezWZVOVuwvTHxjGI9ehOJTr8X
jzTmFkjc2nnaTk4YZODPB0oTks3qbEpdY+5y7V8O4bkk19O2L7TTzTLr8IwkFEze
m2ETMQ3mTOs0NEgymUPnw8m9jG5hVl9gnNrfeYaAhqx+7ekVBL19WLMUtf4F724F
EuvT3Ve1UauJfRm5GAjQF+IKCuTgPxAobEIN2w52F/DmI/2exXxxCHIHWyQS4UCM
Z2K+1Cl21qKSTdEzJ+Iz2Sjn8mRfGo6Q1b8m6NthQQhsGBFZojCx1EPVKalFbUtE
X0puHDTE52ZCGBB4H8gmVJ5s8HAocUvI6+nldhcGFn/pq8ZJWTeAvTw2Z/fFxG9z
U6DzZiRcJ+tVyL130MJvjoTlh/By+PEDycGu462CaJqA3hVcs1psnOLk3aK9LeWU
9sX7RYoD2xKEuY+SzEoCxizuMmHT4bq1ngrkn4qSS4qMru33mTJ/xsBJ3PG0S47v
wNp+25nJ0sbopJ3xpj5e7K9KCIpI9Y4HyIdTN0oz81TM1ezu4mqOkhXVcYfa3QYX
+DtrDSXq8OLt2XhpC8/e1S3DzjF05cudhFKDhsfN0RtY2OxS7aUWwM7S66rANMvE
t+ZWBwoS33+agRd3XBvfxxEaxhc6DSJxKiKBw1e72h5fuQEMLd8B5DPrfvSe2gi2
bZKiV/8PfQUMffpwkl3ReGLhe4CprnD+/5aShJ4dzsZTBBpJiDfdUHC9kHFKOdlP
xG6pbsx8vDapHMTRPUkvXbRhLbjqkEvFO3ba0qkWtaofbGFb0sHXdWaSqsNg3GDT
e7pJ4JU6MniyLZPYXlBq3tMyhzi/P0qHO7bOzCa05rf2jv7rUnKEJqE65pQy1InV
9U9uKZZC0ZB8W6ii3u8u2A2f1n7gepT/MPMFs4XAW/EbfLF45poE/rAiGzPKQgT5
TW5CfWVxJbJ/ZTZ1wZQtNATWgliLIDdSZfMNAy0KxCPulYO2KBiDdJXfBxINF/l8
BOeD00eGtnnwV56rM80SGEfFbfVcMyCVesba8UmdubTjpQBe7zC71B93Kf/RnKJM
FQEE08SnoB7UiXHlrZXai22tTg6osxk5fABn+n1BKPc1w3ENnOYp8YhFKkHXMOJs
+usTXOK7L9sobxLDHeiFizhLTlxC5X9N4yyFCfD76jyw1rorEwTppJPrWTNdJkrT
VohVEV2v/b2Q1OC52bSHoO1m+pdvIk/PTpwIEzxEJtzQg+oTxejsz9AGqOsG52v+
BCrFoYnX8LTSjJGR9soxj+63Dqh9QuQRM4+romQWIV4PKCeiWSHIhJGV+F6oghWO
78k1+hlIKhmfieS60NLiMlpkdr+6vnVRd+5vNK596aWrttmM+7lSzyTVZAL6h136
6jQtefO9zVVF9JOYbatH0tHhyU/hhCq5o/1A1UtZ3EMMczKa26yMPMvxX+MA72Qc
GroXkGCc+6kqsnDSUFv0S1QCjb9C1NBR32I/v33z0h/L8y26CNjefFgDnABADD7x
Giur0i4EmHJqa35hdN37Dbzd60hgUhnZeE7mtraaEU+T0Dd+bBPaHRVEicqBA1hu
89ipt/CBN/TVYqw1s1Q/2nBEe7oK1F8XYcHj/+xvL3PtFLkWPIsDAHNmYGE0fbSP
vBaWE/C4LPVOp7eA7XBX4WN15+X8H7Hs0ERrz0SDuWPvXxvKzb24cOXzmjebfWw+
lHYBz/op0SnYz8UnOIvizc8V5v2P8OXaYuUzQ3GEdl5gR+IP4W+EG/ZmxSa3TcBO
TMRcTbvu6tP2mN83Vc+j2ZBB7GXs/LzfPoA9CtR9CBh5EoyqSjExHdOad4XVRQhb
sJExz7c9GhGkhrUyb8JNtDCU1De/KySBk44EWuX/oaWI0LxbWfZLMlUL755o1bQP
/k67sEosZ66bLRKVTKSE7YlXEjtcKjWi+eThSVa+7PENwwqh4bQf//cHb6bEJFS8
dqvUvJ1yjXMaqYR5eIAyEEq5YMJGcbOPd5LtbP44x53o5ms1nXDNiqHHqNQ4UDiO
MPc/qN4jt4fSqonjWAQgXc454PMz04CjHcDkAcYfWIm9bhCGycXcXODlAj76ViwX
uohYv2uyURHTn4oDckDp2e8vp5XHMeZTAmL/yUTg1X6QXVbBQaaYwGata5VhfC4q
na7aRvAc7MI/miUGmzEgdimRKCQSCIQfLdCooMqe0gUN88yM/UWLYrbHk5iVxwW1
vRNWBb0kzvDICn0ll6S8nKAGOYeCL8lkLTzdPiMjYFTJG+NxOAPLhRr4SPS+FpyO
J3JKPm0uSpPdk3U9sAQDeT/rbAl1JEZ8gLNXoW6Tb3d5+qFXQHKkD9+xJ3jaBFNj
ufp/+/u4vTmXnA5Xch0SCPbrCNpKWl7rm2fasNLJYbypDN6nIrn9ytj9pMPKODQl
cEzVwYHfGHX0nD7/0hJ4N9X81+lfovpI70eyQSCuxXifIyncd+1LqR/WiRd6RAw7
/+Trriq3a7UtcPiDIXxN6SGOWuMN6FpR9DI/13FhEka4akUA4zUfDpZ9kzKyz9Lg
O5OoiRtEcVobVIBIcYRjF2coHu0G4kvHMNhwEmYGqLnOvUog4zf0SnTiDAoI76+C
c4K2EVdj9g+RvwZuvBXga1rn0k/d35TGzdhLgbkig9UDe7uXGE2sgTqKVsoOuqjB
917TfXqDsjw2D1ISma7qbLThORdOXzkvVgDFY84/KBe1TkHVyPxWkwRuq2lMGDMM
oOdx0x2N8j3/e5zOdTGL0A4pN3JAXKSa+j/58IQSdbeJAPxtIw+G+h2KX2JDm6XW
vcUOv9liyMtFfuXf7LMNrZPQsA6f9faQJH1cWO8Tu70qs0e3kqm7g1DzpB9n7HIc
T5haMYgAmqVMM208qkovyVeu+jHxTNB49Uoizge2qOVd2NxrIQB8MyOlg2DEuIla
DCjjCfsqXc/7If7vHNWhFlanv2iw30SHCF7SgC7ls5+PembeXVdqYOv19cqX1YBp
2yAvtDksmzLp+liKv200iLf6ZZJKAw9yfoTQz7B8OUW9zrZeUMWoRDBl96Y1Z/XE
u0BG7aLsyA7CV3laEIZa6WkrlUunc6IEXib2v+Pl88VANhfeQRSs+YZ+B1k668hK
7DlKdgeaY+W1PZ2r0/zBL46VQNgBUQfWFoALHCXHcEqfyCCDhLQaibQ112+WsP6U
72RHpIpX5LDCZEoxpxSjs9CanapSwlyLDvfbW2t261In7aaDZdopqEDBTdfDWMGv
+eOhsRjSdlHzQlRQM/xwAJvEh6zQcVM1fkLJ+J/zRYY8U8KdaO8lcEtyVoqlMmgu
We2Kso2/c9C8OTRRNu+WrhBj+9w5bJ7njFu7tNfkgze+3MC43dFUJMSU3RnBILK6
atVAARJ9uL0TbM7P0N2O7FOYmoB9BybHerVNpYoY+ek8pB+1hd81SuA7aGErhXjw
McutIggCHszFvu9L2ln0IafD+UloVFF+N/NybUpAM6Kd6aUI/7axBDZdsDDdxPDy
pk9DE9SO1r0AWLAwksZrZjXQr3lUWHEJCUpcvQVzc8/nthPiujwZC0K/gIgTNcsW
IPb9gYF2JdiPfFmXfr1eallp50zIiGfvlR7UdqZorvALY2S2+HvikJ1AQgoSWjpY
1Q+Z7i2iiTSTchRDmZBjNnbXdS8gJe2jtvfAz1jSQWIaTjIoY2SZ7eUZcR3PhOdh
spxLIuUTYgq7Y+JBR24wMwr0Z1fpHXXjkcTNUrdWBXo2Pm9iXtw/oYimt2rkgvVN
w0YUhJhILbjo5pE4vpSbDVv2w71yjithi5e0FPTd0s5RGbaKQLd75xMecz0vTN7A
N3OF/lFWiNKdZ1SEguglx2ppzHY70C00CJM8uXrxsbCcJi1/TeUx8sUbWT7ed9PE
KhZcMSZGp7ZTjFxZj+6Q7ZcYWoGWqWJ49OBuDUQXwbgyV7LqAa35hS9EXOlrcWI+
sAwWOBt+OfyUNddzaMDhLZi6LVu9t9ziFvTPPFNpqIGkz9gOJ4FxluyBxEjLxYDK
FFqkY8cbiAsCYJPV4DnTsmAXMXg902ne82k7t8ENhbjst7LNDo6kbGwmgn1TSDUJ
vT1K1P02lmFqFiI4DHQa+UL2gAz57hmFsfHaKUYp5VSZ8Zv80rEZ5L5HYgeVVakJ
HE4iwAbfsGMVS3LjzRuX0iABw5BmeX1wiMTI/Vn0MMpzieF+rGAwLcC9jsLHthFS
jh+Swcm26wOOWEWONcQZ+CWX9v28s86ZE45/j50G5d7zmKjnqXqYBHgSQNau40qb
fSr4TGTLPiJ1duuYdJ+6GvVI0cXp9UwRAeMdyjXo8S4JseaB4fC6r7bbZ1D2J9VM
fwmCdUWzb1qvRVjr+KY/SRmE/HZqoJdKHAWf/uCiP7vSmHsgHlXPIdaW5ghHlQ5i
jadXv3PaDfoM5/8Gjjs45WnN1E3ISoxJohY/ZNiZVylpH4YNeBgFl+aEpd0vBf2/
Uo60g1bdVNWcUqebj0lupOCXLYyRy+ZgNUlSICsHRtd8P6bADeBFRROBj1PZX/SH
jHiQUBSxEkENvk8+CtbU2AOOdnu5BgLby2yrm2hWayWQ6P/10THtK2+Y1R4xEtsE
6Qa/ZL+rrczfe1zs4LuIFd+lAJUz/rjS7TrCrZMkw/UqpGlG7RYwxNiVelxzsY6y
BVh4DoeaOOLyQUNIW5f1BqPmRJI4/GlQOBvNkoR2Zjxq303NH7pWsuf14M/yqo6N
sdllK0Q0lClvGbgd4DPWyiejcsItlKJVR0j5ceGY++UFZW1R6T2bVX1nXOu7b2FR
JT3Gb7QoAiz3tTkJK0pD9T0aWhyNMeQQ3JV3Y6Rm40ihSLtkVFKwFNz+Ip7j9MpI
/0HPaf43xleCweAU7SDwWvCdUfa0q+LS8edlfFY3d2wzgOsu7Abh3XXlMhy9ZNDF
0QEqJOKk9603IksDQuKuR0Yec+LdIH10MBaqUWj3Hf8FXDKnOn2RdX8EM0r562QS
zyxYl38uz56m5Fo8J4J1EcQdqBNZ10Ph4vj7H32KITClRNQ5fmZ4NllLhyXmdm14
WV4uBPOTlwkUaTH/CuWpMu3g2Q8EQbx7400//ScxKb4LhqLLMveBjUDy/9br+QFi
UVUEMCMwaxAt2aPjbKkoVtyLWEzYQZnEjNmx7p5zsEidD94PEBiE85L56UGqjee/
EDMilB5uCdPpqbi3ZHkVN3kgk1P0+aPAua89jB0Zjuzh/glkjPlW3p5lzYc36UoA
rd05cwXT0SRl6TFXbelbYaPRdsMFCCnaYeKfhcufEpxJG5VYpw/nUfoE69C85hn2
7Iicb3MVZrmOQTD/Y6wmFrE19fWsb91FrkTBYP3OX1425OmEniSAfIHekC4v/llh
ZOYun5iKW27NgXMjqAVGy7kKXix3qO7GfU9myAx8ZZkV39c+oXpR6Id6poygn8ZC
EkoCvYZAMgi1JJ4pZACKfKJexJlSrpSMbMBi6hEeDAVwlne428g6yfa/k9OHTxbJ
1InP4HE5I1Iig6aoMgdI4/hO9zAO70W+THzbTIdhbuqjb0FRUgA6udFNHwYnkbdG
LSu+4unAHZR1dgyNW4ju5O3lb6Jjb1r8hxnXwTfEpVSvz1jaS8DGP0MT+dZs7z/m
vZv+dFmm4jQQ2gg5EBQM6dhWM9+fiRK5NrKIgnaumRiLZrVJQgVIIFfBpnJxdokw
wCch80077ReQXqQ3yPQIh/V/KzIfZ9mzI74/md0JHueWvJ5/0f8w4/ChGnVy7H2X
s75tr6QE+u3C6LNDtm1J9QZZiMlUD/rIR31M3UNHN/X7Te6NSqZiIW0YFgA2Resx
XadLli4wHMm8bUa6bdAOc2uDIGENT20Zh0YL0Y4s2bi7MuzYAZOsGm04APLt+xef
AlJaojHDgPSwA3eVw2q9kmN+xhK7tSuP5IzIjEvQDceL28TK5Yn82g85t6eFptW9
BMBSDFwQvZxtUZnjaA4bVdZAMypeTWQI4f1Z7ayflpuyHMjqcXb/h8WON8OMIeIK
UL6g3oWNq7rYhf1fv2oMh9I6zAlfwI9XFisYEX4Ei+eRROf+GVW8E9J0KgQOTgP1
aKA877a9okdggctbHV+jClxn1MrdMR2nnUmQ20bUZ+yu71kgVjCr+gXAU8ulz0Nk
bQbLGqcvnr1QesAWDqY2qZerf3h6jvttDNOTYPCJUY06mdSCTWXjxVbgTKgzbdnU
GRd1ieVv80NVkwuiKjrM9h02svHwMUgvU0izVRUCF7JW6NrhgaBePOI4Zwln82uy
fyE+rcRbutNyeBD5EkFq+lER5xz8BpAPAQ7c9SxskNVi+SihmkGUneOEWJPymYce
5Mk0mK2p5gEM2pFQyj7sV7NbZxKIcvvarAoOmi7Lg5SBaro9SVQOG8AiRwYBSvS6
KhFMjcei1NLPTeGFwqOwB4NrIpecAWPVYk0mBINLx6oyKxFimxPGGXQpKMoq0Gkf
JTVe+5GdntneJCd3E55sYL3VVBO2PcN8DeuykjpSA1ruOMXy7/RhfG31A7j7hHK1
5GLCF/6R7gGjCoFtDWZDTm2OCK6mh1dUvlNwCt5Fw+pq1Wefa/sJMPaFgkQEfGfr
WT76px+TJd1p7n1rbx5PbzkKwMlp9BZQhIIY27K1DcnieJLF6GNPFhhbqD3gK+4v
O8CkV6b9I//MnuE5EM1zngdxnWh0uQsluZu53Lj4EDNY9MIAJyOYeHDriIBKGsLP
ZN6WoKK019ovbiKOoMq17TaLMRv5W87QrZ6NPSa9Y4NDx3bSQxF5qJbrXob1Tdzm
U1lR6a475oCC/bLuSeaNsbcWS/y1WOlkY+hPWbHR/BU0ComgiLJJXSSqcLN0WASm
sZYYs6MSffVHqlDxw2vLIZXqkGmAcYSIlznc2SmHe7BkzITkYSV+mh90XeUYgRnX
keGfxiLB3GMl+Djj6I7s973ov2Xlzd0Hicix1OuN/X1LFJoWGhv6//dfiTSG0CFa
3ttoSRvfpREO1ncJHCb6Tc7i3gkvtBvwkNze0G2osbdXmXwICHnYZR12TuFNq+cx
lkD7dkyoISd3JM1/MUQd1DfiD8pxplaQlpAHmmBlNiwsI5IuHwIXimXBpJ88YpLT
rcQTIyWVBIbaiixw9T5v+Ovfb9+Unq5fL5ZTBLEI6LDB+a9NQCfjYme5a7IHdGHx
ayufsIvjM7xoIT2ncbD3J3ZIYQCqUyTgNeupG1pT6tv7T96q/74i7X9Si3bXm4zY
iibLxlEtga6bqtzn4YT+ZgUy0jc1u9i75rqTM+Cwfnqa79O158hft7G0nOt8vlWu
aJuuF6kfw1W23bf/k9bQ8kVry2egh667Il1B+j20J5QQpakYOb2ZRIb3wadQhKzt
ul3Z2Bx2RAXZ2da7ea2ojaNWI2JpPvnqliiuM0X9Xw3zVtsB3re+QKNOaQcGQ96p
Dtm+tIOi3RLJK5HoaushKE/cFsT6THY2g543SCf4Zbs//Bvk7KGPo8unGsd9Sc8n
dK+4zvwZ/LSiCv+4WS6xqNakfJ7IqXahiODaulPrsxFZKPq4tvf4v35F27VjOJ6a
S1+d8uirxOSONyPi/K9jAXWH7An5DtBkizg+xzcmB/cFuDfvATEI+XSnyVJJD3HO
OCsqjA/ZmQE93O5nYpFEazuqNUKMh9Cjwm3uNKt8drwAxR9KsvymWXnm8UtMSuGy
CB63fBAv1DMZLYWasQ7hsnzddR/LSqc3H8pOLkve+YxC4/rOeH246smO0VSr/8Vx
UHJHWGIWn2gPiSCoghDq1h0zKZUueforUN1Wz5MO5VzIquUxcrl7OjMe6EifFdp+
iqYZn7XtU76f7wVMHA9J3BbHVlz1dE8Yq9JXQJKCaQcT/2mDxuEXW4OoI8llcxLG
fRN3iSRprDkPUDmhwj1mDdbV3qayBf/SMITWorQo+AjuQOH5EUmHomqKgABPKQPr
f7V10qByB6cVT+PaUAdMeJGTRALlUomLMp39xpZygd+mf7KIbTDaLvMI3MEwNoD3
+J9lPrMgiIyKf/Z3CIBXE4Jj0p94/tfBE+nKYFltNuhkJBsRJCCtQBI0q26pUkjt
IWCuvJ8WRegsJsHiQ1a8p9fxdvc0c66HhiKJrosF8VtRF5sBLw56OgNR1NGjt2Rt
UqUaj35jLmAmNJ3KI8+Poa3+belfjVYDLzVM/lhhvw5ND2MCjyy7SamsMKYLC06g
hNprAfXAFkyIrlYO31W8BdNF5Co5k1Oy7lpU/vq7MZxt0BQHy+AaKDHiTXalWUzM
91s0h8qsRB8V1XWYJV2fOd0z+lauhCdVRQvvgRjRmN1cXpPH3sHt6IpaR4uWTPBI
uPYtDi8gsBAsFrTSA9gbTzd1VfpCquoII1mc5EbUIf+Atw5iH6M9Nw/Pc8zGRIM4
zNzvN+M93Eo4pSBdoeBI+LI0edMljE8VlPdN4PKsiP3qIkCTWrUmu9zh6SSGR84u
w0dBqYvK3evYz7rzOpmKFN2jz30+u0UMQNlrKISZTRBUcUqaCxxaB1hexD4k0FBM
4DzRRj1ujh64xsGcrBUBaAjs86rpcjgussrQF1m8WglIwey84Mq18HNgl/aKcQqD
K6QQNRUn/wbH/CRhZZTN3XAuyRwtbfWJt35cKyVaNdjWlMrUNCpLIXGRqeXGA+pb
I8HiMFEGaknmd5igC3r5hd/635l3lMOy/JkUhwicAVfty/uAGmPI/y57f+n00Bbe
Sdt6ca64Yc5AC6YIM72U4BU6WKTBvzknX5XkYHmoXI1WO8K/2Wv9CMsmTNvddcdw
57Ntbm4Ac4/r+qW2EaFpXecTYGEAx1ZyG1oZFrtVQ3Lnr2yQhUSAEe2FYRqfvV4Y
FN4Shq8zvTSdlkb1e4iJG3Ck4toa0wmaCzW/1em05ADmPVSz6P9I60+91SEW7aiE
EmyIyfSFJPD05iK1K7e8sUnbORrMN5yIza8LraiMZ9CHXR9gUSNLKSaxC0TBt26k
3VeT0C80fMWHeBSygKKJT5tQJiR0l1cBfGMLtfpTVC8ALV2G9KZiYYK3WlxMBDf4
QumIH7cC3yUBabmF0PdbxZ0jBsoJXpJ9u2naHNlwkfSf6s0elQGbMMc5lNkM5379
svYCEKs/cysfzphGpaZJ6gbLXHD2bkcVeTyiOKzmVOkWFYnQgA47Pb9yZ/dZBvD2
I9jiZ0RJ88pEBPCeqs2CBAiGkT8pRcE+e18PnNSjj856ibPaFEkezEJAGkqDT67y
vjCFspHPRQ9rFjzWEPz95ZGboWk5HZtrzUq3OtvH4RQAuFWumXnBNAHGKBN64dJk
tR4fvnLC92WjDnTiEGFz2UZNCq7PsMDfxvDdyJkNfC0/E6aIMgrsdshDPu/lFmVH
GaHe/eZYgollFTYf1aOe9MWLkl00YCIJrz2rP2pRDRxwm3mGIr3s+0EYMhaAdxaR
kbKSY12KNImxVPoKFtwdkobcKLy8rQNUO4D0L1VkxTUY+9yukJ4X9Yx6Bfur+Jzq
kOPdTKOo0t9vvxyTTHBAf6qSw4Ay0Lws1zPWzfu1HJ7/W/vMd4OQNSyGT/CKjgBD
69OVrJLeBJIKK7VEp4ACW5/jQ26lOUoBpj5BoTM5Fn5/4qR/ji1HbJxYnrdFe9wE
riA9dxHCAp1dAov++Bh9mExuIJZTo6F8FARYLhLm3JOkdIqs7zXoGqKkg/Q4zk/C
9HBUDi9a/fcUQaU5VzuNOCFCkMWoOOlsT/UlhH2m6cSrWWvDaGmNswlznmwh7IP5
rdnfPaihbjT8pAm4yRNuf258kJXzMR3uipYahNwLdocpNekos/lOYGM4JzKjgidz
NlYRHB8lOwC6Om8BW4pHmqpLxcE+xHItWT1m3drttg2LnpyoBrrADnN/LOpLm9Lt
yX5pqb9Jm5EAJoY8IBRoawql5OoTdV18+SNQOFMlQ+7FstEKW57WRmEpCDwYv7+E
hnXGP1kiidwZqfR2SfsZS7WWZZ65cUDArn8nxf3cKGQWCyhPyVA2nMDT6UHwdUaT
0w+efBQE51yqa94ESeAe81ThOxBdKKmkh3+8fBMiih7nyO67j40WpBK0e/x+vkVb
PaspQH0BHi28a3NmD75NL3yJyjwfZs71LOvK8O8wp7v5Om7wzp+oIWdWga2dpY/R
+abWZ4VxTb60+uk74lEMD89fpFDJB1mlOokvLkSM0CfCdR/kvmI+s1RlY3thlASI
DIaNDpMGOKDiUBXl46l5IfuRxCOsIHWJXTr0VJChrSrdDXmOGPYP8Vsj/Ovz8zSd
6I3vXzpjiRO+JtUcQ9ObEK/rJxh79UZZ9zIOCH5qdXFYQ1ocqqJGK8WDqR+3ahP+
VjIRaiLr32kGnjTTZnwdGHWWpyBjqE7DaOfXXyRGrJFN184a4QS+kGXNwt4GGCIn
y8zP+DkHGTlawdwXPzfdx+D5DgKXngZOOPSc+fCx1Yf847DuOxNmkQ95CZCSf9xd
O1skYja6pAeweaLQkN+GimsOCC6l31PMSq36D/cWYJ719zlbmEc8OVIvdfBskEOo
u1j2E1oxQ8gjVOUy1YUFzsjV1ePZqbdQoRsa3wC8pbBIQtR6X618WccuQKvKCWrL
v27fOiKB1BJbtMZglqmnBE6YOVlSVfynrB3kL5LejMuCjYdPPgwZJ7WTvD2qjaKr
A8CJVGs1aH4CGozRqJDBjlvVqyZ9LhmtYSoeAL5iZfEjSnuwva2o0vRHh3OCLtoq
X/pilrDRWzSFdzz4X9mYjVEdukl8AZDD50KmXRtL51miL98Qvme5X7lPid6mk7nm
tJcfSPU9heGVq+u3hplseFJJ3JEk8maUTUD+1NXZKROSPWv8r9Z78C9b033jy9lG
fs/OnUlKBS3CnKLolZShTpTxwfcJK1r1xqmV5ktsZZx+unrUV+y5BcMLkbUJqxx+
d0/SauIKIC1PcevcU0tYHqkucZb1KQqSasxCORVRH3JZaWq+F1juRHc9qMEL3aM1
Y/vuGMbo5NdpV+p79BvcnYW2AYlqO4VYNhix2SRLrMOKvx8OLiGD4k5+nrefRM9d
SqLSgEUGJetEKeKd8M/higF5JTa+5CQukABuMGl3sxlI0DzOVO6Mqixf0HUXXBge
dT/cQ05UbOnodxcBnOrTcXJOfA4tCP2hUfbQlHwqwdk309mdTulbYQhhKkRRq0lk
Soz2HrX0pxx6diZBuG1ShI/8nGdZ9GJYfuQ8I/wwtoq6K1BrOwtjvTVhgxppmhm9
UCLL+jcorhafbJUPgyydVF5cGx0B8XCGdF69UwS5+5ci4OXZSjgYP+Poeoau/ubf
fnPqxftdDb6GhH1Mgt1ncuqjdKS/rQ23uGEZFz8Hx81KEM7+vllcBRVzPzhmPRU7
trFqkSlA0dtV4mB5iC42VzcOO3VTsNp1Q92sqyvgaaMtPLaowZga5rtIjkZQEpL6
xag31CyDam59DsHp35vOEFXvr+g825crezC5bhGzvRWumLkHfwjFTlKMco4wshcu
kOYQ21ryR/BBYGqdO0b3ksqBHFai3cva4CMudzUEkdDoEwVy6y1EJ27zTKds2ErZ
nmEr+qDphAVx3JbRyJAt+Zf6rtp2glx7ugGNhmimOJUUBPiut87ZqZmCxAaU4KdF
WGrsssLGDpEZ0TngJffba5sIAxPGIEBaKUzunwP2Y63RMGRG1S7+9LmYSVlWIBAl
Ve0egNNWvlBbALn7efbxSVCzl/V6q3CKYciXj1pzAiDHzXL+TgavFehKZSQvUedL
ViDygfgNM0dBET5zHUOK1+Se3KfpTPsZMKq5gqj/2oPWTDNRD89irqST3iCzJSPa
ASTNqwsnycbo4UqFj0/bqBt1rDynCL3Vo3Zc4uHcqO89knLUBRv7OvQq2tH4W3G3
IUqaboAuNTyv4qT1EmIW6vMDbY/ilPKhUCo6ddjf9IEtj2oRhpWLKD+fYoUhA5O+
tNZhZS0eeBgendmlmSLTk6RBzlKDW26MxrYUEnJriThXG+IMNJ7aOKuc+fz9hLAH
9RzssXiwkhNK9hPZJ22gV9zbNlR+1Kl/VYYwH3VHkfRrSOXlx/Y1bLCMH3Y48wq5
0OkXRomDXHSx7jTFg+u9HPJMAbSevpg3FzGgLQTxUxgxq/L5Hu3vbL4eQKl6tghL
cEZP7WPcuO1F8JgtWU8OZLfQxdxPbOHuIaBguto0i8Muzvy/PeVHcg6XCzqjC9u0
eyMc7tFHkwqQsrUNRXpfd3Yg8Ma4k/5Ydxf//SKazOudJND9EIXkFz7Ep+NTSzFA
UMEu/NE9T0PfeghE3FZoe8IACEVZUeY4bhEvRYFm8UA4t43AancrKQcD9TrsOkS6
aICUMHbTEyM9yoV/cHVVrM89eZEmB3Y5Nf90EfcTXF5RRwQQSrhjAH3CZHuLF1LX
2ZwdV4SaWvgYXnv/ynJiuXu/5reMQsDvvV4Jdd+95uSFl+SPZF9uWvQbnKiVNwCd
HYAF6l59fB2677NajL50guBp+8iOmgf9eWQ0b4ENqzZz2H0E4ourIp/VqkmDh508
TySar74KUNI8g8L4WvoAen1kVpfw07BZNZkBVsyMTJuoOEmCGIbd2oIkT35ElhKE
hCmTRXEY9MTLo+N2SFwn4niKXgADfu2sVMA3v8rmaBnVzuoaSHnZXmAlDDvwxS5q
S+bQd+cfKGd4pMxcRotuB4RkXrQdF4Wn/bqIQ0unUIA9AD5/gXRbKboEkH5mJslB
I3lCpMiznFkoXz+WWTZ5A7U/Xq9vVqJJshKlt5SwhFrk2Ebs5Ssg/Tdl+0TPTlYU
wG/Dx2Oxb3G3XDzxvNYENEfB8NltswCBS6jNXEuxUMwgE04hMqJdkrQr7w0bCtWw
9jNDo6TBWNTlN1lgWEZaj3/ePUEpY5DWug953QKeen7EXuYiIbVCV2Y276/NkYF2
NlslcS23qkitpO4JwpK0OYqgknAjZZJ5iaKGbqbnHQtOcBwtcBRvh472bGQ3uEFr
9a++Bc8E+7kn57UDf2x2NQm+f9KNfwe8j/zPWKlxMjKBwz+xmWwbYnKHoEWjfIRm
uU9bqXnklfId9ObhWKACWgNQHCjkO8qW1kU3AwmZPS0LyBkmgozj0Ke4OlonaX1m
Fg1wqvF47dgbmBqw0+ZzPCTAQ5jZFCWjNTj7uon49yQ3hUIW98uGuHZHzC+FGKgr
Pb4GI1LTj2GTIVbNa9FMO+96NXKXGIZUS/jKDmXrHCOIGZ9QAqeTK2uWTjmdNnqQ
RHiqybeVN12KCSeKS3PI+sge/eJfWtFW9PZbB0gKAlzg0w54EvGqJ+DQtfWk0EYz
usCrQJQdChuQlOh4a+GRvYe4lP/nzo4J6kIRBdC5KjmVfEJihl2q3XbDoGII/Vjb
lNk6Oy05N4AcJgn4lBidFdtFW9Zf5GA49LPW3KtRJprQKd/PGa/sR1SmwFgYwRyb
p8jBC04VhT3f1v4SM1dNx2NfNpN5OUl56d96ORdSII6cMrpu9anKqgzU3pJoTADd
53dCXFFGVYC3JRFcJjj+NcZJ8CZQ2GDr34vyV31YywxR+yeyKVdX7ZlifUT4LxQr
cOE0gMFUckJf4jcJNyp6caXRoLwHpKvoEXdI7gpt5zkQlBUndbS8lyMoVXuhzxhW
UtPMRiDGdU4l8UvuOvrSuXfBC6ADjilrjZyp/P/+Niy+Ft0ivCRWSlQ94Dm2rtG2
KeD/m69YvDs8EQZdNEyYcBV8E8iIVipwOHGOs1eAavaToeXIHoHbfNk1nqqS0bRC
8u+xJfugQaEHWUdzqrcwZBVVg1GES/KI4gaU6u3vJ+jz0iPOWJRQrwVVtY6pINEQ
GcMx8HyI7PNqCZ0tA17B+7oNUT7KYb89eWTkgwUFCs51KtdaZnpgzYjhdIN/FPfl
9kGm2w0hu08c1T0nCIA9fe95ZVF/tRlFY+y7zQ3KIFve5OVeG59YLad/Pva/dNuv
9obiD0+eonu/lyDVMDZ1rNlFC6wou1jWCqKLU3kNrJi7veBULgPd5caIAZ1gDpYY
MLzbYIu6H9wcQgswo4Zw1MZ34ZuUrxPDmySY0zt++GtzdfZDeEkHEauV1NoJxePM
dK3QeqC6tyDJMYJp3woAE+T791cFFemT2KdVLNCeNemBy7I1lTi6VsDaje58XfCO
pYDOwf/2XHdxj9iOXCHKtR4SieXFiv3M7nmjiaPcZ6ZDnp4N1xFtoshg7b2KJUbu
r7CyZN87ATf9kO4sNeqZE9mnJOvXkXtpz7MRbpTO8vno7LqCAFcCNrKbmQAkp0KA
vxk2Kp7mRfF8dgrbvDgjYt4SWdgvm9xJcUf2vCqrslJlOqtIGqKhMlc33oCHP+en
iDEp7bprkyLYg6wwOY+0BvvZVQS1OVITIkMjxePz9OXtrzfAwe52JxUmLUjGxjM1
LRzX8mD2QDpXTf0c/7ktXkyJL9ZhodZ/zpnxIHCOQ4q9spLkKQzphNOQATWx43pj
4aWrPsLIc97avyrIRactZIBrAITtYFciLC7gFAGWRC7VlajV8A8+W8nXeoTYpmRw
zKm6AiYHNmz4lpm+KbZRzLPoZh0fOCKJ9TfS0/P6CAo7aVploWiFJw9puSAGx5nq
6JDNi9J//rPgOOc1zNpf/FI9A2DGgq75PKDFGCucKowdFSMHuNye4vWCbrt84dLR
0xm2ee3450ZulCr8cMpGh+rK7k6p6WpajyQsgMIHOzXMrCfHfk02dVhOqB6ObgAl
+bWsos16kDxVGrZzo1jVM5QlNfiM0UrvSRrefcTNaLTUYV7L5Q3BQqS6t4EWoaU8
xtQt8QAxFyEguU+Z5EP7/8hO9Ep5UPCt42TpK7eBx3E44zy8sFAE3Xkte+9kXv7G
T+y8uK6YJLN7Mw0jWsFlU18EUM3Ppnu2pC05d4kFjWbQKn0BQkW06Y88wjCSMWiB
bFGS457YPAO9b3USKpbYG0bKedksBZZkjK6XQFpsF2F1skm4y8rJYRGYK0MoIvFB
DUgYmdf249+GIr2YXb48QSma6vPyXJRlFRNi1nCz4xN5f+BrgcbSZTjZjWKl2P60
NtDk44hdqZifWAjsyOAS7w20zLZs5ULTFvO1+oXXHFF6lOsyh47eEr4e39XPA5+r
jVywcOO0ECHrlcyG1yamuWf3GBj6PG1zpLAbfQ7BBKYbOqqL/Erxy8ZNDkuasrMl
7Re7kgF9O4aa+U3zB638VdDNOmRmUvwTmYKvyi8Krs8IdWFF9IfKbLRw99CKSl9t
4QGiJl6CRI8m6Upu6ug2juKJSRKznw2vlmOC+olvdDGGJ0s9ep0AMZO/Rsw3P2gL
Ukfrz5kU9CeUXX2U56Oav0ZyNa5arKt21RjKQQvBSDPX0ZsxWaTcktPTpf3QONlD
xYBMODud9I5ZjWgG25gu3EIoADAQpqGG1B80lme+8MRcn0FhYTbSuRV7LwKTebqT
JjjpPbX7xc5/Adw9k7Gaus0G9cpUzuUc1u0NFMES0R8d/Aj9DY8E0JENVl/DBSOH
wKmHA5NFPhESoLcwZFleiSv06rBY7rRZA7rSI1JwPesECN9j2H7aEbfIFbEq3wZz
a4G1Gd06ECTvK7zWM0rX9tWPv2wO5zBy6i45wYqQj5FtrPFbCPDTmcGlMilxlFV6
uwTsnYBQSd2YbwFAJtXRbh14CVpt0fTcNgaNTeGMhZOFt7zq3S9wFM/MHjq3hk68
57ptqg2JOe/LaxvwtMOgy+c/E33AyM/tmip/J14T1VlNEJraa1UELkstyaRkfzlo
kbspWR5hat2+ii5UnbPzamVujh3a0voAmNt3MdRY7F8W8aqTAo/ArCMaZ17mwRQu
U1hicfJrS/5yNkJn/lfSu9D1DqRbyrI6m8xvPQapo5ocUQP43JFpuadYTdimpW+w
KduSzB14gt+j+JS0jGOwMmr0AqpqGrVWs1p3sZv90qj2ZVAvlWNP+Tweak30kdjZ
gTFlfwfOu5bUpu0P/1RHfFrTVDVYkQdqwUe+p29BLiXbuQBFteGWTkVGWCCHWblz
sJQvmKRvImkvkYDU3sD1aGyjkWKzhKat1v6fHA2FTu+qMs9Y/cjewEtRAnSJCs4m
LiAsBhqttfvYtI/ZMhG0nzS7IQ43CiIFz1oLU3qjhPOSK8CUMqWYUbyjaYQrNtpn
UsTqVrDmGu72GIPBAwqqUJwsrK2EtD2sPIHUr1Cy7kG3Y2JOKfxzkDI57YWnO4q4
nnh3q+/X+A+bVk4mYrj9+KVv2d0BWTTUSCPd8e+/IpMkFLyGeU82PD3B4QTOUIBh
NPgxLnwBHYJWzQyAw/i9S4GXdKMeLQhcTaH8aDHtnPbprUsiy03//uRObaH3J3pp
fBMOVZ4ri845sSHvqcIN8kbhxMZ7Y6qw+Bz/Am3Y63ZUIzerAVJ9ij0IRtGyVifD
XtmRDqeInPBhicuDhHw7/YShNnv1Q2HR3UJSj2ykBayJ9OGhZSNgUn11JEq8UqNV
G73Ob24iNQ/nuZWBOyjs+aRawwULXOTvv4TUeP/B1nLhpTLcAJ7eeRxs2cyVwmA4
bmYjiWVYXmJw2fTeGC2xsDquc9WGho+u7ESiqEOdxpEznQUET4E0M7wWokgychN8
Hs6p6mF3egXlOvwyfSoGLrW6wg4mJ/Jtt3Cfvf56NYA8ThzE//BmBYj9ZaSpBpuf
r6Rjm0aDlJhD+g4SMyPDc6wyDnZ5xYnMqvJCPXt19N2AdyRHpG4nEur2kNNP4huu
83rv3gLIWKhsgPsAFB+035aNe88n36GWMsVpG+ONiJOHJbEA1foVypmzRXiNVrnh
cm8KPyJRnuue7lwU3cODMkb5jf9tUa4qzfez8YF/huOicGGsXRcY2R4fMks+rzqP
iDJneM/hOYLXeDQiaK6sMX4oH+YI7cRpU/d7q9jqQKxzTkN6FPNf3rFmiHrAcqK8
79YRhaLhQaURPKLaI1CvQHX45/+FpGJ+FB/NEhvwb85OGBDlDDi1fqMhuMZC/U5W
1FibRAOXWekyOLnUXk4wc02L1r07FvxskGnG4fxyWwkrK1ya+ppHGQnPJkDl7IU8
a/N8qJ95DfQtcuRm3JxkaWa60NPeY2OfkryJEG2SwbgRc9/ASBug2w/BmyG+7YEQ
t7KeNf34PnI+eIfvFtvmNkVXdwh035tNCp+B8FlxqPe/kV3mLsH52fubqRjX2ofv
Rf3uvY69rmiec0Jhp7vSIpRmlte5caC6R/r+LxbuIA1xR504dfbzubuMCJK8jpHf
pnokqs7de/30yRUDn2H60gApfX6dKxh+HI8CE8CBwGhllCMfLSt9HN4qWEgw3Q2P
UXIbS0JoVRJKQGnJ/mM/mqIXDHr4CWosxj4BYvQel5EHm28sT3KQMqn1CUyKW0N7
KiHzs0ikTM3AJOSYUJznXy8sDLgLtBqpY/JQ/F1FRS+PFUmNebWvVIijKEWQe1oY
XHKMYHuZ/HLs+85jLH+uey5DgNo0q5EKsDKsiuMmnQf9L5cmm2Xnr4Gl6vdtqWju
gtTVmb4Q+L/QOALCbLpIHO7YhmC+DauFnhICOPCxClxOxCIBLVUVrXzWtDUPFuDI
1rS0KUtOblZPIp4mi5A5d0RfMVrR7yZKtczv31K/grxtkABMNk/LrUDtyiS1ZaNr
vkKMS9jB1CLmVSBzTyNeDLnXZLA4xbO4XRpkMPoQbOR2eWOyGR1d2ugdzeuNuaJv
paDIvAudp8nTdNEBg0zU2rx2dpyCha+K4sCHgJkc7/cn7zB+re4FlS/6zbuPlyoC
ym2A2Jsh7ZTYkjBO1p4kyHi2nVlhv+PoJASOwopuE5MmUy+qXEDqhrlcSvn7tr8e
oNs3/R8Trbdcs3bcBPPhicYXq1FCHvhQzy2WP3oLt633NxHtVyyXmofGN9mOSXLU
BthjHZ31iolbVIOiLXypqYupKKHuavbeY/qywYAUif8nvztPe+7fXFOVj7D/OOFw
5UaMpvUvT2GfDygZKzzzaTN9nM3RSw8egq8WxkK0tX0rmx6/i4Jc6/Tq9JHFH04N
r9JQhW1gXZXilX2LhS4a+v+R5cF4ttd1ZPGQmay+4yNz9bJWykCnREX+SRwpj2UH
BsAHN5HDZURHj7pFo5ekReCFBdqx78rQ56Oia92RvYJtSqfX0CgMeyj2kJPKJM98
wunyJgl2bynmD22rFRBR5LZZihUsR2leQnnPOjbsjCRV/4YkjBE8VBUudX2ySibN
Z2fxVsDnkyil10aAYS0hCPuiu6Jn3jePJegxSYn4mf1lHaJkYJ6ce8bhtyAvdyaW
kBorvcw9vmmTUFlBdlRoJzYulL3fzMvyM+eo2rE1M6oTvnHzsG+ud5LIpn3hrIAX
sKbug6GbUb4xXtchw6qw3YyFZ4rP/UYb9WSBoTiuTa70QrKu8kuhbjpj9OoPEL8G
mDS1bhGVcJzMdDxQRCzt39L/NDR5hGw4BKrov1CQPpzQ17X/i7Ub7MXW5n9P+CaL
IWXTAIHYdJk8mqvi1wzoW0Nne0DSrjx7cdABwm08qWQ1e1SECQdJcXZkbp+3ga2N
W0xi4FZberQfWajSHRRwMbo73e1zeSsUS1eU/JF3eRHNVmY3T3WVDHLBE+iBliuY
Nodv5ubXWJ2dRTZfm0vDJo9W1x80Gu3twtF6+9AjI2/uOQoybDxmT7sTZQThRkI1
+Wp/LnIPXYqkUMn5dXagppzzuvpJYE8Xw7RCICNUhwNo0mMgKJZ+REc/aghQ8rov
OgPzU+Kqb0racB8O7OxJW8J6o4g5Zuv+cV4shTmxqOisKdEiHE+LdJF7ezsa0WhA
3xIhkxO2Eo9xgnH6mpy6mCNC2nsws5tv2P4HOU/880Zv8DXilA/kvTG5qJZS0Kve
+StwQkMP7EdrjnD55tL6EKByXKY8JQGKMWk5p00mgEeTdIPcdmZ54Pq2xWPA4aGH
paYuhzEUxPU4+hqBONGYrjtyEZ1YHI9cdUxWZuErxh+BUyk9+RdiHjtx0zLCXZk6
uZ25Mv3wLZk6Iy28m+NUukWGXKdZxdZk6ccaOEsQzetUE5yMalJEaWbi7SF1yRpO
e02SuGml3TJp66e9OzWYcBFMTQRKYpd/D0tgDoOSAgheT/gv7ZRvAgXEtoBv34vU
E+le8pCinnl+fQBLtZwdcSdpEgRFe3/1Wj/Gib7p8lXuqP0biof7LYrshF15IDyH
vv+ZGU1MvT082JBn0cHys3tRPE2hUUOxXSztxGbZPZmHA012S7QvDDO5YdqNm+j8
RphJABe6PVKCuWudRWDrouPrRJ+ePcS24cvCfE5DhammTNCsuh3A4LS7fqIM04Fe
lvR0kYbmNVD8QdJ77tR3JR2Og8ofvPzlXFz2yJemdVHuEDlLdXVxDZWbty/KcIk0
eESFt1bgBx2I0ktZIl4Ly0jV8T1u/TgdeLoumWoZWG+9eXQX8n8YXwnRd44oEOmu
abQW62fGEuVhDSBfi87TQ6ObGu2BhOH+9u+/W6Z5Pe6awfW8FVtO9aQ/8tF3NTe5
7qn1bDTz+rKXCqCbI/kPhwKsIXVKk8vwCNdNp4KrE2pu2Ovp0rPjOKCvOy4rA/ar
078bBOKjaAfpw4ELQ6WRVpjPBvaWfn9Z32TOQf/jy1wBsJbbr47FuU46u0n7g85T
5f7wxpAmfDznksHwLjwPc+fFCak8Wh7X7Ud4I8M8ruNbTZd7LFyn5tfGvDvFcvvT
O0FJ3/oPEVm6POkjyRIXewFuYsjH+3qo/tbmXHF1+plUF0kew1/I54w/krctiI3L
/LVhGpa7X25qTxpix+HopP6fGOpBugu05YrdAI6DZ/mtQrYYplF6B5E2W7qVFY2z
8YOhuZdw2li90qAOBtFqvNYSnBap/RsWpbOcW/WtQ1nEFEDnJrcxzIQDdVhEF+U3
s0ZKOVeAYCLhv/h/QhNkeUPn+6nK54Md6e8TkvzQnBzAhcj1uPVUvGIB1lvkaURb
uKzfhbhowYlMM/YRLyI7nLFdcWNg0N+3GhkT9ic510EUhEj7fHF9ARmgUT2J573H
WjNDpfi6XD83Vq61x6Iqqbdf5T1yn09WxAlZb6/f/MPVaxV0LM9hPu/vbfxOMoWY
jo3xcaW3cDeQIEIwcL8mH/34IWHsAjDpmqMvMFGv/qrpBXa2UivA+i+fg5bt0zsM
ruLJep83O7v10Me8rGMAM9to7QNOkh/4io5hYV51S43vKlgvg+JM5+4zq1o+gmny
BHE7ywZfgYceYIBtLBia8WWMvMR8J1vkQJgrMIyo3Si8loBisfzVeeWcnva9reYv
Np/fdf0WO6t46d3yuSzLCwDsNS6EIgP9etLTgTv9ak5xrbG0ehCROuC9H8wUR2Wo
EQXEXjPVFM+gTzfOw4GOf18VDK7xXWMVMtT2G5z9K8xUwqvYByk0LBf9hZxLRciJ
8u/YMfDDGoDuEjiSTeFRTE3DELmEYCMmds4ZGpbM2zmsYuU1PLsWZxuahMi+vujD
7azTLHfgP8SJbCfc39Zkb0IpCxXARyxEBKzj/nqIIzT/YzBQY8YawRdx4i33BUsd
MemkiSaBjfwMjbq16Ezj6bjoc+iDlYn4C5L5lJ/kVzZYarWIwm6JeSfelCfT49g5
DUsFApEqjQCAmoWYkuCDz5sFuAzJWNYi1Uq+IPiof4ZxyX2G0SoPcMkkZv1mF3OP
HtdV4rrQUnPnXGPBv2hB/wXddBRdoGMGrOkUNXaAUPhXw/3vJbOEU++E+gVhA9iO
KXGBP2W7og4n7bTVhNHU0FSASUbCUj2YuWVGSpJSVN8hTbPTC3HbY2HoCE4UZLCg
gkSfwp8oMo70O4qdl2YuFGsOJBRyufRIz+xpRNhvDHN2Xj02DldHKncByOCrLVAm
s03L7u6CZoLFqM/fEtHE69rUv5DwU9GVn0rbRYTbXg9KKybi8aMLYccEQmz0KZUw
C/ZqejucIjJzQobJyycoTRJ9Yf6I4eiDb9nC/k7AwG6Kg35h3NJEafUdnRipQ3xn
Dt8eKhYOgbMxBpC7efEVl1NzdI0JnluRQGtJMdMbU4vqTUKrZetOUk36cUgd2cY2
O8AqR4z20ebBpaFfd1lzv0IjCHdlms4pBKObbaCFvKAx2ZGNbVw4kdfrd5bqvbyL
gXlKwn2EveB+/scLUm1CtZUpmJEJp3y1ynpK1aQIoE1/UVIcB+BLnmaiTWN2khuO
YfigzueB9u3OqsFjX0NdL+xoDJ1+Z1HExz6UdPEWjkuMcV29HR6/tBr2+v8A4/UP
2nSQvcW3u/FHQXUKYrYbj3DZkUevQiTNg3okWqWo54fFYCGNmCqkMhlVBKjJ8Zk3
1+iOtMl+Yv4UyX5cCPSiZ2ajJJFcPLGoepM/r7KoKl3SRmXSWlf/B0EMESM8DvDF
vY2hnMMrWeRkwG1slxPxmnWp1Cp0XjCHvqh1cLI3poMGqOwY0Vv41wBVVT8YgKsS
OZ6kvc+zUO/1Yg3HIAcOyUJhztizoAZcEqi31iNOzx7mTJLcshWCPjqXb70iXaBr
rgtWkn8f7CdEs9iVyof9x7fXDTp4RNQ0KVJ/RWBJVG3e00Z93uDU4aqTXWLhyrjt
YNtnr7rH1xJLlvJ7gvxG3iDRnxfVb1mw80QFoBfYFSBUMohrnZdKrRIUuibuKjEw
Ao5hzxe09CjX041USQ0Aa1p0WbR7MTnseu8BFITo1v6Hi/6f6A5uNPXyIqVB8oPc
7pZBQEFfKD8zGeuubXqm/o8N+yuooYWlxHZi5ighsJ6fphoUCFYH4KwHwsPPEhG3
UOwRRHHi88vjaRGJgIjEOGKGsnfA7Z3UiRas/H1qIA1eWGvn2kAzMgVacbvcj5oY
IwFMv5W+pMhiwJk+9JYctx5maszme2izkFheMJiPgBDOvRv7qswh03SLVw32QrP3
HXNyaS9IMGq0gSQ4r2HevNzry1evpQInL9qZdmhj2AHzceui2c7WEWffdMdx4R6J
UvvH11JZYpRTY5SAmnwKuRobj6VHpqqM1SEs6RwDkt/ZNz6BGGt3CJZ7JAOPrAJg
oZBU7U/VkUUBIvvSDRc5ry1QGpvINvLPciL2UFwy0Rr+Rm9tyuPR2PsvZbPOh2Nw
q+HSS/bARAk7AxphL1SPeH/WkvkU+vE7zUvrMagh7x9DIKmvXB+GeTjr525EZift
X+US4arNXqbDK1pqC8XUgWiGfd49hFDCcSS0lwq9/Pugwb1uFc+NBPjFtS1sUm29
NUfabFJ2dQQCty99AdrBcn8TEbBMbBQSHbP8/favm3gPMKZ46wohMXqIFZP4LxWH
sCkQKmIUb943nBOZ2OSDGwFJYa6ezCOwNrOOfxRpny8/bmeWC/XiHHcQxx2bISrk
ZvKbie/q93dKkxBnb8rkiYAUjPA8QuDAkkGaKh9CFBCoNSjB99/CWo3N8UnRiPhm
vS8GhTD9EA5pZiypr15becKuDfynVogxB/TEranzm2WK8aN/I2svLKiQSK5ZUhEu
VMXkqwu/j1GlpLsCtO+L6062/sBpASXA53gIkmKzTtnBXkoDFG4PM705QE4rFBhJ
bESSTDoQlgS6Qpz260jGCbXsSZvJEUR5S9a499BjW6WeKy7poyC9aySSK8Zh+2np
7XGlACBdsN/RuPDThYZgFc4yWNAPEt6i0MIaHGU2oFVM8iG9hw/ll+NoRPsYb7xp
gVOTszRJneti2LscddKi2i3vrlWeM1Ek1ReQMsm7hU4Ov+nJ2+iHiIfW3S8k6N2+
olwxM7J7R8RB3BBCrWfGRl++Cn64bHApTER69+IWFdZTER5HdT4zwzXq4M0Ax8B5
JmgCnaxBCuc/VcVG91oVZjEqbstzkHZjSnsXX3PrS/eeUVsmWekyjmf4eS3iUiHY
NADJge7n6aW/d7iyWIBVpqe1r0Qr/95tByAjpdF7lmqPAkX8VQTSApMENncqPv6c
42+4J8KMtHQzJ2WE43aKF5ESkRSaqpDj98m5baCJZdZv/dQvFtLWwDORSuFAaIsY
1JbNBubDoUzQdrxWHxhCZMsiL5QqqU3tPLoOpI6we6szFqyDi0CjUy9DNYu8JLUT
Y5+P9BUAihjeaI8C9D++hxePMOoAvunEYbrvAcYYjmdJtNtb4K1p23z+un2ez+oX
n7pYuQjUfMVmnvlpHBn6OUoCLNJjIYVNmP7z27m20qnzyyx4dNZMtucdPpQf0H96
cgOHOhgAtDQhsiHMauItwq/qCerSqX8gw6Vls05ElVXepuVEmTMOYL91qgLl5iHy
fsfkKZHphEWuUZANDn9fB5eS02eLbq37vT8qzYAncJnZZ0F2IdRQXsfI5dxxyPdN
0FK3kwZgfYvi9lNcqoqLY22KBIBz7WqTKfRxAfNNLIPNQR+L/gPOhpTZeTYFacLn
0FWyuVVtnqVWmkaLio+lg0t0xLvMtKhdo2NvS9JFwavtakx1JXm3jIA6FK7jvuo0
d0/JtrPlNPS5/SJQmIk+7Ow/wb956Mo3LVJbsXBTOyofb+BmRo0ALcsPaTE986K8
1G6Ge06k7e5VXWnMFYC3N4aUaS0UYnX7+8aNbGRWlI3CVOQhxmi+hL0GjriJr5V3
Gr/JD6fgcHV6yF3bBpfr2S5zaJij85dB45LSCVsDnO57QdATo1jLSR2gL/BwWzsW
Eez5H4kehGCF+9cHw8ZGGIAaurQRa1I/GZ3E8tXVfmF/yYHInZRjqOvziGMR+ZkO
rJ+AUaHsgmu5sLzGMzCvzfy8SeZqA3Fg/obIGIXnB1aAH7g9Vgq/kbuEkSMqC5tw
YbKnsMsZqg+44Po6g0Z5ajyH96bCxN8LibDQg9t7SZEBBPYXGDUwg8KglnF0ulTr
9GDn/BHqkJUf6EltaJvG8tDVrN0HGbLbMEcS6c+cNraUF+08yLLizCkwt1KgDPr7
nZgF6JHqV6Jh1m/XCsZCAIPQhcbS9Qqsqr3RGlH04ZrX7zHcUdlyUqjptIIuIj2C
tfIdsupXHYJLRMH65JSWCKgPyqvLP1iWgYd0hEA3UYkdnhrCjKaZNP2h5Wec2nfm
xzk/uojSkEfjLlr6oT4EBeb0VpHhvFS6gWYWTJ4QEVg0nxRSZKv38o+OpBiszhUb
FmqJCM65nSAZQjLD8fx8bym5H+yORHurgxPQjdTEQ+mXJt0oOyakSOdglDiugbDO
9dBT+JndNLOjqwibfojR4eHDeYYha3nAocahcgQ4m+dasLOrMrhbhHJKVXahHl+W
z++Thp/EgY4pcVKuTfjhhPI3D3dHhCkPz1nBORNGe+DFIxoRmOMvPzXtcqHVzAQM
GWuyiWgMa7fHn1EMFaTdiHQ8WP75m1ih57aIAC2KGShHcQUhKkE5A5/Y6F7n/bZQ
+rmdh1AUBoxNIT9sLgzW9ZTZDs4OIMG5kh2LVrf+fw+w+mxRSLzTkq3aQ8SqTtkB
QgNO3nR3fJWDQCGPdzzH707pxljONKM6WpvoBfkW4lKG3Dk4rufGN/RkEymdnZ1m
sHKtQ0fdsgMMIR/RIMTSq0iLr5cQYePvDbtOD2bntOElC3J63006bplM/3tHgEy9
Dbj/G4VeKCjdJWWR8tslvFqHLoSH4VFzj0f2OoNMZJssFuAr1xX9C6nwPRJNrgt4
I5Uz9DzolHT5RTJbuyCg6QZmQm+8Ay0MRngmXQSV3ju6q4eP2iZo8kfjheRpw1W9
lyFqCpZAqrsws4M8dTyJzoAN6fRY2rVRIUJvv/HO/YPonAefbb8KV5VKppCKHmx9
obS5Zl1BQ4QWEKw5HXn9LETRv7lq4bw8nZSeVixBQ/Vg+bF2K2anHgv9749OBdp1
ZNQTVlSi5PXn1NZX5lsN4KVbwpVh867E2rvjMTqokCFoQBh0CUr8V6xrtJvbsxtq
0qPrR90Q8jc64yKI1iyRFvqIxIl6QUFXabOJzv+wOHb+muGNkSKhxLp5YBPh1ZFY
MjkRdX518N3V4VTrnwt012afcJdTGwl7PTcq6XGPZFfaIkTywtsfnI4DvibZLqzX
Kwzb6Yackd5L37Dcx2WZw/Tqxl3QyXQGpejFFp+9D1HGM8UOW+SgHdwPOcBUuBU9
BJ8RJ81c/kL2FTyyLOMNnwPXCcmRAFOqpY+TGLZnOwUxWjJDzWFYK17YOXbuVQl6
t/0GXENtUtLqy/hORBg5LQ0+T37hiIt9CMiX9xuEHHPCIZNaLeuI8sKUnEv8/uGh
O2xDGeZUxKGqbuMmC7WYBWCBCrgC2Etzw4utA2BF9MsI22qYypzIS/HwSrvSfCcn
ymrpny5NT6jB+F9dz/GByHJIwo8tXNOhCfivxjumUyg1WPX6bM9BZ+615htzyF9/
kmhY+/e8jp9XBST/ItoOZKxA895GPvYvZXWQG4fdKxDv/z4oqOFUSuuoyQpl3Zt8
8UJXyfRnGKwB+iwlvbCN8wQ9AjChjUJ64NNYDQk3qX/4Hnmk/328u5NGRmpMULpG
/SbdcAern9ryoPkc3/gt95HqxNxjBaeSU6o1siGUDiS9R7K0ZAXAUJG1ZC2RM+vU
CI7+38JwLLYTwpwMmoMCy6g5VsO/1bhS8f/bg6MCUNLM5MABqiG8fkGEMS1QUVd6
y3aS9Tkdto6ilyzmWDI90COaZZ8U2e4TiEgup8mQL5vUfP9FS5qD7Ow0H1XfO8Wo
fS4Zd9MMoKwlPICchHJMb8OURxplWqt4f3Jn1qA6Cb0c3qcgNYXW9O85L8a8WGOE
IMKvf5hzuzrBCpoL9squYpN1X2VDTwGWNSf///Q6f5J9EnLES3ZEDKQfLdeB1/IH
Qz2XRjB/4GXNBmZBD6ewdkDUUdGRcvvmwfm1pEfp7HenPVaXTDEaYOemdKSEltdQ
sWZvr3eZimi9UiO87yGZbM0MZk3BYHNXA8LBUH1SBlQRF2imDA3ElGHhXMxjqpjO
4H/B5TQAoQXX2ZGNDEyb3NhQkt1DzDx0Vo3FMG81k6ZchZ0r0mH+GqvOjkUoA4nv
pLuNSQh+Z+Wu6LHM7AadTi3jRY20KDIY6jZZjR2wsC3KMpKxopUmmgY7q2SPJA34
hQRQxt7BL+rtz9XHW49LI2yEBg59qgx/3i71PEPdw9hq6zsFIyNSQKozgTCoSXbd
LcsJ0tuzHEXoG46lyWSR/5wPX6zoAItB/phHN32PjTSN/O4jpq+wnN/z/S/o7fXr
DTRDqazUZRZ7acKjEUJfHnq9E48OVAUydVn7dlFjsrx6qtuQeCFYvma3NMwpnB8B
RN33am0G7JSImPSPEWk+iVtbxIQm1O2l3IfR+MOfNnTz5/eQpsJE7aORi6M1uRr9
0YxQKitqVNS52sOsZWzF7d6PRAQwE/APIoV/YJCXR1pts0XiYgsBGT8xwVZnXhL3
w7Zu3cQWtT0YNEeyr+6csBf348lGYJr/9Un8J05zkgYSF/l0n2WaKU2k+M96K88l
9ZGY2pgGC8WaBHLim28ZPXOq+bnfV1wXis9LeWaf/XXj36Z4VM9sPqYIgWhxBNNU
dEv4CVXevXIpOUNzI3T6D17+036nnLPf8IHqZjrbXn3f861Z3nM0ct8Nljufplw4
bA+M6nQ40VydJyiCUyfURLHgHeb61Hbz6O5uZK41Bxz+GeQlL5CLoOV68G+m6OsZ
LiAAC50uJp3Ss5vMy9pfSG8p0n9Vw1KirZ0IQHj9/dq2ScFWrabV6EMc4sYKpQ4p
pQeL2nlw25IZMVK8QYBy+P6tGIa+xgvDuLZxqzy8UinNc6Ge+NXM70xDxW20Aak4
jop7ukd8Rn7UuWIyzMxLJNUf60sDiUyU6qmZBCkVmcsZe9iqr8z1t42/2PKbJwVJ
pr+D+vQxxoiBsaYQ6zUtlEnKc4qywZlS5smF6Ont5H1nuUz8QqJTdRZzgcXncVsK
VAomER1ukwgqbWWRZeT7Tyb1tR3r9/OFw+V9pA1KrQZKviDErFneiEW1Ip+T/Y92
p2SUY/EWGJP67vyl9q97V4ZhGgEAKFJm0F1NArHFx+FeaQdw/nGgx1Y45mqN6Piv
HVCHVLO3nZclFzbX5jQu9j8Luta1PUZeIWqtvLxDq+FHhUhPVRzPNY61A2GtGti2
7aFvlmmKtdf1dBVlB/BF0PQ3+mTgC/6FL/dc4gsMCSnP8ALqJ1xJXq5AdpluhKe4
E6UEkmebbhfGSpIHBfqLUeR95vB763ivZTXNZ00EkJ6apRnuTkd9dfOxYPZFW/7v
r+5n58jeT8r+ucnDt7/XgawNeb3iwVEEQ/BIL2J4JDpVztVZ/xZoPASiJc2LRcW+
OJL7ATxQ4BuaI4/gm4w8zemeZMfYa8/BvCbFfg4K+hc8cS9/t6l0zw+kaxiWqr39
r08eLB7z/PeyV+mvTnQGtkCqQfjsSIJCGdM3s0TykYvhKVi0QgACT2C6Lt+mH9iL
aJfBxOrWfjkk21ly7I6HElHlujVV1ih71kEl3Hy/DLPOpRfuM6vaP1sffYqa0dCZ
QCQ/XCisvWJQCWBcT1nnj1F0wkluRLg/s+ikj2+j1Frr7ULc1OXLSt2akCw9AbeI
PbTIKvB15dxYNx0Lv+ZOtUEBmqM8uemey6e0F9eIIOeSokOoU2nYdS6gKevF6rvl
Ieq7d75GknyZ/QKR1gskP4NYbQ6spALu9x6lkSWdj1PIsSJKClPhqYEreE8gWaTa
dNggYW2xPQXf26NChYeocfd7W+IlmaQTgv3qC9IoquCxhoUxkEsHXzbKXqCl7wY3
u1KLuvkuIf9MVw5y6OUT6BftKAN2Z2GcQ6zitP4Q4bRTuN97Gnszt+yunIHxBGKB
a9/c2Myaz6k27Qjzgfq5tCFFRL6NKSIjFkQAkm65DJdCocyjabhCce+xoOWgg7NW
kL+0xRG76xSFb2AFM0BeNcRtSh2+pg+80TMBALIoeAmdKfhmBKXIQmrSA+1HTryQ
wk+GwneUPpQ5I5koJMYjVRpBY3IAhoEzeXyNeE6YvNRbmTXdmUyh270pBVMun96t
VFN/jtOzcO5hVBBttcRyLMSogZyPcA6hpR3oNkigA2NQ+vCSZ0DS2FJYhUPvl/dZ
7+niRCJQDbgdfAmicQK8kf+KkffgRgl+F8rfnJmpskywwazM5rkUYJyEHd8pq5gW
9CSXHxY7B9jQuii/oVmsS0+QXa2NN+XVjMh+xKNv4RE4beJYXckGS90oG5iwL7c+
Vw/TFP78CZuvDPIU5307NJAnW65A84RNdxO9G8FBFAsUuwG7dJTKesyo0hi3Edcm
aun6NyaD6EvD5AUqqJllo1JhWoZRHlPU2yPvqjiZlk9teUFTgZ53CP1IsY+huJei
XOgXpPM8ugXIgkniSUmtA3eY0ODeZ2A8vM/1E/azbiYCQKsBMkf3i17314AIZf7j
VswJrogIzsoH3u0/TT8UciQDhU/8iGHX3tWgMy+Ds0GHQbEMaSTtE7BIVUGiF7F3
VhMhymsJq3UNMIdCKqxG00EpPzAY/dBMpuOLCgqJG7z5ZVap54YjOxYNDyzzG88c
MoBbdutV5qcqDF0WAWKtzk61U5Z/AK9tg3CCH+Qex3TTYLu9VoaE3MaqKAT8S5+3
R43ha0/uJGiVn2TGe9I9xRT/ykoScLGi4bxpe4rLB5SBLxqYRV4lFpdXuGtFhUTQ
TIlkboNHHJe0PKeLrk4vfjJ+YiH0Km+JI/QfZesJ0XdW7+4w/tOwYFc4LQuXa5QN
LgkByV5bN78hLL+cuoV/Nij4VEbICh+fQPJ/tAYppNirKktx7Zl+PM42RGgaaGLH
D3CKSGek1MbqcCMxLFJQx0ZPR8yiNRdpJspt9SAzqn/ZBUXfs+v7ibdUTG/Fv/6+
hIY4Iu9Wcst9D/iub7UZ+q1lVJELqdPIYuqmfg20j7l8RTvY+S3nsNftBIXXw/CD
rva+8EQwbq0FEcFE+RtR9I7ZzZsM0Zz57mTMuD/nu/mkdzs8uaPP96A51eWNfHNI
uMSzfFJ0Z7OJZPjP9DHYAaowp+/ZW1/x3E667dJ9pLO19ROpRViP+Ssp1PJ8EbK5
X2ih/x1A30RlF2RdbCSsXhskZplnZ2fT3Hjp+ReX+6wVYvXdf8+70XYZXC1quhqI
3QVB9Ja76zZT34LisKbv5G8+kuTMLO+OKychpqjj70nEcmmXefHA3qndQLAKYpvm
aSSUhjVXBC9U3xSRvJ9CS/z/O6THzZa0z8TuDL3C26i3ebpN9D/NMOglWljRJTGF
rEVS7F2B8E69Gh/80fe/UTMMECdFjMytACPg1eV7PntQlShLEmZgm+FOP9ptCTVs
A+rNG0V9j09I197ZaaTlNhF0eEtjRiDf77+b95pteKKf9NjhhSQcpULQAjAnDjv1
8+Grh+8a6PoM9uguJjnXENdr52jbQpjF6YhNIrmnW1/cVn8pAK2EUJIBma53et4K
UUTtUEGy+yzzKGxUdSgX/626wKun1/zM/0LxggKNPINdzMvk3dumSmrc9BnBuEIE
lHxlh/l8yi18RBKn64kfCkAkHn5pwAuVaaUzW9myCkOn8vSRg8C2p/zmtv/kiJm7
4rrJ+QfXhKN/zhQ+wwtboA5a1H9XDtM1KKiE6wxbQcfT58eNfoXZOOkjN+P7zzpy
nYq/IFZg8J8ZcRHoFU8lmHNPS/R4MboqwEKYvJhIJMI1rV45wwa9mYtmkA1Eyy8Z
PlCcbVSPd4UYCmFdsmiMXyoZsuxvv7w8eP02+9ut0tWkDixsOuHwmZtm7XVgSnm5
1k3QvOEhdKqPkcNnsvj3rjSE89VVTUjj9YgW6BEvcgRfaypy9bcuq0FrttfKdXAI
BN3DnLXpELhuoVNCp2kz85UsiebVGqDcaJ1Be1xy3ZiNgzY2hNpGa0id14iryzBm
ta7tuko61p+48etxLQag27EmMGs9/F0ZADg06ohh+BUdhlBMBgELR1XfoESoN1O3
KAQIQ8kMbS9y69TwtM+9fFRPdXvlQdjdm61M8z0RZzvNpbr6LAK8uAfGq8GSv8oi
NLxAZVPZAl5Nut5r+lImX38Ki8FQso6XAcaJqr6UiVJ+p3Qno4yBkOcJAyanBNCF
1FE18eHBiOex2HnCfluxXZksW6ibo98F6xrU2ter9WqadIgjI2JnrfWDzNSfGsWZ
zZz3a6MzDVi/Pr5FKtZIv8WhtHBH2bWC6i2w6nD2nEtzueuIo0KjwnWembFO3l6j
5DOiEejjQk6b7a7zFr4b4UTWQJEqt4hXLrDo+h+cZi6pXtqoR2m36zdW9GpuR53b
57IrT5y5WMFhqJeAFAzslsjScVC54NQFihokAi9OXUzf74asdPw6IZNxBv6qje6k
wY6T1eqvzfECDTMqPw7UwZjJemJcgCtXxeN7LbpUp0xC8q3LkjawGB9zIYmNQMqZ
GM1OJvbubPhY7BZkPRhKYmYbyA0V0ou/vOuCPoD6LTywmKoHTd+AUwExY5iwvcdi
1Ik1Ty2dzdeaVjg4yo+c/W0zvFt9mcgs7zDMJQu2GF6gE6hzECl1QARA+Gt9P/EX
GGHkJXu5jIct6lJCuxpXKRtUnCXagS36010TlPpbPktF67hdJAduT5AlCwG4zJei
EyzN7aM9F5MXGnel0Q7rShAWB6zduqj7Bcx6TNMhFmVbwWCLZmqf0XdJxC4dY8sQ
IZ1UrPEGCnLskVhbF0MEz+kOQGpmT1MiaY5eaf4BkjGJzK0yNw2NdrPAT7oS1zq8
yVTQreJZRBtRkgy40twWgGIASwbA+EW02vlHeDKM5yFBibDZ5UbS4kfHMY67ZfsL
ade0srjOZHDWwRDty4gf8i/javucgFvDh7gMAHmdvvT7ZAGZq2TgeLPkSO4Ykrq9
0ZOLIZu5l8sWssawAfDLUDhhKhSmX0s8u2d+4TotZQcw+xQCw/apcMuew0j8yiYE
EGzzl8TrguQV7ue6QCyubtXc1If2OUg5l6BXuL53FuVclPcIi+HJxtmGX32f1jyg
ZVBI9jEhYqI4dOjuXj8mQhD2H9Ge5P9Ngw02zArN6C+Cz9x99oPBgHSWJwjNZS2E
T71B5usZ3msSpMdm5ohRVFVuctDoLfDSJw3p2teWh7W8Amfi2t+R0Z5jBaPQTPoE
rvBNFVft7PfQFj1pZrbhBhVDRYfUeY6HoHJoHTWVgYBjSBu3Nx7KxyXQfkrGvTzm
cZGp6ihfReHIqqeM6oX9fNjN6fx+SOLRaGZnXG530zXaJ+LnrpzbKApJXTWJDF7X
g2HSBgL/OFC7ihtSGKl+eQ3lcSTpk9w28qDGvIFk2exJl/w/XlMCGk0U4cU0DAjw
hmU6NxxRBbrPPLmzuuaB+a0OMZq3uR94csKfur9p5wEXX7FsQ9RQDdKAHhPPgnsi
lsiNqYIPldVIjm2Bx9esV331wekPAwLXO6Ms1Cl/Xo+gMMcNDBbnQ9377BWc5uVL
QBEs3Lpsfd0uFQ5Xpv32w9Y59NuhjLG0BiELdH7bFe5JkDmDMnBWqkcHhtomccoQ
FkjqGy2Q45TqZ1w3JhcvTqQjdK+ll/rP7m9tGs//C6pxQo1P+xHFRf54xPpbbb6W
2q2TBa0H5oT/msmwDB/UPaepMSvOiuFHFVT5Y9JjTatjHhzq8wB06jCngCEOtGvz
i9xLeLjZ/26Iz1KVOhNKWFIh5ntPtK2W9/ciJO++97BGePBHM38HqZe+P2oPawpD
wez8MI+fOvlKPdLXrLE6r4U+ZmE1vf4SWn8pRJPM05hLquXBmk0SEbTrNI+63kEL
SHuF2D39tupleZZuh1y3RXdq2QuMNLbOaCSxwqDcv9vhB8jDgBkS9xQM3sM/Bo0Z
By+WPk1L6ShFElUAFBcU9QjX9WpuZ91MOPkMmMoHVxfBO3Xgkl7OwwoTuK3q/8TY
0L+O3owleRtgokye5Uf1E9z5WG5O/YA3bLw6IVIe6FQgQh+RNxF5b8X8QhGpNRzo
Lrqkuu0WwM9gf1ReacmM8duAK9D6CH41bCoaSKsrNBOwUJw4QmuukgA831g0d3N6
steniqAGj4KCk9d4XLzsTzLhHzoTPddK1WqUJCJrIbT+75y1aPVxYkrmSgXj869g
DRSYE77fNHrwCOTnByj+iIbTVK3+kKGBm4tPNot+0CQBj52BFudZHWgrxcHIb1Sv
lJL/jlQ8fa0sQVBsrzEYL8OS5ZFs7i/0z/I4dcKC0f//nqOqGaZL6tPJr2lPd6wK
x3l/QifWn85ljIX2Q+zu8bkb8TNp9G8IKk1M0Q8NCjI9Uu7dIVyz4SQAfmUYL9F1
P4KL/QtLqcIrqrYJyqbskXVyt6FsPNbbnEy7Ttx9M0MHjZdb3nsJ6RMHbgnSK6Xm
VZr3bkhlDKEZsiZ0b2mv0SJ1fosdeM7cfH2XEo+k1YxuvfGtIVtFmGpNIUbKSljG
IwBr6ahMgu/lt4sJS3QK3iMxkBrONULGupL5Uek1lVfcuJ27wU9AlsSRsPvEI8hB
pW1kAzLxhnXzXTYlItu1f4z0uWEoPO0cUVse1AFfYWtGYtI5yv7MeIOb9qNEdor8
5mt4bz56oI62K2xc2Nps2a/kcCKIuy8GVSpHStSDSkvbVM6MWmJzhKdgt51cF5y2
kPyjV134tcJvIysLl+5O34R92NVxr/9dxKviUp0AiDp//oKXoqKl2+mV5PXKK0wY
m1AdOavYhDjOQ6R6Vbvpf/0RNqc0m+l0EDtEphquP2Tpdq4HdNEgzreeJyx13oDE
5yUg0bMrILO8c+GGfdXvFAztAFm2eaSQ/k7rzoaE7B4e2dw260uIi6Ch4xzIZh+r
XjV/hiqr7lncaMY7iEU+wjSWMZxUo+sjvmXwfbD22s4+5nYnZxkiDORYnduixBPO
EFJ8+3akLTFfz0hkE7eGdy7VDVP5Gq7k/CYuseKGJ5yFMjU+CvC4EzSIbq5g6TIW
rHf42VDsBnZkredGIvChw5SmUquomxM0G87xD2cqQGHYyCWPoa7oFu5jFnegub+b
FxSu2GNPJQJDfhDKabhIFSx0kuuFOAy+02isfYLoJzhc0wPRG76uZ7GKPjwvCNX7
5km1A3bHZuXW2/bt5zdmgEeDxevKFvFSwDBPh0ykDdr9pkP8tpvq+mxxGkgFyJdl
vUpN8FrjDvsQLPR5jTq7dNUZpMchU1qhrZ0wiSfDjSxkeUjRVEZCbCr8J8Qpgh96
6q85qirsU8IOdVKltcbqbzIN2zKcunwvlYgeBkzRPyaIt2zsU48uOedfdPbmEC5P
vfhi3SJ2Q9TCI+XyNPLu77ZGEAm0UF0Y2Jb2HYo5WFroUu5w+QjZxpD+nwLq8HUq
QxD53oYTbUP2+3pYqhXtP3pWSdHjqsrk/yKVAwTDGccDfsy0n69rQUfiPe7XH3d8
2Itjo9E+cqp/StGci6+dPskmhGc/2lEGYKIOoB6g22rKwYkw3CYXgUVxPn31dV58
m6SD5gcyMOTdQ20k8gtE/Dm0Z7hi1Fhb6l/07rR/zfw725Ui83g8MK9knmv7BahS
rEFwSuRXU4kUkZNHW2ZJah/nAv4k7E3dt1BAag/8cjYDTC3JBP+RJRzzXYJwfXtR
lA50x7pr/FLRDPOeKKAHNCh6fWSeid8rQEU1PgcU+rylJB7qvRIMhgGJNjLVdmmF
8OlxQIz9yiiPDp9vbspYmIgOV+O4A8Ph/iykTPQNVLpN1tumss5qIhSpKWt4d/Vt
01j0zJ0OF8lufQjpR16ZKYjnUV2zMk17ocSC0q3U1GgLIVolZyPTyimTe82rN6xt
EiKbEzwOSzjVbPkGosNzsFuubvMgxRtoQuFG5RPxI6ogFcNrkdEZxbcrxK52VlmW
6nfOnVuNhbo77Vnw1K5M+oBkX/r/lfZKYqlkeSVi1tPxghBDJwDZ+Vznd9r9U8cM
hxSeUskXs15azAxEkQBUxSL0Y/RpXc18nKVa32jbY7Ocjw3de95sp69UvjVfhcW5
/NnGf6IEyioah/emfJI+dlKe26gNNehnPl6d9ERHhGn7oWBxfn9Svu/06rs1iGBc
EHo++0av/+kvAytpeX6/wH+nlLN1UQY9LEcqVW0CLkY03TOdEh+cbBNJhNUNWAxU
RFN/jx1z+77Wl+7ayKWLYAs6xGMgHYyO84QnwxojuMyfyOB/BoI4PYFurzUTF2qi
CBFtMMh7PKHoQk6pkzD39cPHxgHQo45tGn7sZ507vMxstq8/H/B9G+nWpwdyO76I
PNiEqNvrrk09jJ7fpaaMipNhCaxCjAwPgdWF/n/KSa3Bc6TuKwpNI4AXQoadR0bO
6r2a9rWzzSflUUOo+FtGkX9XPzvzoRE/9SHl7+P1jcKU7BToljl243dREjPD84ES
/EhreBg9zrAL5Py3VdAmsYAcg0jTnZ5yJgGAarAImIKgb9BwCEZQFcFClEcX2qTL
dMpBhDQxQlqM0siJLjNBwDERlVCMlJ4YDa2pBQPo1ie4uVaHForQzkq2+30I8mzB
Kt+2Bh9/k/JTOO+VGk80q3iZxqecSaJF7ekZ9FjLi7AMU/UAkXS1OT/nRTYxWxcQ
XVh01PBeZdEPVeKqGIZIPUrtb8BOPrJqOaczRvjM+s8ndlSb0ReQtiHcCl3E+cEP
5uFMORmY45IVqQlXE1DwPXyd3pR/x8RUTDJVzPCpJSoP0pqoZlRlSrpccEQ6uNtL
P/U78wcpuBRzNKy0+ryt+yJ0PbcTZHpKm3QEn4b+fGKNR3URhxSs2FhwmigF2Mnj
oPRCpAX2FsyxpQiTrr0uFrJoDhl92DgsgYK3sYOrIEKgJztyhyWwvoWO+zf1qBw5
PKP0bYbXft2lfMI7KgdbfzlYZ67j0PI49NybaNNra1VYQH3JMti/+zCtrgMG0wTH
AisWiza352UvrHyKdPL76nyrrUqWViRR/LhiwfCCL75JPMTE00KDEQJDHDeZ6QAr
eJu7xJ8qDrdKcQQzwo5eIGcAqGgXsUPzDGI7mHA+HrN0KTC5bZylgZzgx/3ZK8yd
oXWay8HS3BE275IyCFYipWIjodiIb4mNjsqMSZFu1pxmsD60pJ4WBxSD4hmlrBoC
MguvkgcJ35buntXuOTc/wYNGlIimI2rsovUVQA7gmNL1wu1+lHKmDFCH1EyK7mDw
uI5GNSlUcCTlIVS5pcMJ0tjZ8vqGAkolNOqlW75n6VDfVKW8J5+M8X3KXS/6qBsI
tl35KWa6MgNaLXDCK1/n9UORwIRdmLpxLQ+0Riulu5BKl+OGiGC30s0eIJzWDUm4
H0I/cFH3UIQCJDhRcrq3ZfpiTE6q7c4u8DXh0i6FMxPsZE7yT5VoPK85O2q4ZE7k
BGfcUUHw8ao5nnfNs25fsEEgKtbXZFghOwD0XfgU0d1IxiTZsnbQVLscBPKIAnXk
OcOpMX7wO7yLJs3ENVcrzdnyo92IjTzEZ1O60DHSEjdkyByB1JlAydo5ZwyFZIaE
tFsXc2QMdqC74Cwgf75VZCktQ2Em8E0qjXjTJve+04t+P7n0vB/d4P23lHnpdDDD
4PYR7G/uCYxBKRtM55FRQQlaE1hzDb4O2mg89c6DIgsyHNAzM9ZSVuydYrbKir3N
M8Z8k4okCX1SAFLY2gAGa49l8HfnJ0H0mrgbpC/xgqK55bQzEK5oI9QLnWz3PIkH
IOMMXITZQETViQ3mftDgjpWbbmCfEbIkv2cvY405lwqkaXEj1X7Sd9t9W32odPyv
OSvBAT60Lrb/CBkfgrDV1sML+kxOJVkbwVe/vPU74w6CorSSspI9br5SIFgEBcns
8TuPNB5xHLz+LwOmOOUE0ESlLg+ixVJ/rd8VRxMnkrjGiWDJrl+V0+wa5nUSVy9I
c2gVjBEmJciZUbd+ZJZYIHji/uEQdOlKuAdHwggZItpZldSKyWZe8C5c6fL3WXLC
5i1IB8AyfIRv+uwQlaht1lralJ0MQ+8oW4tHFSwi+GnSNwtz7kSl520QsJH7iUNc
DstolU/syOGc3k+AbLjACuKOIZTdMO7lhCgPpc7Uv/gMDNO9N8KFT3RcmgDP5cgs
KL33xjQxcecYg39Y72JxSAEdcV9oN2aimJxFEgGLqeZYFSKveAHSFWN6ljiPtSTD
b05yZ6uxJUUv9kDUoRrxQsGK8486YFKNEy4rSAUzTPnkaILhsg8qu+dwdDhKvZye
BvYBtpj2OFFZKVgnzTSjS+qUZzhUjzlGcca/WxNGIOHwEvGp7CNb+oijVaR53SEm
dwPyMjnUDFNgXfUKBCyzGiel1sflWdIF5VKT2VbGzqkEfKTZrQ1ezBid8z9qYi1t
Rzh0Ks+0Wd3O1BWt2fSjplYhOHcYvNW+B5+dhN4CH3LIQl4iiok8agddmMEC1Hxm
cxQf4nRzVDhzPd9e1gU0oAY+cadMFtVfSdK8x8xxu0mF2THAvwq5fbgM+qrli06G
qoWVHB571ncrZxC1mkvchdwe3QZaw/1mQycqpiWoxw6HSA78IsUGiKVsjvgz0pmc
z2lmSh8eeYkqErPbYBLiZeYsCPmlzHtUgepXi3s1EhWYiHx/aKSaWevdqbHjUnFv
`pragma protect end_protected
