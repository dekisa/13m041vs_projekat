-- system.vhd

-- Generated using ACDS version 17.0 602

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity system;

architecture rtl of system is
	component system_cpu0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(14 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(14 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_cpu0;

	component system_cpu0_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_cpu0_jtag_uart;

	component system_cpu0_ocm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component system_cpu0_ocm;

	component data_gen is
		port (
			clk             : in  std_logic                     := 'X';             -- clk
			reset           : in  std_logic                     := 'X';             -- reset
			bus_address     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			bus_read        : in  std_logic                     := 'X';             -- read
			bus_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			bus_write       : in  std_logic                     := 'X';             -- write
			bus_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			bus_waitrequest : out std_logic;                                        -- waitrequest
			irq             : out std_logic                                         -- irq
		);
	end component data_gen;

	component system_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component system_pll_0;

	component system_mm_interconnect_0 is
		port (
			pll_0_outclk0_clk                            : in  std_logic                     := 'X';             -- clk
			cpu0_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			cpu0_data_master_address                     : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			cpu0_data_master_waitrequest                 : out std_logic;                                        -- waitrequest
			cpu0_data_master_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu0_data_master_read                        : in  std_logic                     := 'X';             -- read
			cpu0_data_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			cpu0_data_master_readdatavalid               : out std_logic;                                        -- readdatavalid
			cpu0_data_master_write                       : in  std_logic                     := 'X';             -- write
			cpu0_data_master_writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu0_data_master_debugaccess                 : in  std_logic                     := 'X';             -- debugaccess
			cpu0_instruction_master_address              : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			cpu0_instruction_master_waitrequest          : out std_logic;                                        -- waitrequest
			cpu0_instruction_master_read                 : in  std_logic                     := 'X';             -- read
			cpu0_instruction_master_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			cpu0_instruction_master_readdatavalid        : out std_logic;                                        -- readdatavalid
			cpu0_debug_mem_slave_address                 : out std_logic_vector(8 downto 0);                     -- address
			cpu0_debug_mem_slave_write                   : out std_logic;                                        -- write
			cpu0_debug_mem_slave_read                    : out std_logic;                                        -- read
			cpu0_debug_mem_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu0_debug_mem_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			cpu0_debug_mem_slave_byteenable              : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu0_debug_mem_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			cpu0_debug_mem_slave_debugaccess             : out std_logic;                                        -- debugaccess
			cpu0_jtag_uart_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			cpu0_jtag_uart_avalon_jtag_slave_write       : out std_logic;                                        -- write
			cpu0_jtag_uart_avalon_jtag_slave_read        : out std_logic;                                        -- read
			cpu0_jtag_uart_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu0_jtag_uart_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			cpu0_jtag_uart_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			cpu0_jtag_uart_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			cpu0_ocm_s1_address                          : out std_logic_vector(10 downto 0);                    -- address
			cpu0_ocm_s1_write                            : out std_logic;                                        -- write
			cpu0_ocm_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu0_ocm_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			cpu0_ocm_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu0_ocm_s1_chipselect                       : out std_logic;                                        -- chipselect
			cpu0_ocm_s1_clken                            : out std_logic;                                        -- clken
			datagen_bus_address                          : out std_logic_vector(7 downto 0);                     -- address
			datagen_bus_write                            : out std_logic;                                        -- write
			datagen_bus_read                             : out std_logic;                                        -- read
			datagen_bus_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			datagen_bus_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			datagen_bus_waitrequest                      : in  std_logic                     := 'X'              -- waitrequest
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_001;

	signal pll_0_outclk0_clk                                                  : std_logic;                     -- pll_0:outclk_0 -> [cpu0:clk, cpu0_jtag_uart:clk, cpu0_ocm:clk, datagen:clk, irq_mapper:clk, mm_interconnect_0:pll_0_outclk0_clk, rst_controller:clk]
	signal cpu0_data_master_readdata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu0_data_master_readdata -> cpu0:d_readdata
	signal cpu0_data_master_waitrequest                                       : std_logic;                     -- mm_interconnect_0:cpu0_data_master_waitrequest -> cpu0:d_waitrequest
	signal cpu0_data_master_debugaccess                                       : std_logic;                     -- cpu0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu0_data_master_debugaccess
	signal cpu0_data_master_address                                           : std_logic_vector(14 downto 0); -- cpu0:d_address -> mm_interconnect_0:cpu0_data_master_address
	signal cpu0_data_master_byteenable                                        : std_logic_vector(3 downto 0);  -- cpu0:d_byteenable -> mm_interconnect_0:cpu0_data_master_byteenable
	signal cpu0_data_master_read                                              : std_logic;                     -- cpu0:d_read -> mm_interconnect_0:cpu0_data_master_read
	signal cpu0_data_master_readdatavalid                                     : std_logic;                     -- mm_interconnect_0:cpu0_data_master_readdatavalid -> cpu0:d_readdatavalid
	signal cpu0_data_master_write                                             : std_logic;                     -- cpu0:d_write -> mm_interconnect_0:cpu0_data_master_write
	signal cpu0_data_master_writedata                                         : std_logic_vector(31 downto 0); -- cpu0:d_writedata -> mm_interconnect_0:cpu0_data_master_writedata
	signal cpu0_instruction_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu0_instruction_master_readdata -> cpu0:i_readdata
	signal cpu0_instruction_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:cpu0_instruction_master_waitrequest -> cpu0:i_waitrequest
	signal cpu0_instruction_master_address                                    : std_logic_vector(14 downto 0); -- cpu0:i_address -> mm_interconnect_0:cpu0_instruction_master_address
	signal cpu0_instruction_master_read                                       : std_logic;                     -- cpu0:i_read -> mm_interconnect_0:cpu0_instruction_master_read
	signal cpu0_instruction_master_readdatavalid                              : std_logic;                     -- mm_interconnect_0:cpu0_instruction_master_readdatavalid -> cpu0:i_readdatavalid
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:cpu0_jtag_uart_avalon_jtag_slave_chipselect -> cpu0_jtag_uart:av_chipselect
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- cpu0_jtag_uart:av_readdata -> mm_interconnect_0:cpu0_jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- cpu0_jtag_uart:av_waitrequest -> mm_interconnect_0:cpu0_jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:cpu0_jtag_uart_avalon_jtag_slave_address -> cpu0_jtag_uart:av_address
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:cpu0_jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:cpu0_jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu0_jtag_uart_avalon_jtag_slave_writedata -> cpu0_jtag_uart:av_writedata
	signal mm_interconnect_0_datagen_bus_readdata                             : std_logic_vector(31 downto 0); -- datagen:bus_readdata -> mm_interconnect_0:datagen_bus_readdata
	signal mm_interconnect_0_datagen_bus_waitrequest                          : std_logic;                     -- datagen:bus_waitrequest -> mm_interconnect_0:datagen_bus_waitrequest
	signal mm_interconnect_0_datagen_bus_address                              : std_logic_vector(7 downto 0);  -- mm_interconnect_0:datagen_bus_address -> datagen:bus_address
	signal mm_interconnect_0_datagen_bus_read                                 : std_logic;                     -- mm_interconnect_0:datagen_bus_read -> datagen:bus_read
	signal mm_interconnect_0_datagen_bus_write                                : std_logic;                     -- mm_interconnect_0:datagen_bus_write -> datagen:bus_write
	signal mm_interconnect_0_datagen_bus_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:datagen_bus_writedata -> datagen:bus_writedata
	signal mm_interconnect_0_cpu0_debug_mem_slave_readdata                    : std_logic_vector(31 downto 0); -- cpu0:debug_mem_slave_readdata -> mm_interconnect_0:cpu0_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu0_debug_mem_slave_waitrequest                 : std_logic;                     -- cpu0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu0_debug_mem_slave_debugaccess                 : std_logic;                     -- mm_interconnect_0:cpu0_debug_mem_slave_debugaccess -> cpu0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu0_debug_mem_slave_address                     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu0_debug_mem_slave_address -> cpu0:debug_mem_slave_address
	signal mm_interconnect_0_cpu0_debug_mem_slave_read                        : std_logic;                     -- mm_interconnect_0:cpu0_debug_mem_slave_read -> cpu0:debug_mem_slave_read
	signal mm_interconnect_0_cpu0_debug_mem_slave_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu0_debug_mem_slave_byteenable -> cpu0:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu0_debug_mem_slave_write                       : std_logic;                     -- mm_interconnect_0:cpu0_debug_mem_slave_write -> cpu0:debug_mem_slave_write
	signal mm_interconnect_0_cpu0_debug_mem_slave_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu0_debug_mem_slave_writedata -> cpu0:debug_mem_slave_writedata
	signal mm_interconnect_0_cpu0_ocm_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:cpu0_ocm_s1_chipselect -> cpu0_ocm:chipselect
	signal mm_interconnect_0_cpu0_ocm_s1_readdata                             : std_logic_vector(31 downto 0); -- cpu0_ocm:readdata -> mm_interconnect_0:cpu0_ocm_s1_readdata
	signal mm_interconnect_0_cpu0_ocm_s1_address                              : std_logic_vector(10 downto 0); -- mm_interconnect_0:cpu0_ocm_s1_address -> cpu0_ocm:address
	signal mm_interconnect_0_cpu0_ocm_s1_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu0_ocm_s1_byteenable -> cpu0_ocm:byteenable
	signal mm_interconnect_0_cpu0_ocm_s1_write                                : std_logic;                     -- mm_interconnect_0:cpu0_ocm_s1_write -> cpu0_ocm:write
	signal mm_interconnect_0_cpu0_ocm_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu0_ocm_s1_writedata -> cpu0_ocm:writedata
	signal mm_interconnect_0_cpu0_ocm_s1_clken                                : std_logic;                     -- mm_interconnect_0:cpu0_ocm_s1_clken -> cpu0_ocm:clken
	signal irq_mapper_receiver0_irq                                           : std_logic;                     -- datagen:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                           : std_logic;                     -- cpu0_jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal cpu0_irq_irq                                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu0:irq
	signal rst_controller_reset_out_reset                                     : std_logic;                     -- rst_controller:reset_out -> [cpu0_ocm:reset, datagen:reset, irq_mapper:reset, mm_interconnect_0:cpu0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                 : std_logic;                     -- rst_controller:reset_req -> [cpu0:reset_req, cpu0_ocm:reset_req, rst_translator:reset_req_in]
	signal cpu0_debug_reset_request_reset                                     : std_logic;                     -- cpu0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                                 : std_logic;                     -- rst_controller_001:reset_out -> pll_0:rst
	signal reset_reset_n_ports_inv                                            : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_read:inv -> cpu0_jtag_uart:av_read_n
	signal mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_write:inv -> cpu0_jtag_uart:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu0:reset_n, cpu0_jtag_uart:rst_n]

begin

	cpu0 : component system_cpu0
		port map (
			clk                                 => pll_0_outclk0_clk,                                  --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,           --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                 --                          .reset_req
			d_address                           => cpu0_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu0_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu0_data_master_read,                              --                          .read
			d_readdata                          => cpu0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu0_data_master_write,                             --                          .write
			d_writedata                         => cpu0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu0_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu0_instruction_master_read,                       --                          .read
			i_readdata                          => cpu0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                -- custom_instruction_master.readra
		);

	cpu0_jtag_uart : component system_cpu0_jtag_uart
		port map (
			clk            => pll_0_outclk0_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                           --             reset.reset_n
			av_chipselect  => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                            --               irq.irq
		);

	cpu0_ocm : component system_cpu0_ocm
		port map (
			clk        => pll_0_outclk0_clk,                        --   clk1.clk
			address    => mm_interconnect_0_cpu0_ocm_s1_address,    --     s1.address
			clken      => mm_interconnect_0_cpu0_ocm_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_cpu0_ocm_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_cpu0_ocm_s1_write,      --       .write
			readdata   => mm_interconnect_0_cpu0_ocm_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_cpu0_ocm_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_cpu0_ocm_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,           -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,       --       .reset_req
			freeze     => '0'                                       -- (terminated)
		);

	datagen : component data_gen
		port map (
			clk             => pll_0_outclk0_clk,                         --            clock.clk
			reset           => rst_controller_reset_out_reset,            --            reset.reset
			bus_address     => mm_interconnect_0_datagen_bus_address,     --              bus.address
			bus_read        => mm_interconnect_0_datagen_bus_read,        --                 .read
			bus_readdata    => mm_interconnect_0_datagen_bus_readdata,    --                 .readdata
			bus_write       => mm_interconnect_0_datagen_bus_write,       --                 .write
			bus_writedata   => mm_interconnect_0_datagen_bus_writedata,   --                 .writedata
			bus_waitrequest => mm_interconnect_0_datagen_bus_waitrequest, --                 .waitrequest
			irq             => irq_mapper_receiver0_irq                   -- interrupt_sender.irq
		);

	pll_0 : component system_pll_0
		port map (
			refclk   => clk_clk,                            --  refclk.clk
			rst      => rst_controller_001_reset_out_reset, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,                  -- outclk0.clk
			locked   => open                                -- (terminated)
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			pll_0_outclk0_clk                            => pll_0_outclk0_clk,                                              --                    pll_0_outclk0.clk
			cpu0_reset_reset_bridge_in_reset_reset       => rst_controller_reset_out_reset,                                 -- cpu0_reset_reset_bridge_in_reset.reset
			cpu0_data_master_address                     => cpu0_data_master_address,                                       --                 cpu0_data_master.address
			cpu0_data_master_waitrequest                 => cpu0_data_master_waitrequest,                                   --                                 .waitrequest
			cpu0_data_master_byteenable                  => cpu0_data_master_byteenable,                                    --                                 .byteenable
			cpu0_data_master_read                        => cpu0_data_master_read,                                          --                                 .read
			cpu0_data_master_readdata                    => cpu0_data_master_readdata,                                      --                                 .readdata
			cpu0_data_master_readdatavalid               => cpu0_data_master_readdatavalid,                                 --                                 .readdatavalid
			cpu0_data_master_write                       => cpu0_data_master_write,                                         --                                 .write
			cpu0_data_master_writedata                   => cpu0_data_master_writedata,                                     --                                 .writedata
			cpu0_data_master_debugaccess                 => cpu0_data_master_debugaccess,                                   --                                 .debugaccess
			cpu0_instruction_master_address              => cpu0_instruction_master_address,                                --          cpu0_instruction_master.address
			cpu0_instruction_master_waitrequest          => cpu0_instruction_master_waitrequest,                            --                                 .waitrequest
			cpu0_instruction_master_read                 => cpu0_instruction_master_read,                                   --                                 .read
			cpu0_instruction_master_readdata             => cpu0_instruction_master_readdata,                               --                                 .readdata
			cpu0_instruction_master_readdatavalid        => cpu0_instruction_master_readdatavalid,                          --                                 .readdatavalid
			cpu0_debug_mem_slave_address                 => mm_interconnect_0_cpu0_debug_mem_slave_address,                 --             cpu0_debug_mem_slave.address
			cpu0_debug_mem_slave_write                   => mm_interconnect_0_cpu0_debug_mem_slave_write,                   --                                 .write
			cpu0_debug_mem_slave_read                    => mm_interconnect_0_cpu0_debug_mem_slave_read,                    --                                 .read
			cpu0_debug_mem_slave_readdata                => mm_interconnect_0_cpu0_debug_mem_slave_readdata,                --                                 .readdata
			cpu0_debug_mem_slave_writedata               => mm_interconnect_0_cpu0_debug_mem_slave_writedata,               --                                 .writedata
			cpu0_debug_mem_slave_byteenable              => mm_interconnect_0_cpu0_debug_mem_slave_byteenable,              --                                 .byteenable
			cpu0_debug_mem_slave_waitrequest             => mm_interconnect_0_cpu0_debug_mem_slave_waitrequest,             --                                 .waitrequest
			cpu0_debug_mem_slave_debugaccess             => mm_interconnect_0_cpu0_debug_mem_slave_debugaccess,             --                                 .debugaccess
			cpu0_jtag_uart_avalon_jtag_slave_address     => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_address,     -- cpu0_jtag_uart_avalon_jtag_slave.address
			cpu0_jtag_uart_avalon_jtag_slave_write       => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_write,       --                                 .write
			cpu0_jtag_uart_avalon_jtag_slave_read        => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_read,        --                                 .read
			cpu0_jtag_uart_avalon_jtag_slave_readdata    => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_readdata,    --                                 .readdata
			cpu0_jtag_uart_avalon_jtag_slave_writedata   => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_writedata,   --                                 .writedata
			cpu0_jtag_uart_avalon_jtag_slave_waitrequest => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_waitrequest, --                                 .waitrequest
			cpu0_jtag_uart_avalon_jtag_slave_chipselect  => mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_chipselect,  --                                 .chipselect
			cpu0_ocm_s1_address                          => mm_interconnect_0_cpu0_ocm_s1_address,                          --                      cpu0_ocm_s1.address
			cpu0_ocm_s1_write                            => mm_interconnect_0_cpu0_ocm_s1_write,                            --                                 .write
			cpu0_ocm_s1_readdata                         => mm_interconnect_0_cpu0_ocm_s1_readdata,                         --                                 .readdata
			cpu0_ocm_s1_writedata                        => mm_interconnect_0_cpu0_ocm_s1_writedata,                        --                                 .writedata
			cpu0_ocm_s1_byteenable                       => mm_interconnect_0_cpu0_ocm_s1_byteenable,                       --                                 .byteenable
			cpu0_ocm_s1_chipselect                       => mm_interconnect_0_cpu0_ocm_s1_chipselect,                       --                                 .chipselect
			cpu0_ocm_s1_clken                            => mm_interconnect_0_cpu0_ocm_s1_clken,                            --                                 .clken
			datagen_bus_address                          => mm_interconnect_0_datagen_bus_address,                          --                      datagen_bus.address
			datagen_bus_write                            => mm_interconnect_0_datagen_bus_write,                            --                                 .write
			datagen_bus_read                             => mm_interconnect_0_datagen_bus_read,                             --                                 .read
			datagen_bus_readdata                         => mm_interconnect_0_datagen_bus_readdata,                         --                                 .readdata
			datagen_bus_writedata                        => mm_interconnect_0_datagen_bus_writedata,                        --                                 .writedata
			datagen_bus_waitrequest                      => mm_interconnect_0_datagen_bus_waitrequest                       --                                 .waitrequest
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => pll_0_outclk0_clk,              --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu0_irq_irq                    --    sender.irq
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu0_debug_reset_request_reset,     -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu0_debug_reset_request_reset,     -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_cpu0_jtag_uart_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of system
