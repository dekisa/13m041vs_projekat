��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&|J� ��
#P�}i�X�>^�m _�lNf9B�]0#Nd$El�0.� UW&��*=�%�N1�zITDR3��0@��� f��;Vee�s��ő���'k]��u��>т���e�$	����G�����l��,��ǯ��	��Z���(ͪN�y��j�P��Q�������aϛ���0��up~�B�V(�3ɬ�����	3���7%a5c�^�/k�,�����a�)0)����Q|
ɻ��¨$l0㛳>���{���i̤ǔI3|`��9*��lK���Z�7�O�-�%�
è��.w?S`�{�)\T�逥2;v���WVlɖ��R�z=%E�׌�,�MK��x3#*i��bE�z�b+z�����0f!����$$A�"���zE����G�DήuZ(��6��Ĭq�$fDh�2<p�����+wG�q;USr|�3z2���V�}�8��J�Ʒ$��^�@\o�Q!GI"G��9�6��@s�bF������9��̗w����H������5c���ױ0��&];��䑂�5Z��.�D4��@ͱ0�������ֻt@��kȓc	�ċ��=rc�?�e����p����(:���nFY������@�k֌����e$�����S0c�UݍF��7:א�S��]����y��&�P��F�L�3���4ql�㶙�*�x��������"�g���Peо���I�<��Jb��;�wo�C]���`��E͇�f��͙�&�{I��fזe���OyI	����֜?���V�o�8��a�!6}�ݲ�h�jU;?ë��0*ȴZA�t6<P��wk	�2WO�����RF�m���ʯ��h$}�(4�0`��׶�U��r�Z�m4P�Y���6�G�� S�4�P�{�0�̷4��O��v�s�hB��EdE4���ȟ��5tZ|EX�6Ӡ~� �z���h�z��b@��!�'�T�EX���0ހ���{�X6�xoy�>�*ſrU[�@��-��j(�=x�2U&�B�T)�tzb��dr=VU����h��s��
���Z�)���5�)�y�;�����t���_��ܙ��\o�@Uq�ـkr}.�6*H�e� �3�V'�cr�_���L��iz�ku�w�T*��g�7�uf@��;g�F��C��ۓ7�����'#�Mu��P�x)b�<�s��`ۦ����jԌ�j{�p���@�����H���ׯ�b�����ϡj�e��
�i��ň>LE���0�3b��� A��=E�%�X{�	u�2.��g��p��.qYj[���<������sa�F��G]kYcD`G`��q�����mnj��h��?�5�#�crK?As6s8�kO�UM�|q��_Q�T3eZЭ�x���PZQ�ǫS8ד�Y��N��9��e�"*��3����gt<����ed-��t�F��Q�
c��8y ��Q���ON�/_q��H
9���2��F�a��ιc{-N�*r�N��ng�86��G����d�s9�^R���U������t��P3i���_W��?��M3~�H�q����ug������_
B�)Wy��.��O������(}�!�-f{0�~t��RH&����J�{�����y�[v��ϝq�����6��]w*�t�D4p��!��uq	p-D��)�*���ʗ�&*�f��dÌ���� 1,���8t���*��H�S�J���W?'gs�`)Hz-�T\� [G�����5wwv��R7��T
��˽5�HѶ!I;���W�rw4w�ik�*�$V��9l��R�豌�κ�S�"6����
�l�����FzR>"w1h�o!����"�[ �^st�
��,�4����We���m�I�I���e���#R* i�]�:����饬�UZ��g}Aġ��-S�׬�^��7Q�9%n�A�nG��m�˙)���(�ꇻ{'���Qlu�[����-YD��}k�� 1�9I1�oጿ��e��4�I�M���)��z ��)�C²@� ���s��y������1���P��/�f8���_���#��q�f�ݾ0Dd��:��I\��/Y���Y»ٶ��e�Q}J,�R�C0��[J��+��qX�M#��@��kuh$���!+^�O�tc�Apd_ȧ�滧���J�rJ5����U�׏���*�p�	������B����a��ߣ��Ł��>"�Ih�p*�#Ȟ���#C�p�0FEI�䨯
�s[Qre��p٘4��0�Q�)�$�Y�=
�m��I���(�r�����S_����J��oHgҗ,
�uL����ݳ+o��s�5�NMAR�|�;7����PC?���&�(l�<���r�m���<���tk��9�)\r�{�#$ ҟk�M� e��8�*�����	R�D`#��$O�q���6��N%��+%�c�quj]m��8�� [ƌ�!�����뚯a|��:]��D��������������� �r2��L�ɵ�j�.P�l�{��dx`"�Y?�'�����;Y�;]���&� ��}��&�(5Q{ ���Y����p|�iī��`��؇��*J/H�6��P�M:��!rX(�;������"��'yxPkk�����ͻkQ�'�~-
�E�h�&��Y�}���4�<��x��J�����汒MEU_+������3��e��/���b�8�<�1A����
��>7�� e��-����ir+#:�^*�'�?1��{R�W
��$�8�hEdŉ��{W�/�k���]���b6q�:|�F�W�C@,� ���u0s�VBQ�9�P�_�n$�W�5_X�~��z��I�"����k���q3�b]ի��b��Z��j�'m$��"��J��=b����y[�uJm�x&`�9�΢��=��T��4/�K9|��P}eJ}W�E�a�}Ucӭ�m�%s�����_V�4�О=4�l@`f}���`m�����<{C����_��Td���v3]$��sC�4���v3�Q'�؟m*D���	���n�-��&xxpߛ���"��-��nÑ�͎�&!B��Xp��=gp�$Q
�O�!��iVr����D?�V��B,��oN%�.�ԥ!����N
`w7����8m�+�6E�x�7��.7��� 1�@.��p�iJ�-���	��k��[*uE��ʺ�PY�*c�Slb�	^8ua���,26����,���N�!�G���r�ij ^�sɛ늭�کށ��S�f�]>`�/��x�+�/mr�?L�o�b�W2�]��M�$�\|�Н)"���K�N�L�kR#��%�
�[�Js�pж���rc�тAǣݜ���t|)�Z>��|~���q�8�B�YX;��X��چ��[�T��c��w�8"�o7� �h,cq^F�t�Y5�Q�9.�"Ž��i� .����>)%��gJJpd�þ���h���ڽ��'9q�MѰ��4���^ȅ�=M)�����P<��P�.\x��T����I
)�>�^�x��R��@�q���3�bWiW�~���������t�!~��������.�.�;C�}��iO��Ёr~�"��	^�=�Л�����V��XЎ6F�1��j�}TGWW��5��.�����F�/ib�ۺo��KUo�� %Of{/�v�V�q|�g���3�}-c�cR9Q�h��+���~F�������^��\f	3�V���~����R��%1v����=o.��P=���}	V�X��� ��ZD�p�\&X��N(�
Ǆ�R�a��e�R��h����� �wW1
��`Q(��0*��ijA�PK{,T�l�`f;kU�=XR�D�Z2 ��>	�ޥC�3(`V|fxk���:ѕ+����H�EA�KX��?b�<(�=1�9��#���`��|���|
�aB �W��c��� �<�f��l�W���C%m"Ts�Mt�0ի&�ed�\�ms��+���Ђ�>���㍳�10���*v?����1F�I~��u�YI�:�])D�y�超p��?�Z�I����&�9��q:e�daeaDVr0M9xz�j|0�q�R�N�VU[��$k������xX�ǩ+��.��1�˕��a#Pu{zW!�J���5��{�0{�#'��Fz�
,��ꕉ�-E`�L�� -��Ŝ�!~4ޠ`�
<:^�-�bݢ�㦄�Lt�Vj�2Xxfv��ZۂZj��}����˯���L���S�f�4�緘J����w'�w��^%}ʁ�>�*en���=�l��/5�z�V� bȸ_�3�C�bR�����ӌHv��;'���lڶ�xA�;]��1Dъ��:���Հ�ǛkW`�|_�>��G����5{�T��|A];�[��~[S��Y�B�@��ؖ
�GOҽ���r^�ݪ��+��$�p����05�Guҋoy}S~�#�D�,p�nwo��7(W���[�5Q�.m����J(�p>�B��P���h0���}m�29�OYIF� E;΁Z��{��851Ӛ@(��b��^7�PkJ".Mr�����]t�ڴ9(%���	�B-�ă}�a�VxC�c4�GB��+�R���%"�T��i]���:��4�d����)�mw�QB������{�O�iX��ջ�I7���FV$IJ�Y�t2H,����H]��������st��d��g��=H�_��J��u�~�a�C;�l�%�j���3	�Z�yN	ۀ��a�֑��5P��q��{��"<�T�����O}�m-ш��R���ڱHyb�k3i�fƨ����N��}�²D7�o��Xc>7� ���츘J35ìB���� ��0�?Ě�)=�f����4���}��Z�BL��j�{��6mّK��O����9��&�.�^#p0�)�-�l���=t��Oѥ6���8H~b�,�a��O���
EO��L�SeT$_Ӽ�q8E�Z@(�^���Ϻ����\���B9a���!ȿݡw�?���������*�L�d�t17�gD>�C˪�[^yw�aa��B�m�o�,�'縭P֖	���b+���ir�9pqh�/�2���^�?�[������6yg��a��	nߣ
���XV.�'ZR���:�/*��x��,:�(g#_'��2"J����c�8ֹ{S���|��'o�_�7��|�#�ԗ�uef��e�@`q�o�����1�9Oz��-u�6�K�r�ѷ��z��V�-}��1��z,"�~ll�QF���k�MB�z���Y?�̖Y)��Zn��4����l!姡9��P2^�1X[�&���
-����B\�� g�̊�}v��ߤܪ�9V�].�U�3����Zխ�8����&e{����E/Se�?��f��ӹ�I�Cؚ��j�Z(]���7;s2	s�5�u�V2U8���iM�\�K��Y�o����ͨ�蓪��Vu��ݓ�S�Vj��+1�nV�G�1�&��b/�2���+�:�d�U^�/��/��"l���K��B7����M��j�FCfʱ���i9�T��ˈW�I}2������I� ���/.T��iq��\�Ez���j<�F�>��C	����2��/My���bW�nK;�W�t$H���(���=q�]>\�u��5ͧ]�Nw?���Rֹ��&�ta1���'���}���;�M��i.��YX*k���M�����Uc�ʁ�osw$�)��}�Ũ�r.F��G�Ջf#O��a���&7B,[ڜ�s�]�9J��xךExY���Iֿ�Vg7u�|�3h؞�}�U27$p�9XYH˴�LDv�#�\�eH�OZ��$.%�6���|���}�cF�Q���X��36�a�<��Q@�l�B-��. ΪQTM��$MW,�-����h	(��L�%�>�Q�x�y�7H럏I�vT������ܮ�u�62�@����*v,,�^��Z�r�laPO�(��l��z����n�_��l�b�����������?�)"���z4�D�|3�M�������ĸ��=�v�������F�^�ƫ��D���M�K�`\�� �'�?f۟O���� ʁJx�_v�y��eՓ�w�����d1���*}ې\U�y����T����7�p�;��*=4������e�e��޻7��-ܨ,�P�5���e �#,�s���������kUIb���Z���%�r{*h���^�2N����>L�E��Uj�x:o�8�k���Ǽ=�0#��i��%%���3�a4��B��}�e�G��tX]�os	-M�7��� "�G^Xñ���a[��Q��<����J�&z���?8��e�tlZ�E��P%%ch��yH�a܄��v(��
����������iǷ�6;��~*�(tO�.n���X]4���S
<爸C�(�oS��6�J�?���\�b��%�}����Vb�'���ɲ��5�]�8����5��֓�����pr��8V�_�B����7�U�uW98(�S:̣��"p��,��|)D���������+˘���Sc78���Q�lh�^D�DJ"���ן�lDr����ur���5w�Բ͜Y�n<���E5��]ȝ/=��ό���F�����Ib'��ѽx��g�]�F_$�}]\������:=#a[	�(��Pl%[��	����ew=�f^�ub���Nl�P���D���q�+�L�QD�d23��a�y�D�T|�D��(��r��Jz>�d��(�!
�MR[�z�2��P�b�[iy�#!�ȍ?I�[�&��&�C�?��j�>���P� ����z�#��;��A�b�J�s�^{v�.�͋h�+k�Q3ț��6,؈ݝ�H����ա
Dwp�CE������L��$hs��u�����@HژY�̘?��k��>M��~����bpp�3�:u�%�}V��Gֈ����UX~nW4�X�DI�<��t8b�e&��,~@����gV	>���Ң1�S��S��];|���Ot�-�f0׹��
�m�C�%�i��b�i&����IPCܵ�:}�s�ǂ��>>��pn�l�7t�P뗝D,���
�7�t�ki��4�ǝ��s���{"d�L��g3���{�V%B6Ğ0�q�%.�U���+����cEʦ$��(��@VߚLNl�ۏ2茟Əa��zJ�r0.��2ϒXL�=��`�yqꂜ�`o:�,C����kz�8`]�M������e���5n�u�1z�23)�^�k�Vz�D�0R�5����.ȃFqlN@T�ޥGf�+�K���Ɠ��t�c<C\1w�d��Z� \9�6<��V�����F�ky㽯'��M�%*SS% ȓ@�S��9�^6Id㏓�}"ξ��w�l����������&·G 0J�K)B��k�<�Þv�JNc���������C��#�B3P���N3��yu?����$8��jv&��taT0�&���^�"|�2g��=j�ֿ��vEZ6~:�vS��ϧ���7礴�S1%R�A1SB���8������U���.n�|�i��O�'��;f*/�2E�%ii3�n��V0�&�i�?Ћ�J�QT6#��bF!�k��)�L�����w�]�h�ϥ�Աy�uaQ��%(zagьWu����R�����!^t��]���;L�۴ӰR��w"��8AВ���b�%(��Ij�R�"(�`�I:��,K5�=���+�(�k�(Z�}g��	����X�S�:R4E,D4�dͪ(�%��sl��D*����DQ�]5�E��,w������u�	��ݮ%��h���U[g7�q	&�`�ܡ_�%R*��o���'��k	#QC}�n�!G�
2�3� �~D6pt}<K0�P��8L[i��/�>[�6�.�{�˔��H��e��Z�j<�Z,������J�ύ�)�mVf���>H���v��`��T&=���yE���&<HV��e�?�Q�����:���M��J��A�( ,ّ��舖����lC^l�S�H��a{�{�|�#ߔ��.j���{uX�+%���w_+��Ǖ#���? ���� -�0�1����~|�3$ey����b����Lsҕ�yc2���E	��8���,a�LܯFJ$��b|�۱�5*�����������=�r�M;韀��C��q�����.{�2N0��y*4烗g-�KSc6\�'b��U?�% 4��8ur�|GL�:�;�Lu^˰f��_ώ��$J{���?K�5�b�W�����p�D/̤�]$n{�I�fz��Cf���.���W��ƛoZ��|�`�7[�rr*�v� ��a�ʫ^%�=��o^���dw�RnTJ��G�8�x����ق%��s����r�f=i�ԙLHl��A�6�� ~�<f4e��x����b��)D���n��P�/M�hm�hr%)E�8S���E<:ᵃ��Q���!׹~q������4p	Z�+��m"��Q��|���i��JEOZ�*�~�Q�RABu��������3}G�Ȥ�5B�
��	���9b���ȴf���,ĴK�S�M���˗��|;=+��ĪϢ�b�_��_�q�e]$�-���lÙ�G�d~�B��ou�����yj�K����:�vzˍ�qP��m�;��\z%+B�d�̓��lb������{U�pQ"��;��n-����[��'AϽ�يCie��*i5�xz?�5z�LJV�f6ɘ��o�r��퍧]3���3�n�q�Z��vx��S���}�B�6�
e�����Sd��Z��m-��f�����[�䩝Oyz���#�^� ��z�x�&�i�빉0�ǯ`�#� 焐�͍i�'>�[x�b��L����I�>SBᕐ�3�����5^�VW]ϊC~�,\����I[$��ը=0i �h�ﾏ[���ۅ�+6$:z:O�έy����4uh����oD�~��������Zp��X�7��^�gY��Y��4;���4�~��֥lY:-	5S|�0J����� 1@�b�4;�V�O�+��<�51���e>��wΓ����ɸ��೥�+�� -f�dO��l���*QH�`�`d����0T$���r�
}���)�!t�!�?�ΛP�؅a���t���|��=I����{<:��=�n�٢�s*,]J7!s`��0�7�~O]4��}ob���9eR{�B�G���\�~bt30����aeQ��[�f �wJ�UF��f�u����j�EIW��-}��Iͅ��a"R��$�P���<4�3A@��r{hdNI�k7qV����C�s�^ޅ3��b��M��*3����$i��:�Z��(�R�	����	��5K�`�5O�(���;U�3�%Y��'�6ã�M��l��;ᕜ