��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���jl�7�x�֫����_��aoY��?#��#�r�m�"R^F�(hb=��pt$��e[5�v� ��n{L�x����o�x�+@wM�ca冐堏����D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[��Z�2���Q'
o'+��
	�����wsN(�z��ݶ"��b:�ގH���܎�&��l
�3�O��kw�*���yKK?Z}�K�L尐f�l�G�0F����Of>��8�-�@?����Z&�������3]�C%M�F�������L��'�&��SxUޫ���
�s��E��ȷ�o�{������e��݌[�s0���ض����..prsð,d殚l�I(���"WGIR��]�6�2Y����)���eaW�o����*+���4�?^. Z�sM��_�%�|xJ8b�
��ӝl�b�����s�m���U6�[���'q-z���Q,F;�88�s�V�Ҋ�R�l󝚇�i�B���E�G�䋚�@� �b��O`<ѽYdC�׼����[��\���d(��'�:��h49�i��%�eԴ�>��^1U��=[�xkA� ��u��/�i�!$�g�F��O!|�Ff1�gƸ���!��?�v	�!x*�g��*@6C��U=�σ4���%D��R��s�x����";���*�#f_i�M^v.�d�`*h�T��4ٜ+�߭��ܻ2G�Ðڊ��n�����y��\v���ת������}���͒�o�V:�5�J&Q,�R�5b�y�/A��ҥ�Kݟu� �a���k�{�H��������!n-�NA�8$OI�����5|�J�#0��������ճ��'� ��>������F���9�������d��h�%����Y�QO9RG��V���=M�����	���Q��b��8�;�]��95T���h�ӭ!�#~�}�h�-�� u�O�#Ms&bD�a��d��B|��P����U44E�;�!|���+�7��֯=���/c��Y�����695�Pe�	H�pq�]o��<�&��K�9�} A�kL¾�_@��]����p��c6��`:$�b�ٽ��d��ɟk��m.�w��Y>�BD$	G��ih�V�t�F��s�m'��(�ӳ�,��w���_�0-E�*�kAQ
����o�#Y�,��N�v�}���y��1�q-U:�`��{�'����hGQ�*3�{����hpy�S�/Y�=^g�����D� V|"=��u������&[L�*.���j;R_����)
�Ϟm�6B���x��!����{qFK�׎���}�J��x�P��يĎM���J���T�z� �W���E]����?���z�# ��Ie��%-��]� �ah2z>�(�z�@�E�i�f>/jk��6(�9gH�3�ϴ͒r�Q�����D@�(Ij'L��WQ����zc�k�����jp��G>�̓��.A�vN�7�Q�F�r������d�!Y��~��5��,t�o�gB�O:���˾���(���>I<�q,��_B�Ѳ�Z��Z���Ҕ{�{h�f��Y7�B� q��WTp䥭���y��_#�nK#`�+��ws�	gz�!9�����x���#����%��F����%R�:<��4*�ˆ$Л��
H7�=���@H\�����7����u�Ǧ�G�:ݛ_���k�x������A��'|�{?z�z.�5�<�R�>�9QP/сa��Yru(�㯥�l��A��s�m�Hu5G�?�o���F�n�M��g�X����M��}������gq~�+�L���&P�4���b��_I)�M�LJ�����*�{^��w�U#V!<*�78�++��y�);B����gC�?��9=E{�}�$�Byݏ�'��>fC���Yh�7���<.�x�=�5,M��~�ހ���o�=|k�
��,��F�Ĩ�DB��.1���Ҫ�M�L��'�������ꯙ`�\{y!�ډ��g}�N���>A��oзhlF5��}��G|Y�1�G%E�g�{�e7�V��#0�]H�_�k�"�̽:��8�$�a6c*aq%3��Y�r���qӀO�(��V�����kKXg�b9���p���g��|�g�:�(�m��Q�{�~�N��� ����UU|�1b�Ha�EHd����}�|�	kPt� Sf ���)9�!�B�v~'jX ��`���6	��8���gB��&�i�՞w��K���T.W:�J�,�6�2U�x��H��˺��7�DS'��\�!�Ag����[O�gތv4k�P��*�����@�|{0^.Eo�3׈�&�k��n��h�=�ǉ��S3!C�^�'a�K3�?71�p�U���}L�7k��ټB�6ô�~�V�奷r�����ԯ���؜Ғ�׊��u�#IO�gd(M�1���� *���=����y�ci`�u�L.��!w�HuC����q�c�t/P�_�1Xr���=��ݙb-�����|m�H��@�3��5TN��gH�Ox�3�s��L#���ٝ�+��B��+yҎ�0'�G�"�$���T))Q��D�����r�V)d�:��quBi��1�o���>��^�aTzug�g��-���}*�h&n>���l��l��A\��_vjUS�̪��D�9�+ծ�>���-2Cn2Ĺ�hϠ��u��ɻ���3�r&p��N�r$�I��{o ��,tOm�;��ANV���.��:�x��l���_ ��)��y�}0��RV�js�	�MY�׋�jU�'�n��T%��
�mR΃�D�̏VD*�f=�L�w���d�,�����L+�D[�/>ϟX��"{�v��%�2���A����Ġ�-"T��|��-+vd�A.Ǽ"K����fh7�6x9�eH�l�gh�!3��x�8."��������*��U�=�am�2($���s�
�����:�͘�����L�-��|�~�Rbm�(�fԅ\-=�H}/�ujy�o��'V��B3�G:��Q����G��Jҧ�;�4#�s�l���<�xN��]�+_�w����l*�Z�m4zm��7�_I=.�0f.u�d%\�[Wki�ϗX�>����d�ʒt�M�6�����p玊�_?>\W@���C�8p����4��'=)η�4�pte�5��x$1nk�64,��'<�D��sn�Q�v(�u��}���T�y.{��S�~_�̨��wv�f/���*��ǰ�04#wt{l��7G,~0������~�����E8Y)�5ɸ�OCu���R�)�h�譌u�r�J	��\�_�6�^�e���m	�|�`<�颍���-LXحY�F!Y�����ϱP�C���~pCF��4���ܛ��6C�)���b�]��ɛ�QP�P�xЂ�`Bɘ��Nګ�,gS2r�';��N/�����7g|��,j�S������.�v4
"���tؖ�Cr��P�tP�Q�w�&��|]�����Le���I��.�X�>Fja�6��K �5`�O�>�dQ�	)}��SzT��.�#i����r��LW���e-YL�-c1c���(�0�W�Ǔ��K�O|A�П�k��P��(5�>�KE�j������w �	�&�`>�	 ��9�>��ۂT��~%'��Z�Jؕ�:��r�u87G3��� �g"��]�����Y��� ��8���癋��ܕ��a#u�R�Ǹ-`f���l�����$@�>���cU;�[�;�-bD���TL-($��?ϧ�?�>&~�q2�f�y=�R��,�=���Z4d���K���!Cq�Rsf:�bpJ��8m����>akB)�0E�;L�MP ��t!�4P{��~f�8B��_�M�W��?�PB���샔�0a�ԓ��*��CU��	yڏ!u�G�d��l���Gi`�	]��I���B���N��;xm-Y�'=ۜ;��x�u	�yt*C#X]�H�����r9�4ߒ ��N7��,�rs�O�I�Bm�z@O<�[<u��§~�4�`Q�*c����[ $��!���+��g�o&���류J����.��Ը���0�}�x�Yd��٦�![�s�V�nz�z�n�� ks�,�w4�IЅ�S���Kn�=���#F---�|f�X�3�t��Yyٲ�']�e`��U����iǡ��:}0}�3:

O����m��Ey�����U�H��@F�s�����<��s(��l+v�?v���� ��/b̬���ǝH�L�r���]}���i�Q��!T��	�����T'7՞E꒶��,��4q�*�Xk�PD2���w�t���- a.��"�!w�Ԃz�A J�<}�Ag���!���s�Ʈ�Ӏ���o9�г�έ��1
�{lSA�M����������/�U5�Oڙ5QE �19B�&"-<�)˄���
���*�oM��ʂ����~x2痚�!^c��(Ņ�܏� ��q�� �n�7�;�0�D]-d9�6�.s�o�����2�����������u�kA*��2�oh�_�l*�4+�ZG�$-ey�e[��ˮ��5W���wQǅ�#"�4a�+UHa���1z�����F��./���j��]�S� �:;�]Ŏ�3h�\D�n�X1 ߁�3��b���u:^�5|���2mP�r_upt�.����RZP��T��z�P���P��.(�~Bkێ��.�}���Ek,��4-�����p%���"�H��[$�W��հn3���·���/��S�F\�ȘN&��F�T�x6��NH{#m>���]S��+ An�������zp�P�yD3)��"�K��a�/�K.%�T���1�;�e��%�4�ʉ79��-1��?a]�q ���ݖ�^}�_4>�i����� PO�����R���V�Nu�8%�{#�栭���d��[�ʲV<St�	�rMh�U���}�z��\�PUR�C_��t��t�_�^Z���� ��)6W��P��DPe�K�I&�Q ��}I9�,�v�U+�mG���D[a�ÿh�/|�ӴN�ru�ۃc�	g@la	n`A~r w��`*$���[x��}GN=F�	$�-�-�_F��_?,Q�͠Oɚ1�Yn�iFL�����������0ڇ���_V�,@�s�)
�\c�Ą�V���]7�����.��g�j+��xw�v4���Ƌh�*>`ώ�q�;ê��|�7M�`�y�cN��A���k����~N@�"ˊi����-ĩ_7P��lG�˻dn4,�z��E�J�x� ��0��g�%����%�W�n��%�쬀��PnNY��א��R@��(�4xN��gX�\l���,v� �x�7_�>A�����X.7/�Z6������k��gie�-�A��S]�����<�K�d�]�ShA��|h��8����|����X؎'HN���s���-+M9�Iz��d(��Q<]�ᛊ���?S�l'j^#pȘ�5$��Lr�Sp��KE��l�,k{N}�����%�[�@�T�g�[�)���uvS�����:R�<�����ta*� ��m�m�0@neT�q��̔JS��'S��ۃ�iW���q`�mT�Ga����s	�e��<�����Eh�!�ܰ�k̲>8��2m0la�^2p�%���f�C�{κ�A���O�
:�+{n~�HG����r�a� �vB�6w+�k�1�"��>���;�	\����wP>g�{Xr�0�*���"-��l�5dL��PpW[f�:J[��EKI���E��&�t�:�G���>�8J�y\�c�~ۓ��O�W�SlUj�X��G4u���*����l'�4�Q��PA=�B����%[���i`>���yϘ���h�u��l�>0x5!�������J�NO�u/��5r�e����kD�B�n@N	�U9��0�Y�'�=3���|�k��W����&� s#� �.$�Lk���3�@���6fvZ�3T�3��L����(�ؿ�m��{k��G��ϑ}���+����[]u�ՈȊ�e/�	D�D�똼e��~nQ*SC�O��0 �)�m[U�Z��(��f6�c�>�@`o1;lr���+Ȭ5���\�F?>�UP�fY��W�%�L�^�}��ߨ`�f�\"��5$̷t�+�	[����O!��k^�?�[z�K�ï'�[�����W�F�K���)��:�@Q����h��Fgg� '�9X�A	CӴ�����#���$�k�� �v�� 5aI��U�*�(�hϬ�	�N�0�wxѥ���E�&��(O|�o@C>x����jT��0���=(!�|h�|�rY��< ����O:{���q����CK�$M��j����@�V0��MP��4\����t��е6k\��R�_F'f��]/_:��w���/�j�$v}��[);Z	�����q֫3^�3u�?����܌�_�w����]��+���,?���O�tc8$� g�h]S��K5Vz��H�c�.���'"�v�waR~,�!W�ڄ�0��¶���Gu���Ip�jQ��#ўq+Ԛ/�<%7ߡ�>��>������2���;���M-1TS��'����*����]AY�a���[c�G�D���yJ�.U�)4Ͻ5G�A�d�6	ܮQ����j�M�we1A8�򛽰P� ;:�ޞ�$�R1S�C>����6����a�Eew���C���ޕ�q^,͛s%�Vm��6R�D�,������:�sB_w�z���1��ED�Rm[��.���^�.�at��d��ڦ��/d�	�h�ėj���Ōl�ը����#hu�( n�Q���� �y�G�%�t�M���b���Y�QѨ%r�cX�Z���c��D��L*"�����|��������4NZe�/p��t8�olT/.w��sO���Ƥ�q�p�#֯jͼ�Ht�3��6��8�y�����s�Y����5Y���R4�+_g���'4�����b����+b�;�S���B��l���5�:�`֍\����@�@��(��,%��W�2]�W��0�n�pX����t�c���uT�a�]F�l�"-/3"2�t,z���Sv��|�>	}+�	V�Ū`)�T�mJ|�S�u�+��{8��2:��L�����]�"�	�2zh�E��#\��������k5�:i�Hl���I�{�i�2�O�㡜az�8:_��%.>�v"����񄦸�N��m�n6�t&ORn�|c�}H��p���o�uPV��,����ބ���f�4a_��r�}��в�)�Q���!���OOJ��*�V��$����B�2p�(!k:.y��#V)\/��l*��э�H���8�C(qg����v��Fe_I0[�Xf�r����BLCh�+��kI�{.$w^}�=�ڎNy����`�!>7V��?`������k3#GL��v��)=#�ҸY��݈&
��Nx��<ȵ\8cjloi������x۹��y+��Ue�\�Tch��ܘ+?,%�I�8���jP}�$:��R���1��a�f}-I�F�u<��I���sw�| �-��^��b"a����c �U"�kq�)�I����}�z�l�ja�*�_���g�mE�U� �Tw��|А>4�v��*�;����y(���_�ܾ��,���������5\�ڪ�9�C��o�*�f��%�ީ����<��Cg��ǝ��y����s�C�鯓�����3"����X��}}�z������ ^�uj�C��AT/vށ%}���W]L�q���A; '"�;c����d؝��IW�g�Da�m��a�����w�i4�7�R��&Vs��3W�PF4�UzW��ed@�2���IĎ�n:�n�=�L�J�u�~��}�H@���|����vU��F�^�'�qs:�W�L��y�t�!�1I����[��,�P�o-�q�5=�;p�5=�>8��l�$���sɄ��떽,��㙣�(X��D�'8�߰S���L[�=Բ6�@\�S��D{=j�t%s�g���f�׎n���ݴ�����H�1����j�븷c��o,�.9Eõ��e����vxg�:�-d������.��QE��xk��t��^�sD4�ҡ����#^H�����f�BH�RD
��:�X6����yw�m�ꄷ�f�웟
vb����`�OG�
n�����k��k�n42��"��P�����ÎH�^r;�/N$)��$-Q���,�O՜�\�7 �(�3�`��O���0#��;��9�w�z�b�U�R�G-���xnɪ7��{���E@`-�ܖ��o�}�v����6���j�z�W���>����LA��r����L������Ԕ���Kvȋ��b/��4���4x��_v d�Ed��wo�T����pb�2j0'=V�I�-���?{w�}5y��x��~���dq�!�W`aG;iG���)PL¶��\�'�7�i�ހ��h����Dɑ�ez*+m+��X'l��\��
�?s���-�:����^�K�u��U����m���� �
���k��?s"�v��~�,u��w����4StG4�P@���CEfm{K\�_�5��TY�V�p�����o7_#I�~��^�����.�LDןk���L=9����0��3�=8��=��i%R�k�� �J�կs� �U�!DZ!�æU��YG�`��6�u��C��*ihU7�k7�Jn&0�� �(��P~
�9���W`x�/�0��6b��a]�x�>?��)�X���0S��`S/�6�ϼF���1.�SJD�ʾ�	]Uϲ��6���R�����ƣ~�/����S����X���k�r��)-D�D�y���^]�%L�F�J���J����>��9���Ϳ>)C�����z�t�,����M��� 0�cq������@��(�yaQؔ�`��:[��x��*b�4�l� ��K7�K�No<�������妺/N����tJ�4�/��RL���&�:�|�4M����e_);�)����Zд BK���H��id]�G��ʑSM��5�?��Gk��:�$�u�e�)�Ƭ�Z_�bh���^_��s$i�7ѡi�i����}��# .��p�e����'��#����y�5��C����p����$�*�o��ҭ�AN��u+�ȶ`����:�pu~{p^on���f����ǢΏ�=υGZ?gV�*���f��!�,���pוmo�����h�ޅ��KN�g!��c�x�n0$R ���{���2?ݫ�/��,���Kb{�Z^����Jv��0 �y#�R�s�oRk��f	��k��ͳ����I���LK^��G�.�WϬ*����O��A@:1�M[���@DԌ ��@���5!Y��
�����d��>���6[�<X�����8�lJ����$��SN�Ŋo6���{��춹�&��Х��!�"#��[l��_`�aF��=�w6#Q�1��;����N��߳"�cp��z��'_��|Am��A^l�wy2.��+nfF�M���BM��}C"�R�+T�mbt>w�8[���/�"h���T~s���dh/DttO�I��>vgKG�Zo��%B���R���⏥�R��Z#�,L:��};~��!�������;ʰ�n%k�OY#ù�@1͢�G��҃S@'��v3��ޘD�|'dgg����雠܊����(h��Q���]����1��v�X���];���ؘ<=�i�����p"R�5�Jѕ��C���ǌ#��tГ�7ٴ��B����D��ҰZLb�9�w�=��V�$/��8�*L~���ڢ��n�S��=�	h�Ԡ���+y�᪦'��e�,�W6�.�E���sdu�8O^���y۴\��O���>�!��t�2��&��Ym��Y����T�Vk��Q c4a��@ˑ�)
MN��P��4�����xa�'^�ӻ��te{p=��
W)�)�`Yn4���G���ĚL�$��Qݳh���cCf ��6ą��)L�l�e�/�&sEl�dtIF����O|W�Ҥb�T�Ğ��j&E���aؗ���դ��H��h#An����@�ā�cn�ג��0\.D	���	���$��dk�QpO�v}�w��i����-w)['�z`��j�P0�8����
i�F/�������nAgo�L"g�r:��<�c��I۹�Ơ�Rv�0=&l~���w~���t<x~�G�����{M#�S�>]�}q��� P/�]�ݶ�w�?�?���TH���_r�{B�c��	d�����X�#� ot,�[�ZX�;�Y��D���rV�JC�6�A�7cX���~e#�倝]��78u�J�gD�C��[G�����җ�҇d	Ĕ�_�_K���A�^\+�)�A/E+�$�$VX/b>���pY,�ط�2 ��&�:��䕷T���@'*�pa��t�h� �Ԑ�����b@��P�JY�q����j�
[�d����waR�3���&ߐ��!���R�@'L�^� ��.���������t�|V���ƍ.��d�Kp�wM�6�<;��38Qk^N����Hh����ٰ���Pc��6
]=�EE�I�wX���{|7��i�5�m���Չ�%��,�_�d�ZG��ٜ6�(b�e�Z���>�D�DE�S��I�Z�;��6�Q�Kx7]![�3��4���i��r d������%7ެ9��ะ��T���Sc �s�0��l4cB�Hɗ��U��B׫9�{� �����YF�Λ��K6�F$?��_Fp��������r{Hl��Jo���2�!kȵk�h�w�c�6��;=x`�Rd���q[��d\i�Zm��kFb�+�'tQ��ز�t��v�
�!!:!A�}8G75⤩��<heq��^�%0��Xf�-�GM�r�N�n�WO�v��kŜ����(�[
mRO��QW�EC�Mi����"�<X(�6�;w_�d�[TL�*C~FDi�䐨���8{���(V^"�9�}0��$v/z��c��L5���ʢ��l9��x<G}.t����i5���^my׮W@U1���� �L�`dP=�\+�� :��z����K)�GL�8{�k�%�2�qa#=F� �q�,��� r4��|�f\1ǲ��'YS�)�v��j	.le��k�o �޺H��U�8����(o�5aD��*��ܢ�Ʊ�O1zw�S�Сx���a�)�:N����i�!#َ�T���n-���8ד�	JL��wLD�����˦�G���UV�/������X����(�Q��v���	F�'b>�-銴�{fu��V�3�I#2�5Qί(�Ȍ����y0�b8��x�_�o��gw�
�V<4�K����eD6�+��K[k�-p#<>,�z��S�踽�6K��ѽ��pq��Y��S�F.p~�ֿ���رpLQ	OZ�u�/(�N7یC>���L<ŗmcg�V���>�_���l������,���H�[r��~'�6�9`�f�s�~ר�+sIJ��u--��E��4��lH&T��w�B��D���԰�+:c�l��e,$U��3x�����'��Uz�CS�n�w��K��.���F��1Bpɼ��";�Ft�@+ҧΊطmL�@�ZD̾&Pޑ	x���6�`؂w�m���:xW��q��U3?�9�=ZI�o}Ī9#��T�!d��?����eP#�%����yk<�!�Qf�[�w%_�D1�E������u�(;ঈ��r}#d����E�5�
��<G;��	���K��{N_v�Yf樲�a��㖰fҵ���{~��U��
��G
j��u�T�<C�Ź|�(@1v!�c�A,T_M�VN��z���s��d�� R�d~eX$G�P����z�#!�G�o780A4�1�V��A�v���D}^��zE6nu��n�f��*5�F$NOdds�[b��p�æ��.��N�p�ߚFz�۹
C%�M�8��0�(�D~�s��tM�|d������@����B����h��0�e��=��Rơ�x��E����z�ۡp�+[;@����'i�r�����܉��;�!�D�?���Z����p�fЀ	z��w�:��(����C��-h��r����ln���,��>e�N��C��m��f�+ �����E�_��h�Z�PQ����8�A =�?���p�-x�0���(�|�ھ�i��X�D�����J�zJ�s��a�B Ȟ�痢Eh�c�7�r�aSa�.{���d���;�Xr6B��Fw�<b2A,fQm4��Nơ�Hl�4��+�6�����<4��o��Fw�����/Oξm^7�l%2SC&��w��s}\�Ϲ6�w��!�ɴn��z��-R�9�_Bk_?o?�iQc�4�7�#N��N��Y��H�A͓���ސ�!	fL���|����� �$CJσ�c�+�qS�%�|`>c� ��]])����v� "&�Xf����bb�@+�W��A �y�^Y���#��xc$�>����"*�X�ug,@����/5�Dz������(�r�h!��m��\��:��V�x!�p���zI�5�o҈e]ĤZ�reXwיa�~���mV�"��D��[���H������ڛK��va<�~(ء?�w|�#tڅ�|8�lA9�T�����z�/��+lU�nb⍅�e���d䭯nF];џ�"H�%��<�榆��I���"�0���7~8T+�(���ӢsO�q��S 0�������~���]��6MHɡ}jp�T9Ͻ��K�\a������8BK��`���k��0sH���R���,�8�NB���Q$Ve�N�Y��<��C���+��� =���wa� -��^Wb����
�v����U��#�Zk�����)׳Ud���#�ObQ5.�2���#��Ƨǩ�#j6�.w����/F�lPx��Q�}�J�;+3��� ML�و�$��/�p&E��M�8[G�/^R%�Y�8�#�9C�jb��V+F��+�T(t"0����
�v�x*���2����[Aep+���'2�o#6����d��a6�m�X����Qؑ�+=�X�.?�B�C�N<5��?�ַ/�i�=�4��[��~�Y�L$ЗX��ߎ�_���8��s��gY5)��3	���At(֟Z���]'���)�uN�)~d�wL�O��Z{(��C��I�Pc�#��i��,���uKb8b��Y��꽥ݧ�ms|����׎-��7�$��2��	C�
wpaK��B�Ġ���r�e���-	(�����ɩt>!���'"�ޚu8n� �R�}���?�!��t�pW :�+R�d����ӹ�Yg{����ܥo/��R��#n:~�F���dsUW��ӄ����|$x2���1m]��ڇ�����	���=3�7�[a_x��Fj4��D42 Vw?y/p�݊��I-�hk��{dh�]D���x�����"d�f'Gu*�g�N� =0�c��G*zG���N������a�C�f7ۣ����0���Ch�}bSnв��s�ɔ �t��~��lV��=��-q��y�3���ft�,���6ւ��w+�E3�e��7���k.{:0Z73��FL����@�>Z-px�=��n��H<H�ߡ�t=m��(�^�WxX�o:�6��/�3�15���U�!
�؈\x���'.x��A�g����Ptȴ\q�|�v��eì�`��d��t�����&R�uc,�.m����	Gv8fH��5Q�$V �N@s���K����B�,�x�C����Τ��d𙒣|���	��ފ����|M�m*���cm��E���L��j��x9,�Z,�	>���
�V�)�J/y���a��Y�M��]��/���2N�o<G7ϧF���l�jvU��r��
�ML��k�JQ�)K
+1;�O��'��t_�=�ɏ*�/���Tǆ����o�#b�@O���)���։G#i 7.d��R]q���#!np���V�7Z�m0I����������T.3f��>�Ґ���ޞ�V�׳`���9���(`.|eW�F��urԝ/cz��4OY���n��hO�v�Amٌͼ�u5�8�rG!�/W$����!Q���2\h�3���t�������.������7�S���nr���^6���@Wܾ��%H[����f"����кv(�To�]��wz�'b��Aلm��"@�:
h�6��R��rx���(���:��R���'?\����K�Gݴ�ux��ג12���p3}�r�����4Ak�[-~�OX����V��טI�3���J]�`��/4��������qGx{a.�e�Bf%ZT?��� ����O	(c�w��K�<�'�z���E}��V�� �d�%'nON�r�ם��5?��[��lv�m�9�4'��Id��+�p�m���� �G�u�"�H4L�,��6Ӻ/���چ�
4tL\�Lxr�(m�h=� ��ɭ�"4��������<�Dz$b�Y>���;%W�s�Nۚ�Ԁ[����^�d�������b'Y���g��}�_�u��z�45-<�0�:����T�y�%���e/O8�Q��Nkv�"����=?�����	xU����8%
��Ԭ0(�;.��K�����8v׾�p�W��7��������8��ǒ�p�L���y�Jc�7��;fH:d����9m��"���%c�uxZ�[��舍�[�yT�R�n.}����*�2��'-�I���-��
:N\����l%,�y��-.tϯWv
�Zѱ��eq#6r��-'7"�D��@i�w�ﶖ��)|���g5�ǵ7�݌ʪ����ߦ�E�Z���ۑ�����Y�:��Q�g�8�f��/LV`�[�L�\oOqQ#���ǥx�@D%eF�a������y0�?�/�%�7'�E��Zk�dG��7�t���k/�Aw���ӥ�K�(8�Ai	ƹћ��ݼt�tԻ��C@��W��實���82.��M����癙����T��%g��P��(���+%�~����7���Q4,N�x�aK`i�Q��;�B�#\j��Ջ�Ft'�rO ���]?�����c}\�7x|5��(�j�9
� �"�Cu��Лq�C&y����A!��S�&��۪/�ŢYA����Cˆ������n��E�L���z�`��"�>��Q6IH:��c��E�a&���g���D�؝W�W��:K���	��sa���`��=��WP3��M ��s���_�o�F�� E�O�>]������"�s��6��e4�QU̐5I���&���I�!*CE!/�2XG!��]0E���%njY'���"�ƒ+S�vf�=* ���kBWL�0YZ��q�����b������0<i+=�х�x�?��]�	�Ǫ"$�v,q��?����mV���Q�R,���L�K�W�B=N�i��II��\��N&�Y�B���~��Fw ���-�l���VLړB�������	�w�^�0L�
s���������m]�%v۵;]�.0x|@;m)!-��Pڄ�ٵ�,����NR�* ��"��*Dn͟��KG�[�8[��S��ю�!�3H0nbD��N/��']s�:lk��w��#�	�D�Cٗ�1�9���0�M4��~�"���CP�#x`y�(����h�� �n��-�o��Y~`>9e@�k�D�_7�D`��X�ߟՁ�b�v�qgQ�ؚ�z'?K��vE����1+�� ��렄R�!4-��+�����~�
T��q��h�A{.�3Y(�¢v�n � �`󨼻�c���5$�(� 8��z��h�%`Y��Զ>���[�G��i�����M��O�8���ů���\���ey斶��.���Q���n��Н����-֩�3���������'�0���q��z��]!Q���׀gF��u�m�N[��$�Tj��L5T&[a�4�Y��#�wx��9������$ �}�Ĳ��k�©�����¯D8��u��D	��M������1<�=Ȭ>�՘*e���R�B�U�mλ��&PG���5Q����}�%^�n��P�}�7�<įr�KmcͿ���,�K�������,KW���kO���eJLφD��J>���&5d*����(�s��T�����p�vnQ��t�+i
�j��ݹ�Tb�\n�^=eY0�
��ˊ��ye0������2�/,j��h�ٵOo��!eR�2'�%W��]�ўj��g�����x�@ـ��b����K��x+������J���'¦O�U� `~�1C�Ȭ �3*�,$ ;�Y��"Hv����b� �o���}�[ɦ�b�~����#$�]�����*RG�f	H�l���|��������v�������
@�|8��,Ģ&t
�
@�1�;H��V���!�#��g�����-��D���_��7�j�M�_�G��PP3�Ko��!X*���gkx;�n&ԙ�������ޥY�S(�uO�6p,��'��������鹢���k�5'�O���&'s�Zb��\��Q�(��*t�]�v���Fl��Y��lMJ�A�[���Ġw\��tV������uP�~�p��ٜ��áS����n?���G2Š�w�ts�� �=!����V�e't�Z��$���i�����v�b�u�z=���N�6���x%{����`Gѻ�W�S�1_�{�␪b���$M��}�ԯ�V�/��1�d8�+;vL�\����^��ܰ�?
>m؆w��W9���V��P���0Bb|������zs�k"e�W�&H�m9 ��[��n�q�"�������(���9Z�i�bQ=��z�ؒuTx~;(Nُ�K�D�}jw͊R�����!BZЉā���� Y�=[%?̟!A)l�%�> ��B]��>#ww��^�Vx�	y��X�Ѷ3���BP�j�����̫{�4��Vਪl����������_��$����m��/^RH�8ƺ�2LT��|U�a�\�k��C�t8�Ѵڥ1�R��߽5��;�[�5���[�o�9�hː�O3Ej~8���|�BěKjnQ3El7��0��F�F�78\<��b*��PO/D��8�,�(��=7w�;`&��V��*�Wm��� ���3h��o s=ts���:[���~$ ��_��ik��p5��CUܼ)��3�}aq�^��t��?�	��j�?��`�Q@k�!���'�yۘޱ_��h�a_����<G��f/;
���>
�Q�Ym�4����bb�/�R�B��{:�4�%Q�'er�%,�n����U7NF��)�0tkW��%·�#����G����v��۫��=r0����m��ã�����Ln�a�`����N�jV��܄Lf�2)ì��k4~ �`f��S�ƨ�`'�I��PK��.q�r�Y�DB�T��@l���p�K]8풢	��5ފ$L���E ���H������ey�QJ#|.x�3�8>3[
�`��ۙǈ��d��}l=tn
w���t�x�6Z�s2�Hq�� �C)�	� �KB'O�3tr\A:7�m����K�z��O�����׆�5� Y���^��O��3����	���/�����	��kj&�'y��,ѠPim�>����247e� ೢnC*3�5�q"6�(a�ig��P�L�у�K_W�s���;�mʘ��5_�0<�ka��痞j��X	MB�w3m���o�h���Q�gUЯu��1so!w�� }FY�s �b@�*��#Dj�$ Ӗ�����{�.����&"m����)YҰ��&�}�c�=%��ֺ�9򿜸!g"U��%�^j�o�|��E��Ti;��s{�ġ��j}��Ѽb���p.D妩��g9��39#k��I��±�<ݭ�+���؃�2jDn�;��${���k�k?���3�6p�ς�=zy0���y���1��h2?���)���J	?%Z�����!<�A2 ?���p|u;��T�L�:�"9O���pm �U��iK06��&%���HV0JS~@��Nr��]�)�,�Uz������xe��Zo��.5�������Di��m�k�]�'�Nx~�9U�ߞ0����K=�l�_H���������A�+�~+�*I�c���d�eO7b�wr���{8�dmp���,�6�P�������t�O���Vhͩ����!lق3���J��F�ߟ.�b�(��cBڢS�%�5{@T�/��:�Q�,�P�O�:��ԇ��Ca����v��N!e�Mb�}6 /B�%��~��*o奯i�m�h8��;�]�6�l4d�
*��x���6}�r�ｽ�S��;m�k:F�|�aRAs�-�t�~��kKap�H.B��4�ZN��T�!��2�t�P�!�����߽�[4�z=`���M,�?�ՠ�j�m9OUjކ�S�*S�)C���Q���<4�����D\%���F���0��VZF���k�Y�?5�m��� �mby�?�rl_S�ͼy�[m��0�(���c}\w���S����&���"����)�
�Q��!q��ak��BVn 5�U8w@����L�D6Z��s \��KU�m�+t =h_����*0�Vz�x�K�n�����~x"[*�W�m>.�Ω������L��̴�Q�ޔ��nWd��|
2%��*.��"3���d���D�s��Tn!#���^�}�S�u�_�s&c@D���x�_v����%�e��B�𓬱bx=E�ExB�Q��A��˰H+T�\����m�y��)VM��nr��Ъ�))F��b��GVHɗC%LM2P�^�������F����]��8�V�X�=@�3տ�mʡ�G#dbP�~a�i���ϝ���\���]������~�8:�-� 4F��>�����䝕=E+�.�2٧Aպ�%<=�gt�2\���5��X����uy��KJ��OFe��ifG{]JXi*��q��J���F����
�/xz��Ua�O��O��L5����z�x�)�)�!T�7��Z$����Y7�t���s��h�yu��,
�Or1��^��k�X��8�9Ƽ�Sv��'�9�c�������@�N�F��C�._���Q��H�]-��o{�0m���B��K$�ssmh�ƹ�������b+�C����!3�;C�#EY^��]ҳe"�m�k��F�\w&��1��a��:zF^�dm^D�o�]��@�oC�?^:*	��pQ�姗�
�yv�Ikh,��!T���e_���`��`��zfCyXU�����3�X?�%�V� r��f� ��T�3A���,��kTYF��=)�D�7��L/g~�^-�l���M�C�Yr0���IEm����%dL������Q�����z�D�P�fGaw��s��m֦��*"Ѹ��xi
ȫ�N�!��]2 ���Ne�4����Ƙ�Ͷ��>�I��IX���8����ۖ�Nɬ��uҞQj���RwfK�к[m�5���Ŭ#��.�`4 xo�ܣ!�\�F4$�$\F���Xa��>��C(�*�Yݧ~ByZ�&e������}�P�2:-]+�yUq�d����a.O�I��yN�����5)<2��Nd��������k�����$t���C��d��b�@'4��])��	/`2�fۭ�0�E==��`����f~�Ž�B��X�0M�C�v��Bb9,/P�Q��Lrֺ���Y}�+��r�?�o�/�N*�M�m̮vt���M������g-��Ey��7�,h������PZ�fo�՜�O���x�2���f����uN��S�������k����g	�;�mZ�ؗ��x|!Ց�����S1��7Ҝ�N�;�l��"ء���/����ZފW�%�Xf)�ˆ��6I���[,Zl���lL$�W|20��1|��mj� xϷQ��Пg)��X� ��~�'��a�Ma�&����Y�+G��	���{K�W��6��v,�l�
�U�9�3_z��+9�
��5-�:�l�4�Q)PU�i�or��=�){0{�h�7K^0@�m��k�9��6>Y3JK<L�*ʇ���A �@Y%�I��0WQ�q	��Fk*6BԬ�L`;����5���2����G�>ݵ�O���w�����|�L��Za���R�z���yDӵw�|��{����$�֚��Ox��#'�Ib�B��t!��w_9HH��?G�0� ��%x� pq�*�:�5�x��2MB�� �z1��04�ric���	j+L�bHg�����dp���-����t�+HL�x�5p0�[(�c�+Z���`���)�Y�B���̫��ӇN�v,pE��4��}�`�9���ˤ��*�a���CW�{ƴ�"�`$��霴����{��� ŪY��7W��{�1Ax��L���p�z-��Y��،P�h���D���z��$ APe9��\�$2�������65�9�R�K����N����[ȑ����}��B{�(�w�e^<zh�����XA&�F�ۓ�*t��R6M�^�7�5Z����$�}��V֏���]�����Х����]~
�/����OuCı�i�NF+D�QG��oF�&Q�*{��g��3ef���_�E�D��\c2pQ�e�^d��'i(j"œ�v-���En���ny�J�b`	�
:�C��L�x�ڊ�	�͓x�F�{:�wx��Y�RB�v�	��JDxeU��`,cE4��j�CP�ps�F+KR��l�ӽ���D���{��ʆ�1�BQ����1t9���i��$��Ꮐ�^ҍ �xk��2=ÚUHrZ5�r���0�I��� ��_Y�s2_���B��ů�Y�Y��
����~ʝ�,o�ˇ�B�Y�����Zy�U�Fy2 �.(��Fv��cɛ/��Y7}�;����_�8N���g��b���R(D�����ug���w�iP_��ر�w�O/�-Ad�ֻ{��e�'���˥�� �&�":���N4�� ��	����d����}���<o�ng������`���g1�pԚ��c�V�u!B�o�w���0�{ж˯ D�Ŝɬ��dJ��Į�IkTz4�8��G�]aFn��hX���作ޕq+Dr��l��'�>=`�1�:M�?b��Ȋ�W�U�)�"[C��؅hV�A��i��22�q\rm�A`x�Km1���C<��O���I]?R�4"��S���X�ȵ��e�Y7ѹ��Zi<!tྱ��A���4�P'"�n��X�&VH��k��a[�f&��D�n��#>HJ�qK�|B܉�,%�
��K�GBh��b!��h��BY��}\]|`�&@�ǥ�.ô�0%�t�2�+|�@mݮv�pNSP&����p��e1�EW�=8�����/�1��f��b|��FB� �}�T,��ԝHl��×��v�]������Lx� ��'[����ne|m�=�^�C�G�A.#�l6+H�;|-��)c��.@�-���n��!o3Ĕ�$ibj�e����c5�-U�����YL�t�>B���N�7�$̖n?b���U[���0�r4杒Q��������PY��uϖ��`��v�>ގW��Xi_BDPԠ��L�ʧB�8꒲K�=N�h���"�^!4����$���7V��/N�,�L�~�UUq�K	���I�V�������a��Z<�W�:+c2ܠ��k�N<�6��7x���Rh�01Ƀҟu�t%�wNR��n7���B��9��/���ə��lͽ&܊�T1
b=1W���>�<�S�!T h�fZą{��2ݢ++;�m���'X���h��������q�d�y�m�X�����D٬ �<�
��#f)7?#���>�ŕ_�>����&U����tWS�������1�9f2I���:��O��q�,�Z�4m��u ��(����e�� �S�K����!��D���m�%�Ql|L�TA�xCv�	_�ZU�!$�a�(志�9H����PmAk����* �	��bj��`Y�q�������n�w��N��ƒJe�H������_��<��i]����l�{�!�%�t���C �#��h���nRG��g�+�m���D������Z��;8��^�UY&�+��i�PPjbx�:ߐ���9ȼ��<��d��5�S;�X��Z~W�0/�ޣ9廴 ���W��M�3���"�7�`��qP�n�Gې,����ۥ��_� ��|�$|��*�3T��H5����1�\G W�.iv���Z-�hoT(_8^V���LG�v����G��CS��߀�*]IA+����EB�F�p���;�̷���TO�,2�&S	�ғE�Y!N8�������ӭ�w��^*g7#�Ms-c��UO�B빂�&\o%�)�w�}�/1jj%�d��m3�`3Ɇ���'/�s�s��JYN��Rм�U S��Z��;��d)m啟�ҿ� ##�}�|��E�s8�[�A{:+�~���σ��
��$jb�r��ڽ<��K��J�U~���6�IOa�a�hz��8hk���XAel��1�kT~#[�`Qn���Ң�}�S�a<�^$	�!���Ɖj�������w�=&~z�f9��-�T�J(���	\�d�!�Fv�3��A5r���R�Ke�:�.��"�� ��y��8�&��v85�Hqc�;թ`%��X�%�A2�S<�_x��e��)�<�_~1O����	ui��z=���������{
�:�c��&��V��[���zD�)FE����Yw�JAU��o���_�!�����"���[�0|I-�ū��۸�JGٟ��=N}�ơǃ7���/��3���Ӏzj�5�����9h���	~6���V�OQ���-V�3�A�-�j�!.hn�1 9�>�5���������Zk^7�[�m�>��g�x�һ���|ǎOH�wqzPz�MUc(��om�Ӆ�:i:�������خ�"�>$3�(K��goO�e���C=�����!ó:����1
S�zt��2��2��������x`�FXb<L�G~/�����E�|X�l��5f�K�v�[[����O�~�ٙo�E�"�N(��ĵ��d֙�txJۈo����L콳�y�aP�7yS	!0(R�+4`����R��5����2D����'�E��5���S�E�5H���]-����[������$��wAS����-����	FйZ���wĎ̷&�+����$��b�֎���,��3e\�Z=�����79���> �m�h=�ãS� ψ���ф�^��t�[5��{�6=6>-1�#�M5��Ʉ���g���I:�z��"I]m��?SG�w���ʉ^%�� �Z5����霮�oBr�e�����6#�3������x	�� ~+���8��"d{7*�;ˌ��$bZ�K�ۯ`�; �i��u����X�η���|�6�/�D�08�]h�v�XR�S�b&�I����"ut��}����}���1�B�Z=k���j�4����r]���7�zY`��ys �1��Hi�l�AM�q����7݂/���[�=�JR�P�NO�.pS�s�a�����x���9�%��T�%}������S� 7�݇]�ɗ>�����[-�<ɩ] �^���ޮB q�ŷ�q�yf�=H������8�x�';B�A�Y�1�)u�,���I��k�iT��D�)�ƪh�x�׷2�W��-/e���2,�>�uC�5�ߑG�#ЁgҞ�P:�����Gl�����;��E�na���G��/������Hmw]��d)(�b"d.��!0��ʋ���x�
�Z8�Sv���QVmᎬ��'Lo{C3�%r;������ٸ/����&���1x��Ѱ��Tg ��w	1���������PC�,΄8�E0gʒ|B����Q2�$.ǀ~��k�Q�O,t�x۩r���Rd��[�A$�zoE"�K��-�� ��M`1�4$�9H�KY�$4a�0I#�y�T��Ka�4���:�c@�� �����^cO5!��O�"{k.��^��D2X�ʯ�/�"�{e�l&&�t��+�J����|s�H������
�
��zӓJ�(۳���B2_���U�|��u���aBt���b��؟����*,���oP����mhV(遭��G��<J����H���~��������Wзmb���Ed	�:�KD���J��@��&Oo����W��Y������ *�4���{��D���b@:C�߃s����d�aȻ�c�y�e���n�Q"'hj-M�X���q�	��\�����g�O��w���JO;��z
��N�A�1E��e
k��}�de�~��t�B(㍄KA�Vo��cm���
�"O�:�?����z��L_�c
��>i�?w+<���\TH#i.$l�Sjq�>�Y�D�[���p�;��qA�<
M����q!Y�����]5Og��}C�Ş��I��C��V�� #4O��%~N�Q��-9�����P�"ÓS���j�kM���nw[H���R�D��ؠ�,a��0�6tt��A��s ��i�Y�C���a]���󄦠� =D��� eƺ�:"�����2�gI PREFc�N�m�F����/���ǈ4v�t�v@A6i�o��cɒ���[����Vr�nK�U�(s��h��<GU32w8�h�D/�A���0fO�}��i��]�mn}�蒕����� �	��ك����_{&��(&�̫��'$�kxP�;���D�!g�#�F����3>03�&��egi���Ԇ"C R�ۥ����m�2��Ğ4�����xKە���׷��Cip�$]P�� �K�[�b^���<��!�{Cؼ!9vs n7����T�tC�4,9n���u���xz�_6��	��@���h�y�t�LE CBO��}����!�%
�!�bNQL�g&�
�2qo�5��>Q�l'�����L���
Sr�4��爳UI�qׄMǒNqg����v7KW,Cl��_!�>�4��S�����C�/�1l���!��TLvN\3�\�K�
P�U�l��6�|�Z���4���y$t�������uh��%%�Fg�:l�t��DO�@�1�;�Ϧ\�9�)Es���[ŮNd��,1l�fр�����0���t�!<y	�e��S�Ä�@��es�h���?��i�t��9� �YXL��MfB3�K)��U9�����\�'�L��-��#��d�E me̡K�2�Q��C6����x�Hqc+��Ni�Ǟ�*Z#l�{*�.	b>��Z�@f�*Cf�,��Z��U
��I2�G�=�f�ٴn�A$�6�Q�v/�
�lm%/�1G)��tU�y~��|AQ"3�}9l�CD��0�䛴@܆{��z����[�i+3g�a��7��`Z*����+
�}��e<��QF4r@� wr��Ȑ:ho�UM�a�-�`���ɚ�V�Z�I2ֱ�DǑ	
��Ɉ�"�x����S�����+���t�?����K�el�m��"�������-�2~s�>���,E��xܛ���C�\�E�Rw��N��|;%	��cx�Z��0���5� ��Z�"��ޱ�z0�8��Z�	��h�w�80q�'*=�G���u��?;��X��g���R٣��~�N��aq��Ds�D�	G�����~$�X��Y�h`F$}�n���?BFN�!f?0�M@!�\����WS�L(}��B�Ze�eg�����c7�P�1��N��CL����г��g_����b�q{~Ĉ�8���'�}�S������/#mR���Zm8�L�i�aX&�&�Z##=�}&/�]�l.ڝ<�Ub�<G?~7�dd"��\
*qB.��	n҇��;���SǨy��� �rt"�{o̠�i��Z�U�J���B�`����,��-���� }�`�l��D�ߎ`��`LpO�R��N��� +v��U�����g�~�5_�J�����O��������H�����h�N~�U�qG�v2�F�X:uI�9-�a����#����[���j�L�������?L�*?dƝ�?��acgN��)��#e<\��%ȗ'	�pܾ��h�����^낝_<�Va�,��} mt�0���V*L�l��e���}���}`U�霈��8s�F�n��%z��KL�>��k����k�Ӭ�>m�JIڰkaL�? ��q��U=ތ&����S��?��R�� ���R���b���oIC�N��ׂ���댿�'�\HCA*�I��Փ2�-�{-ɣ6�1����F��2e}��� !��T����`�؞몚�]�>һ!�8�]����P��7���1��mlۮ��+J2~[�9�4�9��;�4�R���ƕ #h1�:y#�ŭ �YQ\�3�:֦O��Ja�m�囓 &/�=̌�q����e�T��)U��%{P�@�*�J�䅞�� �9�ƊU�T�����PI�������n3�E�'9ևjk���u�8.�W�l���V�3���{ˆ�-$/�F�W�]��@��8inpU��G�Eb@-���[ C �;R:�u��VB�Qքi�Ê���e6��n�F/񴌐o����s[�{e��9v@��?����T�(���**3W�R8&�h���I?����g�l�+?���mm��,˖��;ߜ:L#�98�w~���9����fgN�a�GԪ �a>��h�G��8��������/�JP��	+x��*�A>n)�
��@]T�v�F��a	6�I2�z�9��5�\��09��-�Oْ
�Nܠ9��g�^�֛���a�^}]�8�,�F)�V��8�	�o��O�^��,K�U�p���#������9T�ϩ��E��.޶$����fE/B��/t��_��J��8��=!A�KީO=�U�ǼRi��h8��~3��6���ŀ��<=���;�����:!�Iٲtdy�f�97�N��v�I�х�4�X�4=Cd���ux�C�8٥�^7�6�z_�{��w����xm|�*��[�C՟ߢ6�1�7Vq�QX���g�HQl�O��c<n����?|��8s�F_G�a�v�>��'6�e�	^8˰�q*�؞	�vv�H�؇�h�J�ٰ/���>���S�]f�XE�]�>�*$G^;�;E����oܬ�,PN�M1��aX��KI��K�?��'B[Zp�:���:>���N�;מ�~(#��v/�*g�,߶8L'/�@���^4A�ׁ��4~2��H,�3ԙt��8��7�����C�j�J3�B����3S��* Ú������0�<0)%��)��Sp4�6��׻
����y~��+�ޓ�oY�����^T�@�E8��mt:2���ʅ�X�8Un*���?9���cT�����w��{���)C���_"f/�ο�,el"ↂ[�Dhge�K/���*Uj ��w��*�n]��R�9���K�IH��.^PȷQ���I��
��}i��n1�?_3`���U��r0��޹:
ŷQ�Y:��S�3�@!�'�ruǙ���wy|���/Յ��ʘ)���eM��T��ˋ�D����G��H�J~sg^� �p�v5����V�~��FEK ��@Id���7"�#�@�i<����L6%�ω*�f�֐�B|7*�}�?�Q�`����ҭ���Ŝ��U���N�@����&�N,l�y����:�`qxT�g�lI�&a� kʩ� S9�XpceCs�{��Z�`ٗ�@'����3=L�J�G�if]�!c�C(nqR%us�ħ���+��e��|�|�៴wǵa�>2��^�M0el?g>ő��,��f�١Գů�'4���z��ȿf�`���{��[|��Pu
.�@0�2�먨�36�Ak���}pDB}�V2�4���'HsuQ�<��$�y>3�n��x���cq�8�J;{9dWI��<��{�B �p>�:�z���`KB�d.�l6�go�Q�A��Czmq���fZv~�{��k�.����:z
��J�\�<���\��kL�=2ZZ���8&"�:��
Oᴲuף�M�+T����:���-�/�r+ݜ6��6�w3h�Y�@��]������)���|�.�!GZontG�`j�M~d�o�sr�j@A�HP<y��-��̣���~#�c.0>���E���m�P'E��×!��&Lx��*� ,Cm�0�8Iֱ<x�	�~��Ag�\�þ�;+�+F�M�_2�*g�?��#��z凸.�G@�e�n�7���^���[���-�!��:��$&�䱫�lu2����(?�w�����wXuatG�Z���>I�y\(|�d�x��m��u�L�XZD�44pׁ)>��s�ņ�`{X��(������c�u,��'�X8�����i������&߯��q�*F+ڲ
Z���;Ț����M��/ƛ�O�����Ҷd�)OL6���"�l�$�@b0�H�8��dH�20��́����̒L볙_I:�- ������'�i�>"m<�K��|ŷ,q]���pp���^ؠ�`�zDWa�\,�QLG�"����re Ѻ���J�<�&�c���iPI�ftE'a?�'[�l�j��	Xz�"�h �������I�BB�p���yD,��mvy&��XQ�X-,x~f��Y��/��<{�3�=�?��(CŃ�9����β�'�)����0n������;+�8������Xl��:�3?vʡUXGp?7�Ϛ���%����C��,1��w|"����f�ˍ���UB?1P<������{�]O' 7�d��_�م뤡׆��j��m��ҍ�^�� �gWӛVv
�D��D�>n���!c��zu �	̤�6ab�Q}[�����ca��ma1KG�����sq�X�^Z��Z�3�=j<�{4�g���t�M���[���&륄?�O� �:�)��Q���J��
���f�s�W�E2�i� m��"�1��F���^�l[?[��e���5�./'�ag8&�qz�����mGo�����䯸@���)M�<�r=lJ���,������ ���¿��n?�8��$�/i�I������,$-}���H9r�� h&� �����!r�	[�ąE�W�j�d8|u
���!�D\1�4P�쪉��{Ĭ�V���\u��SfK�&���2�EH� _f���̦�X��zi������跨
2/K�$Q��f�[���l{��s�'��`NB� G�=�	��p0���q�C�j��ƾ�妊��=��Ѓ9� Zz'V�T՛�hk)�)T~Pٺ�F=&��}�u6<,e�;��i�ֲD@-�t�Cp�|j�C���/�Ğ�@㋛A�^''7Y����θwHO���pR�^��ID�º�gƊ}�I�-����O^�:H�O�ӫO
)=���ٚ��JW�j�>�[���B*DEz�^� ��tp�mQ��w�Z��eE�v�����nL�u�C��ANV����frG1i��e��"�؆��1�$�i��$0��V۱�*OΒ��ˑ^��{(�c�Blm�h���N�1ݣ�Ϻ�P1����*
����m
�U>���I��u���q;̎S����\�X�yj�(�U��yJ���_���igw���Z"�L�E��d��\���*��̷��&�G>ZSI�>#yqVE��� ����*�e"�N1��Ǉ+�o�y�Sۢ�Y��/����857�֮Maހ̶+�����W+���˵�}���E��v�
KVks���vC�8	�}y)�.m�������]�/����"�����O1a0�ym| k��!�����r��<��F�I0�IW��dyf��uEu�/�"��Ù��}���.X��[C�� e�jM����q�^�>����P���u��d^i�V�Y�Pze��ɻJ�xk�vvl~|dMQr ��D҂�J��>�Y�T�Y���dKn54=w,�Z��jJ�Δ�Ҫ{�2�-U�7������y#�sh�
X`�l�Ɯ�=ҵg���V�j}.�V��������c�z���K8̼�m}_�и�v
�a[���ۘ��!r{���� �M!5�O״;�o���j_��@�N�����R0���ƪS+�a��Û����܆H�z������R���7�m(2��h�m�d�l��,S1���T�H:	���0�~r�ˇ2[�U�����U'�J�{A�����J�K�;�ܩ�S~n���~I���)��#���;��W2q�x	���kνwOSB<"��Y�E��?m��-`՘9�rk��MTڧә��)S����f�_M����x5d
Ct�,�:����o���<5~@�<^��#���fE�3Cc�"�n�7!�`��m���WǨ�>�&fz��W��+������C�I�hM�iZ���y���!){��d�H���%mk���I9�v**K7x=fљж����RFn��ZxzX��T�pK>��O	�ז
�|w�h	M�W7�����Q8�)�Ѹ1����f���Ik���Y�������U�����\����/@}���|K��qˡv�Y[�# *(�@0wm_������]~#[b4��5�����IY����#X@�1�z��}c���.��F�A�#�I! &��F���M+$P�h��(i,j@0R��	�i޳(U����::׾FX*�/!��υ�!��]�����>u�͕�w!��ơ�a!��+�ԗO��;V&�X�YP\�b\����W���+�v�U����;|�=��-z���-,�&�@�}��
i{T�vmӒ̲B6sM���$n@bu�HUYtC{�(�3.�y�LH#��̀	�ZY�
8g�0X��އ:�oG8d�'�Ȳb�眺��qۇk��xXA#$���y�~�E<���O,��1�`�g"�)�>�Z�cӁf&nz�3T���:M��d�ͺ8�x=��_6[9�e[>㋔/����/�*�e�y8�׻=he��mQ�4����.�v�0�z=��y��Q����>��_�B��wg���Kz����@Y%����9
�F֟, ɝ>\���v�@��I�N�N+�m�t�l/t��Vj�FcV�͆��(d�����D�Hd���tߋK`���۹e��Hޕ�n��T���2~�U���*���
R���#R�;:N^�/��$��k��dbΝ��}��s+����,$L<�C�N@5Rm�?�ّv,цG�hQ�qy�I�W�^{���@�=�a��� �F֮�y@��I_���4��l���b �Z���Co���:f�-V�<��h�X)h&6������bBbc~��Ǟ���?���rt^*@��l���{}ZB���M5e��������j��k��K�`�s����d]�\R][�	q�x�:u�ݢ��.��G���dW��6��u~ )����r��PkY>v{�w*tU0W0U����B�0M�g��	TN߽ǥbPJwCˁ�ڞBa���o�.����@wԗE��:���8
�9I���˗Q^�}���k���8���v���R���ְ�")��@v���W$�2|���^��z��p��~9Jv�s8����-�F] ΥN�V���YCT���p���ݗ�����_���� �Oz�W���k�'�����VI}�[�5\��ʇm���(y�Ԑ��"�t�����5y�,��Ľש���UIms�{��@�9��˹$��6�ڻ�!����m`eA���\�jeC�������!�N��k��4��O�~��y���U�:o�Q��x"�w��0
$�w�-hh�?��ގ�����9�ֱ�,}[Y�o��$���H+���շi�`!���%��1Y9q0E��5+��z�#\�lg�*��)�	E������^� �I]Oar�`��'"l�a���4��E<05�J�{�(��k`���W�AM�� ��O�x����D����3J�g�=��{�N4��z�ޓ^z�
�td`��+>9�T�@�!DTN2�rF�T�֩�		��i�S��c\��2=Y�M���0|��l�m;�DG���1n�Hv��!^�F��,�U[��g3N�欶��j׈�aY�+���0#q�ŌxԐ<z/�{Y��q��|�g.����=�����	r��aR���$�2�K&�7�V��Y�v�V2x?��Jn�^�.���]Y���fZY�t[���kQ� �����-GF��K M�s/�N��˃���x���:�}���+�l�����𑚠�����n��|@�5����'����S��-�e
H�&���}��ϳ��N.�!�t������N�KX�oH��;�g߼"0'5��CES����
8� t�wW1}w��L�I��'wH�Z������7��}A�U�ӓଠ���_�E�<�y�@�J�6��,�[-�4�g^�z���Q��K�ϖU��i��ߚIX�����-���`��!1�b4�/��������6�P�U�?��t�l�4�S��{��̛��Ϭ��A�v�[2����W�X�4�x����rҬA���Cc�3�0��'�*zM'�I���ŢF��;�4 T����$�Ằ@�ŵ!���^�ڬ#�`���Ц�B�\�ö�q��7K��M�y��&vf&J/Z�O��30ʺ����P6X,TS�Ñ�+��gON5e�T�V@����"�Zađ�$e�K/����[��Y���* u��Պ�4[Q�<��G�TJ���D�pJ��3]��EڽU���L���ط�u�^��
����e���<첌1�&����>W��,��{ڙ���s�N�S	j��z�/5WG�Ey�V��!8�d`cgv��e%��{0g�Ks$%�*�e�鴺�_���!���8�W�p�i@o�"D�B�cV�73�=� ��T+�7��<<��&Ȩݝ���g�W�9�0УI�Z8�@/��{x�Pj0�5�J��b����I�DTe����]�9&�>V��u�~�X�?�	���l�j�-, S��MR>�������tֱ���`�}�dӹ�J�3mN�ӲC�^�pz^%�uKsً/��H������AQX9* �
�"�s\"���\�l�ڧ
�����Z�5]���
�&謴�r.Ŀ�vD8��q���5U��	 �V�R��|�[^�g��NQ��2���\L��6����n��%��u���
��B�`d�R�$vk�x<_�B[��*�]�~93�-�A����o����1��7�z������MmRqa��#Ƨ����3q����D����BR��;��eW���
8h�m��A1�;���T�,�i7���=-�ʞE*�z���� ���4��9m �Ȍ@>����j$�x�=�<��oc5:��S����X���l�!�Пo��>\���ɡ���2�\k�����y�,�(Gk�(�M������QL�6y侾�HN��@�w�y�{=�����64����l���� �A2̮;N��'_ٓ��)��6���O%NK�J)���E#��?P��|I��.�k`� A�|#[A0K�}+��٫%�R�b�Y֌���f���ᛔ��Rl�Qt���a:Ψݓ)
��ڣi��v�S�����t�bw����]�7�9���vNmx���|(�M͉�! ,�zk?�Z� �5���Ԍ4_�����^M��Y�.䊛��*�oi�`�4��tEY���o��-�jQp�u\gR���:K��;n���-D/�c@4 B���eOt)��W�0��!쬄��p�� �$I�3x� ��ῼ��<��Ą��=������!J0�6�o�q�`�a�Y����V���a�˩9��*yrH2GLy�e�Ai�8����ל�����;	��a�Q�:�¥�-�&�(|W�n�r���������S�w�O�"��t� S'\/���s_�5J�f�#�� ����O �5K�����
 ��J|��d>��x*��+i�7~�:��!x&�5P�G5��J1R�8��'(`\Y��_�-��'��,<H!���"���i��wJs�tK��r%��U�Kj<G�jӆ��Yr�ۜQ��\���y��W<�Vi�U��=d"��Y��7�rN�p�=W�����X�c����ЂM��$���a��Y��Ζ�&m1\ӟ��;�J��"cq��r�_��E��S�J6�J7��8�;�"�x�!���ϴ�?�%�ٓ�|�Y��u�@'H��hz!ܱ ĥi��tt�;�m4��X�p�J�;ϗ�"#��	K�"�W�R
�ŋ�{��w�u}m���^���
d�.�BՃ�n+���6�}���I����5�J���.���Ҩ�l��{�m��O�$ei%�dT�\�@��k�&B�~� fJq����ٰ�P�v�5�2����{�QS�Ѓj��U`�iv�^I�Q���
<�4��3p�g���6yl��45 B5rd��^�%�]F�͒�荷�l�e9��4b�/�T�̑\<Xs�I��#��hqH�#�w�:j���b./Ű��˟�w��*���EW=Gr�8.t�^���*>/@XB�IeS.ԗl�KZ��By�W��5��� ��6+�Pz�l8EܳXD���T����h>e����GB좼@�I�"}aja(�T]{��3��u�Q49^8�{��wd��UI���_*��8?��߉5�c����dz����&�㷥_�r٤Eʫ1�b(ȳ#������]q��ܶ�����_���o|�'�`�HiPn!��|o*����cݚ�=E���:�H>��5�=�*oD�$���rQgz���|�u��ː<$�wW�`4���}�_�L)
����Q�%�:DhY��?��^�Z�CN���V]�LJ�т�[A�\���[��X�FA8����'o��x蒧��7=L�*��v.�� rs[��T��t�s.�<;}�&���nc\4f�U{�Phf�e:��.(�=!ܥ�IL'reC�σ.Ln�Ms��b:vY�z�E��t��T���,����z��W%�X:�E$=��c�¡2���k�P�-ُ�@�7���/����0�l@R�MgͶ�a��u���qq�)r�4_Yu��T�ue�a��U������˞���h�5�Oؖ;�XB�5[l�#�e�o���8?c��*A���Q�zth���BƧ"V��H6�Ҡ�"�Pؾ �J�����_¤}�F��E�=(�ʖ(Ho�bz�0�1vv��/a*��?�G�L�$0����RX�!��gS˸]��9�hj����jar��t�1�7,Y�c���9�5z(�	3E�p7��҄Yijܹ�h7Q������W�֣_2�,��M<dKdi,|a^pRI��AU����˘�I/��ɍt'���Gv�Z��#80&��P}���+K�����#=u�|�#�8H�;ٿ�7T���=r��/S<뤲���:�#�.B.�/���m%�.��|)f�Y�������P����1W�7�IV��=��}��(�D��Z���������랍���<)�Zy!T�x͔p�y������Uy���H���ti��2gJF%�~Y���"_[���`�߉� Ie'�ǋ��ߜ���h�A!��Ѿ����&�X�L �Y|7,#���Oa�������=`�5k�\`��*ˉ�$�}�����ҺAF(�"ū������j;猇$"�-;Fy�z�h�A>�{�UV��<�$�;$���~luʹ��۳=y�4�Q{Rj��X��m�����e� �l;��<�)��x��z#řB��j������Y��,ߦ��];�����:S��F]��9O�	�U� 섪xK���5�c`�!a����o�g65�8j�����d�����?�mT��#@�$��BN��-��*���k�R�W�UWBq!���;��&��4�srF�	&b��kmZ�I��>�1��(x����^^�0��
�^P�����'��q+w��{3zE�<�/�����q����^�4";�勸��ɏ�+]���2үL���oݍY�h���ꄴe�IXv�gt������QƲ�/��6ןn�Bi�%>Vђ0�I��E�|�(��~�9-�7�L���>v���i��(ιftxIɜiAO#��Z�U4hc�l�,�\˻;����)���VqPs�K�����v�R�I��왐~��D���Y;6��ơ#ˠ�\��5H���\=QB�Eˆِ�$�w�R:< �2�C�ŉ�~_�ɤ_EW�	=�j�X���*�߮��i�X0�.G��F��������̃�;O�ס!{t�1M$���f;���E�n!}���_��%{_�}g�ˋTg��}<дM?�  �]D��$�O�ƿ�E�xfuk�٘�� nc��S��4H12�vȇ�[i���2��|�x�ъ9C�?U  سv�	��̺���?�+��r��V��UK�W��d�%�I����G���7{��z���5�	�(�w�,R��~�*8�/n�J�;���{���1�\P�}�>������*���K��韽��u���I��r��"��Q�Y:��=��>j>yx'f�g��s��a�/=��)�Q�<W�%I�����"����j��eɋ V�^%V+Uk�����.�a�X��� 8cX��:	��&⺴H�ST�
��)5u�5v����^~�Sy�fB-]NH�K$��5Ԟ$�c -�_��A�}��	��xW��P����˫C�B*K2R���h�Y��0�ָo6���v����o|�#��P!�G6�;����K���pWc��6���c7����,;b��jp��#�x/fӅUu}���	���+ObZ�[߉����#/�|�D �k���n"V!V4�e=�C��>�	B��pp}e
�w���w��3���2���9U���7��b��T��~ɤ��(4�Ri�!���YN�%��7��J)���}�n ѕ3���n;��a�9q�R)Y�@旀�����aL�)*��MN�]v-��\t/jh!	�O_+�7����+`�%��XR��Sx�n<s\RX�Rt�uŷ���%]ł����ƅ�&����>J����h1�W����e6'?v֢�E3z�k�ő����v�z����=�ֆ�0����\�)�O0sV������8T��\«t�a'���!�����3	 x+��qbk�m�O#�Ih�S�`�=;z���J��9����>$�;5�)�[���E��]�[�g�t�h}��6<L����g����@��o��F��s���!?q�u�$���d��.+�~$���he�'�1��^0��kjSw�$���O�'k�:@�>�����ˡ��-���œL�0��C�g�ܧt�PD�h�& $3��m��I6��=#��G�)��]e�6�%�ͽ��"#~�H<-��ߊ�\BiZ���N<��X6*U� xu٘�"�Gt���c	����Vh�޹*��B�s>��Yz��"׼e�ss;w�)3�J�_�&bʞԊ���e�~6��i0UU�-m�UqJ��0�p�UP�b8N��]cFP��f�I��ozf�J��=}�ՠ���@khY뼈c�_��KʽM^`Rו���	E���ǌ���Db]�9��=�G�Z>�%�T��tT.:��wl�3�\�o�H�	j
����ʞa��C�?y;<X���SΔ��c�TXUOv�F#���5m
��} d"b��W 1N���-��Ȉ�@jN�E����%*�jA5��/�FE�<U���M��h/&J����BO�(���T:Z�,R��B�M5��
�Ai�v ԯ)r��l�L�3I
t�YM��h�q�O�W[	�>�����h��d�r���~��s9�@�<%sesy�d�-3F8��W��U����#����@�~_�L6p��%�8�CsWY܁-K��/Rn�S3A��ͻ�nHy^O�ҺN�U� ��k�Rq xM�g! �l�<9t-X"g�p
��iZ� ��o����W?5��<�F�q9��_d��޽���?��ěwZ�d�I����-�ƶ�^dC�qHj��U�ev�����-��=}ozv8E�����w=�(tP�͋�d_�� �f�;�9��X�G!di�b��@��[֊�
��L����HK��;9�Y��˪��&W<g-�zL^v���^Fm��TA�YNw�p���d��Q�g�M�sXE[�������{� [��O�Ic�-��<�4:�����m��/B<H[^N?5�׊�Z<�pf�]�Ԓ��|��z��B��i]�i����
�Y
��Gl��2���p����?�~4-}�b��?�\ꭸÈ5��}����S��1��olVTG�M��B 5�}��-8�ݏ����ա]�V[�̮�:B�⮱;8����%\f�];J=D���k�$�ܠ�uE6����+����vL�4�YV�kG��*� @M���Zi]������z��B�mPn���R�O/d����"g��k6��e���-��팔�'�X���@7\T��+��-��8�!zm1m��|���]��I��N�j�R�x�x~����=�2��wB����Җ;ޖYh���F��҇�K�m��ݿ�W�ܓ�?E�Ç>�G[@k��r&��m�M�4��ݣ�Z�o�&��p�J����u��<|j�,�Yȍ�AFbI�#Vp��_�:�8���2[:��ݿw�\@7���ej�ȆT�1�J�����h��!sw��-@�S�hj}�o�
�o����rFG�"���М&�/���kψ����ev��G*{�˂90N�+��+J'�+w��9�#��D�7�*�u,�:��M��2����;��fO������#� _U�қ7?�Bi�m��4��}�	@����ygn��)�h�(7�-@�<�k����j�&���e�J�5�u����ܭ�����u7S�֔���B`;�j	s!<m�[�
9��E�]���泮�����BG���qŶ�ts��r���)��r�w�9,D����,\��}ձ�f�+2��"����Z�.�*��EWO�f%�a��v)�`y���_v?�㔆M�(�r$�(d��,��&������_�շ�po����PA^��xƗ����LN�z�cC�"�߸9����n<rpK����ZVqH��S�k˳�l�ZIN����AG���2F�*�9QNz/i�+���p.o�SF�|�{���T���Y���
Xo�$Q�W������v�ݾ��?��޵4?����#��== ����u}{S�o�[.�+�x'J!R�����͡s��G�*�����T_=]/|��w�aA�j��оw���2����5�K�S��*XX:$���$j�|��`\']���#w!��V��SԄ��1ۢ�*���Y�Kmn#�(9eK�ڐ���W�c_�OYł��G@A������ֹo-Y�S�����|�
�B*����bqֺi����i3e��`���~��-I��m��}�g@�&���7�kW�v�\�%���E�R�zg��AE:�`Yn��ڐ痌 B�ܯ��9�9���b�z�M����o���!UI�Y[���T��?u�ju?j�Ρ��\�*���"χ�#����"�@8�,Ϸ��tN@?�ΡJ;mV3�%!u����X�:o��P�D{��{���F��L�Y�|�U�wcf�Q�GXiV�M�96��L�\Wzv���A�/x����D��8����q6������N�Z��7([�~T�2��#�&���u��j?E�����@*t�����]QVuFwc��jK�~K@�� ^��ܧ��0�B	-B00�N�0$�2��l���nK}� �`=ϣ3���/B�/P���]g���ى�>��@�ԛ�Ex���Z��M�o%pfVG�"*h�6�wH#������g+�������^���WοR^և�,E��y�����eJ|��#�(�W3J�����P����fe~���)?�+�k6EOl"��f���J3���3>�ރ�z�=pf?��G��l�n�iD��О����C�(��Ο���l�7F�'�-^��~@;���\��#(T�vSxD:���ʤ
��� �b���e��-C�n8�s�b���}�̸1㟳����)���qJL?6C�52 ��9n1��Rʀ����W�LlXަ�kIQ���l����(QW�ŷZ�x��͔ay
���u/r�n��MaN��ϔ�AY1}^פ<\x�������T;o�V�_*8�~m�^ȑb���D����>���F�x���I�!��ԫ��	�úضL�����������G{tbAtsc��?p4�uxF�sb��΍<~�z���&���fҙÖ*cޭ1�k[Z��1,�F��/C���'�W^qa��-X��V=�:}�(�.�E�\�#����єՠ�i�u2�%d�Aq�$#l�x���L�;�a��D�[�&��r�$g=���h�ߐ*�bL�P0'̪�ɱeN)z�G���M6��k��V�Ew�9n�B���I+;∷Gp���	��O��2�d҇\��d�W�7+*J�{j�;iY�^�Kf��U�p�����e�t�Ʊ��
Hl�e��|��l@�nװvQ�z�Eԏ�?6E����n�c�8h��شh)�k�[#�� ��9z/��O�յ�w���+�P9��V�B]�2�-C��X3��l�4���2�_� a��,��:�������k���L���*�����Ggq6����ma�A��
�p�M��=�Ɂ�b�7A(�7Q}ܯ����K��yE��TQ�g��<ZPU� }�W[�);h��`X1!�Z�]�U\AG6�R�����o�*i��+���J�k�W���Y�5���?�$>sm�s����x�*�<76���'+A���Z�������_�)n3��3�R�Ayr
73F^uF~�\�����]?���-�t�^Q��*�n�+��z�����ȁ�d��";x�X[�� ^o��c��%�?��[xS�r��ջ<6�AG_�3n�o")}�f�;�Z�t�;/�yw5Ֆ[����}^N���W��w�aC�����̊>.g1�JǸh^��g����ӣ���a��H�}��4�X�*.�}KE���@=|"z�b���k�ב�Ɨ��K#�{BG�-�t�J��~�}�F5��1�M�@�1�s9
��dށ>9�K7im��#���oCw�H�ܗ�h���&�u߬��CЛ�-%9���Ѻ�u�ը�>���^�6�FP`��ϡ���]J��)��~l�˹��(-��J�7]���u��'M�R?j����M�	[`�H3��J����,u1�b����ͪ�� -�ȣ1't�N�יq1Hu2�O&
H��n�Z@��T����쌦`�?�k����]EZ�m{ʗF�5n�τjQ���$������t�y���Z*�N�{mGqJ_���F�����%�u���� f�N����Xn�Y���lF�jP;�c]}�b$�þ:�a�F�s�:G��u@�?���P���{VZq7\;BD�t�~?��)W�m�.���I]�+�W���S���~��ɭp&q	k�SC}e��elS^'�̬��6�ׅ(y��-@dۙ}bt���k�ٴO����Vi/��:X��!�%�2;P�0X�|\�O� ����'���1`����7,|�:�t��a�n�:�<N�~��댯|g}��e�>/������u\D-�O�׊e�u����V^
�|�1�'��2V�m���!�>(�.��h��S��|�ˁn�9��f�����=�[�{:��Ʋ?����:�0����b�7T~[	��9�"���Nֳ��h