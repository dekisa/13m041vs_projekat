// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Pf62NNGvoMwTk88JGy91PBi58MyRvdp9SeJGtDj5qspVJgaIezXrx+y7QGZZm3ZRFUNVgvVH6Ru3
0lhQ0rxKT1KC9yFNhQPesRDSZU1gWFWmICCAMLR0Cz+hu2aeSqnoV3Ga/WcFMyHwKvcOCYfJ+jWk
rF5gxHiiAQ/VZvWVE5598GqWs/7a2lOCHCpQ1iOd/LozmdpUhLdfM0nwEQNU6ENAQeurFwDwWwVZ
gU9Xl126PRoABfBoeFxf+3lOiSUiCsNAo4BdpUih3Pt37h+Qy4IsnOj/af+FkeGRGyOToh64JF3C
plDSlLqKrObarPk/L8Uti+ztx8K/qaZp1VkdCg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2096)
HeCHlUA3qOV6DvBxEvA+v/ktcnrbzEiFT07638A/vOATXZHXD4nw1Dd3aIGMFI751pv3RSPSUzta
nP3nSjO9B9tbW89GCxZonmZFlnTiG/88D40W5vRaqbf8jxQZFzOJZbqEc7EEANm70Rb+ht+zC0pp
gHhWAw8uxin9odUGJLJuinhocT/Qg6m9tnGOcGqKudV90W10nhDkmto4tJJVavq0hID975APn+Gy
4wkQc8JykxE1E1kblNTJBCD8LVPnjqnRqO5YqoPttp4pmhjcrIyzYIouSSdvfrDGfuqAD8Wv2rNL
h5UnTCQDASOuT/p9M8wO31QwXsDNDo+YLzIk0AsPNb5rsqPcMLt4Zy19r7/4vgNt7sjzgy7C4+9w
7O9mgTaCqR8pNdFGtXQq/nnwstyn69m083836CF0rPmC6IPyJ4OqkvTjQ7qcYTjPCd4jNzETsd3R
z6SSgSOtyeS5XIOtHDJigVNo5M5tJATZzPr40lG8mhvJS53ZJNAZCxEz867jstSaGGuDesuOkZwb
n5vyy/O0MPuK6KcANTjq7XjpSurceIGIfHCm4ZKZdRL7mYXLNZLILByK5DSQjxo6gvaA64LThQ8D
vNHgKhhcE2WZlw87oWmOrbi4ro99QW7YeVN0Zn9OBi3LMnmEHp1xM2mRtFjGVufREk+FMIubquAF
OuzHM7o6RqFo7JsKhFUnMkKEnE6JDIdYZL/ELhnYdqBjjFJHm1vyg9BgJHR/QjEFMMP+lkqYFZ7u
qK/qGrr9sV4/4n1ime2svy3VzN80QaX+f/ZbFXDgpxJmzv+oIZieUbTQI24utwACAfeJ6rXuLWot
ejrGs5RJOZ/iy7TLWjMpu4swBCTKLRvLhatMbu2a84WjbOxZERkEaoOIe16eiD3KkgdbbAtAcbKl
TbdTTzHFgk6B7d8Cv82SrhsIxU2YbxMOCWhbBtI+0SzkLccc+Cqh5p0Xecf5rXWqhoZkwZdUF4LI
u4SjqdFKpnoEVfDWFkmpwZ86U8uFKjGn/+xz1rsR5qp3Mr5kHvE+zKQorYKzdFn9nHUKRGAMpRCU
zhSc+cfkL4Q+LBS7mcSUS0PR1M3tYeoqFpPGOBbHlhP/lL6TKgs61yHHNi8ATCtqGYmyEiGYcYV9
LkPLTGtZW2CVM67YyTJiZzH7kGWfgkDFuw67j7B0oh8SO48jW5qV1Lqu/HXef+8ml9sq9lRTR9Hq
Pw897BcP+Z1l5dL9SRK/Pj9ZXGMprhBkYftV6x2mWYEuhK5FY8TPCHeEhhVZqGbjV9K9kqQMw8PN
O/Q4hz1l3o4/eSEx3tSC2MRUz9OodONeqPj+ydBKLQe6hbQVhEggjuLEcCchZ9zLZhSuKNSGczI4
ZcqowjA0yU0P7huKYb42QwXvOgYoswBKm6wa2uh7sOCosciqLZg0lc1NSEok/1W6F5b/KrhWFaX7
OWXZqaXt0UtrCeOTVvBHYOubwpAibYhXfNKEJ4t5rIg2ekmtY8PIvZD6c9Qu0VQTs9z+fXq044Gm
8VlE+ee3XXcwgiDXNWqdCJ3nlVAkUuK1ndDXedBu5OV8mNCMtu5gqjzF2osjeKo90lYsLC6FMWEs
PsN1+v8t6Ih6wHFEmnAzkNgagRHcHVAduDOUx0F3FJIqE4PmZPVB3Ll81Wf0ljOdCgJSib7kxpGb
LfHkaujhLlaUozSD8S4MvOPqZ2+hWhMgkDyoepM45/Ma5TEATGJSEVdjA36BZVPptoiScwZqQkta
V6aEPAkdJ5KUJEpYIwBSjwmBGDFVkazsPZ1Nd7K1S5KwNpORcMKjsRaJOcknUhssZ4wYmkuEvCnu
6rgwLbHqLcu2zbOfJb6Q4NVpBLKtWvyVyfvBbnW1+r8Qf387kAsD4GRGx3yEQ6nfd4S2yYi+/H9q
lqoZuwwYFaqnCB/iYh96a+5dPlNDeuCTNQLg6eFh2ZWe3eFGuV5A4PuVtc+ctEjFZCPaZEc9QOYW
8yjKCpgJXmOJEuuGRJjUblYEmtt/IHgkvFuKIYFRb8A/iZy4RCJ+apwmoth7KjIbDpNUwZGKYa0Q
ABvQoe+pLs0jTWx/4BxLD5xdjeUVmSZ6klTEBScrT1jq3e5KJUTocX27JR1jSphqEw23sj5jZTHc
X7sw+LO+FMXAd7cEAL7EzyA7I18uKE+D45wvYUn3IDukvwZgFgsD3lKfTRPNwY25WfdikxEV2S6i
gqdpVDpJMphvvLZdh9C2Pw76jmZkNmk/g56mLRTwRVNGKArZ3VSW42hgBAv2fsWpj9KAc6C+szdD
/rXCD0oLS1UU02P6Ejn25ccClkmLZn93pqH2pVOubu1nf5tuXfDNNHkrb67VyOJNa49wRtFB86Bz
QvBD/pPhw9Op9EO6lKbmU1TB+cmnl12k9ju+NWxU9AhoGs+uHdYSUxQVdXxafALNXg16q/vAv8cE
FvMzez5ZJXUebN0sWN/eez98lpVrTgE2/zgMjBntPjB/66D8kGu+sOS57c+f+ZSEXa9CtfUmU59M
NcMNGk9M1u8Tfy2KtjiMjChz9MU2Uf2mMDQnsPLYbVsmbGlyOPeT/J8I+bfHkjVy7nQxdh/kQZza
qj0ULNWXkin+KmywuEO9r2u1kPo/KHCH6YpL6lknyRuLcCmQ5YvwHEPB2slTaIB4pyZuOpD83vb7
nWHnks9Lj/optd8j19o10M40SYn6UWo7yyQx64cRyMDRcGE5oQK6vaPkXdENsqRUNZWg51P4PExb
M3qGjXU8OPHIPdr11+bIq6/Q5JjdYJRNvVfQDf+bBjeYAKsYK7XFsDl86K4=
`pragma protect end_protected
