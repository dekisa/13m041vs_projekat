// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:16 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d5wcToutGT5/PrdJfzuDRUGIX+RAqL9+4mmK/HjmP/WiIHnx29iqP21kkPcaCm/C
at+PUfja91kA9AE1kFfvDWeErHmManNFKpJoSw2+bNbnHSrN0+GKmzE+0Iovpsv8
pjSuDW1V1fbla9A/x68huPpW/nZ7pJkDn25cy1kDhdg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25200)
KiStu7HvSIboLS+Fj6Ybf6cv9BT+SNQxY4j6u3a+u1X3nrPBxi64RwWw9Pz4PmXu
O5EFBhlLkkAILJvRdCfJkdAiZxxOnZ9c7l943U8LJlqpkfRsj91DnEKLjG8b2fQ9
QFfQSgABwqrHrENNIrbbtHXNbVJL/FhcKN/9yqcIrK2O/3aU4tLWzc/6XFi9kVl2
vAepsxtnVHrFOBqW9oUO/2Hc3P2HuyviNE+JQjzz67ZZ2R1twGOrdVYBXSJY3BDA
u8comO+eCOgrLq5XzLvmqkA82zQZofvGdbv9JDsf/ZIGFyZ8JN0Hmar+QenXzANU
cLFOw3NScAxzMvFp5Kho8jq8ndrpX1WgQ75S/ctyjkqeDwM9zYmTbroFkF/MxH3Z
ufGjBNfwyn2+8qKZ7C2EQ1qGf1CE+iN80bSCPJZH55RY8JrEBI+pTmnX6hc+R7hi
Xih5RVEiNTCRTqxEWtCNhdFBT2Ik6CFh1fTDYbkHG6h3x3NSqhNEODlzUk5j+thZ
gGFaI0ovNf1i5JHpMG2G4aGyFnLMvp3N2GNtgKFqH6ovf/OuiW9c+L1JFbVPqGbG
QP4nwOU9Y7aCrBwf5xfBbaP38OwwhkwO2veAxWQt6EZi9h82cO+2NYrhQ/AUCZFF
mGWqpsHw2icKg5HrArnwyH3agnAdkMlXOS5D/oXRUqaKVDSTphGjk8bFb08hJLAf
0Z6T0uLJwYr4lb47JSW/mIhHue8Kx0JXRzETYvA8/POoX0Qo6KKPkBSIWL3vfllM
23U87QI8HYWoGz79MUlRvZT+MOvDya9lq55CdgT2J/9hgLwMWaXaCBETlPSFBf0d
QqncCqzCPnbkUtgQ3lxWAii0vnZHJ4G3Wxekt8zeGRV07jIk/rvN93XE0fq7IbJa
fxefvvZdiVN6RZ0iaXS3wsZkdcNuaMMjZduIP4zmz2JI17qaJmJGGwA15wyWcC2I
A77OMyV9lW29V/dxR0nfUQphXvRHLnbNO8gazqByEcEy0Jy5uGZnqc/CSMoR4LIl
JT9jcdAhsSRH3uGNYFqMxL5jqMWoLqv6pGsEwblPwUqQeTIt1FyHKTBF+fu1XXmB
sFZZcyGniYafLzhgvbsZ+Brj2kClgsAhdpwhcDFY61fChuh5VKQtYcMZ60pQBVWX
4cbH9L83TYZR4v/sYTvnSNPig6Zvqc2UfnY00jNfV1Eng188xoQahS7JJPuhvsWY
2k4+KfQEYY4CXZ21V/pOQVkqLEOCPhsrF1oMwy9u65u8sk0EZcZ2h8EuHTh8UC0a
XIDiwiAjx2M/ZlhzYXD2A6Rj+n2eSvhry210JvqIrVVYCJGWer7tGnh5rO/lwByz
5MRERG+aDxgSiNKSQHpwzM49N1A68Jx/k5jX83MRBk9ljwy/yHKjJatKbCbuPTNb
DVTqKatWjfguO/OAnCzysj84EbMHVn6sWD+mjtaRqv5p75Uzke9tcjlWfLcRW0lE
tQJnQ44hM2v190Rden0AGIypYsBk8EewjF7LOo6or0Deg1p98IIsZhS/0etXNXBX
YZdsRSDYE2kg1k7IAZ5KRYqQVeWxAwI+cVbcYyozKf4r35gQOLppDLAMMuIWD6Z+
kkzBI9FtdXgrZgVJ8QD4Br4EKyFBvL3xGOamMVjTVgwfCBJAMbcY+8DChdiBrZhO
vSs0Fjy312Li43++yJTmq+OSibd98K+fK5WiQ7n9h45bH+v2+k/S+qbtGG0iLkwR
7qYBpF8iQiDX9h+I2wS4ooRfSGViPn83q7iPi6t1LunUgZYdRzCbY1fLo1EbH5/B
nKrihloPBEjdW48PtMLOysqGNfyeuOeu3+oBNPpuvCPCO5X4T7sRbyBcxe/SVVi9
pM2DE8axy1qcBuj00wr+d0hO9TDLyClbHa1JStbE2UV+TY0U3C8Q2NXom48m8ggh
vK1/SLy2TCWwdzCMBeDW1qg0iyLRPWrBjz99EBXUAwZYi01jJZ+oRGc5EBMrx6Ie
03YXMJUCRblhMUtlOMZzxg6HFNPf95CndHBBsobh7cxXfVgQVgjkXCIU0L5mOYUA
lef5BhTYhMWmKTmPnfAGeNfxv1DtRWyRfdPnVGVc3LbRwruoR2OQmxlnLZLYO3st
jmWqR0rPG7yRBonZvn6+MqVHaIyqgf6GyKcWIbU6fS4sX55mDOzh4VtksJFeXX/6
lplwQ9c9fFRS+iy2RgZHFj939LGmSJE+45kbnBFaVDanvgsl00pxDZqu8p+HeJpa
xjcxcqobxkuxtQL9+dmp+pf18nyAWOz+HZp4wsiuzzm9fW65XJSMvhDdg3BrjsiN
Nzr1rtCbnFcouxyXIqkV3ORqejOd5rvqbGGrXV62ii5DfuQOzG5uT530QDD74KrP
8UlerHk5OpcYdovFVHBnVLFvCceFpwGZnEKaNQP+zzffAefqknGthcRJ5QgMal7O
RawGLR+gKMAm4exWEF2cY5diSTNe9yxK+xLqRhZRYYY0o0Te4G+JSmsYhqAqC8ur
gAHs2HXcwuYaqx7KH/Sj9nH26WYz0xa9kscKT6PLuG1mo0r+KQwzwJnrkF3NkVDx
6pWAnOlnIxY749TuqrPpM/d8Cggd0EulJEby+74mm52Ucu6mWCwS2QDFatbA3rk/
BJhBFSaBmyTusmhV90egiQKFQ2jYNezqssulErxC3zdfS1Hty8ltKbPBBeELeTAK
dGsODz65XHyHae5MlXQuBc3WuwxFfJM4YkZT9H+baCFs93lt+5geNyjcQp+fNxpb
hecqsAia7NswJsKxgtK1ESzsid0gCGiuHUJoxvQB3VH6NtkWDeZYPF2YTneyzouF
R5pWXUccg8j2nJhMgGz6HSnMItYxGGSilbm4ZSGzUpbOoHk6TmmkRc1xtXbf3j4g
I3BX2b5xE5z4S+W2O2RUg5HnKnNZjTZTCDcLUSbS9nr3NJEWhYEhqJpiHZmVi2WT
L/YrSCqbwc9g1oyRljytuKeEhepMb8Yg0SpchLG7PLAw3ZmL9ILBWJi1ZxpOPhJF
KyvzwxUYgo2tZX1nvkxkhuJ3FzsaiwTT8ZDIW6qIywnJWERVmyQgk00CAKdYTtOc
XoDZ1Y60bFfTrQRvRhLTpg0FhH7gel/7m3G7RBOtgDllfxoSKJp8rSi0qAS8EAFz
OF2TY+8YUB8QZ/5fzoCCnKAyH2paq6efT00PlvFjzER49aJBmOSoVg+bHH6EVUDD
oZiuznsldf5XjoyErlugEFo8Bex6WCURKAac615GDtuLW8RdLnbTkCmm3ar3Ioxb
jYDA5iSgttWKoOTQPJrhim9a7sLHJRyvo/owMAmL7QNJ49RFEPmtQfixhAD8ZaIL
P0RgE6H8N1nxJ70qjIZHTRJhgMIERNHMEsrPTYtkuFC3POKJnbJPRk5q06XC+3SH
/PfUzu9bp8latAeiH3T3zImmNtLwkFP185fox8LxjfLAGYxQgD6eEeHuRFIlS8Cu
1c+B7tEI3Zfr37HaAG2v13hQvxDhvDLsQm8Zf1q1dvXPY8yMREMTF0pSxUWU6wXt
LVpVLLiZtUv/riChbIKKTGlJa2Zin2q+uDIR2StPC9zk1c8PLizZEMWC5grRpifz
epqWtf/YDW8yo3S+Olnn2/Z8LV7+JFasFD1JxHEb12e2HkKg77WKe28uJWAjzzaA
kUX9MAcyaGWxiCK/vL/pBOp78QKtQ4mzv0oQZqvJW9Xu5spjFYEfMroA8+mXqwQC
/Cn2zDrpyLsx0q3+aP1aYVsG1cwG/MAi/E4QQN7zgH44btLBpt1X8b+0fycBJWl3
q/3EnVdzhuRQsa3aDedj/7NSAfwduHqKK1iCEUx+jkGbZjmmfgjiyOHVUq2StkcW
a87bBb6dryRp5qqwBJvYslyb9JVSG97Wmx/PuhZJaSu6aMnmOUKMymTrWrvGinfU
+qOwUK6cs2nwTTr/guqG08cBTHFsqQezIIRvW6jB3HTxer2XQVFsTDj4gxjibC/b
08KDv+AN/22lhJkRu4pEwhvOxRDGfUBO+4rCz/TB0oItirut1nr+UFciXOnnbFDu
jdMzoplL7pPMN6S/iuCjibNSymrEc8p/oj5JIyoQu1/rTPvxg5eT8uUMQeWDz2Ot
prFnDTAAcQpQIVNyzByrJ/TuePRWQ0RdVm3pTui4t8m47amDFQ7cKA+ed+2LfZ91
W5vYk+Pyx9j2h0XAiRUYm21S6AuhIsajfy8dtrqSCnT+dTQJxtMPINLYzc6u1VcG
fYusQG8q58mMiKAELDFGnoyvAF2DULvSptk7Ody7Xqq0IDz9NSYSv4uBc5MO7Z4L
ePK/FoagJBZJNul8lWfMCUmpp+XgR5WCrn+chIaseD5qSBBOHrXMJ85OpHrri/o6
FicPPcxiORzoXqpT26Y++MuP6hbE0S7TCmPlSQXRqwrseAO4cb9LU2kSmGJgidQy
In2GPnI54B6XIXz51t4iBUczEWLu7JVkA5P8HxngUWxBoRRW8eF4qJHdXDUr7f/t
JqM3aTqf3ZU7GMVXtz4Ifb00np9FJP6K/A61MJ1hiQy3thP6qPKUGk7XGn7SH/7G
WzRK17g/s6+mG8EwCakJ1aPKNJe3o11MPOrQNFhSOUcluE302rudzh+3C8hvffgo
SRHHqRvYp+Rhl4BgV8JRC21KklTj6YiHca5hU37cfPvO0R1VmiAbgF0PVu+ZH+4R
Nb+Jsom0OouA2Fn1phGvzXqEFmzubV7/KBBI09DgEDPNXbJnutLj+mDGxEnFDBDY
l5wg34YmVMhjpsZwXEVlZQi5LK+3JiEB76LJxBgZE77sikejrW87LdqSb1dYDTqC
gBuoFTriKf0W0bMxnVoaBGSOy042Lsycgdok3SYROWSNFr2aHXWppXow2KO+ghy6
S1MYyMhoovOqnuFAo+iLhMrZONhduR2Ep8VvTb+f947EZAzNmhVCv+4P9xKNl7EG
bY0fn7mOe+602wUOwbs99WP1I0j8t3Z1oy0frEvQYKEehkZttOxr1/qBGzzz1X4a
f26m8+kSTWshbt98hEsSlLOH6tg2KsPmfdRf1SlitZy5DM5JTGTMn53Hok3fy/To
Bm7x2sQzkB/snORzDt0/gPTDiZXNqh6dtpChDhk8JYOlcnUI+FXO50qctJ/OBDl2
UKpxD8NAXQHRc/4Q5EM1VuvSkQuXMwvIHjjXihiQEMggnEyzn77AE49JlxaoSnQv
CP/lHVVqvSRwwsCwASC9q5RWAm2f/s8ZHjAKMuGm4t5Hji0IBXN/dP76ih1yleM6
Uq5y8LmaHOiPU8KZ9+IVaASsrf/wTsUw3dcC2mjJoTIxuTZ/r8+xky1edU5gv7p+
3l16GnRwM9oEFEgSaC2rSJPizl3SGzhiQzemvAwqAOFgI3v4RPUNK27DTlIIeHR1
hKqGcx9OgDI1h87/M29NGShRbtB1RFgYbidbhqczeS4zs54OnadH7RbM9AgcVu5K
+L19eHqgCF0/FB61NnvcLnLv4h0uLqMTAphOIsIagEVfY3nXxwPnZ6xKdcIFi6MV
kf8JoxMGtZoSR07mWnDwuosbCBAtmonElMpTkrfEtNzvLukcmdfP0ee/OWxcHV63
sEXb0Sxhhn6NwLFlFwdY/GF6blwNp385NIgxZiV59FkSMAoz4APK5DA/dFAgwTFY
HzNXj5g8puR9agjjhVQ3oy0kDdor2FYTJgnLxaagQXf0K3AV8nXfQx9Q6MIS57tZ
85pOWeYGkE7URN8VbFjhq/uCVbyDKsrv/YxffPnc8OSfSTFb1s2+gBk0sSwhcuK5
QB36YDJ9H2KpcE3eQI5F0EiPnXrRT31CVpilBL0q5mk4QAfg5CJG7T8mcZ5iKIJY
Cf5Dm7KA4y7cjfOeNepk5IFRigizDKOyfj2R2bHgpF8hPQeenS5+C4IyBET1amwz
kNZfPZPqsOQFcQkTLkB8wO2qwAj/Chm60o5/L69gm36KXSn88y54v0BeJNjWzg/o
b3RDGgs62sZNU3/C5i+Z1NGlku0C7g8x6H3tPEDBweD1hLfurvuWWXnaLZ9ptSbb
BVsYiG0XazShifZDxQ5lNd/7CxuBeYwdWBlxFnEfe3lvLiaEqORKc6cevyoUgL47
UlyzDJcvhLotTFgdiBAkbLwr8oG391wSY+aN381+J/lIaUoTyM3gsUlQ27h5U4cc
mzigv4AmQgAwCkq3Xl98j4MeIIMEYX0t4E9ilFv9ismHWUTWDiBEAxugPWPEw3W/
EBNhPKmU35i1WEyyCCyavHGqN9APvU85I/uhF4iYDzSl1BV3Fdwm7LAZ797Il2qQ
HETAStn+my01vlkDeXAqOGhqhrpAOi5wiTBwngzayAWbJ+qqsK0hjjn6QiMQOudU
3FkWn1ibYxEdvCIKo32KqlfFUgop0wglhqc5FqqikG9SARI/xthcz+5yw8aknLzQ
T4BNoeMN/acHxypYdY8pVPvXb91EZF1He2JrWzFk/qFTsRujFplX23NNe1pukJ7s
KW8DOXz2e77VzyHoPEFJKoBW4973dC5HRMgwEMZRfSfwU72U0OzDhAkfMxkifXVW
pZHeGlrs8DeR4JHt+iH8oeVTrMueSzsyhZkmN+zWlmL1kp+t3mj/IwUr7+Hfoknu
RwasLhjSAZvJq/aDMM0qgsqDxsXAN9Bx9RKrMBKWtCiYq83dS2QbPYy73yZEkHNU
yrhwuiLxj2tC+GBNiXzFbT+sQf9DEKgKmXmSyHcoCRDSQyVZHiqLS74XLM9pu/cr
INlIyG4tsy1IRJjkvJ7PC5HSkROYR/nNOs9J17QVJR3zWmcIX6vwVbQ7krEIQcm4
7d+r5tZ3nddTwlzre8C2uI6ayE+e8FW6vmHIayXjgDyoI/fnnKuSEouMiesw9rcQ
lDlEo/DNEgTQ6QXm0zo1+0svFTDbxogc0UY+GBd5gdkRLoqWgScRTXfXOGZhpa7o
OZ3qz65L6hEEZA+nwCwDdKrroHqwtsV/tOd2Y6WEntrumESxch+IhI7vs1PlE/Hj
5KON1zBQJEcLYcd2Zi/K1nERa4fl02l1GtofZiZOdUZkXmZasY6KRdsq4R0fngeK
buZO7O+/AigPkoYsmd+DpVYn/KtFJ9Iyr0EZ/Kf9WmtTzO0CadgSqwNYRzB/tltO
RIckmkO3WBrk6jupdUbt6M5wf0tKmbbe9wKyjxFFWoRIVmGB1AqkFGJZgeamJP0S
cMrEJfI+AWyXUbF3i53mZvPxO4apimnNohIcIPCjSNvzhCvGc7UhUACbICIioCB/
kdQvc56ud6Mred/yGy32QXWhWzvCZ573qBzMgNf63NIoENRc0i3dOsaeKG9khVpb
GpibQi4PJt2u3nRJIjZAnXI2bHd+ML4hP6LzLm/8YtTcGJEw1KffqspWeP8JtwYC
3ap4uCsek9VrkdM/AQSs8XBtY/hSFiqFVKZTrJmedZf/gfxPmeXpGTk1qycZmwui
oqdY3me7KT1INy/4hO8sOOl1PD/x8gvFMhrlPp+mIRajVqnVJsHbirg1Al9Z7k99
UjWwSHkQmfeU0YHn12JlIa6160KjSJXFXPUpKKzRFxuM7N54R8ydNtw2YkdhIuGN
/w1Pk92hSDz42YwiTFiBvRyi9CJ3iUXwBsY7iIIiRuv82scFUkkwBhfPmqYmAn8/
7oGsdzAMKoCmecVqMns0gl0rYUhnjZXcvWaJMeIFMQyxAJlslOCn5qUdxd/xuN7b
2+bw0o88i+nGyFvtKiGZ5W5sO/vjJpMTErt22zkCkyodXpd/VNRx0K0Wb7BndIh2
TNIJ/4XvOFHK6dpujJF2Nj3HcGq38OrlUfpYhmagOfHyFTgzt6UnFthB5g0NKALX
00mMjDN1XcleSmpz3Scsd/d8HgkL/3+OQAas3Gl7r/CAqKc3cOjfgvq1i5ZdGf8L
MvtOe1G3tX0IQuAC9V2j+xiS6dUn7/3qhrwZkoT+CMNLjkSzSRnQPcVnSct6b5lU
Kyu7s/JLgxRi5Rr+b0p5e+Zqfww+jbTwwRZxgbmn/Hsy4vwwu56rQSyiQ5kSfloF
Xo8dMd7n/pCLKVTsvAEozxlCtCrwSqYIE0VrJa6fP/eexuk7tU6Z2TzbnJ+i3DOM
suaMlnq/3u+yf+kUZUxS7X1G71gGXnequNHPx1RFio+kOldrA7aOYWQS8PEwcSmk
PjU7CL7EeumHt05AlZTXGi07rbE3eJ/lu3Kdm7r+LZ9CAVC6aILhCaWf1oh6+ftr
QNY6gtwfHQPgnEgqzuI3RJNRxvzeGVuhSBu7xUv4n//E09mMkSA2muAiH/NfYHci
3gBXq3/h0ccALcWFB441MqRXhkqy1cjg7InvXQtUDDk8rhdqt5VnST90YJolKsuu
ra108gK+ifoc7ivOYF9KkfYlUdHj5Y86PxMY7YPcFhHizO3tgR4Kwl+D7qoBE3mK
C5XcIXuoG55Ca3+l1vIcicx6Y19FJt4naGprX8aB7lft+XDSqRxGC5ESlwLXbApB
m3UcWC1W0MuFyMFo11yfrtT+DY3yL1upKvm45MEFhDAAO00g7N+Skv3MEk6RlRww
YV5hOHB0lp40DOwd9xE2pBVSTECjDJpVbsZQaEMQ16EYNZgsCtyFqntC4UjQdBto
HAVvMzZZs9JXEPOwjpvqLbKsAG+IP6DSzRdCDZ2Tt2aD9EVIMS3femtK8fFVvCog
MuCMJHku3crohUIptNBka7+5Wln4Ld5rWtO1RtgrNbTSCZJyjVjxPXocChHbFrYa
+YD8p+3852Ps4igujfyFVYoL3vBfEbsF6xNFBnau790qA28uD62iz2o4ZHqoOTpn
igTLgvm6w9Ol2eQf3TLQM+AVDGSQy5qwjfAKtxaBX39ZQVXEpxANDbNi/cbz4AGy
cw4AVjQJLUPGbpRLGJZmQRRtLnxNWaSCbK7HE7kNdv8R2+5fODvIuEXe8Ie4/IV+
qtjWaBCMxUh/nd6RnvJUAhMOsj2CRUf66V2Bx9XIsQFZ5htE6y4rDenVuKHXJJzu
HZLgRfXmLWGlFjwn3Bn2yj01M9haAoGaFxxzI2HsMMllU1wEW3X8HJfvZXggi55q
7cbgRTesbgwKVkIP+okIYqQ/pQYkRfWPi5CI45jg5F7HkAxp+swC4f3qotgXn4Qx
9vXa6iVZHI23hDujEg104kI/pMXQanfu+r3HWsDPnOExqLV4Zc0vfwqbEWOBC78J
l2j3Ao9Xw/glj1bbK7M5JUZ5+bYz7ItPL206n4IYlAtiB9XOWSbjW9iTTntOf2DS
RUwssWWb/nbD/vtRXO2SZ34myDMCiJjg1Zbr16zarEYfo9qPViCntIV7BR0mQPyG
cz15YUTo5WEfuZa2/cqaMhHfOCLa6xwdBcbIhSzLF5+kWdI9PhvA7mDKW09Mpt3k
yYLhEn/Ok3PFYVDTRlOtWI7R6pXYhLJKibklU8BekUaEyYK3fWxUCWB779HyM56d
rvsE1R+ki8ypKTDvLP9iDaythXAwh712SRE984BMRmGl1i2lTLOmQ/Xc7cab4AIG
8nExHuZWy9F8a6Qh5qvtCguBW99luIkgkWQb3w5IuW8zTc4ceKY4kzDfq/CU9F5A
0y9kyMX96EQJzLIZoDg6QWtD5zMQblFIWCyZllwkdQ+6XIjQGXcrIKnm1Xm1JCEL
wIixVXENA0woy+c7PL0CGBelxvdBUvUoQOrKsuMNWA5ERU6MbN6/pit17uTeTsX3
kbUoIJqbhLLhfoY1LWkzTsLGy1sploZ7B46GONFCR1Bgyo6Pu4BOfVLWEOF7hAC3
1l4ra0xMXLvSDlK1byPDBq34uybihB1f7ij7JjMojToU7Abza425U+m62AQ31bxV
CrxT+CbEBxnFstsDl5neEi2y97oDZcPqZDI7AOZHM2lJrqZh9mgoe7Ir8s2Ygn8f
6lbsIWqKGF4qK+YJCajNmhuBAxFYU3GWwfD8ezMCxWLJzWG9GmPVSEFCKUxJQz4Z
GEIMDX6zKkwysuIhXHssm/53gHCjyQ+nI/fw18vx4WSSo3JKdo7cFm+80iaMj3+8
aAKYdP38tMOgKY18bigGGCB2heB1+u0mUC17zQQ0+R/y2DA0w/Vw9IaS+OIDyZg1
I7JnGmHMAzXwmhYTUVYo8+qFb/AigQ/6Kq+VLSvVA2msFlfsL7IjdrfOLx85r52R
UtnNW8PbyTQQRR3xIJaPcfo+KLYU+4OTYXw+xw5TAsEDl+x8m6rGLy76bUjIopft
6HQaOZ+B8LgURkfIacHBVPNSUSp9h929euaN+T7cDz5dD9lL4zsrHkDXeHj6VLKk
Xjvy2V8IVKGbR8FrLAV8bDnka6FGlIUbTZg5HOnq//RnbNjIv1iSP90ScX8PUdC6
WToTjx6Wi9TcQ5CLcPrDD4bzV+jbmr8RxfJMUO8CbMnrwsBhTOV9fh70phWF/9FE
GQ0c9CYJZ7NKFE4olvErngs9sA8sTYglp47B8PQP0uIn9bZSQmvNt01NXdsHnbI8
Yb/0S+fYElyZLPEX07zpw4YFfK8JcCJcoax0blGOehxZyYIIF6JZG7trtyGroicW
VJLtGmjhzFj/QPchvgFon5J9+5UwW38Re5p0k6SA3ULNyfY39brsza2dihIsxz3M
3hxGNM1DsD5Mk8jUnjToVkwKf6z8gV2Bx4Pk83eoDaOk15havOhJxh4M2M9wQ+w4
ck9MdmCysZFpN1BN627KQUUmTfXhH6bustFXVW6Pmbk4d5ErfazEchv2kb04likt
bI6ye+y4nU2+3JmQ6oxT8dZMRXMekTA7FFznt8PYTIjVHNxLg9gOv4STMH5BHc4V
s1yRqYAWTuD4ifOH4y12hTDvahuVywRccfoflZNneOKQnZz6wFx2Un215urp1k16
YeicW+lMOEp+L92r4C+u1E6GQSBkdU8goYzDPwMmy/Hdc1pwtKuU9wvQZ740y++Z
nzMEyFYsxdkcZrqGyC9WiTFEFSHm4c2oNzl5GhxS1/dF+otlJFpWz9IRfESqz1zj
QJcftwIvSxOOjrYAAxGhZZRDmAZN0poeBmd9CzAVFih5I9oDJEwL8xZqJDRmn9hO
X09L+cOikugktMbvrhjjccxIaEngoReN4UAGQUNJ+SPV3sE5ZBgdC77YB/3+bqV4
tfkcnrgPR7wLZcBzKcIYG6V9zVuKcguBR2V6Fc2DgAU0U0lEsuP9S135Q1K+dNQT
26OAe2/sYcr3eV3uPTFRRgU5GECJ6L1hasO8HZ/sS7kidU95Vq4iiMogbcLy0EBQ
i5+xYiONl0dmPLTmgBiouCKNsXyBnYIo56NXSHvNPKVchI4zNvy8RpK4ZY2CJqEs
DG/kA7eoD+V9/T/jnIs7LuBPyWXLZTq/8SALpiuaShjDOM6K0QIJBAIrgbb59mLu
mGN/B6Z1hvAw7zH+7rvuZ5Zv6/CbiF/LUvBJCotCXvDpLKwBrmOXbwkLi65/Nlrt
pfiUMa/QAenaVxUwuJSANsal0koStwoKs2FZDGrV1zx8WbAEvwXbT84/rs07la6Q
f1ur/z976TsER9CiysbH3QaL3ETgyxOb7MZGlOYy1GwR2K/FLQUZYqmc9f2V033E
p4lM3Q0FnB44kRzUP208sT909rjKJAiIu4jivSEIj9horDigoioWOzg8YouqxGs7
+B3MtjXPlfsnjSJpD70aILBnHzyvRvs8M2SIGoJLhYxwavhIkFGmbe775LI1LCgN
xB/kA3eLjyH8PaOMh9eBulRkQvnajXhRlDBlDsjZMlmjjwY4oljNyii82tqrS7Ff
buCnXI8kWaivIELV6RldwuZXxGwfDFoP7e/EmadebKSxfgb3+uFvrGGH6+TNDw5o
dLG2Ab3bFZEOazrld8aQTygdrqUba6baL4wdtGo64543iS1OARBPTTsBSbgVlmO9
SyY5SWO26lGphgGjsnspjkqv2RDRBJZZdOvOC3mdLu2vhmzGYAtlxuk4gMf0YLvA
FofZUaQeSZwpqbybNCouRwUEkquMK2VdycAw9QrbUNDelqZ7mLICWfdqviwYEKei
xrQCeXcRVc9i85nF/yvIx6+vHY/2cz/FhLCxu0dnWOcivkJGwAFCeJDbkJB/PI6w
SksNNG2k8UGDPfGX2SIO50VqL9p8YLAIZuKzvhdKm4a0OIbdDGN5Sh6ArhtbVF2e
DZ65NMcTnyrmwdqsjFlZB7ozc7P2uQc6ojBYUDboctybEmWmsRk0Zd3gZtknXSyv
ZXLWGQDaJtNoz8m6u9IDJDRfTmOpnxpQ803jevgJdXpOW9ljH6YBpU7uyEnE9QhK
fT0LWKEWZezWSi8ITbsJ20Qe9Ivu5CawaBdGm7E69GquW0qVNurgnRVJHtVxMru7
8TnVmD21GxKAX8kwoYn2GTEgQlqapDBBMS/eA2nWxEiqUzq0HorEPOwjCUP4xksI
GfkigDCKMzB6+ff8IMCFtFWH5fhtd+oK2SArHeZYu+BqUwmavphEONSa1infRyXD
HyEbco0Yx3Hr6M242Bc0hukVP34Rq2q0RzNtOYp+RYPMuOVvcarrZO1KYff5NV1f
Jbg5CYBS1QKb2z/3eUfbSBHeGUEinQvFz5o8g9euTXNrlSRBaNWVNBO/BLeIji54
xHDlbTKBMkYbyNbXkwybFBnSwKnGhCSr2AM5GmUU3E/lGmiTWpj865RxKNDMXO1c
dhGb+m1qp9KwymbgzSHhpbdNGu24/xjoF8gaHn9iit9t6oZ0KsyGgvdepNI9LSD+
B+ISzCcYBPV6f/pSWpoP4kB+SxGXVYlc9PbZKhpGIcmIdzilFVXhKQTuf2KMhBF/
vMbcLJ011fBjq4xUKU1dNq5N1Z7hA+0yFmA+oJDjITH/D1Toz25eKxL7ZuTc1+Ji
H5O6C8QytbTDd121Yc9fGT5VWsZxlo11zSTNXAzk7H+yjj+R4BVvC9QYwXEDfshh
Urp+9Rp2tW9O9M8uZJUFktS8CmaVekT74HHNOKd3ZAx3TOgZRcMSP3eBebmOg0+H
OmaIjMDNIQYM9mBDRccufq4WUubx0aMy6yuPVJag2ZD1602MoWkltk6pYvR2dfCZ
HsrwkttbMJdiHUQ9ryJyutYAEuBdefkN7XvAE3F6Ntgss7BLEtcQCsGqec8mlQRH
+3LdPChymobEg/XgvaEuhiexNPAFgOZ8z1GY6n/TDR0uN3yeaiOrBPLIA2araj74
Wors8O9mcLJ3ii77p4ABDcPZ106rpKCzXm6O0p1CTz01FTWSdFzb/kLcLTi1Qvx2
Nfwa1kIRtKaN852cylylW8X76/owsRLG54NG3MS2h5M/sWQj9ZpdzZz7O0lMEWbe
GnilCLrkpOl2s17zqkhon6N8mxji5MVYj8K2F9DLHJV08I+voDFsjG/S473oHkEW
8wJbHVmFDkrUUEmQzuxGcp3Y55aKb5BeCyHg30jeiNDDscPUuS3pX+i/48BzW3JS
OLXi5FSFjeq4xn7bHe+JuUTPjs5xxuoM9Cw2hQn1E3fLTLFMczkQfLS+1JGhj9Vy
3fOgu+6S31u0ZJt26TDWFA6YEFmM5ukhPYXxASpbMgBFv+3Ol186p9DfRhwuQSvW
mYGuA4x5ThW1yoQvYbd0jVsltEB4zn6LGMNf3OITkU09VgRkS47ZzcK/+9zQz719
Ex8+g3SLAQPHLp+DIJ9ulpVKZShWhiEXx98aYMeKvbbplS66Bdz37BtWZCwWdyHa
tAZV1GIRRUZ3cCbG/+EFbs7OTFNXFFL9774ZP/JPSfY78hHfnXmOaC97ypLxU9/9
Ps9tKTqJpBiMgxl+XL523vIlq0V7kb+PF21DnTXhFPic3r8fZwVP8/m+BEO2YzMD
pTIaemkVd4QBvOaszB9uIywiGz4EceXZomRnzAoSh+Ziey9x+9CPSBU3s7rFKwB9
5Q241cSFgVQKcVLPCbBrCmb2WBSrM+PYBrZTX/IM2l+nqj6s86U68E75RzXdqqcf
qDgsso4hbWNuGSnKhye/gRIHm5nLs4syoxyISsGA8nKfdcewPrhdCRS+wubdSv6P
XH6WA0JulzDDb/6vyobf5gpwF5hvQU9+Jv19NYby5SAvPsmkeVdn5py1smrPgdXF
8pMsn5dwClDekLVmkspTb9d9gD4rHfbVvkFyGxU+zZGMj9S3GYxtjk4+yCui4UTo
/LWti0X+Sg2TA7TqZcpHqZtyV3gxFLkeJZ0+G/tbRQXecfxcwey8cGa0sJ/mu3gx
+OtnkxuFfLBiYkpqh0eC4hTFkWctkprovPZfPfWcJL2xhZ8T8N3StsG65x5hmTSj
QuqsLr7EYXmdUmXjTmAgEIVK/9fWbKOJVqMcRAVmz5Mn3Hma2frDpZLiO2ogUQAe
POr7Qve45mvMQEaQzI6j3y7fbXl2sKVMoRQXAlp4yeCvPgcasjoaQDjg9+4YbWc4
xC26Hw5Bdv1Kxho4S11n1AUJWCpEL2UtQo06SkJz6ZnI9Y0vxc2HOVTUgW7ki3Ym
B8HM7u5UK7u+AVzvIhfxWFW9gxhhNiT67CbxB4kkN47eOGm6M/4crOEEMs1t8TMR
ZfamAjmjnwbFshzkegNYB3c6Hkm7A+MOUZBdY9oi4q1OOHakLdZewxc7aiShxfFO
vOzNDiN/BnlHK8jrz9v3H3/ofgYrLz2tCHrakwXJsv+uB7mpIvxULVDn2mRfG5u0
512DwHzztXgNoBHwGLrWto1CdLXUgrTO15oyY9+z06AjywpYdhozlwR9ayJmX+G4
LUte0uFB2H3kONE+TOmdCWq8pQGqAoVkvAxRNi42K5qbZ1rvApEyLWvNLpvu/bnp
Vxiv04oK/BImgUWyIJ7XLkCwTcOZievepd81fwI+6FXH2Gcp6dZcGPte+mNyVXrK
MiXdTDeDLkyjwUmW0/iJNwViOH8w4ZpJeEGtGPaBE6l5VB+5c5PaL8z2LQCBDdbK
V5Xb4ljtqArDOBEOtRhf6sYIklHXQL+6WV5SbBFlcvqEyMZj0ynwLiZX8taTVRuF
lt9tFAG6IFvlhQN5h5Vnad1xJjnAbmUgMgji4EY89+/jqlDeALbi4DzZslkOzSks
RRts7Yx7xD3DBMXOggjEcP12dkmqb1JCt0gc6Wn62g2njbJYj7/WplCepuhaGeHO
tBePsWTyUzIC3aIy0EIh0f5RWU+ej7DOYyA8Ti8x/y+my1rcqICtRq/vH0+obaB+
nGGIMsaWx96sECQRp48cL5tuB2rfBGflLUD9n4XrCxp4hstD8qxvXwFwAyLzngUR
PijnQpZQbfz4tFIz8IhIznVSxav1c30kaG/t+n7K7zM4JSOXb7XtM2i0yw7YVKrB
gcT4sXyv++1cKysK1RlmwWLvxwHT+D6l5RtHB6bFx4JBEJQl0aJ5wD/92wiJ519f
5AokM48VJxq//wLwbHIy3GDJrlt2hKxBLdGqgKI8sB9htF+pRPsZZiqDhAHy2ywu
K8IOpAwJ0WbOT/MDTnJs3yyyD9NYSZuswd22NVrwdUIXHYpfzvhg+266sY8Afngd
+05DSFuJQl75e9gMkyiWU632Ib1xt/KwsMad4pWHUkoVPVh140fOrziUypwsFS9N
nSHVWsfD8nwQHizPeAzrNj73pCc0XYoamRmvhc4zfvxzr1kfM5xr+2Wu8AXl+O/2
fZqoULtkTHx8wQRwjPA8ZHnO9+Ok2psiG5GS1gSiICzPIKnV+6IdvdOyTKLM0dSN
utbYQZR7pOES9uhVdbTCVG8si6RGSh9ioZDvEN7yjF2E9kQu+zg9d8bhyf0Jnrqz
aFdK67YvnuqKW/QRjCRj09ln7is8AaRG8K2Iu9XtNQriAPmFczeCLxveynhM+bIo
DZ/3284XvwNtQqgMzZKskuiNRcdmfiLdTifd3AV8JbFrlH1TjZ5sedOUrpa7yQFc
boiku1dsZpX5Rgaaod/GkhyvhIbToOGeXdvcSylnE3vA3ZhEog0VUj9nCUQT10SC
qC5O02t2wstUAOv9UuXMA+VEekcB0GFBNK0jCJ5u9eMBFESCu6Vwur0M6co5myDF
rewm6DSJg7DYETsnOFoOLCqQILVB4cbpLyx49Y6MHK7HzVdnsbvueZ6BudXo8uOq
JbW6CAQeIxTzD31uaXH1TQ9Nrab4hsBQAusscHiqtMwuM+Gs4WGv+8SPGEf/sdLw
gzH4T2AznSWFJdwY9MfN04lYtJwLvRS/ENWBlMX3pLcqKM2j+tDCuDdZmCvAiNGG
Dy3QIHsOL3KaGUPL40u6VeEb5tnDSPUnNl5NSBc9otpATb1rnbPaPiJZwr+Z6kwO
/N2JmNSqXuBWIIoVBe/U6sUjz6tsPLX0LRDLJL+Mk3YHIccldLZwZJUdCbVx6Mrq
RPtdiOLmQZtD4mXaTQHsSozir/qSZQ8yJR0RtXkzvyIe63hAvUFGBl6iuo81qJZ8
xzYSYh+zobkibK2W78+cgIuMTkGjwjEiNfIrAGCJIuYjNCWSkW4B/s2szdt6Ulat
Q0jaUQlDkdd5HlxYWBQhiDZvERI9TZpNIKyzPU6j39aywtbU9L7pFT+BrQgUVK58
qhkU+NdDhTyOviCwbUjF9ESWXD7qZV1TQhE4EdQVX6g4NwAIUtVVfwYCJ3xYHiA8
IU2njnbHipKAvqNgy7Eks4tMKMtWcboGdelOWTzPpsFOf7o8OCglBw2ERMjHxo2D
sfjhvMf2HXIdPD5euo5QhuHjoaQK0GRwaHpDxZSRERcuFQs7Ik5HHar+w15Kej5W
aLbW4mzPHSlJehG3lIujyGv4cjuqo8dTwHpEFLt8+LtL/kIIm6OxrO5k5AHVBOjX
AtPsHMVBvupg05Ks1WuEG/vd6o3Avt5lv7OvEe+aggnlEtkp6+OVmAqvvW6U9yum
lQvNCy+QQfSaHYMWQAjD0CkPJLEanvU63SZdP1f7O0LkekdahBY+gahRZXgHY+uk
bRxPQP735NLbz5eONoRZ+0tXe8vdYr5GNcaXolhicPgyjPJf8JKBaqLq00fbZ4KN
yR4U3EElnC+J+BVHaVFbZKksMcj3zlyTxA+cwShRcVfTnm8IaGYknrCdcHtclFUm
pA+PH5ptk7Y4iTPe26WiW1bBlkPtjdfYv+xXlQtHUR3dRr02I3g8A+S59idRZoBT
hpe9PpWi7eSXBlQr9FSA4E1D70SanhTj6SgajLSD0hf7bMbeadb9LshzD+F6Zy6v
e9z3AqCXHpuBmBpyVfSsb0jgsTUz775Gkfxi4OYjwEKl8UrwDqztWaOZ7b3EXiZd
dVDM141cDtgB65lQWICgCOvjaVxk+vcvctnNRTrsHOp3Z3VxeX6XSaZh4VOSPXWG
IEV1dLGhyWyuRYkyOdkqMjNRjYniFQ9UeMoW2RzIo2sge8eiGsFtuLJgOKqGEhaO
Ijv/R6dm8+I0CsMrqmobdwRtjGjUfexYLhxM3ZeilCo9sOTrGdBRFNvED0Mo5QxK
Qh7rW2iZ12in/paoBrNU+Ys6Md5URy4tIx8tkgrcEITzNC5ooP5IEMGiJFTmVlxA
k5kZwIGaZe5kJKpBxDuGbglk4gMgFt/sPBR2GElprdMVqOwkvAiAqk02vRplybBh
I6bCkC0d5bogCtKb+2+SGQXbyoZaFSU5bMBFbvOMBMlizEyCOdHvTmDHBg1A0g9F
mJniDxASbNPNYNAqB3ymEiDxGcIibwbnJ1odgXvaQAqwZlX292gMe2ddWTbUEn0a
4BtZ3M3y5Q2haH7XixUY/xZUuwk9PtuGiPFBhp1NllLVWXlGtSGHoTRsbvai3Pzm
EzYYd/uI52QdhmUrb1PiQn9RPX0Hr+bD94pItsYMfEhkn+raFlUFk6rUo4klpOpI
KOfc9caU/MCIPAZvrM9T6QO67e9mxJPlFLHH6b0YfRwyZ/JESPG0i/vfenKT8CCP
fbJL6sRF0cApSA28/T08zdXjmxzUDNqmBqXS4gTKaNnDuJoM28IcsfotVzhVyPnT
bW62qxEW5OTSz4vEbozHC4JmAWeAKe2jNOplSO6si/rMeYzUQih/s344kox/a35v
UbXMcoanqktGcIfwh5EY+Ss0bcc3wslRvOiR2n0rmvouY+k0ugA4HQxR2rmMSNj6
CDDoslnoHgqK0RJDVYtkUf5wAkyk+RiJFfKfIgPGWGvEUGIEgbg8/z/MKe4UhPGZ
p94HRyZkb4psA9IjzOHKZ6f5CgaWs/AUVWXrhyk/QcXzy9KhFwRdi8fWOBqKbRJS
LPNuch8FU/KRGQ0DND0KfaFb4ZZC8loxUMNFe5GsA+ykrB4Rik9hbRf9aP02506i
8U1pSCweFpBRQMvDg9uv1MN3gTuNEI3At2M/hGowGLW74w1Jb7klslYMN5E2PW13
IYyG5fD8yPWdp6KH++pbh70xHUhtqwFurRqiYyWIiZV3SbvXdn8pkBOLf9PZTajp
vkjChHVdU31PXuI9eXPpD6PYF+Qft/wCkyWs+3kPkYWky4CRiwPoDEKurVOgTvQf
u3pzvREClKHc2QowJxcDiYRJQsjhkMJBGrrdCVo4oZgSinK4a2W6HxDODLgxlueg
a8/5wMaEObV9L1YvlFXnwtwlpwcgDrQ/Cb+oNHi4soxheKN35CkdVpyism0/OT0+
LeIGNGXk96ku9tpVrNfOAQPrXGBRlwl4cNkVvvVyPOztx0x4Gx6S1jWFUkbkiqZ9
VODkNlYTi5Pk1EHtPFmcZG+E2eq0ld8kmrDMfUIeCa6O+tDSDNC0PtavC5eiDL0H
3nqQlqh77aYOHyFykPZBAAlsCCS+EsHN13NZ08887EWpXoND8ldEQE/ZkEFW6Pj9
pelIh3OOZgAnmCkaAttpVgQYiDzvoUdgDs8r5nrcmihDFDh18n2ty0MENl3XR8uK
fHRahLYDVohLQW5olKDSIabcr7S50UowTW4rdINYg59LWsrl2BamoHUlLXP3zARJ
PAvKIWHUtUMEf/33ogZnN5Y+OMBuXEi6nGUagvhUtlX5OkmTHT7SzPSK1FQpiVtc
FEOEApSr1LezxvHmRdMDHhV9e3U2bwcSdwTLIqGq/oI1HH8b3onx+rFSHbjW7NWb
jFApeLQRa3FaesEDZVEAQXOdsnoYEYgbgDfSNkvMC0Kbrochrt94tn39yjZa/PZA
lSEEgfb4qsmrVyl3+PxHPfkg39siaI/FO/Pr6P4Mh7g2bviAyIWaBIfbDAtWuU76
6FdjaXVtOlFEgTRriFAS+ncUAUrR+nMrH84uuw+FCZpLW6dbSp+EXVKodUQI48HQ
OiqiFWoE/oVb0LX73cTlvZV9QYC/1h1DxSr28QHQ8e2XhgGTdPpKLAL4AfbWKSSB
soh48XpcA7wWks0j8+eYVuxBJ1cZHevhe3MjYSPNqaDbmIC8K34ke7gAe/nnVEZZ
43Pzf1533Ytn+Yzmf8x6iKGaJFqL2mW6741eoQEvuDVBnZxkCO3dl3zDsBCH7y2X
BBgUGfAXgAsE82IZvu4oTW3A9cwVKn8iZ9fvFFndikSTVVrlbxlNYJmAedkGBZOG
dZws4AhlAZQTmVeE7K4ogiwpm5DexVpX/ZUo70JVQ65aJBWfJtnckl8um8Wyk4bH
t+sDgN+2auSXdo3fGAIwnqQi3sgLcdzKcZkj++8x/QG6C5rQFPLNRbY65YKbDFK+
VdGOh+YZSUxe7Sx9dkxluObs+axMiX5OM2P6VXd+V2v5Ond3hJ+Je/IWXNrbtT7k
6R+kbLHSMcO4j2qu+02+Im7wtTW3mw1eGiOKp1gm3ZGRlqR7W+3wD3D1lVt5xQR+
jjL2lhWy4JNe+AggeDLF4mK7pGrCL8oRUZlaJUpEIH9XnpSo1X1Pik/EmTZafwNp
x74BFPmjxC8tAT89jQKVbgkXdhSCX9u01HMHHMOBLodXEGl06XRPt6hHpj9CO5nH
KtqPa5oPT6iKaBbRyJn5TwI1adgHZxIga8uwNYGPvZkMwPW/WIhBM6tuPpNH7r6B
Xqp6CemkLDsIPr/6Gkt32qBdOI8TH3Spw3tS3ckm/CLtmj1WwcMNFnzFrh8ka6zO
/g5VkTQSXOa1wn/GZKs93fVRRGZ9Nk8k067/L9S1ntN9nnRZtKM9mL4tOZuf5P3r
uLHYqSGXjZRXQFX4yqaELhSu/1hUEVv8oTQXRWmeRGvDXHUArOEBgzA55rD3hAJA
fzLwX17zg2NI1/7QdZB6uI8sJ3bDIBy4HkRYTGmnk/wuC/IRmMiyruBaFj5NoQ59
htSztT/czpCxrV7Ep4xVdWhz6wDQcAR/a9ZFK1DXHfaWTZDM+P5h73K+2O7XZGKm
taAxIqXH/W2U73npRkW9W9s0Pu6MuspMPe/hTQZ4GakGlU6pYs1fQThjriHt/nFF
/O87s+MbjDC8M6hVpNc+HXB0TIiViHIeYMzBGPlCZP5iiBwOUPxYpbnlcrU9q/mY
V6yxqmWjCF+4ciHbNT4P+TXGkmYYSx+uizFE/AwxR8ByF5605NGeHk1Q+Z3a169Z
2JoaWvREk/PPUE/JwEYurmKY2g1H6PpZGHa1xyfolaCdMg4CNRyNPrzey/zpxb+S
r0GBREzQlv5nhPk9oi/nyn2aMlqJXSN6wXvj+IVQW90eMDBBSJ6/TYVr+Q2l9Aa5
BswipaXUUri1UKuEOeZjvpsJuTM4ugAr9adrcNl81ISESfrOiIry9SsYpJbWGfwb
8u5FdHjcRK2+4VyJ6T4ZEJeCxzJghEbAQOczUD64zN3+6E1q+imfjdN9x5zwUONN
Ed5nULovmr2+dl9X1EK5lUOahCZAToLKeMgRG1/476NQ3HVK7c3HzPYuJ7Kq++G5
H7I5XiWiMfejYYMglyz0lkz/ZiArGjTuS9ATvtJrZTRyTzD6tK/l5prPEMFd0WUR
kSR7P8rgFwPZUma/aHFrBmyFKICs7C+8+3f847SuiXCZ9vQBCT/rFb6YiP6+s9ff
yrm3HeluF9F6Nw0jA6AyavYGsP7SaVsZw6WIA+9Cvf5SUjllZEOB5tRT1RCLi6Ff
aATbQEEsI3iirkoIny0lbBdpyrgHpj7gx38tHgeSAlU8ynpUQOF/SYeUF5eEujc1
X9RkqScVyF753HADf4ynHIzlt7lAfPFGfksiVz5mq7j1pesjiGtK2n7OgkenraF7
YQ0VV3c9n9+8vd3A8mtKSw8ofBz5TBYlaNQcALBkrHpuOaUv9ut7gvniFghyKPBm
8B7LHd5+FLAJWdYA+GP6uTmRMvITsrVKXyKLFPeaL7Z4FXJlgNhFyPsPRR8rygm9
rVfY1PGDJK3y1cLuydB63KZbD1nRucB9pdWdESFdh7ZkQpajpQknZaelAN70aWiB
QYPWwBKd+1ofCkV2tuUUsvuCOV5Ho4mE/rjsMtWziq4UosAnDw8NV1DyyAJcPvuq
OOMLm/pw76tVDL/WOiJfAK90GHzUZBrv4aAyFTY4G8/4+cL2vDhNCC88G1MNTbWz
YTJ04Kl9xXVH35hlkFFAOI/8FvrsYAk9quDQUPdK9o17QLk9u0bTnfGYE0usCd9h
yoqKsloX8sYSqHaoCqWgvX/fNFlHy5gpfMgOz/d80fiYPUD6rYiibz+r0HnlYO2s
RVw3tkFgdmxpPw2OhzlTglWvLDDx5HuG3LAeT/4nVueQc6aGoMlKyT3zqgDZZRK4
81osKfBIeHgR8mfrLXtcT+Rb92S16mEo54xQheE5hr6vZraEger3OnSsYK90F7N2
9QBg01vabAcFQpQCt5G3IUfEfueEFbpiwWzwUqIPfsCpCEXnEK5Qb0PJXyFxAc5/
jUa9ci64FLZEoVepd5fGLQSYXDFD/IgYqfIQn4zgoZVxvzTUQ5ciZZ8HM5ChnE2i
9+um9+y3bI/IYqnKNn4yMF+wmgy1i4OpVei4Wm+ZdB3VehlYqM81ESLroJbOfxOe
99PYAG88WT4W8IjlYiajiBiEic5Wu3koq8X2ncgKuHvTNWB5yHl+LUcG91nH8LKj
cBgBJBqVh66eZtYcN2XTS276EwuT/lBTynHluF6i2c6rWznOIfzy3/IXHbd1mhT2
hbOOKEBevfXTLqJ1AAHLxn/Q4m7VN/GTu353gcBu6qTGdzotD6kPgDke/jR2uaWk
lEquNFi6vi6Z537KS2gt6xpvbux6GzyRogpSxKzB6OmfTUnPbbgCk0ObZPOCp0Ou
Bmg9FO5vl2uYDz+7HOqK2mbgZm6Sfjnsb5qbpYM7TKXNoPbYK0OoSSP3Awzoyc1G
/mgDea76g+6mEI1b3FEbj28vcn9jz4os37kgtVfmM7PIZPxgJrXcvvH3JgASxu+O
tAa1CqC/GWDcESerYuHiyGFPvLgzETmg/0Ap7PnuWh/O2ijGzN5lV6WAJ3mYhFDh
MrJ8SYMQ2+41H3BfudkWilkzkQ1bKYfWrkFU0CrLzAACxEOdg37alCyaKcAfHzMZ
pz67adRYAKlHcbZiA7JAwpsYURxGYQAnnkmhWjM2Z1UERZwnSD2Weo3INksbJzmt
6k3F99NZ3ZXlOgD3bZURTzB1RQOiHm8se4paJ+r5dhCUJSmdzOiyxBX9V+3wS5dX
H3m3S5JY/slxHFFd56rO0et/w63vH/YGYSuyhLZ4feRX4HlA203l8ueDmSfWyy9/
Ofy7uiWwqy7TR7ABLunCvxZEne7ihHdCr1Zn7d3jTQ5lNaAbFuBisFiZhSdQgpPB
7d2OQp8sIG8IhuqUWhFpW7S24Vq04wzUqlPff8jIeR7ly42Ja6FrMx6dnSS85gxC
GkF4SQxHRgZHdFDzQNRzgfYqc1hqI/9/6KB0Q/UjHexlLryISOPEBK59jgESiWq0
tickFaJK8AAg5g65xzz0qm8HM9MwUY7gCfNV/JHQDTwPWPdY8DIeGTa0i9lLhgE9
fO0RMlRQNE4JnP9s94gw1Vf3NAOXU7+xP3nU2vvn+G6JADhbxNjkol5c7urmv/ud
d4CiEMhAwwc6qeN50hjEjoBeYTX6UqE4O28PUz7y47qkgU8YhQQ7eLJgIba+QWWJ
m/NVJr1jWlcA+qkE8KuMtuTjNv8z8SkEvmlFfKeKDM3U0HCZzsIyexGv4n6CDIxl
s503W3OL7BcdFJIpc1YD2tBnkpH98LldNnFDLnZAZoRVxloqrNLMbLJK8lvPYx++
PEbewrE6Ku0cDqsPO7PjUp5GTgtTmwyP1oDESp45bEW2Pr5p5Jzb5WXUtOEnSIds
WHyvwDXmUrPeSm8Mq3tmPQZ/1BLJwEafF4stmoTp+DgtN3giT21uOqcUxhm6RoZJ
eG9HBjEiODDlMUP33tzVfCtrQv8eNdgIxnBQFhJBLpiQbbpoq+OK240XpoWB5oyg
w1vmFTUfeL6Vla0fW5sAlDMFK7bPE2khg60cwg55AljBXs1KS8VOGxzaPj3rZWrM
Y+5lJpF/HIepyrdWcVjleNSWo5FfJluw7MdxkQzTbdbGJrQGUeXYGgDGtOEPJGnE
hwr801TKzXsrzC7KDiLeYOIpSGiA4rLO2bAp8BAwYv5P8J7u7+Zn0eG20zIf4jc+
Vbrge2rhWf10QxyB14jN0Co9yrqgxMTJiGjx6QdiO0cKnMv9ZU8KaN04oqltl8AK
o25/OAY6wue4D+HCkJY715h9WCb3H92WjVPQ6FXDvpFCIIAMV6ICkbSLwZHNxQEI
JXEUcPUlt6yjci4bpGaEqcGWf5BAVfB4/X1eG11UyPSSFAQGHmne8P/kGME9BmT7
+z/bbCtVU/PuF2x0g9qfbFKbd3oGnqXKULIKIvCYPdtd8NWRVxk1mCuojSN60G2w
Wp/nDfuJKd0GnCrhlhQLRG33d06nOb+kc2ljXXGG2zECqubaQcldxA403B8SnoBP
v4DqcnHx3B6IYmBHLrumsdbLiNv4XSCduuJx+j1+Ts9TLmr/i+Ygu0vIVR3jlLxT
5w+bli86tSncixP9snE4rAXh043gb3l9QEQygT7BppxYntYnZ9XE3/4Dhf4U3hwj
3J780/pl3IA6WcpQhFldjiVz/2YZJR8/noYVRdUN29+tIzldcIb27pbuHNBvhs/+
9V9ACrlc/FieHtTlqEFEEIlnuzTlItl2HJeezEDIjcUKEc6gYOhkVfD+SXCQ2YP9
GNxnIcNbXvNxfe4Cd1GA8jFovRQ3lmmLbmcTWZ9vNHQCncD0U0vfEjqNqYqcVjhX
UodI/V0+UlJZu/qKJvHVpo49vb80WG3ZTObglqgcq6ZDB5vtIqDi7XMlnodUlvjI
n7KfzqK5/pWQ1ETK+EL7X2g8QXOXVF2dQ8UV1Ry8N8OA/4vb4imUqVNSJGIG+sha
4ggoRLnPwQ1xCj8zes6KsrGcKqtXkOOVIP4SWJByL+6Ua2iRw7mPlJqAoLuDp61Y
1jXTuHAhNZ3HlNKAXjjiR1mBl3ldPuiLHt5IoKExNy9dKfVaaMVm3Td4TJlhdTSC
YroFygRB1G3/PxiRDLO7dCftqi3USKZBOSXCFsHX3MH3jm5G416shDS6LL+9QnbE
ElvhlEfO+QjA/L2EiQ4fzyC1XO1dEWG3P94a7k9fA2Tmotr02FYZTCYIkd2ynws4
6CTpkzDBRa5bbY5GmZNPGkzE65uc4/hL483d9IloIlUdiyNy6LU8kKtOyNjUv4RE
6KBEyY83lKnSuG9YOtrjhebwlZEV/HHDjKu8eKCh4H8nY2jEa4qDUePhwEvcHpak
B9DufUbsuOywQWBliEFJK3/prP/scodBpzGAxibG3yt32H50i6oJhvX5pzXycotq
5l3K31RUS8x3vSpDYRdikwJFgCGzq/ZsTRGuVXf0sRh2aeEwSgpvZCNRSV5czS5/
CoRNpqMfoiEWf9R5tU3AeAmmr+Wlhsc3NW05pIvjt8NclNsrj5KcqlCo9NRp3/1d
CNFaqSZVfWRRQ1IAWsAeiyhVKxpuonJJVamcRLm798ZM4YjTKgiQgspYnFe5C7MV
7rWNq7eKPwPVgf6O2HU3DKagYUQmgETojv1+bX1o47P8fKKhVrw/vyaGqH/88AJb
AIscKRCwKX+LR1/kOn70lNl5iafBA+L7kz6yZpQyBs8s8D3uLoe7cMVpcGervQJM
uf2X+QG9iMUQyjTxeRACur7KNGANsgRKmBJC/ATKv/GLo3GN3VE8eN4gUDLSk30r
7IyIo0KILaCfAqssfXQUxgOZOnSfBpwDVkepJGGlMpnroDefBkBla4eGsAGnPbDX
67pkD4oTsjuw+PiDq1scUKJWET560r2KcMHs/FCOuun3lOMH7xKQBX5p2YAqa1Ql
I3BVHKlLMu3BZhMM3QkyDfBks/IlA+ItVrTKXADngh3pumFE96fZad0I8sOWm3l4
Ti0KbxThEXxJHwS2b/A0ChLLShsP4IIzcaH1O0r+TrJdjkS+R48PGWzaK6IXeB2Y
YnIAr4u0KmfniLSQrsg9uMuOTQBnPbzSzxddogCm+7hPZldKWFz1ZRezOGbNy8/c
IVEjqmIBRhiqXR50S+XLmAM+aY2x3xaAEdhDHg73uu9py7b0XvFKEVYJGYYHSEx4
2RkPRFhkfD3injHnPoCgjc9wHGBxla3+E2+wp642yXHzycDDQFGi5C7ujXMQh8pj
4nPf/wpG7GZe+XbC3m8QcIK+oz+0fJxRDzqdrxagBcgsim3d4nqPvy2wNgygynC1
I93yifGIGuUl3ZrkzEtW0lReEPyHRKdp3gr7FzPK2bYr9VPCxZfNeoz7LAWK4Jq4
1v7t5j8S6Ac/mYCqMSXGi9bMv/BirYdMtANMiR4RtwPivXwxxlJ1zlBA+zZRRaeG
GM/n4ccsNV32QrKAin7tbuCGf3okH47M3nTR5poi7I3aPdDRW38UJJlEokHU9OwT
EyD0xkOLsP3kDLE8TdGZFeZRY2ezOWw6t0g1NOW6XZAgoMZx7yRL9sM2PZZGTOBN
J/fc8JaZD3W2cxepyOsKA1zj6/9Yw1F9EOpOaxmZgHzKAPf+ITx+oKxVr69CbbRg
na+cRWzN5a5q/ub2XJXWys9kENVoLMYsCOidz5UGuXC42xzLok8Je6fJxo8b5q39
h24iZad6g3QEP1Mq7+9jZmX/+PwdY2/0iJL8BRzADeEujiICC1i7E6JTZoVcdZcs
Y5vRweWriNrnBKybuj6/1qC+2S4BWFz5H8K5qDUYodI37jc6lfm+bPFcKTKzudqW
7eA8ZDFpkv/HkL5wIVLntckvFn5xWJ/XM0AylS6s6ZHmlCSwvLRiyIZ4v3evM1fD
VzgMU5rMNl5DbVWd5CIlsOFD6xKTQcNBC28+khkwciXkDY+AJli9FcR3/qrlyifh
cAXovrxlybusfGwlmdEnFE6rMJzONzWaPpriGEhlIdAVpg4OrF4ESauyjWCmssHx
wzsZQXrDdX7BYFBbXIgduYmcfqgDfcodWUus2QHGCI2qeJkVl9FlptfLUBrgH/Ct
tGkLvjaRiuDQWCoG6uyuKmJsztKrgiK/oUpv5CN62xzPes/I8FoPBwoZoefgcLjT
mqUQ7aKpDQq64UoZspxoD5NaUP26dZTWgXwQcDR+6jH6o6RGcjdmpiGPl/w39y2V
FGDoDUONWbCOpp7eKsYXWR5aSuAXa8FfgT5ONoQ9iBr/ITkiXYg/3JhscnZuoowb
wPtCmma5fsl0PqjfgFasakpBnkOftkiRIQV1TC5QPZ3T7AtWO6XM/U4re8kEG/77
VLfZq6IDZCXyLm9GVV+ZozYKHbotNlKWsiItTObDzTvJKPBYp284y2bnefC/PdrC
g62R3Rnr5iIPstKDJtjJ+M/mWZYpJ8NP+MdbTcUmMqItK9madcdXA5xLW5jL4DpV
tX4o59txEi9M7iycXnZeTQg7934nEK54LU7ePD7/mhACv36oAA8ZRx3+vaTzhpKc
JRVfx8C8UrwBh6MlNT0usd3EJImd3TqIOJ+JXFUqjoadEYBnUSLm0+K3mk9n1SDD
Z3hbn63f5r2pvGkTOD9HWtr5bT9+5RyzfblL8oV1jGgXS6gZdF/GIx/rKNvdrytv
6qKpQb1Hau9FAT9t8Oa11PdOgFRYTDbKQtw1+2gfMKRuY2xJrSx5lb/SFsrXQtpv
wR47x8Is34qg3ZfX6Ufe+EfktDHIv5zYC2eH6wScXJTl6y9/B7G+d4EorJnkfKDy
IGX1jWuP9xFiC2XNP4c7hv8nfa+s1hDhtu1TywU+ZHmWL6e/LccvoWIksTwn2jzd
fcxvIjnbEhe1LNqmHPw5/NlSZi40mVAwX9ktnaYmgmOr3yLsEdFvC6wPKCCZlJ9J
IQohwgOskDoZ1bSe+6p4q3aint1xEM0j9OiynFestlcKMm5nFfkAf4Joih18zFZE
YqLJfVwsALfroMO5G8T94W7qGdo3t5h8RrjfuvU2KsVWjOlm5eKqwo7bskPqNYjA
mm6k6ezCc5eIvJinxMv0PCW1zb6ixrhBCLIiZVHfIj3KWARKJLLPCdpwp0KhZF6l
TGIc8I4q83RJV0Aq8vxhDTxFsLtZLu/lYuRjXJ/35puzsnYdOHSflSDd6mZZVqm4
pEH+1tGVuyX7VZw05xiGjvgqsOCHVbdyTZxL8xe4bSK9OnArqSoy5SNi2izkh1vG
b802LKqrJxGOZpIw76ItRPXDJbQn1qkUx7Up7IB+3MYVHf4/P3ndjVtaG+DE3O6l
R73Rzs1WLdkYS0DeHw8JmHmWX06ZoWt/wVuXxvV2xsctBK/2uXga2flYmGrYhGwG
G1M5sDQtJ0CMYRPianWpuzfGLXixFSwJQLk6Hxos9GJ+FejB7iKWDxRCH+0VwNRr
THFJQgXOhkKbhkfZYf0kjyDcFm+ORe7MsPDYEqp45fwS9yynNFSKv98jzJrKi20p
MoXtFUJm0642WKt9h5YpWOjkFLNfNngXPbaFRnH6ZOShPQ/3n1G/vgPuPg2FSid2
oPJboR2HZ9/kcpKoyr3wQfd3Y0/19Oa/k5pbvAd3D1Sjfts7BxW6YULVVrqsYAaM
EQ9CH/q3FTZqpkWm68BFHTERi+jQhTw7BpvwgfwojTC64jNC2aBAu0fM+v6frsVS
SVlmA8avHfc95zmuCSOj5apjhHZlSP3yLTI6lN11E9pheU4wmkf9e0hSTO4ebEz8
0udWzaDf8WfAu5Yh1oU7nJrq6HJCqBwgKLrhJN4p1SBjVk1CJd65z7dErDyHy3cQ
QoihKwEUdNpztVBHQh7Pro5YHOQBBLkcxJ8UONsOFErPlm+YKBNRghHx9nfwIQ4j
t8D/bUoHUE2jqOtc8s/AlT5QXDXr5ft8G7wOC9OAkqlwWNjPjkObhfPMvjvJm3Yq
9k2M2B4VWZUOKrMTUYpUEbxSE9JM9MTjC6eF+bnLZT18UlaqMwMZMsLmuPH9Vr7+
PygEk6ocxytbJtgWWd9gp1clnh/qjkZO2xzz9Jwql4nMYIMDxg1bcOMlfQzRRZXG
9LUEtNvy8cz1Uj+FBnfJUrXVFCy4M9BRDbwX/Ba6EtP9Re1S49/ZGaprmZEEPEgL
EN2QctVJ7fhX/RKj0Nt6e2xWZQfXrBa20G3JA1BaByqQaf4izebZSAY7yc6RaLkJ
YjVd8WT8uYnzBU5R+JN/EXgUHu+3qniHU6Fp2sODPNTyJdIOj09LBmQJpn/tj4B2
UDY0vTJqjTAqMyu8TnYSBDHgXQXa+wPks8PMNGfMtBsPa4iYtXfCppHOpwxDaxI2
qY4oOobslrisRP7AhsSXO13Br349NBOiEeCdWCjap0bYBDMhDmNVaMERq0ADXzgI
Rz/mjKpdjE7kzdvKtCV6PuhoC6SSLIDTbRhxaVL9pRvZtHaVtxKMvi3qTknor1Q9
mcnnIl1RLprGKceOfqgLP1oMpDeMuD/jTz9Sb0HTFkp45PMHgpouhidWVw5XUnkH
L9Xv43mbK8KFaEaa7BMIj5Rqpd2dSOiDMBYwhM4t6QSd0CeIWKLC7NFV27O37Dgf
67RZVVOQG115UjKnjhXl+k6jXWNtZcftwGHSgGYzjSyvY7f+/q1wCokVtyD13kcx
xTINKysoRF2+Lcs8ULutl/5+bM2GkZk0lHlxAQ1heTQv/48FOBBre2k0rLjjNrgP
U9M+D0HLkXfUEX+/NKG+JgyhSFnItnK9N+4XvsPkcMSdn1DvV2PbVG9JO1iPDr38
jP/weM6GQTMkJm/6kB+3UcI+SgCouwATJyk0QWgp0cgcsMjV83Wkn2MHtOzMuLlb
aoh6bYwafh3lY7cZ8pKJEB+sbo4Ohr2AkbyCWxf+ndiWChQsYN6eZdhz5OVCNXGW
lXuYySOB6jFXlujouVbYN5AqoPDk4xRD6beGThgvehgerhzg3oXoQ03LQrxxNwiO
cqJDuLtOXJH9t8FQ3k1IgOPPp5uuiSV1iVlTGNZ2G0E2eYsMTsyaambg09D/C5al
6vdETz+sTXobAHmyw3EiqORi2A7ufgilMC2KAJPAeYWKq1fNNkNIU6tABlj+HX32
KfxocuxgZg5NOsI1hZNbMIMkmrvTrr3SniR3oCA+/mA8edcGR/WXLuh2BhbtKjvk
ykKGeLTyqxNsTGpid1zXxNeLKN2Hy420ihXqeOZKC76oKfks+XNwuEhIDuI/LBcH
mrGRuBMI8MBO+9P1rX+TsL7Hs+ewTOPxJFPSEwnq4+4GhtXxskJdAX0mwvENvq3w
nEtuOimgHNhBaaB+0xOZ5UX6AK8yjK1RD+jgXUFoES4qYlLNmnMndKnH3kZ+DPC+
PxHDKpPgOgNu81pEaSkVctL296Yr6TBol0FU22x6WNqIq7lJ8Tr1R7na4kyHwh/Q
bYp4xoaOVLthOqP3nmxRGSu8HWbrGw0WyZyAgFp5VaQxfZvpg+wHUAATnBYhw0iQ
RxElfXjXg169YNqy1LpcVCUJNN5BDBoxsywIpmn6zB+SqBrbi34RSBM4ZZgbdtHf
ZjOWdlXxP+pHKwHr80OBKUIveL0Aem4uqcVbVee2czmWnT1TEFSq398SPtwP7L/D
acUhqtvEgfAD0auGK4xj31Fj93TBUZFk9m7+2KUZh7kDSC04qXF1mQkBcCu0ARLW
yPl/F2D78We85Pu9reveWYFsWQ1HTk4zqkR8Ge4wANqRR0rrSKLKDS+HuGIQZ1jF
Xa+pUIOksjMMsG154Aaqrlox6knxj3vZrzgQwUCBCtXln9cISsZY3WDsir+gg3QY
7ef+k3GjK5CyQmScOYBBRqrSlFxyBYJYI884H9rPaf8aF+ewMmAip2bfQX3BTkGu
YkAm18RYMWqO5eN1ekSdlddUPcDLc1/xqJvXSs3qbg5DQOuTL2sKT/HyTp2SzPA3
3ZSA9nMbbHNKysQQ3BDa43aUPHSAz9yPjnmnBGYroDWCKUQX/l+ktR9hijo/4ViX
kNfH+PbGSEwgo43rJBG8VLdZi/04iJ96zVBZYHdUj4mRvzmYrQZylFRISvEkRUyZ
dRVPn1t5O5gCFh9UXeIa0lGlMRzXPUUXBO51YMR4IzoEXdteS63Tq+9Kb9b6Oa1G
drg/ZR51fL3YwPTFXFADfu/QxTAtICIL6KJWdNyffeMMNwUJg/0WEngFuE9GFJ85
HZnusXh680DDN4OhdDEDh9BdY6c/PhuHh0bN+c3mX5wYMCvpduWsEKiMZc+pljH0
PUvDLvggELj0OjaIAdzidL29txn5A0kudKudYyfpfJMFZfGIiDEs6xCuCGouFoWc
Btye2Pe8cjojl3F1UYHmIsjneUAk3ii+gqNMhQhH/S5dBVBpI7XuSf1qd/EUTFBO
gLiymf+vabIjJLE4aglaRLiirpPTE+EjWw/LqitmSqGvu6YhNYutPu0XkaOBmOdq
UCj2VDnA94vEl86ab85xhgKoj4ZAhKTGE2aXp5tWcDbwoiSixJzpqSK1hHVkaxGk
M4Rbe93IOLnLdeSaoP9vk4ZmqSlIZWMzmPSXL9A5fQzllTn3Up0Rmf2W3DryCb6D
DiOCgdpEacey97bG+W+LKVHpqO1omN862J4S/y1oDUFiyrCQ14ev57r6Q47Gn8QA
fjHwSsGsnRIw0adDrFGBMP6Xo/p0OLR0coOQoYKZBfH5N1T0S4Wpn2T/ySyFuQZN
Ym/zhFGP2xgrKU2MCWKkI5e/tIIkYnmUTIzTRwSYXPA29yc2m6VD1SGTlbeX2hAd
u6MFUAqFNbsupIqxUJYuJMOA6pmELQ2M2y1R1/GyQGEOPrB7IpyLF7hCQg7/kiz5
piOXELxbQ9/deBojMhasZhysNsxYAPZZ4lcwTbWulvvleHcxXQDDUkYmiGswtz0y
+3kGzorpjgA6p9lEZdTfknRl7mG9gEJduqcvHYcLooPjuCQgJ1gbLmV1DoBzecZ+
/oPF2Gom0rRtEC6Vq2LY2fyDMaIDcLBjvU32DeKmQG93535CWKWD3HpWE9hDr4cF
DhIaeKWHF6vMCX5Kh/kbJd5K/IFNUq1Hdq58Ixhwd9kZ6JovqvVha4T2yK486Qd4
ZPDfy2fuJXxRDhTf/Vsbw+lTVLgbyHo7gxHOhVBf8fCLlY8OSOaF9n3vAgZCW9HF
762LyQ7oCImtz78iGI3u6va2m9BItZcLr0kAwmAIM4Xcpdn6gctYLvqJZ4wPT8X4
c6Js0tYgpXiyvFVlgasgJNy1D2o4usRtWe9F1eEV2tzsbKvc52XYLwxtH0YbWsvt
sKQvaZFy2TaJtd2U67dDbMrjSQXFDlN708enqLyQwLllT6S07UiQJIM81g/t4gfb
R/ERAoPU7QJEA9dOp4FM3ZxjT+h1i44VWU/TVIC4x7wiyK45rSYirJ5km45gQIzT
7hVreJi5SZAbxCq1GKcRtEwZoiqneutw7814i9Z0qc2+47/2n19yyoRrictTbqth
Alp2yUaTTR/Qss3cypGrBUfEbM4eaLpVxE0M3MnCSceR+cWZ6DYPq6CKQKXV37Sm
Ow5yLi8qoSgCYKpRF6KbyshdKVkByuiGK/YI0f/8A6EUYw3Jrtmm/PlRegX51Jdj
+aRe9CQnRt3WUnZKFOx7JB73oXc1YeXgIGAVftheD+F3p/4cxiUXoNkk2p7J7OAW
6lwPWP07kog0HtB8YmCMVw2YWZi/H/10NFVwBInziWc5dw0Wfpqvx1dyCA1vlDUW
hgL0o/bj+/v22/X2Dxl5v3vlPtZ310xRHRGu4yuia4T1QxI4zgnjevAFWsR3bNDL
G6d5DPTkyKzAYhb33gqT9+1gv2gVfKbd9G99rLW+mBC4b2/1Gz7truDhHAfDaSTn
kQDVGO1p1LXk1sDwnLllxcItOgLGxxbmmP/ziNlGaBJVeErgWYhiCRamAtqCARLQ
xKR0rUgY7kYsvwkEopUDSQ/BDJxdkfa4jrNAR9EcglorF0NtR0w4YtkWIdXWXZ8f
B6Mx8kgDGXo4xZth3X9qiTAQm4UP3GzS4EeRXAr7tIEPQboc2DuygQtUQl5ZhMOe
+gLpMfsDWsPLpI3DJeA6oJkbsBc0hJ2N+OB6OyapkEHtykC4vY8PQTx226qAvtPL
7bm4vwgKHAY0kMg+H3VnaFSTyhRdYkgXaNFE4SXx4AjF1LlZK8o/kEwBDLTKaWDr
qJ8C1muIdihVMKK7VrxceM6Nwy8O/P2wc3FKkvFoHZoMO2Yw7Fyce13XalpDZt4o
89YmKPbBY8Lb51fmY2/l8UD24W4BcKaKNlG84ObHwXjw/LoxB5oA46crIClXWXCX
mLztb40Z4PSj060kGiWMMNNXpD16ekpreRGOW+d/dLA1x97apo2GboyJFFOHFASV
L9gIghb54xqt2dnfRRH+P4kPjv4GiYdUsRq4opHaTBeVIPLzWOKP53Y79/aARS8R
Z2zaoF4SsMvXDxPxZaG08q/7AoX1Xp4MH0EIzm0kuxNhi08Q1luPjEu5hJVGL347
3umMj5camqfAUun1z7StKOJ0KfmXtVqUQMWXbicWQTsmixpLuVMvFuyDl5oFVc24
5jQ5eX5swWoNC9eAWaJT6+iHz0P2G3/CpwfEWCHEg1hQRwj0p1tFlQfl7SkcEwUd
FTxlrjxaayj9yYenUfb6tMeHEaXklN4PhDY0NYJLzTNkjLPWr0SfRTrgNRs1hkaq
WMABgvuvJzeuYlOt0eK1Y7uuwsXfBJj1Qxycq6QECvBTYAjabZU4l5ip3eosodfb
UynAg4m8+Gw0Rfr1pA70ZibF8M5GoBuV9iHjT3Faer+CqXspi8/MzmCmV6PMc8HI
xxA1rI6U+oexmMfQ2jw+aXTkGwDlhcLZzk11S913XXsf9mF4GpxIsZwcKuZF0rhJ
DIduRuSGlk//6/y9CaRD++feg4h3EC81B77OXAR81zdmpHziHDCKAJ6DKZvSMAjf
ZXM1KfgvgY3eqgJ6SYQC5lL4jrmjp+rsSFPi/y/k6SeQ1iZxcF5pk799g7HaROq4
R5F5WeJx9yoaksD1gKYKKG3wjMD2ysr5iXMuQyY6PedO32BXjE/aOr7SOUPoDQhw
5ed/hel1oBkHWkw3n2q0IQFcioT5oepxL1Yq/MWncYf6E1N9Vuazb8sIxJ7zSEyt
whcWKbC2zAi7PT5AeoB0Sv4zpq364xcC3URLqoiFyFB9bxTuMnbCzuZvFgtEmPo/
in0zSQu8TLAgBmfIso8kw0AvYmfVVgg9ndBbTI7h9NecSYy1q2kQkozwNJfRVfYs
WduRh6NnnTZiJ9aDDs3SOKD5hc88nORseMtqvCoYKv7og/QGRGM9BqXko31RaGUP
QxMqxZjR+yGh39wHPEqAKWUAkZ6UQDGZ4F+kJJSBFzguDOiLNcNM0kiU1W4F/wHG
hbRZUWZ9CuP/wzu72KD1+YseupS2l70Z84FIwszsIWEtdXbORpKRNfrnwKZMMC23
`pragma protect end_protected
