��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���jl�7�x�֫����_��aoY��?#��#�r�m�"R^F�(hb=��pt$��e[5�v� ��n{L�x����o�x�+@wM�ca冐堏����D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ��q�I�`�c��A6�c���Ӵ0Z�w�A��ENG��%D��!y���G�&�B��)���U�<?�Kŗ�������^@�����pX:g����,�~\�a�B7&��ݣ�4�A��@Ɔv�OӘ�XG�(Em��N*�Ӏ���4�>��9d)���&�^ώ�td��6�?H^�jce�p�6��J��B\ч}W���C|vz�T,��[�-b��$z�~K��7�}QXS-���6�G���`V���-���]V�6]eIi�Yt��V6�����Oi'��9;;J�z�^�fl����B�|Cp��\>�ۯ@}��rSڃ_0;e�ո҂�l��j E!]׈׷J�CL��v�T���u�|=P*��dT�r�V5��?�N�c/6�!\������Ҋe���/�k�e"눺�S����.����f������פW�BB2�03$�D��ǯP�+NU�e����DB�3�YW�wʨ8!(юn.�������B�?_�x���$���� ��4���k����{����}L7�!y#�E���L`�DΏ�sα!rLn�������z��:�s��xn��>�<<e'��{�Ǚ�X�^ȼ����3,��i�0iJ��/t��q�|2������TX�4�#��X�Ф���1F�ҏ��D��{��w�ܽ��G����8rgVg���e�+��S�sۜ�̩�뮣��V��x�ڤ�>m��d~ɥP
�u�4�'��e7�6��k~^���Jo�?�kq킃��R��.�r�%�Ť�V���SA�N�8�=�D5&�����L�m�g�s:� e��/3��J}��Ķ>�ޛ~��j;�'�5��?���%���^�%���.".n��mc��ƪ�B��������+Oux����>���Ԧ�i��D��կ�d��C����.ݍ�7�;��� ��K�YX������xA!x����-�//8(��-9k�c����MK�eA	��D��M,�#7����S����v�sBU�b+,�I��8�q״aG�rEoR�����;}`�6��֜��p�E�5V9cf���܀>�K���' �w���|�)����+��2���ir�9� l"���]�H��1ҽ�-8�,ՙ۔��oso񁓠pw�X��N�����+�51�ԜZKݸ6Ԕ�_���>�娐D��b`���@�jr��!4I5>���C�h��G��\�R���\_�I�Oq:P��AJi��t @�\T>�T�z�2�t�c0ɣ��s
�������-�����쑒�e��Ռ#����Lg���n�χ��lW쬀�"��_Nܪ)ڼg�O�һASÆ������P��QF�Od�� �쨰`�뛅�X�5�c7�:�O!^���MO;B�����rv�?:��W~�7lRa��X���U-�8���[&'�_��ɢ��`	�v�s�i�<� �TQ��P��\�W�*RÓ-�2�!�YH��ݵ\BM���9]I��gR2�*Yf�3�։�C�c`�r��;���FHr/��-��j�Hx�>Y�ͤ�_�>K��q1�]?1�ƪ_��?v�"���<!|�����NL)a�r����yH�=�o�?.�l��cG���a-�p�6��me�q�u>(�Bc�BIi�g׻���.��^U��c��� ���8�ݏ+�y˶�jUn���+�t�ľ�y��?�)+`5���Fcv�+��j)���@ȋ�>�����6������bơ�	���S�7X[�������������-˝���3��{怜t*����m��^�ԙNi�J^�#=�\8�\�Y�'�pR��쉭<Wx�����1�J*YGԌ��ףkɿq_�ߝ�$x¸vYU���F��v��&�	w�}��i$��ӫy�U���H(���:���Kk��h�G��0q�����6'ýc
���C��6I���j)�
�l�����x�����Y�vٓ�$#��|X��eE�)�iV5��Z�3GK#��n�uI<��I��$�+9V�m�c���9����=X��(��Ք$D�K����	.D�����_ep�R-d�*�>h��AFmM���/�T�v�������r��B�,�rb^K_e�.㆘��SUE�"q��w$cn`��c�.�EA3Z,��p?f�h�Lt1�HY8}�%�|���P�rC�ޮt �+c^>��#�72��P�+~�.H����l*X�����J��D(������fUz@�Z��B��u@6�5�e��&d2ië��"�� *�d�.���n ����D[EX{`ΟTs/��IXܹ�|��r�����p�7����yT'9��h���5��䖅�Ԅ0>u�������A|�����HlTg��k�n��S�8�����������V��	��>N
8(B�vN�\��ia2���i��6���Kb�8NOq@�^i�?��ˇ��忼wkI�Zm.���k)�a�f�u��VP|o�J��Ӿ��i���I9�}��^����~�Bwq�G��,qy��C��G���1qiĖ��B�g������7-O��wl}e��>A؇xx�b~e��$΄HW���1G�r���k&�3&���;?�T��/�|��ޛ
�W��S���l8�_��~����k]:+u�]�=�@Y�5�ٚs ���ђ�ک_7>6[r~��V>J���nM�NH�*�Kȫ�bBQ�l��Ԅ!kwF�u�����˛-�Q2�"s��엥���'Zꫬ������V7^b�� �k��T���������+���6"P3�u�v.�����F*�P��,u�`�d�����4��*�x�
Ѥ�ɾ3捠���4*Q"��#\}�B����(:�	� ɢ_S�Z�	6S H��K��+�zEn
Ǣ{�={h헵�c8pATl6�Qd ;MN���R�k�(�(�'�A�J�Ps�p��*N�ⅨQγ�mo=hf�LM\q�w����X��/��w���Q�'�5x��	^z�Z��2m�g�46��˜�"��Y��F]�o$�Rb����֫���2A����������+ؾ�m��ݘ]P�u;�V��
��ɾ��axݐ]*[~��ٌ�r�g@��������X.���(�,��%�V��ڵ#�LǍ�'D�|��Z��̎6�E��[�:���a��[	���߾�w�p�	�?�:昖�K���l�R�C��U�ݭX�U"�"���9��)����e��^�oXN�	��W۾����Z�1�'F�<-��K"�*B�f������(%�'�g�p7�/���Z����(���KB���\x�KJ%��T�mK����@�bv;C���N �m�])ͦ���%����q�V)El�Ca-��FR!�b�@o��G�'�*�G[a4V���{�|�N^2I��g�:��Bx0m۔}�t�0����AOI,�z� �������4�*߁T',�������+��ď�����C�z�S���)�����ߞr~�I�i�s���d�L��.�K|��i�C���u�W�8�׸W,�������|Vks�bN�l�D� D�Ц���ɓ��Z37�L:>cYo��#Fy^x�3�N۝����8M��T�z�H]in��XT5��2 Sm��z�f�.|4���%j��`Ӥ��M�a���fl��৙�Z��Y��b��'?z[<}ZH9ģ�*��A]63`<�Zc_bU��0��]!u�~y��Tx�'C���F�W9̣�2����b-mp\g�'�.��W=��:��N��nA�/�y�F��E�
��ؠM�����z�X����j�Y8��b����l<<��c�R�j"Υ\���8��%WZ�hV����d�����l��F�M�	��}����#�N֝ǦplCT�~,��Xrp�b��b�����F�%��*G��b���i�����#\S��F��-�5��g�_�Q�2���3w�-�\<�C� g3v�����g1��A�Z���]�#���B13"�����"L���u'�PB����o/�S�xIq�@�^Kj�xC���pW>=�sDFj��:;�s�_u.V����S٠�c1��&+��/��u��M�	�?�Bwi?��Oĉ�0�pJ��ٓb���K��1�ѩ�蝧�4�re��b�kh��P�$���ł�o�d+��:<�o%�L#_�Ğy�ͻk'�7qM��{,1*�/�ۍp�Fc�ډ	O|]� �7;�d�Q��|�=���NP���^&�s�e�h^�x���Q
t 9Cu٤�}^X� `n����3�� z�����;ڎ%H��d|�?��;_ۆ�.F���B$��<9��S=sSg�X����>	WϬ��4d�c-��le�'!%jU����}�uCtc�|�Ux��]~��S��a�~Y ���pt�)���r��4�&���F��� `A.0�ĩ$¿4����)І7�J���C����λ��t�7Q�`C%.ڠ��Fxq^��t�p��V�E�i�'ۖ��|4�{�g�q�u����)�`E��>�p�<�T�L�,^��b���-���)O�t� ΄��:�������tZf��"ۃ�{u�(�x�/�	�{\�+�����I�f��T!��y��2ڀ�z'mЊ�(W��.��M�e�ⰊpZW}��׈W�P�k|����G�����3����n�.ϝ�P�� ]�0�]��u�.@���w��FI�7�eC|��}��zD.D/���A�I���Q�%_�՜	@1�W]�)OBs���'�	:���ݕ�O�o���ŀ7G#/t��y���d�)���Lx�I��U�"�5Ǔ����J.]�W�ʡ��Q��49�1pvz��'r��W�[ �+e��y7Z�M�cf�7���uc����53�f�I���%��b�_�Y`>;�H���h�� ��ɞ��0W[�ӡfv�]X�D���$�A{<z<�/$��x�+ފ�]a?�s����6��B�|vh&���6�I	�*v8�z�9+`j�a�]�k��]�'���UE�ȓ�U�Q Z���@ ��%��ӊ�E��0��Ic�l��(k�l<f˘U�84֏�"{���*p�����Un������G26?3Ɓ�:���5�t��2�MH@0&�R\֍�2�H��ko���q��nnF@C�����ve���&�u�Xy�A���ufA��A�Zl9���*(RFZ�N<���2����քnc��I�^���3��a����YX'�G�l��.��G�t����&xrw�2��=�N�W�Y>-Z��!x�D�4T�g��2s��C �X�9u�sbY�Q�t'%�b��	L�ms�C��S���v��H����ߚ�
FP{u�F�ܱ�2���db[�2�*������mwSvRqpi�W� O�US�$A��	�[���:�f�9D�oI�L�ʚ�Z�lo�^L�ӵ����aZ.��f��W#1�~P�i*_�g��*'\G��U��G�g�j���%��ZM4F?�Yxĳ����^���U�&C�t����xXꗯ����g���fϦ���]!���{�b� �����ҏ�ٳEq T9H�N�@�W���ঢ়5�9����ej�҂m]֗_�ǚ�D��FV!���̢7�����@��Y-�$Յ�6�Q�8Ic?7�mSn��bf4����oJ��fӂ'4�����P8���孬U������Ϗ�_ly�r9�y�Dboa�aQ{��}�'�3��!Rc�I$kѨ����e���ƿ�n�!6���N�V�<��=,M{'{-�H��N�����P��։4U��~��
��F�"�Y�ʣ` ]M����}�LWq�<�u{��f��˕ٿP��ȑ�����R?��5�89X�'5sC(�x����Y��h|��g�EZ�?���_�����5����]p�3���Q��D!gi��U���aE���8I��-̙�%������+��y bWlD�y�O���M�N|&8H�R_x�_v~���p��m���v�����C��v~"��#r?�c^1���N�N�l�l�җ���C���ohl����_�Ϣ�(�_"�(�1��O�,�$1���zA���ڰ"�N8���3>�8�]�u�4���a������t�V1i}�!`_4�q�u�՜�4)�{���� C$���O��|����$7Ọ$^�l3��.tX{�#G���k��2�E��Z{��)����p���/��Q���-=�Oأ��,rZ@������-��)�v7�}ee����i/��XM�3����U̻�z���?�B�n+On3Œ7���̊����;|�#e�7O��n׳�G'�u�uGw�5cd�������S;(A���ؑ��{j�~E��p5t$�Y�@���%��\�c��e�"�_J�����c^�PC����yo�2�E�P"(�����Ü�
���+���W�_��Ǡ�~Q������c)��E�A�n�[NyR�K�C�m�#�b�q�p��
f��;=��'S��!K�[��_����QA�_mk�Z!B��-�S���l]i��_la��t8O�˖�W�2�*��$`w��x�`%D���,9t�(6��B�V�t��h����6Y���z� �Z&�v��|��7�1�����]�(��9I��4_�� �@�e���3�ÅR6�ˡ7��̟��С���S��/`�l�Q�)a
~V���5��`0��`���" ���2u��O�u�	�_W���#��Wz���3�-��ǥ�j�	sw��_?f��Kv�:!��q�092���
��S8��"��'☹v3|m/�g���hDV�ZL�^D����p�n�uI��0}��Y�L�=��.yu�B�y��82|����"\����@���Ktx��$ҲӃ��m��'8����:}iO��"D�g2�����h'�Is[�p����w�P}�j����y�ͷY �T��/���eI-�D�pfI��8��.�O���`�UG�W��5Ӹ]����)�|A���.��s����wY�=��f�x4�6�l"f(<��qdW�q)Ta���ꃚ8\�p��n���[3� ��E,�Q֔'*�	$e�g�	�Ԛ/9�j
_�B}[��d�l�����`�dƧ��z�����2Q����G6Gp|��pe.U3�Q�
���T(_M�6��, a��D?؟�[d|�uZ���T�׷�H�:6@��s�ӴI���n��Xh8^8�3_�6Q��e��VT���m)��'⊵�&�E�g8mt�R��N�$��'�yϣj�����s��ے��R��8�|�ݟۑԼ�X�d��\��M��4�Q)��J�!��a`��ِ|���qR06SX�簣���?�>V���s��O�a����s7}�>���6�RR4,��E�Yhcj�N
�/�2@y�w.7Kx�1�(Y0Rv�I~� �F7w���7"���ހN�?'������gB�ם5'�8����)s�c^�;b�\5��gYUۤa+��a!�gW(&��<��6�=JP0�$�%x�LU`v�
"�c�-G�#��Vl����/ہ���͈ҋlzǦ���'�!���'��P$���.���thHm��c�Y��к��h�T�$��Y�),���UlF�ʌ���J�<69> ����_�W���BK�����@�^N'���,R{E
��Rua�Q����N�£���o9bU˔�/�PP��5|�z�?��N���N���z9O�y� ��'�����%�~y�t�w)F�g�&��nr��?�w6ʘ�B�۰��V6odZ�I?ۉZ�3Ns���-���u7���K^'QЌ��\��Ae��*��B �u�SY�F�V�L�YF'�=��q��@mr�v���1L���"Sw�С�6Ĩ�O�p��M�	 8�~%$I���4�D?��~{i�DX
=hxW�K-.=�A�Ʌ�^��f3EM��S���x�6��q���ml_\UG�Uh����	��l0\�jtE�p��|�m�g��D��2���|3|wϦ����Ɂ�Atʂ�iU���m���m�RtO��"�P籿ʯio���f��֧�YF�U��U� 5�TsƁ����X��k�#|�G_��]����)e�!;ژ��fqG������:�����rR7���Ƣ�+(a�/�30�]HR��LI���Y��J;�2�aP��AL̼p���,yj!HfS�8V��'������ex͵"�խ�����벃�ZSE�SS���+ �z�d�n�J3Q�qJ@��@y��;���z��B넱��B\o������ӿ�c����F/�B�>9���15O�2�W	��Ul�I�.��~����� �A��`[�Ѿ���f�tF�-��p��4&��<SnB2ۊϯ���P�k�G�2^8 ��&w`L_F\Qw�δ�y�r��In�i�^�P?�W�C"�Ҍ�I�%}�X�h�0Ӈ3#�b�'�Ģ
ÿa��3^���-��6V_�Y��AI���y9�(��HJ5��xa�4Ů�鳥��'����)�R�⩮E�A��l5�|.cG���K&sQ�����`j��%#~ 6lCo&8�dzީi��N3Ts���J��c��N��ȜZcb� +�®3o��K4DP�oZ� �V�����)�?+F�$.�=����2��)����˞�ݽ��OX��C<�7�������t`J6�	�&�1�3kG����7bK�����r���2W��	m��*<kw��� ��P�c;���p�.�U�lN�_�z�M���P����1�8�1��?�/@+�o��Ϗ��ףu����B���;�"�qfT8P#I��Qq�sM%�J���(<h�Hޓ��c����Z݉K�R}�S&e$�{?9�Qm��6 C�{h�+�+��z��������c���/|�Fv�#^��.��J>yww�a��-���}YۖU_ݫ�/��	蚀��{���g�՟F)�/*fJ�R��r���	�P�/��ztE����9��k>��;"0:c���AU�
������FP'8�!T3�w�B�To/�$ �g�j��3��8�s��Ol]�#�<�����r�����vi|������|U��;���q�� ;��!h�ݬ�T��M^(�����f�^J�31���a�\�r����T?塆6'��;�v����j@<���m��ˌH\_��p�|�d��6|G!ѓ=�o�+-;���l��ߑk-1A��V��iY�JH_`�ݨ�?]�5t�c��NH���oI�5���Q�k�4cn�(zG��Xr�\���D�G[.o��!�ʛ��h��[�_*�|���Sđc�k[̢.�-��m[�:�`��!����L����뱂Lt�>�N:F��E�;&�h������:�l�M�`����Nw��c�d
��20���y��S�tKY��~��s��	ϑ���qذU�2�NnSS��	�ŎU�WEA��Ԝ�z���S����	Kd� �UE��&���#��(�xj{����U�$�D�ğ#Rx,��K�8��󠦜ѫ���&oe�9&�?��d9;��x���q���f%�h?���0 �w�@8D���d�L|�q�ء����@g�Q ;���ܬ�
����Mg�#0I��L��1�M�!�� ��I⛾:V�9��d����C��{�<�m���rz�ϳ��R�?2� 'X�ΠmV�I�,]��w��0܉R�+&ҵ��-�냂�X��k|�Xa�@� r�Þ��l��/�m@8��T{�w���3���G���(��,=2d20����V�1�u��ˇ�0s�W+<�3x�9�bնE!��c�nCn˴���dH� Ŭ�IX 5�@RB��9}~:�qF����"JNꜘs02��yŪ�|�2r���z���GȚw�?"���5N�Ot �o�C�tA�$�)�����{��v�B�l�,��u;����E�3����5�u|mdl_��|c�j�WF\�ڮ�iaȢ�*}�8� ud�f�k���rq]&��rJ�'��t)�g"�&�KO6]V��2|����z��y�\�5JiMP��70"xPkT������&>��0�p%'�h��AJ"U횢���.�>q~%��W*{ʒR��[i��,K�+0�'žPv��M����XN�L������NO�pY^s^�Q�0wLyH��K���ȓ�0�����ɕ�d������p���c`@���e�ǩ�C�h��rUL��4�=��͗?�����c�3Y�X\��
�J�����қ>ݾl�G�4"�5*�4� ]bu�����pY�6V�v��� ����K]	0 ��\4���`�7�Z�2�:;�޲�j��Z�%���Ѻ�<�j-Lܪk�%#'����gie�+[���'��2�����m������"Q����*h�#N�>���ji1�5�y�Z���Qx�XD�4z.��Sb8��l��R�m��l���(ד���J.��E�S���6՝���g�46�[)o|��M��� L��`g� zq���ߣ�X䃰3V͑�?���a�4y��Ł:ʎ]4i+����Q��pM%���Y�z}B�#�
��9�\]���`�A�$g���r-<dv�lE�1�f@#�(�@}���W�����݃�h���_��k�a���g9�&`�jJmv5=�ᇊ���m����i��PVQ���щ��?E �E�U��N�3v��m`�n� ����؎׀�dޯT��V=+���3?�N�\��Ƿ|����хX�,8+P���	Z���4I[|�� ��K���!ji�1#o��*Ly�j��l9���/u�0ͭ��Uy��G����|Yj��,�@��x�>` >�b-���{���O���)��+���{�+�	�<F�A��|��I�<��;�5����6H�1lI�+o)j�}����C��C�US�~��	T�����vn�0�'4;��������Xd�uc'�.\�ݍ*�r�bo�1��z8�^8��D�L3mzy�4�]���H��������a]}����acӻ��/���8o����!o�
�y�M�~Q����(�7.�"��V� ���\�*����J���M��<M��w^�o�-Y�����9D��<��I������-���2�[3����׀�Y,�I�K�o�ķ�����c`����Tp�Mm�%��J����AO{��,����0���σ�7pL��J
N�,�ӪŲ��ioȁ�s�m���G�X���xbX6�an/ �|�L!���eݫ4`��Wnh�k��{q*jmѓ�~�6T=�����4�p܎�ka�U�M=O��
s:EGQ��s����6[N�mtB��U���Y�`~L�1��1���3��v���KT$I�sb�꠬,�c.�����O��\t����j
��C����}_� ���&�]I�;���&Ie}��ޏW٫{��`B�E�l�����W��(�/��õPӵ�閅��<}ʨS)�D��O��@/y.tIL"$�b��#}FB <���}7��Al�G�_mh	�Ġ�'ML�&���f<���BD���H�������g�¡Q��m�'��_x3)WPo�F���%�����	��t&> �z��RR$S��*��y��)Bʔ�]���,�J�;�1Sr.��:�ꭧ��
�9P��R�����t����zl	�J���26��������7q{�籿*^]�� �r�t �'^�o�
ʀ������nc/S&�"��k>����6��*���������<�����������2�C5�K<ʘ�b��:10.���5|�~�qѳx�i?�uuS�V���5��J�����;v���q����!Eʏ<�	�f؜�f4b0�bۚ
���@�dVU�OL3!�ǧ.�z��D���Ҡ�T�׸co��.��IϲC��/xA]q#2�!��!�E�t�N�����V�f""[�NF�&>W^R1&*||�#&�O�$*��
81KJ[=Ln�M�'/�r�����_D�2��b{<C�o�ngy٢)B�3�7���5nF�h\t�b`֮�Ѩ??�h�K�f���[ο ˕Z��̞9�5���vӑO��0u�K��36� Q�u���?1�Ѻ��o����eLB8X$�Jf$'b'o��0 �U׽pQ��`�7\��P��>sI�$�|����u��=�����_$�}'��!���A:@d�$[�f�e�|+v���]�3�� ɔdk�{��7C_�G^Ex������S6E���߽Y�eX	���ٲ�:��ă��'�ܝ��Fph�`:}{q$�M�5]=䋶Ժ^xώ��!hݳTs��{n�#ߊX�ц����L��>�o۫xߔv�b}�O�E{��]g�#"�~!�^4R���R:B��������m����>�?M�>��E\�)��y�Yz����y�-��i"�1%L��ܛ�ݩM�}��p�94+S��ՠ �^x��v�!C�2�@9z��I�}g��i.,ĉ¡I�d��Q�S�I	Rt��Đ);���9��6��|?���c���ĖQ�C�
}cvV=�Usu�;TLO�^���!p�
��$R�f��׺�6�.���K�*�3�T�"��׆G�R����@���A�U��+5����\�m(;ܯE�6���� ��������u"_C��.Ӟ~ʺ��Ը��<�'�ac�@���8"�l����4�ȼ�����Xb��f?V�G��hF�ڃA��s����N�Gh!�P�v����ki�&Hh�۰(�O[��g�.a��1;��] �ք��g7��mwZ�p	M���/�$S��(�lp�sF���̐d� !=�����LE�w��)�Aө�q�Y]�	8�vef{�,���&�����uP+-��Z��T���kRm,t��i@ ���-��T��ݮy ���sVY�Jz�b+�%�g��OPdb��j02�n;�fcF����e�F�~��q*2���t�^������]q��c׺�^E^X����(e��j��߮8Ⱥ����S�T���ӇE�3S�w���~W�h�xZ �O��� �����y �S?���!4G j�G�P�����Z(��i�ƳG4,�0?�iPF%�R�;^�f�l��
�����L=��ae��#k5�l'TΧ۩�(��6/H�K����lt�XF`�>ʾ�o���Z�2�d$��5��X���%W�X�JK�r/^kY,Z� �x��c]�.��{��;�^*�	[������0��u5��(i��F.�]�0Q��'
 ����D��QOi_P���<x�"y
-p�A6��F	��@��*t��#�5�6OP��>����s�g�L�i�W��u�&�|� ��x�Υ_�X��4��Z�QF\ڜ�<�^H���bę)6���l�)�G�c��u��iG�Dr	fLUI�	rQ�@��C��خ�%���M4/�25��/N�W����6+�/��נ��T����-s��`?�B���֐4(6�r�j�g��7ezn7LJ%0��/=��áEé�ڐ?�i����j!=@V���X���⾿��e��Dv�T�V��)A}�Ej荥�����j܅>�1T6���o/�`����L��D��?��y�m(�Z�T�[7݄�����d0��;z����t=��o��� "L
�&֜'�9V�<��g���x�� H22���p������q����QS�~*�I	�>���>Mgni��m������w�Q�xN��b����Ob}��ɫ��入N�:����
J�/82. O�(A��C�.�F�h�tߏ.�[���q.<�߽���w�;;�y���fn��ɝ�,,��Z�v�����k��	E]jSK�^(na}�r��) <���Jt��?@@ ����� Ჹ\�6�S�f8#~ȴ:Z��"Ue���t*>��G��>���Ȼ��XA���k�TJ���w�{%S��\�X��S���5�ܕk|�_k�͜�&����-.`��7�����Nl�ErJ6i��~� 	�R1]]�>P�h������SF8�԰"l�X�
o2w�ʭ�Q"e/�J9V3]�9�QE=��H���K�n�Q��^a��I�v���@�^��a���l��m~p=�d�IB	��S��;����RS�,���Ӌ�ӡ�ӈ��sRp�P��!��l�ӛ�-v��=H�~N�{E���y��'���GԾ�b$���K)�OTX�$�06��g�+� �醽iT�9��'�k�r� *N` *	���_o�2�/ �NH~K�RHm��$��F1Z����}�T�jm�n��;�I~z����'���r��U���
=�U���N��I�J#<�QKJj:�᝿�T��k�"�m��<ZpV�i�g.hd���i髜QRP�_�{"�j9��l֕�e!0� R�B++W�'|ߎ�������rGі?�y� �qd�a���`|���C3���G���IC+���ߵ^k�yP ���
�0��f/-��~�'�(�+T�$S���$����7@��������qҲ�-3w�_=~�R�#�jqD���7�@���9j�.�-�!P&���6n9�8lshaI�{��g|L���$�5r$e�z�U�JWi���ϥ-�?� �t�B+�#+�%@, ���H�4'}|8j���=H�Ջ�ƄQ�WV˷В��q������g��Н-��h�W���(��5�"؉ף����)'D:g�&[��;Ɛ���W匱�����O+l#x|4�s�nχK���d���;T^�2g>�ߍ����z�����^�d�)�9,��/ڂIo������4�܊�@�~Et���80��Ӽ��%����o[#>���jң�	�hZ�j%�X)h>,�c�p����U:�C�6I��j��1YG�L�k�5	^U]Z���BCx���q�:�h��JN!8�V���e઀����/lӒ*+�4/h��5�VV�s}X��6L*��Q�5������b��4��J�n�m�U)���
���bA}[� ��t,������X�0��� ���\	t�óQg�kQ׆�DJ]f��Ճ�=�S	:p�ٓ���ʗL"}�}���n�+��k^/9-~�o�&op�M@%���v��3NO�<nU��j��)�:��1��Y��q�8:�uv�)��)�X7�1p�F۟�!�]U�~e4j�wn�o���+x#9�,hԹ�b���s�Cg7����B�h��1<���da��,E�ؿy�7\VnG����#$�p�bۭ6���v��o߁0�r�u-F��j�V���/�c�1;�!U�ϳ��~
�r.57)Bd:���K�D��L{���kY�R�t�ΥI���u��No ��-ܝ]H�Ck�n[R,���s�� �6�S�U��dڱʰ#�����n}��qߊ�?�D�Gw?��-�5��+�ܗS����2��V��<��د��L�`���k/F�`r�?��b����̾�-$��dm�yY��!���Cq����y I~%ծP����M.�a���ehjE�E�����m�c�����|ej�	JD�e�Y�Ԟ�� ��:���܌��s�����1wݑqx��ѱr�A��"�y��N/�R���bvI�+�Z��������y9��� �ڷ�I�r�ԕT~��are���m�sY1Z^��Ԭ=��e���
�u���Q��8}����d!�O>_�1;kW�� *������c�����@�>��b�.�o����1۠F�g�w��.��o��`�b��Ķ�AF�� G#z�w�H�sI�E��w����6�
V7��<� �Q]�h`n�k��c8A�{p�*+���8HT���y�T���m�bj`Au�<]���R�k�\��,l�~��h�j���_�7��U�H44�=�1(V۷Y1�Z0�^s9�(�
C�:I��{��݇ߺ�I�Fn�i����� �5p,��ȴo�ۄ�܂�&*~��/�G�/˹2u���V��ś�P����ܴK����O��T��MɌƐ�R!�	!�~��x�ؚ8"�1��/C兂��#�3P�s��uhZ�W�-oH���W�)�m�%����o@x/hf@Y��}g�;B]��h�Tb��E�O!�Y�'��%�b5��?�����ee@��N� ���E�OZ6�`��<��#M���������Py��nn���ض٪V/�䪥'#%E��S�~l�K�<�$��Tŝ��-�1i;hD�f-{~_�d�S�7q�"sX<���(`oFO��`��v�<�{1W��`�F1�\v��	1D�����h�pY�[�{m�L�����e��H���<�t�� ����ܗ��ˌ���i�P�o�T�7�K�,܉�`��Z��oo�n�W2Fx�H` �J��F�7]���G�'5�zO�����Uy�PׁyG:�	��}��o]!H]�?�!H'�|�Lzw=���� �R���g�U���x��2FPZ��	Ǹ���g���Ȣo�0c�`奄h�Op��|5�H%��Xl��3`�ɛT��BA� ��6	6MQ�-�p��7o�Q�M�}�>A������_u���<�h�]�[[�(����X�I8A��a�}�^�j	/��V�D����#�ʌƥΰr�_�+sjw�pX�nY�5�f�8�x~�AOO'�6��Y
�4_��Ԣ�~Mg��8]��鸹���9_�V�c�፧����.�)E��U��1�/ME�V�5 ��ь���CZ���z���	V�z�Ԟn��_O+�+Xo͘#T���,����iۖ�3�I��������>�1c�)�wѝp��d�@#���W(���UAaߋ�*��ecq2��8 0G�y5b9�3x�_-��aNa��o��n��� JX��$�?�JɉR?!�iD������^�X���}!��Q���V���RS��j�ֹB3 ���/�N/��q32��Pr����ߗ8�l���SVWd����[5
N���nN����I�v
<w����7"J�H"��A ���h�����?ߙ�\Oepn}��5 pRHO�ŕڠߺ�
Ǜ)GX�d��-�_���f���"a�xS�P�E��{Vщ��XK;q�%��y�M&�jl�e>�J���*qR�_y�$�q&�����j�M�#Q��pP����vA�����  �X�C%��Ex"9��<�k��H��=�Ms����F�B�2�� �k(���MT�c{�vM�C���[���2�ge��S�_'��~�Fsy6D	��۲�T<o��<��2�%�ϯ���bYi\���>ǜ���j�Աӕ�x�I�L�
�!+����)�
k��ʭ�TSVpE�^���O��M۱�N�����3:UL�����YP���P�e$��2�E�p��/���e/��@�XZ`���g�.��@{�wvfg��3�"�aa�q@�=�D2c� f)��Y�ÏKջJu��YYy*c����@0��E���s!&����_�I��"y��#�qVF̉n�a��"Lp謏���
}�Jt�hT��X��8/��2��-�����1ii�}_]�8hA����M�Ǫ-`��BU��\�B1��m�f����Sʌ��3���zѐ	�V���Lo��k*ߵ�|b�&����DT��2��D5q����3�h��Id"><���ll�{`��ؾ*ܨ[�h���*'�^$x���<������2���-28�%�~�^���k5Ǆ��y��r\��$І���_�yf3���8Ȇ��]9�H�����1�B��8�s2�9���t<�����Ӕ�ʿ5��P�i�ɼ��I�d�ȉ?�9�ó�hd��8�
��%��a��(�H�)��޵E��!����ۦc��N��� &��H�2�X�O�Z]N(0Z5�N�謒P�E?��o|��h�p`/�[p��36v��}��Y��\�@Q����@����� 7"P�1|q��4l�WMS��l�>?o��
�Q����
�!�GXQL��?W4�O��ԞF�,Bx������A��$�ʴ�oN ��g�#�nH�����'�2�Ϟ,���%�[�	����O%)���r�7��'���y��Nl�']؏q�˝
�DE��EV���
�G5�yXS��P����d�[|'ʓ郲is�Y��<���j��:ss�lm7O�����z:��Mtz|y�����:"6��Hߋz��{���'v,���2�eȡ�Yk��_ ���v�^���#.��Dy(��XwH� o��r��_W:TK�G�y�A��IAh�rx�`o�v���U�də����b�g���p#f��gW�<���U��
����� �s�٫�e](�=WՏ�ק2��F��F��kabt�ty�dYsi�ݏv
����2��d��gpf��TIa��<;JZ�%_�Z��Q�$\*���t��}��珠m��V,�h��+Y�(� �� 8�D&�����ǘ�5�=m0fxP��Dh�V�2�,����Cw'/���sU V
�B���7d)-����r�Er_ìL�#ؽ!�!��5`�]��5��5#ݛj�1�@v����B�Iv�:��C~�`u4=�c�e������j�i�=����.(�M������l��2��QX����`'�@,�9�^���yy֚uGW���:v�٧4L
����`&�ކ� ��ׂm���n�P򯫧J��9|J�!����wjcZ�4���,�-u?�X�j"`3���M�Iǟ���=I���x��+4�ݺ���i��x�W�#�n� �B�A�ʢzf�<ώ�a\b��6C$1�\�g�F?w]��m�D��	aXXf1gG_G2	�N8|V�?D}l��a��T���R���S�*�
�S�Bh���֞����N��ǘVU^^���G[xՐ
����|I�y|O�f'-�,���{���SG���zX���5���o xx��%/�V�?˴֌*fJ˺O�y���I����7;.7ۣ�J��l������qO1V���f��A5��pN�1�myem�iǀ�n���M�H�����/����@Y��_�P�Ő7שw(�c:� �.�P�rgW���f��4.gն*�pQ�����/7���Ѫ�*z������:� ��܁Z�s�㔆�'�s	�C�ӊ�C�gE�Bq�IA�"47�)�"C�MӞߪk�7Ҡ@�J58����G��u
l-)ڕ����32�|>���'R�	��!g���ɫ�m�r���8���1,���k������K%���B���D�+��:���A�D6��1*�.��D|�m��?Z��ђ���,��Mى%�Tp|ٷ��<ŵ`�ؔ��
g�}d��h�ώ����BH���� �P_��D���yͽ"Jd�W	��hA�J ._��iS4�I˧�V��R����q�>��9���˽ZdE�D�����1;��u�����[Ñ$����H/}m�}�]�U*�Ir��[Y��~I߽�J���&/���q"�<:y��o�QD�D�#����}��oZ�w̐�++<�Ȩ�U6�4+He���93���]�j�'���o�S�k�̤�d�g�H�{�	>{(r
̈�5�ʆ� ��[��!k[{6�T%�l��ھ�X�wl"r�*#�@��Ǩ��Ps0A��nf��nt�9��,���f�d� ���fb�T?+6\��ub��Yp���Z#��+T�Gt��OUs�?*C~��j.�t-|�L�D�TH��/G���;(qއ���`6�G�BH�����3ۿUg���ԇ��w{�M�[�ׄ<��
��P~���/�R-�zv����JS?���B�T��`����: %&cf�L�����L�<���v��T3>4M~tjH��7��Bc�� A�Q��J=�x�z'mŽţ)tHl� Ľ;ޒ��T&�b!�������j�˓\�^zRF�,�����TP'I����YBc��V���I	�t�S�ͭ�'	\c(�'T����V�e�,}=������D��۩�mJ��0n��t�����yM�P)��B���J�7�R'ꪆemb~|Yw�i��f8}ǋdvxS���6����m�=�Y��I��@�8�=!&���MM��R�շ���SH0 �K}�v��FB�K���r��G����w�ɕ�U*����?���v�F� ,}�����Oj���țQ G�&���\�W<����"9���ܿ����
�/,�,�<ݘu������AU2˭�QP��p�������8�	�!c	�O½���*���J�E�k�&��2t�PU��׍�'��s�$��uQƤ��(�R�@ֺ�'�\_�H�7W�l8�yB��9(FQ+�n⣆��c����%��'�1q+���L-�l2�P�H&f��%����1d@�c�Y��"?��_D���ˊ]��-��������z���V~G�@�*%QJ�����
#Au���u)����S�3��L���{,8M8�  �U�V�Ϣ��4�>}�w��PW����2�{��M�b�P�J&�>~-�v��~z�Txx-ǝÆ�i.Zp?�h��sC?�\�΀Q��Jպ)�2�
��r襉!nJ�[���[���5*Q�rbO���&)�0؇g:��սr=Fҝ*��ȉ��� �C��ҙ#�,c��ٜ=���!��F~����: _F'�
@�`w�'�=��]�^B	J��vY��O�ht����cE���97V8���W�
rK&I�}��$z����w�>v���{m<=�����;��RU6�
�Ђ�W-i�a�o�]�jl�:�
\�Ϩ�.�׻�	��mZ�F�
���g�_���Z��}�oz�]�RSD�Y�J������5��Bb��-���-pd�%r������}�]�p���-��SI��3��d�ڀ�H�ٰ9_q���!�0�r;����:,K�=�=�+n���F���,P��`H`K$��q�d�nqZe�r�G�������ʃw�:{Hx3���ӷ�ok�P5O���U��F�M�P�-�	���|m@��>�)�ټ��e
E�������o�=ք':�@�bR�.�ԓǃY9k$p����F��i��C�\�ֈ�R�30A�)s����S��/�n���<IU^�ѽE��O�Z���'y�wfO�b^�D�SO	�CMDxB��{N\�A  �6�4m���Ҳ|W���L�����"\��9k.��� �/f�-¡�����4<�ѬF�r��+�>Ks��.p��uz�-�;x#�CzC9��4�����aϠ�,�CM�l�[+��P�X�.3¹�]�ݙ\�*	f�H������C	��TK�����h�ܕ���4IRc���ZתI�<���:���1��#���3a{�?���L�H��'�ȃO-X���3 �Z����Տl����:��K�� �t��a=��Ŕ�p(�;��ď��͡�1Q�$��Z��PJZ�Gi�p�o��}��pj�LzR����ߔ���asҸ���6����+�m��¦}�^,�fZxK����F�)~�$Q%������j��ǰ�g���J[dƴ���)�W�J�%�{�rљl��%�8�քd��O�����Qo(�LYʭ���٘]�"�2Zi�>Z�!_y>3��-�ۺ��[^��MM�%�ҔA�s��ǰM7��a�u�.<R�?K�SLdc��N{�$����_��Ac����0�&�$�sB�aB�Z@�(��߿����U�PD�j��ݯB�{`G5Sj8�Wtu�z�ࣷR������	~V�\���L�q� ���n�OK�cl�H`"�S��e��j�3�Q+���MTC�*�3L�Z����{�}���B\|���脳P��-{fh­q|��?o�eZ<��}�KFZ�(<�N�k]H�?x<�zu�!�Z�?ڍ:������f�\�
ۍ'0Mq��8a,BZx* Γ�˺ Mȓ����p'<Ϩ�Ձ��4���oK}�hĲV��f�_�� �EML������	�6C�-�[���5�b�z���P ����A�o%!J�w��E�qV��~���鸻�t���J���<�e��2x�A�n��>�>K{�][}C��ǯEk'�&В�Qa�q����H�ry�:�~�d���Ag�����L}˛[MƑsl��M�"B�4�,<�k�W��yL�d��3B�|-��&��z�gA3Qy�P���S��� QuK�$u[o�zq���ymh7k�R�WeSe^�O1�-9��*:)�Jtet[|�v̶g�U6S�XpwYD�^��H�1J�Q�R�0��r|��a�	��T�P�^=�,mb�<�䝈�(�����K/U�ͮHq��aDE������Og��jcbˢ[�f��ejg8������]��t��~���i���C�ҍ�hqIE��?�b����<�|	$�;��8����\����w隰ixA��(���	����wu��T�e�Yv���V� HUm�3V����&<KrZ� �7c܄ڿ��X8�M�F9�@�����ܙo��+���_|ib���C�0|*��WA���A>��ϙ���m��1�v�e�Bu��p��+VSP�^��g�]��k��}^�^��e�*n2�(d���\ù�=fu��Ģ%���vn׽�����!e��"sk&�Q��e�7Rp�l<��J���/r�I�<�;E�			�d0M�\�*H@Fl��iĵ�g}�����C▥�h��aS����
D�HClu����4� ��V��W(�oa��� M��
i-7)�|$�MC���
�w�ʳ�^�%ui��O��.;G�/�zg
��$�R>� LסQE���`��崇U�8I������ ���ݼ�i�
�U���;�4�3U@�Y<l��4|�H�����'rV�$>�f�\�:��qx���ܭ}�	ޓ���UA�rd�VR�<~����|����[�p8I�#�*y�G5x�*���1t�Y�m/πM�خs@JO��ka	,3�'��ρ�I�v`��72�P$�鳏�9�	*J�h����y�3#�G�yZR��o��4���ӺgF�*8�����68|3sĿ�]V��[+
�tO�^4�(]��*�ǐ}^�#&Uf��VٸsF���ѡ��b�i��t��a"G�m��?�׌��h���R$�KW������ڤ�ÈD���q֥�R�#aJkٸ2_r���U�~�nzwYytt�\7��xdKg�\�w/�f�NL�|���em�K �rVR�~2/���|�eW��L��nSH���I�`hn*��-����X����O-m�(��fRd����q��ԑ���>S;t�r��~Lz�Ӏ�U9�!%�^��������=��C�c�Ǳ�L1*^�S�ps�p�)[�3��>p	���&1@P.�)��wGJ�"4@v�W��(Y�*�n����f�E��ZEOV�nBU��e�ր,���(����[U�u�a�O�xO�}���Ǆ!t�e�a)�������H50C�90@��_==�/���_
� ���Krw���|���6��@�b1���op|]dщþKぞ��R��ݢFu�.���!���K�]uu�W�LD?��@U<i���<��rG�������u�%'�$#�:��)R�*1�c��Q7C�^�I�5M��]�1���f���+g8������@o���R�|^��@��#ye���0����9��A��w�܁f�N:kiǥ`��Kr�.����e��p!8M�ؤh�mʐ�5���buI�m�9��e%w&��U��ʆ�\_x ��űLdrcl�0��m�q2��,q�@Tuj�
���[�&VA����ߪÚ�GZmROt��M�6|�������i89����8�QB�������$�kȌc�3�z^}�h*�R��Ң���f�g����o, �>�[����U�L�8�b�[�E���Ot�k1�p2�� z�\��q4j���~��C�!�˃��H#[���v�h�E�[�Hq$
���|��р^��7�觨O�@�<̾���af0M����F�b��{o�T[��Jyd6��Od�9/��G->�f��h$6��$Wq�\s�O�Z��!Α�X+��2��J��hDk��
tO��Z)r9H�vQ��P���M*�A�> c�yl]hMqw@�7ڕ�]�r�QM��!EuV�NZxӷ�KDK��}o�5}�'	�꨺�#�'g+�Z���m���'ǯ�c#�<έ=�1l�o\!�½��.�-Y�Y��䝌KX�k�o��P��R�"L��w�wT�~�7A�AM��WMWx#{mwid:�5�k�@v�����t�5�G%�8n	,0�M��<�C_]��f%؅D����|0Ϲ|��/��@�I;(v�y�I��i3��Xk	�v�T,��z����!H�?�Ѿ�gj_j�I�'e��W:����Lx�<#��hIE�Wm��:�!�ӛ:��|��~�����}��2��=#/i���I|*�3����}��u��gؕ���.d���G�>��� m���f݃�����{=�φ����=j��*�����p�
�ٔ?]���e�4��)G�a��;�J*+��.�9��74��[ Vu�Q���h�]�L�Q�PKl�j�_u+��'yv�r��҇Y��~��NLrb|C�Z�����+}U��������װ�)Q��no��$/nS]�<}�t�t����Z]|�yQބ�1gA�e��w�[��5��q��Yw�@� j��4��Ÿ<�l(W�hU�'2����q�&!��]��ůʋi���q!#������-[|K�/�(at<���xF�Ϛf�ۨI���>7�s�C!�Ʒy����I⾈C#X����S�yK��:6���-��ܳ����wh�牿�i��v��/6S���v@�gA�MIj%<$�(6�(Hq|'��acy��dRhĘ<��.�0�`O;���c�k� V=���(Ճ��bF.�Q�m���>���l_�ny�Dܵ+�+q�d��[v��+նB�yk��O��"qb����	#3g@��.��Af���U�Z�~>?0�I]ì�c�ʜ45Oò�տv�ɵ�e� q��*�W����I�G�쇎����ciF1 k&gd�����>nX1��lI|�C�8���2d'���WxC�r�^�o��2.��hN�y]H&P~i��j����]D[I��1��}���`;	�V�S+�؜G����u�,Ce������Q���_Tt��\��Y|G�7/�hQdz6���Bݜ���M����@�� ���k��0��!-�OCl� ��ڀ�5�hq���m�)�O�y�im(�����e��c~m�(G��O+��W��vc�;��:��c-k/�������ɾD�amdF�/Th��phn���*P2���qm����K��܋�˾%���Ǩ[��o�p�0�����ׁZ������|�a�l�T'�}ϭW�܅F�?��.LB�Ü)�
��s���.���]Y�W�V��,��Я"3��w���.�|GE\�C����]�q�^��:�_����5Z7�~J�ߛtJ��SQ��P���*�^1>"�}�z8f4]�?��5������S�t�o,I��1�]	ͽ1�Ţ���皤�X��ؐ%/w��}b�H����+*a7���pâ���<�P�	놫a�b6�S�jg=��¶�$�/�l�J���!�!�|U�>)|�D]-Q�2C"���<�ps�ڴ�RFI�6^�a�$�~�s�N���In� ����K��Ъ�{l��P�C1�mtN.Ʋ��/��^�F��8���0��D*�i��_[8�6(�\�^Ƈ̡����>)45�NOSR���D����3#���ނ� ��n�'>f蕕�k��xtۭ<V<��� 5�������c�/�5-��6��^9CU�ӯ4:b`Jъ����LU�k��b���M�8�յt���93�ҷ�:b`���2�E��a=̽�
c ���l��X��	q����z�wY�j���yR7�0���q�BIX����zA�L�*$ǳ���)\�$�+�!����/lD��Y�(��h��㌀p�^T�ۄƸ��G���W�⺀�O$0�Kd��n�3r�L�m�ն0i�Zn��=t� D�w69�p���������&0�HR����r��������:��o�N0F�J�:8�v�Q�"�h\d"-�6�-��Q�Z��˙�Nn[LmtZ��	bT����:�1T�^.=�BY�Y��C?2���m�K�wW�+��p��!6��W�����bo�O���]N�X@������]x���T�Q����g�y�Q�{5��Rwo���z��#&����D\n�*� �0m���i�y
|(_�D1 ��ދ`���������`5��� ���:�G!\Q^C)����J��sU�Tg�+�?�uE ��#e�f��I��0�	K�ŭ@K�S�R�����Я�2�%�{T���*+n��b�`�d4?Io��G�lѧ7'�tq�%�u�K��b-s����j9��>�̚�e��/Cr�Dy;83�ǶA	� ����i��)\&3���pV�Xμ����0RY�r0��V��w3�V�C�'`>+)x��'[�},0\/Y�T��5��N
��L������+���/��3�o�Z���L,ߡ����6��C�ǆ�r촙�����e���ϩ�[.:�o� ��߬�o;d`b�X-����R҅�@̫)œc�nd���o{a'���Ǚџ��cE�D2�*L���jK�K��H^�����C���P�T�;�ɜ�uw��� 2����
ŗ�r���[���?薟���ZV薏�_�,�A��w�����K��p�u��d���=$��5��o�C�G��=n�'���Z`�����.��q|_��leө��^�E�/�3x@Qޝz�0�ݘ쒛�B�AU3��ݫզ��k�!�TӋ�.�ŖVL��A�%w��Yv�c+�?�1�N!;qM*��Z� �Jmh|\s\����E�&�GS<P-���3��^sd�A��ӳ�)�Y��j�Z�_���\ǼM^m���?z��y�Y8�9�RF��|m��|���A� �����;�����O˜��,�0�KNNjx<K+�ዲ�`/2{@��k�Ʊ��{��,�莹���2x���Wi}��%����tCZy�@�VV�	�$���?�!.x�W��0�U�w���r&���HC��;�g0�qy�b���a"g�C��`���M� ��hG�>S�J�&m��tB���6Dƛ����h ��C�g�:X>��2�ew>5s�O�M�hp���>94w���Ct����R����M����R������su�R�� P:���H"�3h�KQ��jӕa���һ�`y�.���) ����8.�k2L0S������Ľ,��~8��A�W���ڏ�x�!�R�T�5��{�)P'�s�5�c��vT���֩�V9��O�,��_�0g-@�C���Sp"H�꬜���<�[���6M2$y%���5�Q�<��VJ���Z,�������xF����ާ��-��%�^��ڶ{��	��?V
䰏8=� R|O8U=~�k�N�چ�Jst�jD�u?c�=}�q�?��ƢSĤ��)#L��+���r�>p���<F����?p� �i�����U�O)���;uϷ��U�����R=��f�V6��dg\�5Ӕ\�&�⍳UK4��g`�`�+�xm/'�)����f����y�Uֵ�U��Z������@���=n"��ɓ/��c?
{1�p\P�U��M�K�|�r�/��˖�wmҎԒ��G7��N/�,C�ղ;�C��"������Ȁp�J���/�H,���4'M���i�2�L�_e���࿄A��ѿ���Z��B�����ȞO�9C'`����;z�k^�p8U�~�����P�[M��v��Y����SIG^İc>f�Q-����.
��oii?�|�ˁU��P`8	%�S�Eʾ���ޗ�;1�ikl�3^̕����+�4!�������K��ng�����,tM���W���J�	��G��w��挿SV��'<z[��*ˆc���9�����a�`Fx�N�O	�9��#�iVI��m����w�y;5%v�6�@�P	!C�3��K�żt��Gx�^�e{i:�yCh�F!3�s��a�tG^��.����Z^ZNl:��s�k����5N����W�4�5������@4� �����h�[��Q]�'��Ϲ��w��ֻ0�V�0�َ��|�Xs
E��%8��2#�?D^�)j
"Ϲ?�uLi��@��
Z��M*�J����0Yt8E��}����Y��b^0\^���@��Y��G�a��3@pX�����R��J{�����sX�E�h��;�B3��&
Հ��N�:AORbů�\I׌'dD� D>��n�W�P\N�-��={�|�e���"���uK{-�<��Lw^�b�C�9/b<K���طrn�r�Mߦ�\��G{:��:AF�lJ6"UK�gǇQ}'ca��a�%�z���uSh�_:l#�)�;?�	2Rv�S�F����蛒y$7d�\C�<�a�{�}7P���&Ĳ��j�XdLkܟ��n��M���7�"�����7�8�7doR��^�j~C_]�:U����Rl��3�r�b?3�f^)F2�W�cl$���M�� 	}�>��!���G�߻��/kx8&Ӡ�&��F^H��o����A�����0"�B�z�j�O@ ����H��Mn�[��d.լ0DG�S!��A��E�D�l%~<��h������{���^��Z���[Z�t����ۜ��ђ����{Ć%����/��2�Z�f�d���N�]�5���9�Z��2�y�,r>�N��W5�9��ҭ�ƅ꺕R�#�ƛ�I����� ���
�(ڀ&�X��RGߗ�^�(n�G��}(�3���� ����@�a3UEHc8����O�ZM*���?���_�U��2(�Lx0�Z,�[��jK@��t�i�}�k�6���I01�(�{ڷ�_�Cha�g�.Q�"�%Nbj*W�a�ìO �Δ�����=(Q��U��UX�)"9R��p��my�D�R	n�';��'�+��	��|�PJyc�AԵ�ԇ}�5T����*�^w�^N|�|��__�[�j�jԎPYQ�~��U#�6�������i�ƀd	l����HT84��Ņ����u��V�N�E�)酦����g�;�aԪ@� ���Z�ׂ��}lX��/�sw�f��T�(��U��Ə >��l���fB@�מ������RZ(��!
����Q߱���lgp���ރ�6��FIY��7���y�����&�l'�7xa�¯Y��m_o�?�zy��#X�i}k�VK0H��Z�Y�( ��&�A"����I���1I����2���t�_�t�����Q۶k%ֵPH�wqM�� b�m�B8�B�'��Ov�J_������Mݫ86'�Ȭ&�p�h�n��(�4��<5o0#}�y�!�4r�FT;�j��=�f��sq�,Z�Z�ֹ�q�Μ��o��!�P�B� ��t��3��L~mn9�����Oߕ�5Ȣ�T��,^�q~�L "�q��E7�0��e����������|O��i��PV{�#�g��%zd Q��g�F�{_`.t�Lp����w���9�Bĝ��[�}�x�A�'�Z߶R��Ϻ�.��<����9���J�+˞rܿW��QL�@�M�?/'����Ѩ{��n)'���|����I��3��j����
g�����Ä�9@=z	��^��=�c�2à/lQ��'�AX�V�
�Ly(w�(����$�Q<�qF��Ϲ�}	���?�~�_Nk3��C����O�=�:�ҤL)��E;��2l�X�8�3]�0^_�p�	��T��nRYa�U�2���W�����]%�a^�w}��Dh�E<�3Yqhl_Q�#��i��l6o�������X0��n� C���eB,��pC�k#f��5V���3�~08,TD��b ��V����&]*ۘ���Ap'����v�
o��q�"��H ��&k�"_N���ո@	 �+�<{wm�_�B��|�i#�:w���˕���
��⥀��Dׂ��U��7�@�5��"
�d�q�"��(��Ѯ{�������
-Ș�@M��&w/��>u/l)��%�eȐ��y�gz+��2Q������x2�d��b��*�@C�h��M��эcV�V�Gul@~%��A�?R���5`P����c���4J�e�_��]��|w�<�p/8�]����x
�mfv`�,��`66�d�K��GP,<���4H�Z+t����X���5���@��cW�ٍG�	��QI_C���3R�-D���2����&�z��5V]vj
jh������_�Sl2 �*刞��]�8x�2-'./��㱩=����)��j���AS�8fD��ڂ�b�c
GF"��g>�̝RS���a��A�Hӊ&?��� ^�CIH�I�����(y|}�q��_s$ߚٕ�Lv��7����[��t?tÊJ߸����3����È�A�o�j��W4�������|�[,|�/d��a���$7����b|Jr����Uo8%�L!a�w���3?�>j1IPuӳ̵��;q��f�DAE�o��>���[�;K w��K�NV��q��h����yt��(���
��XTs=)�)v�Y�C�$�7�?ݶ��[V��lzeT��"?�ҵ��p񞂻ɜ��P��r����9��D��'Q���[�4��7õ�!|î�%N����c�2�2���a8a�a?�O/wM/{�j�*%��_m3]�����D�����M����<P��?<?��v�W��7���9���)4�4�>QA�'A�o��P����e:�r��.���l�&!%z	��'wҚJal+5i��<`-)�������5vL\V��/C��E(���&&��!�L�_z�o�W�5:�NG��cاSx�h%�U�Pe?$��zx\�׾��K`ه���3>�^�E�)nht�)H������F�p��`�E�پR�Ek���C����8�DσC�%7�bu?~�cc����Io���},<BҒ�[��J6�*S�Y-*�DeU��QX�}�ġ#)�h�Y3]����SO�QE�*0
�b�5��ʤ�-*w�74q��/D�����(̯U8�6w?���HXyEY�M_d��m�o�%i�F�����e��&�V.=���`TcG���?�D}�`�ٜ�k�����?婋�쥍�e�����t�`R�������W��Zk~T�R�-^6J�V��3�� m��R�����!�0�}d@˃�P�q8��Q����ӀV�){���t[���[�g�� g����>�wŕ� �[��?~��������N�╸�S�����X͎��J�@�eQ���b'7Z���-�OXu�19Z9/־�	��ÆJ��4b9���#�"B*,���!�ƈ5��ώ�I�v����B4@�6�˾����/�eq�<�Y#�=󾠥$sD*R(�d�;�"�y8��V�(B�����ap���7Qe�h7��a�r]*\x4K��NN:,FU!tB�
�ϏPp���<�a�XH��9T�J����e���Z$�;BV��סq}�M���G�P�L ��6�Uo���?o�3�3����f���}]�r��O�Dz�Q9�����Ln�˸s^c���@$�f/��k]�O͒v,��F꽳��φ���OQT���SP_d�C�F�w�zD�f���_��Q��Ng=4V��_��!�1HP9��S�J��R�<����20�ɼ��3z��V��0k��wK#q0��I'L��(��Dj���f;x���!�+�s�����pVCk
;u�����L g�Y{�>s@��)j�MK�P&�~����
=��;�M���)��>�\�$�Z��#VD��n��{�D�X{TP�у$1tϯ������.̓����7�f)�%n�~��s���a�H�K߿��n��+M�zz��*�����2����ʭ����P��R��)� ײ�r�����W�;�M��t�߸A����'��=�l��χ��1͢�k'�!�w#~eU�Z����}�׼����%@��@��v:KSɥ���D�}�y���e�o��J \;˽V�%"�#�E, ���|؂=N��9S�$�ל1����f���-��͖�&!�]��|q��x)��H�ҩD_ ���/�0ݮ�(=�z�E�����l�̓)l��
x�����<zec�t*��d~�@�X��d]E��֋p*̓�G��%궎���R0c<���p����d�ؚS/^���+|�ǩ�����|�\{xب�%�ټ AYy��wMeP�sx�m�4ko�����y�ZfQ�cw,q6N���qZ$tXԥ[7R2���T�:�*��+�L�+4$2��MK�JJ�F�����P�Ial�. ���I����1�`,� �Ca%��X�B�_�3�W��&~a8�N^<{fh�<��},��$����ؿ��H���.��z'���y���Wj��i��Ǧ1AY�z�W�g�n+�-	�D��bB��3_}Ē�d� ��7�6|�6��D��L� t >5M>�Vs7|�vۮzk�eD�@e(������S��| �o��B�`��;%~@�QeG��MG-�#Y��n�[�4�Ç�['�i���!O�.уm�.@S�/��݃��ym�v��/� 
�����,�٩cN����f����{A��?�l~dp�${ه�+��\u�� #5ʡ�3<8����<o5K�X�A���&��ܰM���<#�4R)���{�z�^"�f�b5�wz�ZBTu4�x�؉�h"�դ,�H���[s�4��k��MU���>��{��"e����j|�r���=��m%��<E�1���>|�K�;˪�E�n!�獶�jic3t#�v48�I�J��Q^�O��)e�9�؂��.�������´���5��7�m^�~?���O���pReTX��r�����4�V'Mz\r�h�d���"]�>'l%~�� X��Y?f^"Wai��gwBj�C؃l����x���f.<�T>�5n��`RX�RL�i��y��S5��39�(��RH&Uҏ�W£��
}xb�K�=ST��
7�Po\��wH1�>E}�ܢ)06�\w)��<�E	���&8���6#����2�������5e*��������c�5 �G�G�5�-� GZ���
)����<+�{������J��]����LI��w�Fmkx}�E�[�ZW��1䁦5p\z��e�\�K���!�`Y��/��\9G3]���iޓ���>��snj?~(�:t�1��/ށ��]��>m	K<{N����Š��%P?�qg�l�E�d��a�mTԉfY4O��r���Q�!�� JY۶�vO��1��Eq����4�F}�;H(�b��7hR�A�῿��.&����d��tʝ,�J���(�h?��'Q�>��
*��d��6�u�:�O���jfl�Z��:�xx06"�c�u$��X3p��;k����_V.���?��F����� Pu�B�	��I0�K)f5mh�*�U���+c�<l���v��|��&�Eg�v������2eL��s�_v���y8K��S�՗6����k]��n�ib�F��� *��Z-d�هeT>�db�6�X��>������f#}�*8�B�n��G�@��{疆�t�lJ�`�p�s�ߩs��Q���\����� �6*���ؙ{���w���g�?�M�l!҆3�[G�=��)�w��^B<Vh�B/�[0	b�q��h�~3$8̦�R�Tw�oNfN�rt�!53�q�p�N"���wT,�������>O���l����Ky͈~�0'h{��(*SOq?]ںi}X�u)J�I��d���*Ǐv�Y|���M�)H-�x�\'�B@aH�0����<k��^�N}JG-��Z��sm��G����(�UW�[\6���i۪[�ԡ*�b�/|?�LLㄸ,�Ly��Y��7�|��献�j:@p�~VV��%z�(D�f��Aސ�o��nRS�I�B��>8��u�oՐ7v�#Z�����af�CQ�D91��[��A���B���"�v
��˿�Ns`�rܠJ�HքՏ�I�"�o��u���)>���!Ev�U���y- ?���5Y������9|äᖀ�Z�G�4j0�b�=�|��/W��u
�:B����g]�N6޸���=��3��������T�K}:ݿ�~;_��e{J<���
.ہ�����=Y���˅4̺����^Y?bd7h�4��� � K,�8n�;�����a[����� �ͿQ��h=RU�l��$ֱ�%]�ɩ��o8Ϩc�[��&eBw#��Gb������7%9A��v������w�4P�!����w	E)�?������V�t��~�^߹>�ï�Ay��D��.BO��D*I"b�Ψ'�?D�"�߭��}x����B!9	�箧��JW���`���%j
m�F��;��-�n�Xy�1b]��PJ~V
�Hc�����f�nj5l�7ۂ�Xu�k���qX�%�4��{pg$��t��x����B&.=�oCY��0|�7�����B�uN���Q�X�/�O7v5����y��1�'����P5�@�3�Ft!�Y���s3JN�}��j+�E�=c��9��B"�}n}KO;I}���M-t?���9RHt{b#�1!�木�2�m
c�Í_v�J�r�a��.s��= �Q�}�3����$z�?���=���J`*�ݞ�]�m-+��͂Q�s��%������K3v�hd�X��6�/>:�-Y$G�Rݷ��U��V�Fn��gn�����2MA�W�ng�zn,!�oT^���B�#ĝJ� -��6��6�٭�]ݐu_���e��Ὴ ���eӠֳ$�����bO���"���p�<C� �)��Zz�Í�QWq�]��T�ܿr�A%[ίn� ��*�0����W�']L�u��5��u�//2���j�ۿH4	�1i��M�u�I�L���EK���G�q�+B!ה�ρ�z��nF[m�g>^�9]�Ł���o�g��b��$=�-)��@xU�kM����v�A隆���<��&��,��CL�K�eR��L��3�3,�
������m؆� N/���ސR�:���_t1�|�P��r�@��5�a��[-P��L�!	��[�gG�+����Q4�Fԛ�L�ŝ���y�#�Ƞr_�vz�򩎄�8d�՗0���7a���K.�UTB�UB��ӄ2�l�m�ׇ3�K���G��#:�r��tEU�4��@݈��b��}�6l&ZCl� p��`+��&%1B;~�x������s��$)���%h�����cꤠ�3B�.pmN�5��>� �vof���C��VS��?���¼a���uM�e������O&ٴQf���m;� u�>3V;w����B���`�h�`�*3��Hb�C�iTҧ�|P����P��Y#+x�V�{��;��_��G�/�|��/ ������6E�%�d�l_�b3y����Ū����s��J�:���NOjh��ѕ�)^H�9rT���mR+Q�1�<�Zg~?�@2A��8H��]����q�K�������$�^�	"����c���7n�~0gJ�?^�t�}]��pz������r�㛏βS���Arkui��{[
��7��s�Lkkm��l�����f�ν�bϽ7:��@�>��i^�T��K'7�s�؋a�l���d���F������S�ޠe6*��3��m����*rSG^�������t��6e;4T���B߱A���U�ߣ@���5�yj1,ʻ���o} ���ihw����<Oӛ��U=�ZP�6���1��c�Q
�ӳ=�רP�V,�l!���3�����hR���q���@�O'�OVH�|�;��M�Ȁ����uV����B��HNg��6�aq=.��0�	Q;��B{�: ?�n{\����/�dm��B��esG�?-'��]ܼ���%�ߍJ[Ӵ��%��,�?���W=!�S)�g_`u4�����;ֺ���2�X��`�"�)�R��e�]h����L�W�y�&^wp����0�G�����D
�O�7mk�E��Mt�jj�N`�~ ������oۨ��\d�LI��,`�\5.��X��@K�>[?�c3��e�N�G�Ҭ����jñȧ�ѐ}�Z~�]jc19m���b+�Ƥ�L��H�([j��J�`�I��dg?��i*���t
(�<��C�:u4J:�y�����|A4�"�<�g7��O�{��
s"I{oE�b�����bo���|��5�-�60��Q�SO� ��8���։�@(���zK�!� ����ny��p��T�l�!ުȼ݊2M���lҙ�:w$ J���d��wT���A�(�R��<��sGU����f�Ш�i������a�@$�7FC������L�n���)�-j8Jwr��,� 2�1���Ӳ�`�x���b�@XYd�f�̸j3�3���Z�/�����Sљ�xi����NǏ�ҵ�×-E�k������M �����5��aވ�{#߲�i�����@r!.��oYxs[�&[['	K/\1&f�N*�,����O*&�p�U�k�ARyPa�e������B'd�Y��s�ͯ'�8��x<��GR��C���\�d�.N���#��������NSuDD#�"Թ��;��hg�� ��R{�n����W����>4���Y�l����Yd�YL.��C��ƨ>�i�u'�kGi`:24�{O��G��-F,O�qؿ�J����y�ֺ�1#�^�z��*�С_�J�a?�H'
��&�~^
��E�-�Z�19i>���5�H�r3@DQ!m�롽OI��=��3�����"����VN0�.�I
T�d1���Η
������{�XWPUlV�y�#�rMob1��e��>[2�VW�)�8+��)��S���ǟ��1�n��=�H��M�}�i����"���iW-��S��j<�H��S	^P%�]=^b��Ql��k�Z�W����Sl�c�7W]Hb��iKf����4t���j��3�z�;a'ꑓuH�<T�l�Wh�ZJ��S �<Y?�����MD�AO�DľMS(��E�-��S©��d�ݢ(���x!;�>Wܶ��.�<m���{��&vx�3XZ�6:�_������`�Ї+�u�v���_�)Kwvޕ�G�׸�kX��$�㇍�\RiI؂��"����dRV)ĖU���r�߆��%؃�!熼��m&��m�_ܿ!���:�A��J��Ǹb��X���4Z��s��`�Ӿz�#}>q�%��D.���{�;ë�[y�݊�C�˴MbKo�Ĝ��t�a��mx�k�Ͱ�@����tk,oN"L��	�xF��/�3V�tw ���&�f���;�k��ľ�n����S,//_�IyXzY.�9ߍ�w�G�${.��B:��eOp5�W�&=�)��ݱ�>n	I[��ڵvQ����W9(����b��e_ ����W���]�S����T�T�~���!>(��pG#�"���0�G �:�}��8B�j�8�>���#�i]N�x9�tԑ�^B��U��	��)W%��'��ջ �i���mM"�_!�aLcGټ+i �"�����gZ��X��E���k,#��du2n%�f�$IX�N�<�@ȕVb�O�_"T�[Z��u����o���z�LW�!ڨ0�_�^Oz�ҁj�w"�݋�@��WQv�|�R��LNϪ�q��oE����	g%��U}qe��gi�c$�v.>�X�5���������8�Ź�T�G�"ZS\��J2)�o�?������!Ev���wmoAЛ�xuIם�W�ʲ��n�r��۹��FX4�e�vt_Y���
~��wFˁI���suJk��G-��-ϓ�~8̆��'�0$�S�qaM71�#�}�:p�V���7����֡�"��Sz�@�����c�gÂ����qӷ�9`as�U����5R���F\���d=س`�4���}����uY>��ݓ?�)8�ض���\�T< ?V�[Պ!=�}U�lL�م�=�he��r�Qt�~�P��D���M�Nk��Q�ƍC�j6!�O/�#����b*8�u�C���#�+�����x��]����fq����(�VE^j�:م�VuB����x�.~ք�-�F]�j�s�����=��D�<���LEWe�� ��)qLQ-��A�)+��W"��	�~��V�G^Kbs��hDs�巳��i�{�Wx̦���R��7���=��xF w �	���
�� 1��s>�eD�n�#�����q�}�,:�&Ts��X�� b��]��i�+�ۚ<�(D�/�.W���$�jߛ/�&.���r�w�k�D�\�g�i�f&�� L' �,+���������|��@�!룷ޫ�1/?�~Q`]���4�;�tm�=�}����zsn~���߬�W�.�EPi~
�*����jn̿^�?*���_=ׄ���xb�f��M>��4@����4�jӚ�T���\n讖%�Օ�L�4��4W:�7��'�}��~t�F�l�c�?�_BjhxSSv�����h�ֱ"���J���&j¢�����j�����4����=� ��G�CP��t
ZD>^?�InbN'�ż��O&�tO޽S�*R��u���|�� �9�7���⼺�(nn{SP�պ�@��jȊ�9��B�O#,�npH�X �|:y��,�Om;��Wx#fa�2I�����I��[8O���ΤaTT�7�Y�;��C�e2=6��p�Sgb����`�lےB����tr,a�&�k��R�ya�$��q&l��M��*
�X0:�#�g2�Q�xY�z�l�1���!�q�bh9-�7�ǘb���|��A
�A6J��[�kد��ϙ�t&Ԩ�P�©[������-r�M6�XN�%괘�T��94�rz��(�����Q���	|.mϒ��:�P�7�[��P����(�W}"R��pY~�S+�KQ
E���������|Ȅ/���d��iN��v�!�b��Vrc���r�Oj�7��G�A!Ĺ�&o,Y�-�j���`�S���c"�N�w�1���mq���|�����O��ON��Ŭ�3|�F�G�,���W�g]�P\��xx��8����R'ѧ:�Yam1ߒ���4O(�&ZY�UjC
���G�k��w���zeD��ľ�]g@;�*��=��9����%Z�I��B��ҚL�瑇`Pt�CxN��� Y}�9�Z�(E�	�9���){ίI�p�"��+p�۬�#���Vk��S��^���[f&��3��aB��^�� ���ڭ�T��՜�zօ�q�h��8���1v������20�U}&�ы*ZBK�^(�Ԧ��~٬ږ����w.OSX��xs�cx9E�ީ�za<G��JS-!*[ZP��������u���,���TY��Ά%5�*�	 ݉%��4XW�`��R�>�����,�f.�̒�Ȍe>����'Q�X	}��F�@oNd�#��XO��-ݬI\WT�wf�u�1��GV��,����;(����!IS�Ԇ��>��QI>Z��18H}�:
k�7U0����z]�{cń���ћs��?�����s�[/۲�(��{zI��^\gIPP�=�Q�+�A]=S�-H��P0_ۙ�6�k�R,��(_��Cd^$t�W���}�/-����"�	\N����pIe[��ڝLG��%��8����5A�^�h#��d�+.6~�L/y�G�����[�+��ODx�p�Pٯ�^L%��Ͼ�`����oy�+��n�T	���4LXKG	�^A��V�6H-!_��"�;)����ԣ���Len(��:���Va	��1��3	J �J{���~����jM�C���\���z=���t�Y$*�C�8:��@���%#�v��8[�fGR��rEJ��5t��d%Ց�A�G�K�.�З�0m��1JsՆ(-"$�ѯ����4��ׂz�\�y�0F�P�
5�<}V�G��	�sn�PAI!�R�1��_.�0b)Ƕ	��6��>�S�Н"ZW�pbrbΐBַ������{��A��[ ih�0�_�n��Q�e����1�<�B�Y��\�.��gfҔp����4��k���|#��u_Y8o���CcٽSχF��?�
�[��x�<�I{��<�;���z���F%����K;�Z5;4ۣ� Rr���8g�jY���̶=+Ǔ_�r�g1����ı��.T�Lp	��=�	q��g9��&��%�W�'#?��B�@����F�=]fv�>��#�\	3�up|OMztv���c�M�U�����z?=�md��}�t��=�rt�s`X6�~���*o��M��=m�Z96�W >��>'��:?�C>�L"�	����:JT0�ɵM3��o����fy���2�Z]���}Æe-�F���T&��m��_;�}������*�<�}":z!"��ŀ�r�8ϊ5Y=��
2�k����X�B�f"�3.	���:�/����t�K��U�$Rm�C?�"�\��sE�z�t�:�)�\E7˫	Y��D��e�Ds^�q��KOʂnl��Z��	����ȸM�r�����u=����6(�:>9��Y>�1�G*�U���`�l�Ab���`RN�J�HAlocz��wv���ɧ`�(��"\W�
�!<[�9�	y�,?B��U���u������ѳ�-ê��_��=m��R����G�VVx�	�4ރ���S�d ~�}��s�2�)N�x5vf:�� #�䪣��E	�լ*��y�f0ʚq���RLF�a}��H�9� T�+^u>����'ԏуv�'���-��턗Ӫrz�m%�T����`J��Qk���F�Qq,2��Sm(��y�2F�����R]��ӊ@W�%ȥ�S�q�A��o�ѧ��B��)E�k�}Ɣ�fO`�>`ҳ��6� �W����!�㱠ɗ9�ⵕT��6�K��t�-H x��a��ߍ��s�ZH\�z����F��"�G@��e������^hH�3�h�_^'�y����� j�p�*u�����&a��,mI�0���~� ��6�eo�b��)e�݀/Z�%Kw5N�d���n�c�V��f�th�v��f#=����i=8s���$c�]䳣�@���M|��%L�'�upn��y3Uj��D_r72����OV�����c�忇�,#��}�5d�/�Ǣ"�;�t�&�2���_f~7��� |�8��/;%YPa�O�y3��t�~γ�|>�r����;,�+g6O޼��3.���7ղFr�1׼8���U��$9eT�#s�t�HCo���f�Ft�{����;hQ���B ����!�ʏSg�5#RzTb�=R��>���)���!�)�&b���>b��h�ݱ�����\�UV���S[����\W�;�1ZZn1I�T�w �>2|���5!���N	��%�L�M���t�s�Xڮ�tNw���P�XL����;O�L��6ƒ���ʮo=8�������0�-�ܪ4C6d}��O���E&��Ӷr�ҧI����b�����~VN�O��id��)0?����#���L��"Q�p�c�֊���.�1�3K���ZaB���4��=�n5j�J`�|�i�q��֋�&jW?�^�9Ͻ����
�w���*d镜D�00Dz%�����rc|��f+���QUU���<`�E;�b��6k�A^�y{g��Z���\����<e}��W��P���#���;F=lJJe�t���g�]<��gf՗�*(}s��i���ytC��c�鎙&�1�iu��p�yB~�'{�����qD��� ���r�dvd�Y+t�4��-����h�~lQ������7�P/z��w17��ŭr=��*j��#�ώ��s&=،��{���*ܧ�N��6�� �[�R�'o�xg���*u���Hf�a,����-ώt$䬋��Fkᒺ�}��kȤ���;�-�^�$�����lK�+
/�=>���B����p��R3���LU5��c=��IU7�ɋ���=FFq`������Dp춃��}���P�v�`�`G�&�o�{�ic9�����K�iA[H"Q�r��	��f\wBtx:F�ub ��a��\Eo=��8բ����d�S�={5�(�/�L�W�>ۜ�j���4��{^�<C�I��1	K}����?G�)g9|��멿$�ݎ�Vh9j���<q�2�KƪXNN|eu��cQ���gA��SY���bhj����)7�{2�1;30�WDN�}�%w�ߣ�2����1��+����(�~�7:�VE��`C�Q[~s�?�{/
�k-tB����)T*���Q�˔�" �{�ҒqW	1?��Pٯ�WG�-�
p	D�}f��9T�&��j�	ʕ��������w�%F�t
P����gW�T,����M@��뎯ۨ7!)8���@�)�4��!w�2�q��|{rF�}��A3|*=�N0!E@a=d��f�8OL�� � H����[����80GQ�.� �p�="�Aܷ�!�;�?�8-R��:����c�&��+WcZ̏3c�C
�d=�=KЬ��}�ֆ�`�=U�s��R8:]R��!Uah�aAU�h��lL�n��ܵ2�sI�_}���!�V^o����6o)���Ս�B�:c�?�L�R� P�h�U+AL�I���&%y���?)WjdR�R�6 f��*�D�=4��Z8�&y�L��\;b�����4\A��ZL�V�ʓ��>v�������˹iSb����mm�.Q�tr���������=��}�T_���a��a�bH^jU���Ok����������`�;'��m�Sj��}��")��`�C�3���估�+� ?bU�L�β���Fѵ#�B�OJv��m�t�wY���+!��h�^�H���P�=u�����&��{��6��,�u�pdt�v�@�A{s���_���f��~5m��lV���m�mR?������R�u'�5�{���Ј��J4~F-���od���}I�aT�Cf�jw�;Bs��P���X��"��	<}+:b$��<a�%���j�W�@�؀~��)�2�Z(�Z�\��W�t1����w?��GK�`��j��N�����$)�����B����o.�;_4���aw������e�d�fcZ��o;q�A�bŁ<��Q���[L�Uަ������Bf��P�p~Ը�~d�(�7���g{����\�"ʂwq��d�Ɓ��IJ�A��4�R��)S�1m��4e�嶏n��;�v%�0�$6�UF��GvgV�K��ȫ��|ꑫcghB����ږYl��ٳ�<��mϋ�W���-�ě�P$������.X��Ȣ�-�wM�#�H�$���r���adW4g�e�:��z����E��-"�h�w-�(;0�&WXBYo���Rn�r��T���;��g�=3� ru�S��
ʖ�R1���=�Ӊ3�Op����I��א��byM���l/�5!��ۡl��&)����0!�56	��O�FѨ�ьrWߨ��V(~���^��8ӎ���/�`�h�xߡޣO>Q�'�G|Jı�K��p��S�+_�+�$�Ž��se:��WLV�7��3���e��>;�m���r8���j��"j��5)��X���7���+n���۠Gb�fenp�|�����[�=Vt��'`.�g��֧��?zfД}�,� �>��f����(o��e'���X��.I�
e�7*e����� �/��6_�oq��9�ǖ�o�έ�7.׶t�F	�M���In�.���������C��Q�P�-�Í��4W��.���"ߑ�D"_���U��f�?klM�
�R���3��̽��1�M������B��N�_��x r�mE�P�f�A���܂Iyw�_@�=��^gy$%��;�ƼŇ���v��P���ojI
b��=�K�h���W=R�`�ۦ;buD�R��^��͜ޫ���$/��)dv�#'�T	�iUҹ)m^�g�	ԝ��Ǧ��}Q���oUQ[:�>N�홣�Y�s��cz=��#�8�G�VT��N��Y_*1��@�wڐ�(L���Hԧ��h_�J�:P��le�riDV��w;}1�v��RH�@���%�v�j�gQ2�L��Q�p�xb��Iy�n�4VA����+���/u�9�خ��oȐ�����-�^�܈#��q�?NPq!��:�Y0a[�GH��b�9�c,U��Ū��l�+P���ۿ��m��*.�2~jtȾ��\	�"�s~�֣`��\��6�gbw�۟�Q�q-�����9��c�T���e���\:*�p"�����vdfÈ�'6Lw��d��<���8QP0#�j��Z�&a$���NF�tl�]��������kQY�.$Z���P�d1�T��h�]ʪ�0k����bk��������mz42�W{�s�qf>gj;ex����W������%��[�cB<N�wh�#꘶ǣ�J=����r�ɜJl��RC�L[��� cC��X����_� �����h�<��U�w