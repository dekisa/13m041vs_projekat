// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:27 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EIOKk+pRn80AWmz+Y1SuyTgKte5UxlkaHp6iLJfUyh/Jer8kZsKYZLPDVZR893p+
KeJEV+131J2ki7uBlTIfCRIq7sqyJgH836Uf6/TTwQHyu8xys4pFdJ2rGtr78/oY
F2BKv24+qEJ7A86pWfpZxG95xK9TU/8F8yFX+wiNzl4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 110560)
4c2INyh7Io1CHxYsT4+GuyTkO3CPPLvXQGDtVGHOPeu7nQjX4Kpp1+yeuADaR/fF
OpuvrHO4+8jvzAMiOivuDgJPJp2VfsE21Cf+kAXV4hnm+z+2T7NZ1/GY1sCPReTF
0W06hpP6EdoQfGPoA1lOYtErPPVYiXFq2o44lx4sNCivryftOZcIA/xiWAyz/IoT
lDkiy84jTaKRs7TKwOk4/n25k29KtWh7xqLd5xcN4y+9FFlw5PW430fhFHei9Jb6
m3vbWv8czptt3kInZFIW7Oz+MU/VnuEC9QljWHpU4EvDcTbd/2r5J62RERAQ2TWt
CSzoiVRvVwz22Xa2x1hgoQPyTyseXmHSF4GJpwD75zay3nHXrBTXcyoqbhceaFAr
9V94Bo9wXViSAeD4Q/6WadStDfY0jh4rz2WcCEdIBqVbhXTdgrPfH21PAxsqUazY
GL8BwqghdGzGxhZIzNI/FTaTKCZdz7umBeCxsx8oaMITIbPkcEVt4SiLJf0XseEX
8YBmdsPo07cpv9SzMaIrPJqMmD8I3SHe+TV8dXVCdSaiMStcfVAui53bFAEH0mz4
1XPoMbdUkt/Bi5tIdziTSmDLKeaZRvbH0serJo1+Qi9vBbxZsLGFfPON8S1FmPry
xW1/NIPSSo/lsJSpGU5aaXb5H4QzlEGWSrq7VKj2XWP6pck4kXMid9E8++Wfbo2i
jpFIqxLv9CogQzE2Rxt4vvmza5jsWdn1kyIaWXC1C3JsleqV4gFXjkwZUr68KxQ3
BgNCOkdHt7CW1u1JDvnSsbs1MB851o75OScU6Q6j+GZNdWmaKWQ5SWRQD+TzeLDS
elpRC2hz36HZAxLjEPG8FKsrGnH+ZU505WvoAcgEiaiN4AVmkJTBUOmdGmHTEDfo
xPq+GnGE5Zd9b99ZudXu/FKfbkQ2IHvX/KKQwfTaKFW8DqNqURrVGt3UR9gaFqWg
nSWGy/nR5qM1ERBY+/lEqwU+FM0/BD5UifeLPlAADPg+Mlby6nU0rWSzoom6ApsT
BK50JjHWCKjyaaX9ub838nAOJhBRztFUX3L3AnasD3dNjj+yZtrvVa0Om8fkqhcL
2FlN/HJkRe2L9MOrefHUhMdK3jHAvXWpIjdDP79Cj5jEym4q9/XA0PZpPc1gz5NT
RKg+LySU+g0vZ5WzLm+eleGnC5KCp2yt5PPdw2WjMD3GVbPysry1ipwL+9Zr+9uL
8U3B13qz0MuE7z9zN4E/HUaSZzuIQiPHPyU7huZ9R+x9mMzwzQW2/KTabIyPvbDz
59fo8Iz+n9o+3s2usUoAbZDR59QsEFh1K3PGhUp6w16rjwldrl/+uTXcQibRzf8X
z07nqoNleGaTAQ9mZCb7Qt+7K6ABSoWRBCF9YwUuRFWK8/w+raNqaARwo6vUPKq1
T+p60JwFsWfEQk6ZPrv2I+yRPci8SGVJiKOtw9fcHbmAE1uFRS6ACzeaxHxi2bbV
p/gqufqqWifvUX/51h2NSMNy+1RP2TfNqEBI85/YOglNzOZTWZKeCZBGyseFCXX1
8xZUicFpmA9FNPOjITmO3Lhk0njp7botgp5Fbv3OVk0sgFFRGal6VfkzkgBt/ubr
XWFc9QbxZ+Y+ZWTV1qFzQDqWpUtGetnWfB8s0HtfQ6Ra3UBckNfNMHckUOJm2oo6
P+Hf1clKjagsPQc8lSmtGVj+EU4/W7YKuDwHIJSeRqD/Smsq05UVQ7smee23760t
yr78RUMiBM2vNQeXkYmBoOEAxQ2R5Vcp6QrlNt1HZyLpoO2HMKQ+CrfuYJehZKNq
OlEjMpfprw7DMd16oNUYNuddomDFNHhkdCjbamZczMsMwxgCrU65BrPdvoUyQm25
eEam9U9ou35G8V5PBXf6COnMzh0Zck+GcKeLOMqRbyXT+aImiLlEqKOWNWt/o6Yz
+80l15jbpv7lNE/iOsWR69xscyB9q4KjSGM7tkJScv+4Znef9ApYRBES1vD6Rrd0
0ruJSB0xEMvzX8xumjMjw69PgtgeMwruQvoSSWroDYMPNJDlE2WdR4sXs2/5hbue
X4AfMHol8K1P6/h9FHvUwKKPD9R4Cq58lwyWOAN4ZqUGvLhZVGwthwcBejQvEvGx
nQ1jsvMuTbjHDOU5Mzq/nU4iFdLH25vAUYckmMjGZ9cLXNCC7tluqeUGXbnT3MQA
rdNmNWBQVskCihQy+FrMbL4P1ovaXjMKlO7vVW+6bVlkF2t3Decltr+2C+n/mSSm
gMIWB8/J9gidcmPdAx9ROW+cmbwexCSiktyHlUFGfaqLeH+qvl/pCGr7lCeP5Gj/
/CabewclFXUYIsLMGLh29rZGPgLZrDyIZixbVqQQe3RovKLAzap1M/PrAvvivghD
SBmAqqZxWdexUD7LyTop7JQNjOiKLZgz+DW3/6bCO3E7Us5i4uGM/1bzOlFRoxek
ggVJT/Zh7EjMmD4aKNKHm5xI0kGxc/eUnEbwfX2nD9HFDKqY1qI51FftN3JPq8sc
3PK+7uVt+Erx60m0EvZjLaspJfDVdq4h3l19gdD04+3GwI7LogUDsPDij+g8bKr9
Kf9Igcz1pIsg0e3wcNzrUSeT//LNiwD9YYpIJm6QPdnBBQsZUaek8lkDNp+NblOh
armLJILJyS4X9E3yf3r272SsX5zx5wWDPD21+FXr3eFDJCdv9hPZeXOj2ccO6Xx0
VfsuO4syIvLvB09SMvmwKWSFmJxtvdUEMdp8hXzUOzO1rNvGJMj2Ai0hr41wZ71S
RHkFsTCdfNoeLVh+t6g3A0ttpQB08WVq++WDoUW/W7UHKcPf4VJw0j5A9P36SgkL
C86AfLetgiP1kmirPJwBxFT3MMbbwgME9wy2FueiEG/JIVCADIywQa4eaUDTOKzl
eNvUh/irjfVcBowdu4fM4/CLBeozopwvIU04VDLZY4xZq+WrqiIJKnlSf2R/ztB1
jcBPiHr7ti/MENP+AJ2CTIU/HxYO7onzEsPqSqT3ipiCzpa1oLJFyxaSxUjfATjs
UTPjAYq9ev3zGqpy0i56ZqgbOzQyoOn77Ya46d7tCGPyo/x84p5+S9xsPEmdVUq9
5vuaNGjoLV1+3xC18LyZt7I0b0mxHpQ/z3wnDpmlsNpMs54UrDM0TrQ682NLthX1
lNYRO42+0Yf23LttjkAPhFPhdmXZCCq8XVkz8FC5I5CRIVqFLsvpmvtEL1vfsN82
/P1UMTD/xgRrFJmGTVzVcRy3Vx4feim0/7yAGP+A/aw6QQeaUvR/OTg5ygmmbvtC
n5IA4QRm4hx1ElN0OXk1DciFagltTIJtvT4iEe+oHjoXTPoF822TGfDW0zlkQlKH
iRLtbDzPT3Q2sPUW3bBcjGzBE0jRgnQ8lbgjzqu2q/0PUIcBPRM/o7xXmeJENUU2
YviXM35uT6OBoNtBFvZaBi56tvjeGZJTLQXRJfOTut5vnh/ixqkVPixSN+RxMmEw
qX8HnBle5gGe01pbOvU/S9/7HoMbYjAKwy9syYoIL3aaBKcttylnIHAYTqS5feA6
W94FAAKKN9zHPsE3z6xs/i6vcMdzI8WFNsssQKk436FbXjTn/v3fHzEv2fU1hUyo
JiTo8lf/fiEKiat0HZzAa0BoVsmdhnBZg/qBEMBYNpmmnTqpZe6Hbx5wTopRVPm4
OobXzitKn7UBNYUO6nqNFGxRO3OdqzVl7c9guGiJzc7CqOmuqZ0ppM1WfddgB01l
Fd1VoBfyg1Z1DRX+4iVuR6EuL7G3TRgK7a4ddd7QVhojycTOVoI/LV3DOEH6imyl
dsjKYLN6AiuSxpcKFxJ1tlyDeSElS1tRJLQaVffQNHMf6n9CtaupdKInniAwrtMG
qylFa5RAqPQyV+wOZAyf5NEj6rQh/sOnysTsQ5Jw+Yvs5OtzWz4ym8mlFwGF4rGL
PYw5PJaz8kjXMyoyPiW5lxCq/NJsRW8/M5rF6BdgnoKQz48ygnjjDnJ3Nb1ZmBsU
xHT5hmI5wPS88dG/mdap/nyF+Rpl7/HxDwcv2HH82SkY1w+mpkIrxT1QH23tNUFZ
zD/35wxN9UMnzWVaxBGDnAAL9+PAyZE+R+668U5Gid7Euto5q3Xb8R5lknWVSror
U0m7V4wjEeDyLl5WSUXFoLRAXPp45xLcInZYXF55WD1+Ia/zIhBexRYwLrE3S5/8
SIRjv/Lb5dFKqrLyM9abJ0eg9IpoB1wZlmBiQctt7w/2k9ngGAA4LYLPWsWOmffJ
lNfXrfP4mpelCgf3JKSDv5WP+C/nB4sUVeI6nXddzfrzIc8in3Y64XKfdZqcuH1y
uwxDLidxruJSD/GtpreP1apuFfLMvbq/fsib0RDHl2UTd5U6ey/kiMNe7n/XGx/s
MCQEkpO5B0ZoG5ivhcFfXSsiUHhcWAaBaAY8FEMJJz9Tqwma0ANc2+dlEWHIme+9
Na1pSuqu7B6DO87Ss2XoJYdz+j0rOsqkKqHuxxZKFYb8Lgj8Nh481YxyFmQ51WDP
pkcsOqkqsl/lb2SqkMZBK/8Libj6sNsquIB7DGWDZQ8j0QONFL/+ZN9E6aTp74on
IdM0Ib96mDbMlIp7u8jeSpLp8ZVWr4Al/g3RdAr8jcZ7PkW8GgSsYsO8xNZEKgnL
FuZc7KX+aLMNRlQyF3yxZ3AG3h1ljnRGr/pEw45FEBdrvPHmf6jTHJX/48pf3J8X
EdfPqj9DCFZg4HocFjoYUTgsWUVGnXUlsrInZ2lThCwblPSRj5YSHEmsVMTeAtD3
dRBFPR8GkvyfqQRafhykKSiORHgO29RuRvO1C8JPxNsyU8jFkP4TZe6TABw9q4Ul
3gkuFwmOZi11pWmQA/W+ONJxXsBEYAsOPr+UDelLWgO1XY2Cexxwfisj27ZGALNi
4i0BfkMFAiPw0gBvIfRlTClI7Id/1w4MNw1jP4pmsBcmgg5C4pHSioIs1eh/n46o
B45NZotdPqKHmrae0vK8velDWAkmKj581PCP26vdBksQwvnmx7VdKXVEnBf4cKGt
E5+nWAfW3Lcwis1Rd395YnZ8FlmckjYeSt/WPuMDrI55n6aGfBjdl8KMwJ7RKGeR
9c8a1PrnxfuKPfcfi0LGpxxOsbD/J+Mlkmo0ZVfI2LtD6q2YAWLANQv7vQkPlCTJ
Inog/ARtSOn9pzq5+i8GYk/6ojh6jUG9KnUqhghWZ6uiEjw2U1fKchU9SkdOHvYA
usdpZeZKGoqv7jnCNyDJgdGbbj+PCcGDuUjxL7E0c3RsCMMbgM2tC6tTGgl6dmxi
CkUUzuKED2iu4mNKhNalz06gUOeCQcsjsQrUpgAQ7r0NW5owWynYrSnUAGwneWJ0
dsU9lf85Hatx8cuYPYbSN/uItlbM1sT+pQH+uHcLOI88Ai+iAsiMqMo85ShYrixW
aXMt6f7I11ED50QrH+ySXE9hvQ9OmVY/wOxjwC/NYIkXGqujOlxyd/UkX53aAWWv
eOsS5Ll/cnko+bYpeABRnLz8gktfLY8LwaKekUKtxkDkaf7cUcGPUNMAHgPdCUy5
sUgrWtF3Lf694ruXTqMZWyi6EWc/PSc2hDITx3c02jkgUZRZzzTwEtMrY7KmDJ2H
a4JZUOkdv7EOJtA7z2oNjaOptqDMoZ4Ht1br4iDeVmNtVO0K8deVrOv/I/3b/o1N
dcEAkmMKq7kcNBrhC24vz5JkMjuz6lDoj1IFYgWuaMEB/8qbHBUpTghGZ/2PeaTY
LeaFBsLtO8ATZg65muv31oUdECSGP3chz0+LrKvRxhYmcZGuebNwOPppZ6p20/gP
cGYTsQoUUeD1C+1+oraMIVXOf6C5EpI2wwkkO3WGY7YaaZ50gvCZXhXkwmI/n+8m
DcASP37NxUkj7HhDsy3ZAfgjxGejwju1WyGvlXv0ENkoXP1Lmj2EYw+i+61Mdiir
CSaRK9APwM9cTIoPZWHx5Swsp9tLEsXZ67XyWHr5SmfHdCBhzUHRgJoX9KMvqOOQ
WEBpPw7iqcrXWp6ymYjFHd4h++fWOBGzk/oUFZ3ZUOQurcQG8/62N94JKHt2v+ug
Nio20gmXpoYQoqdKMjPvsDugYXG5tc+VjfqqhKfBNZurBvuldQq0Mzj3h6hwVjRg
WM6LJI57hVe8ULS1RKK/Q1YxS14z1mnt6jKIqURgZJHl7+dQiEcfwYJrB4A36UAb
JeCyYiMxp5Wp1Z3DsvbNiRtWj44vQ0MwKpVpNVc/d4tlz23CIr7eKtOVFwzV3+uX
P/pVR264rQ9UMXu/SCWxFj5ENzY1toJ9hqqfzl1vEnkCPrxHM2U2krH/q6HKN1pc
YRnjGG5Or7a4fykOxCpSVGd3DAbcYXk3QzdPf90qNZuQPRYDR1SZGI9MeI9lw7U2
0NPQXdtCGTfbgqZpaSAdCNgJ8imvnWcwhFu70P/kMRJS28adwZliemiDdPkQPM8i
HjfmOWJPXkq/wZUfBopMfbMrxwIptonf8E5bUZ0c9mvgBCo8DxoBOtZ/JKmtJRet
0zUKmdJV9TFqa72iKhc71SsxVmK8Z5YW99sDRsRc/hqtGNsgI7uBp+6mH2oQSv3g
vdcP3GLhYQuyfcTqFLX75GZISnLgBFZUSZpsfw2sLdAnrL1v0Ult1pAhCHVKyz/j
qkwgskfeNfLdzKw2JeN31Qyjo9ZrmAiOBYCTMOUVINbU0bLCi9dR9FomZwtmks6X
PwqmvN/FiOR2724PQAo09yjbu+nSizsiksbi+GHGT3ZjVrUTKK8rzbaK+GwAR9s8
dhL3zVN9xhOW0yWNX/GQKQ0roRo5n9Lr5gLUn6c6SRb8FteUAEHrdWlXQflCkkYb
QIicXG51pM5h0SkzPFad0obxjBR2GKugoLCa8wcNzPI7VLb2di55IO88JJk2K8Tk
7Dp8pXvqJ8UzKOAw7Lbfqc276LNPcCXjFYKgHstwXrpTkgYrqjyTzIIJC9OlZYOP
XOR9DQHtJkSJOFoWo77TMuBI3BGFDp9tDePVPg3w6kuH7T5Yk2DUHExSMNSm1xsc
AsFoDgQ5lqjQKVHXm33YIp3GSxI0IwWB5cj668POBvrTEhWWORBtBOcnKpf5gaV6
1zWsn/Q9jwfUivhFjgquIk26vz66hv+ft4FW59TfDyjXzlH4iV50FEPYtGs+FfCd
T+Fx27Kj0psLypqf6pSPOKpp8vtjKdxGQyJLZl+GhwL4H7jz1HavG4/dPREQt/2Q
mVXl2eeOKLfYMcCLShZsB87FnHNfpghekZUjQyp3oeV0EbNI/InaNcgd4b3c1zdT
5VUgpmxqt4rj9shXNVeUvh72W9bEZDvpmGaTQSpgE4TiDeCrtLVuDmCUrcit5nhY
gY14CxycMXus6xdObChQh4Li0SM5OVYFqeN/JfdSj7s65cZ72FpZJgjBSifauMIW
y2vglSTdtxAbfzccHc/BcTNxW4uWpuR9igl6pO0DPOBcymW/M3PsfEqW6eIp/QTZ
yw9nBkKTL+cRZECP9pMdBcHhvZnxri/CyODifgHUdF7E0Q8gyxgPsbQ1sp9vEC9o
HpA2SQ+1CXR/Ykanj/xcdMBraAA3OC2a9izscYxpnESX6c+3SnyN1MS4VF4Hsl60
GgEM6WwTHIuCnDdvLoJx23umPeTWrJyLGzmlX3iLJ9ATV0mTKtTMT/32yx4WCEN6
C3ZcwEhvKZA5mAqt+2ll51EZlUeJYpOM1nz5/wrylLn8eU+Iy1olj824fBZCgvx9
x5XPXmAcryx0W0c/wuahKY0B1K03kQlxLI/Ym+Vf92OA/E2wb2jfpuTasr3OAND4
RxEQR4YFEkzoKy2AbSYBZkT0FG/I18TTLjRQwFkwKtaFs2Ex1+bZeDdLtC93/QaQ
IiVBzCIcR99oQiu4m9aNnI43eGZUu3MOE15kKvYrwLmV/jiteKbohkKJLPLh+Ybj
iL4Cr6nArrGG4TB+oWmI2m6aMjybcDaYlaYVo/CX/zK+8g678EsB2rkimkWIXFuR
eQ2ripGPGf1xpPphSEuV9BhBvp0UpOy4Rs9KHXrWUGYWcv6mgEKRYZysnk27xGtk
EN3SDVJgJlfOjTU1HtWB9Fl48tVjP9PJiWYlxMpn3lZrOvAHA+kt7hxdFRYXCW5G
Q0E4J2i+hTaAOoZylnAFnZIH7tI/ygiN6BO2Mo2Rgkj2J+PUkWEqjiPnBZv/WaSi
SEARGVaiXMgsRRwesUaURABxQreKFiruPGHA51zRKlQWHNcWNXcJ5CPmnn09qvDI
19LLzHrJTmg94LuYSmVbZyS1VJYR2a03DtE2+7WAUgw46zTvvJcrKFx74B9hdBLe
o82UOIuBxlt9KQvyfh665XMaF6QWUWOdHebyZbJYcIzU7oiMp/C0KYM4YO06BC6q
CanoDbF4zxW2kwAwxlpkFSyVDpi+Y7mM1KrivheH3K4FlLfiEuMtiT8ThwGPfFHI
CGxm8XZaK3rOC83/+vAF3r6DGJOwMlnBL6F6JgPXjN+/Q0LOy+UdJ7OZK/1vwGc1
P7c9HiNBYYkvyvdX9BBNoZ2YWBAvBh5jYzqi4oPTGguUjzi1Hu6ubQL8jXf7E9q6
qn24TuWUceVDda6YUGHAeuymsdi40H2kRlvfByuYN7KW+jDNLDlFs3WCgJYPpAtq
6AnR1oiGiAHRKhAjeyEMxZLumlFLLsCC2kYqQjIF5ZcZi8lbwwB6Ju6YavbiEJdb
Hyz3Iga+hQZK/0zQRouZ1kSdG8dCE2SmOGMnO6EgwozX8Oz/e+VWhsAMd0th7Ugz
kJSbZkVoSvkgUS4l5mru0doc5p1yX1UKul+fkctcrKlPr1mOOho94Af2b20Fj4DM
0q0s+L+vpZni8oYN2bAL9U1ST+gGiyzZmZ+dlomxi/DXUt7+Chmp+IHOQ3D+RWgy
pin+mL7W935Ys5ioMa/STmNrMiS03G0W/OFxhZXd2GGdbP+dL0WdW6oI+fs0BLhO
VBRDTHo/7H3BMS/iPcZNdH3rvJjl2CxGtXL06beFK/9aHxJHBZ/0AcUQvqR7H/cF
AfDn+O31wFwQbMi1lQ3v4FU4wOqNkTsCQjYrTS02e5iEN3+AkGrKuYgNkwpvFhda
6PzHk9B2x8/enyJUIBflU8St4d9XIiOkLRbDVVLUJ8JNQqfuq8HiNdkAvkNUhQFW
wIfUmFCxulLwpo+N8dTfn0GHMee4lPxzXF0YPyGj1lgsGIhYbXV/cQAwhWBbSqGC
7PU1TprMnH+M5CzrffSchKueHnq5WW/OWwv/qcep6hrWw7DOLD+8WmTLCo6Y2D68
Vix7HInspGSos8LwIVNidrKVLJnwVWwTurHI3tZvdtW77bFPEnGXVMlQijWVKJbO
/0Vj7Ks2NRLkS/AgKJjqr3EKQF4mIAt9mhmrDJHmVx3fhCaWKNwcAB3DGiQcCuMa
S9wuLeEQX63MJhJ4TR0hOxbksQHyGrbzpCjXBCo55zGzGJ2ESajy9fgphhP3zWMK
Qjygh32O6zOoigoVb+w2hYwgOi2bFqwf+FRBiqZtu/dG0Bh0HfUZQHRT/mqml5j4
GnpIVT0VufXQ+Qjex2GxcrIci7aPlm5uwrfqwQIe80mn5l4S1yTw+IkhICXSWPKI
Mv96GirsmXt9ONg39CqWZBWNbHzUkfH87pjp0uVIyYYKpC7BIn0RTiynt3fY5A8p
66dfxxm6QEd0tgk0ttCEuv2xyNb5i6aD8ZLjacITGC+X3v7v4eQjBCMVSXi/+8ou
zfuWJdIYakYlF9QxpvzpGUm7f+1RL5V6UQBivSdVirrxjG3WTSG1LXMzQ387nUTn
lU+cjBsx2RKCwZM2/0/BY46cSQFhwBnlnz4zgrpfIZVgXF9Hks3gkllXpefOqSWG
zValfYOCP7eIIjjev+lUiWzAs5RuCVyNUBB9B8kOMIneBwPgg8XuBN3JnL4ax9uE
x/IPiBuaS4Pvp5Hvf+TLpcNHjGElidq5twpQqJWxwKcLceEeTJl4QkxsPpQi8ydJ
tXBlO5Pv4XwxDk3Anfk2LNw9zBXEC7/WqACI1g7mgx/RxBHGIvTFEYxYFEPsYGUU
uvyU+4Xbhuua2FOILJEcs7JX89gSN84cOTLo7mmFV+43nvXgECqSVDCNEHFK8MAm
bLgnW14WDYqwVO33NO8I0+oDZzOdMI2nNPYB11dAFMfiIwG7DoTCJbXHOiBXMINx
LqA1128B/Kvpgc0MllgHKaspYFJwiK0LGLe06WyPE3GGDNVgG7l3W83ePP5e8h9Y
tdGRfwSDuEIYIvm1Js3aVeQ5aAmffNq7RKjuUmUJ6p/QkOGX+lrWp5BMcu+y4PMf
d217GEPiREZIZ5ZtO1S9HGtcOUgvgLNBjS6V+72jtCQTfi3RZLH5irLWQ2WIBxgj
OhO8W9eMZv9oufw9RaKO9PQlCQ1wqt+5/WQDEXFz3cPa72sD8GXqvVk1rY7a81hq
CKi33klNkPTXIsy3Q+tYwo3jGVyfasomnI2xU1v9AAz/Wle9QSXfrWfyumZ/qLoU
+ikBDlGeAV3+M5zTsBOTI7RTnOrZwC0fYClMyEjLyEx/E/AER2gePgzFyNDD3Llz
/7uUi2cbcqUeGTqujGBveAL6N3roAsRyrqCxtk5sUoiCBT67jFtSIwXFdnuSPIIL
5iSsoZQLwQazrKO4eUrcuR2mDLRJFKt8SRfkbg9TcYJICtccNs9DwB4CO6IAi+yk
xNJCAyVqyzi8xP0B2OnTmKyHnxVpjOBr1VmyBE94lu+N1JB9/R0zf7bN4syHlxaR
ynKOmKhStSAB4oAYSThbKbX2HpxPADmKSazf5NoqeYXqS0IQehmR+AMEIhzkjVFU
EDbSNfYkf1LmBxwY6Qd0mcOX46nKcowi8HHWwRw0WHejKzpTuSWgqTPH7eHjBINM
nsMa7QhiCQ2IK28XqgRlrjbAL7fibnezzXSOgxlX9Ujxv+SChhkb1sOx07J4lvCl
wCc+f0oQ8LHIa0IlQATODcJqbLnFaknxLhy3gE1FcQv58ppzOEtMClZUQbZ/n//L
8iFZTb69O7gbcvXzOqATyhp1jyb3fEzsowJ9D8c6nKxTmC0LPET3KsfgU0Rmbi6C
aRQHRhsiV5BUfdnV/M02+rINGJTsdkzSFEFhHbGI3kwmDB2MMjAUt3YQpL4h3pUq
Dq/vq6GIwkKavKZ/aikC0blOJH3a8+Y0rgn850H3pfZgL0/9/yG4fQmL0UeGSjuN
C/l/2QLuDbsJYgCIInyJNYohmfM6JnlYu1RqP0mRatDajJCvCNFwebdW5D2hSLNJ
ngmZ7MXWTjPcKv9eHkbPzAqk6FwaEPZt+qjgWA7DasgmwIAZkKwC++Jnuolpg6Gm
IEMzdsvr2nC8a5ZLJOI2S9MYuRkWJPQyvNy3jZ+hKQZckDcg0Ufi4ZWkKvUkYqhM
KvcTr6zpuDpr3d/S0m+DpMqvYSe13s8Mq5XCxc4Eo9Z/soL2j569++/ajxvP16UP
q2NySiulR8d1gsdLHjc0mGTFADz4pj6gyviZOPzgQ43ZwIcq7OI+xdztfym7GBz0
eQUqLhU2TKreD3HD7tH35Wfk9LS9+F3NDZyRhDsDAtdGV7gMZYNRhwdL7im/1pbj
bjb0Ky0VsX/a+CRrfS56vvgDvJNk/tLE+KltXezVMBARD6Xt91gAIs8NBjo2MsDY
GAAOPYPd9WUa/xAzu09GbgMNgK4Bh7MGZ6bL4P7GqEyTIBoJAOWj/pYJM7zEObNS
HC0XAQjuKgJOqHS8fLqvfx4jFivgj0LonVuQjtFEpNQoMCT5Uw0Duk+sHIKW5sXI
gyA/Vz64HPoEzoI9qGhlitejHWLIGYvmzoEr2nAwZ4BQgrNNs1VIrxk59ke9fVqx
uJjxq8T11vqUv+X/YMsGP2AgxROZ6eQxM4miSAEPpn4eVjp0fFtgfrw9s3MX8RQ+
T6FOAel1+p/inlczmrj6uCB+lbFyhVx8z/IWpDHGE2l/pMspFeYKgL/yPd7TlROW
mdgqJw4wTZKjqHjlbRii60YASmuDC1INZspxxwa2d3Fo3bDIzd6oaar8XXNDAzo9
y0aaZBCdguh5RSJAS246QE10sslYWsFn6T2TpeZpHhKb8pvTzcTiYgdCc0GXq+Eg
5oUe9nUrRWRfQM7lkScc6FrgkzKK7vl1+XABwoPsfscC4RymWnxIa/UfBW7y7+bU
9oqVBm7sWEk7Bcup+3qJxHlbfuswcw0ZWaqqvXpPqOF9AX4jeEGJvrPcoky1gmX9
n2iKS42sF9hqZVxiopAdVKX8ERaAq71BHL/oqWP+fX14f07M/KfQJqcuSbzAJY+Q
NlVNKzle0b0x55QQy6TCp6oUlhGf21e8/lC1PokRllK+H/fIhtJRwAhoGYx+0j9D
iEBo1lTSok1ZChzCcpCGfq6kiedQtBJDVNfypdKs98Om/EkjGDOtmXqb4nm072ZG
BmIKmqx0vkslt7Y7ydGgvMxiltTsdHHMZGkznhPtVJu2sHpTqmIJ0B6iMibC/r91
Qd3qXHrlfNRf8if0qtCFoBO6P73osmmImw3f1/Xjzh3ntjQiGJ/b9WMxxtxyhums
WhIn5f9qpq+jKKkvFH6/adSnLAwB3+Q1BHta6r5S3cnd6W9cX82nihmhMxwrbS+A
nNsJRlXo2UNpo68c0xD1iV0xoNnCw10NyctKKj1uCIPuwH4S53F/vUddP2fGMBc8
ZP+GNBucpXTHef1LV7TxcXTDDsJ/+BQNh3iS4CZs/HRSBz9nRR5uUAYAl+ab+sqp
detJAiBr015lImhbx5tEGy4YapqJeWSRnOM6dn8JRTWdHzc3JcqnuxrY2fnCiu5M
eMAQ2gNbbMli9PV/RJX53EfIAvLQt2bMmlZA7VxY67+3pjH2nQfU7ri/DlRV9XPl
THTNm8mlgo0Iwgi+7wXF3gN8wiCW8fRQCxFWvnv/fxFm7HyEt/tXIKbNBwZX6Ame
Tgl1Q+tKhPjrLe62K6r0rbnwTyUFygqQF5GIcDg5+Hff2BI9jo5e5eQtG8LNtCNC
/auAY98STGAwG5ooLjYs+qiAjYJW2Yy1nJZr5JgmNfj5e0KXfF3LTydwYHwU5y4a
QkAkkwRp0vL0fdbAP38hZbN2n8wvw6CsoLwt1u5UzS5muq0CP5Kcz6TZVq1eEJAP
N6AeTeJ0VW3B+4IgetfYpkC/pJ9w3BrVF5CYiUvjz3WbG9ZYWzyftURNB1+CE1IS
PRtJBeDhizlTnFpXHIUk62SI/9Ra0zOOIuLhPSgwswCTw/VJyIO11z227IfePeE4
fMeDaNdB+OSDv3BPRN4y50chz5TZNHdJLLmeTHG3V2oevxnps8ZS1zI0UnV6GcSJ
AEhl9AIN5CTWFGtvP+MdVvZFD4zPHABweSSxUnrs8v43rbFpGu7+SYNeswldxWD7
b+igNVIfW1J4TIjnwz01TUrYXy/Wi3Mq/9lqh1ADN7p+Ap5oK3HJMRDzW26Sx7fg
R5XvhgC9Tqd1N+58EZqUUAdQkOW1GWw7Y8Iyo4HQIT4LpXedfwBq05snaZF/yRiH
v4klmltMORgeiDRyUgxaoHJcDeMckDKW/9KideSiyeIvSvzp7m17aHXBoOpShysP
taMyNzjCX7ts/jHlv9AhVyq7zNJE9bLMxv29EFUJhyilNLNB1jjobWJ00cPTXFJ0
ZR7DXjledbZdGpXwlnTF3uYEq8r09pSVF5g85DfFK19+x6HWGPbXH9ohTOGpeh5z
SlFiB3Iu60MxfgDMo3wWFX/7VeybeWl7aNnHYYpobu6HPwKwOOY66PRLLGMljY/n
za2nc8/Nfw65O4uIb33X61KzXnsUHlkLtTlKtVBUEL6rwUsU9hQE+J7Hbt57T7LC
FcQqW0V6LQrvhweIxNyysB4RrscAhAmj+hZA81c9CWMH4n5UrTHQ9dGGu3ZDRGN9
U3EAjZ0AHjieLd96XUQNSXMUmh5u7RAvyRKTYZOxICx4ddaEAV8EvduiR49ib6Gg
glLVuXrLgiV6cq15L0/52TeqLmdk7LLcWwqJ188W4ZTtvjuiT2Lzy/Rj7F5aVKuY
WRn3PLUKCQYhc9gBYwqCTMga7OBN8GmnD+8Fy50M4zRwlh4Ud+z9JgK/A9ASN/cA
5jLuGLP/KqelMTkUY62rRu3Zzs4jgSBu30uRcZZAPuUBVZG9kyxvgNX3/YSl73RU
gqcnDHcmkp+kuxaH8UUq/Ja3hP5X8NVqkFrISyxe5akA2mg6LWD1orMU3YyKMdGv
UrwG8m3avHAcWSDipZMi5RDSi/pUzEiAR9To4wCzzFphYbXnWVCOaZsldkE2/BmW
AV4cU0iAHjv9eM2pylO6V2Vf2eLUM+D0dn6JQkkEt4q4RMAQ6cmxq8W6mdrQ7Ra3
njALAJy2HdFlk+L8h9vQkWNq41TrVNW0PKJx6tSDnOcv0GtPYz7loAmpvhJ1//mu
ckF0lMwPP9VJpQDK18MGbZSGJrX9NSnIulBry5L2KDMSOFahJf3QwLWy0ZHGqDWL
XpPcZiqgerxwD8mye8rzUyGB1IlvAbvACzuIaKGgPWxjyMNWI0Pr90JDJuAAKcZi
u3bNM5hIht6wVnh2zsopO7QvrcDdURL78PzpLCecAqLQGq1DBhhcrMTNIm02TIbl
lQGL3ou9JsbyvntDgUexFuOewZL92uC/5r/gJBJx3f+AV2OGhr/1RK/V1s+1+yqv
pKDX2foocUDlVDgZ16ssiW2vFtpMG8mBHWKmsCuo8aDGCSTKr4GkoGvM2uzDqV+y
LTbKJwfqBbkxzCt7i9qYiC9TcEl/GvHj5RVGwhbK7S0FQhazUGrRY4sxNIPHq8nZ
8b1zqzAJ98mho0MsAWpQvaaRvVwb4ozQDffOpD6jY0hh1oCamU0VPdoFLhZwIXDx
VBcEZqy2BEW6Et8zNnQ7q8pk9u8GA3IGdrXYXmCuPOoQJa12wwb91Njf8+lV2WPD
e+XBDI+EOicTys1HupICXswI13WA1QhRj8ZpfN8wN+eoPxjH3F+C6Le0uwxJ/aYH
BGJdSk00lbUb8cnFuQwffxb8r0Nkf4UAPdPha4ET+Q8Hh3FN76Vrn8w+1vXzvXch
nDbkSiwPzUB2qNtXJtEWVJX7ygDUIzcmhTV2dYVvsvMtvu9AK4/+ApTdL8sPx8bW
mAh3n0Yipzpso81gYRlg8uBza7zLeICt2IsoIkrpyDJgq5pjMmQU9WJmebJQubfD
gfN+3zHUFJnN9X7dvKMwC3MJbWQjmonunaIhOVQYFRcQlV2rsXdkxIJk2NBaYn49
erpacuPmdIX+/cSLHH3nU9VFC39Bb/larN5dmKYwYziDG8nz6y5BzMrjBZtjeKcF
WIwCnj9MOqCRS4qEIzSe4YG5tHAGa/d3KjeTT43y8UfvdL9EURgNHzPDLars1iLq
dWW9gL2lrnwSo0uDANDZt5ggU5z2t2MLA6TUmYNNpzmQXKd7kRMs/3xnJC7/vH84
yp8g9h3iX9FFerwxwckhzjUKIVix013LC1sm27JqJICjD5tXfD1Atxi+MmrlbBIG
kd3K0Gsf3xmCBDBQ/LDVwfrNlZT6GhIvg7kQtHqHly59dTAzr2UIDDTb1azUvYkt
GkT9+9H3CbUoWaqsI/EIE4ayFKCyNjGJWAdzPj7BYEKOey+zPWFTnjuwJvM4nweG
R32bVmftJaKfj+NP2hgffLbpHNo/0gumD+Bg6m6gJTz8Wo1Wx2ttEIzYiNqelpTf
5w+m7Hcg4IJiiSDb1u5y8M7zaU1r5lTO0IoUz3pU1jtjdtW0lfsEe+zduMsXDY1o
9I0q5eJEZYZTYD+vGIeVNFyPUmWGb8N+2FyZbD8/vuwCuwSnNbpMzrqlt/WPQLRt
0Lq7ajY3S8StMXupaI6uJ0Mm4QL1rmlNon7uYlrkGeYwqqxA/gGyhKyP3tblyCFE
jscRb4ZasDPzGU6UnNt0tb4LudlpiCbMiLblnnpx64CFCGpdyjXoZYd4jI8E9203
A9J7wzZlRZ4oHA6B2YydjRXLnpVBbm3jr3JFh1BOcLheFkD9tX/xb82oQQJQZWFg
1rYns1y0HKG8x53N7nnyrOOeqx1JyYEVYxBiijzYjeCnDNjKlhuHfcmL9HWeUnLi
BWaR/wtIcF6V/Vu7/t2Lq2A0obcms7FEPDoMy916LqA2N1mWHKTZ11ZTZJitfN8G
ja8lSoEN0PgnoFUG4e1UUW73+ZGaUyyAkT2AuTIy4BlRb8y38xKStj84qaVuP/Fn
hsXSA4e7/r0cfbmVNyqZqgIVaG6qlO0ltq2YfXeJ4uGGXaNCzAzAjBw0eFzr17Pl
n96Nx4uT4y0ptePOA1OAi/WUt+qVLUN59s2QIactYthyTlgzFrcz3/JudB0vbxze
lbI5X1D7SD3sWFbSW0OoMtpdTNOMzhLStA3LZWUQ+YkxatzCqBVXQiZUt7AcOdNG
EB6fMR1a/Bgv3nap3hnla1s9L0N9WCmq9djFGJNcdWfDK1oR9rsJmih/w+/G7+N5
92C9mFS2wj96ShBydA66c9OGB2h1JfrXFOAYnDe9mR2YkN9dm/oFWgvlm76THY92
0OQ5HJH+P2z4wO1V9Fxtt9VIZiw7PBr3EeLV0/pn5ISl503xFXxykgb9ixS2wDEg
sUECgoBg+WhnOivKT8azJFs7upIQLcNz/Pugp/7hEw4hGdAgRNlepvEdGQvGEDTZ
VIWTS5XWhy2MTGXoXGTHPEtVzTSJCUcsqAh18XMpLP0oW/CehHG4ocs4mMD1upKE
LctrjjC06ic3FqTNAZF478c81CAgWoRgrdAvkGt6oD6PCSzXTsMq+PG9vfjTibEK
CluRvII+g28H2UZpKjNudztIDGizdban2N31jdDjePf6753tb/11sZNu/Shlvr19
xbhvdpLS+CmrccSoomqEkWe2uoqWLJk6jjcRI4LmfQZoXG4iIksK8hzSV0AMwxR5
Tl8i6hpr0PaWAMJaP7pTEc3CebtA8fi4FO5vpGnEGGUCuSmCuy5zs3q3tzO8MHIC
ulAn9MNi0Eia1juDqwsIJs1L89cc/4yC69fT0Uw8n89q13BeG3YF3e7c8szyoU93
hAPCDD+OXbIsLXw9eLedymuUaALxRw2zT8Tw+8IVL7adv9iV2tbn2pFG8GifZSHP
pt4K8Rt+8XedYwI/hTTvPosnBUFZ5LRkzU99lA+6hFkJqnkAsGcfts050ciFUzqs
AoKyRr/VbmW3JBeS4Ou5HwGL6Y9wiwBoraW3kiSpUfUh8BFh6Q0zd/lvAxuwDJYT
Kkv+KLW4UVi9397sKfvsAMqriYLhQmHwp24jblEecfO5DbW7mlnoSWyVAsYjbXFE
7f4/8gJMYoX6vFbdQk+87Iq22AyX8dj6ibx5AvYvcl6Ywu/xNLsi0LB2HVjv4rri
ekgTDHI69G2rfiX/jPUmPZz2No6CyErpMuUbJv2X5YSl9CgZgBMiywvpsEovUk/Y
asWamQqTziDyg68NjbQSthtqTOTjPU1E6Ai/a9067mGuyIpZaEjsdlXzPlYOzHqv
drr6XYjeC/z6MF4cM0KtvoMQZfoauPkqBoU3Dm52OBT9wkWzddd4QJQ8IVPYYqbn
fmKio/TXA3HiLgIB9ZTzTH9pE1T1E88K2S6UwIqSvzVSTI1L9NSMKST7Ot/ANT8j
cQjGuyPrwL8HkJEETF6ZoHZu4K8XmHMK/ehYX0lUQsSBBy5fRCMg8wnLUCbvaQWD
GV4g8XuTKDWYEjw4iO5SB6euh3Mm0ExXUJCO3j4DA75sV2ZrceYSK3eL3oryn4wH
nY8o1MDFAvGumH1bT2L5Lw8MHVeNpr1/CoyCHq2vIQ807xTGqv23a/xd4wg4kIyS
EuhHvvs+boU8u6fVPRIQC22gl4d6RNwiqfgrY4hMkJNdTijfnACe1DseALqPHhAS
YUuSMEdRXxJqQg8YeVCIYZyUdksMDiQ/nueCJwRkCn1dAdmvg3rrPecuC0TXI3wm
LHZEm2vfQLUvjumdZ1OjdGF2/ZZL+FGGs1v3jSxIVFKGTHskJ2pAvsQnDKLFhrzn
R/S3k4kcO9S4DlvE8mkrAloG7FS5LxsEJHIsi/uYr97+XxH1RSfEpUqh1Zy+UiaX
yqyjqkiCHThgOCGpxgzos6dSAPXe9V0Uqtgrme71XmqbA2E6sp3eFCRCsRB7PsO4
IRwt2ItFTwcA1rU4glBhCEHsDhAzLTt/Y9Fghpk2rGRyU5c05qA4DlFCqIP9s3pL
5J5tpEQI752bKtNjQYvhVLeeuVMxB6PkjhpxovxqmTMvTthjf0Mm2FHpf8kMxEDZ
a7ymuORcT198v5QN1UFcMWLYXiDzHKRCwGJSN7t6/DA0J5/ZOSYqghX1NUxuDZ5a
DxNXdDjtOLiunhPg6xzgdLiS7m/UUjfdC9kRcKgd6GAGZ0FD+FIx/R+G1YgedgQA
zpZKf0RKFQuKOKhhPBwxq7og5NiBQle2ElPlH/rKC0poIA2K12LsrPpTDQEDFXo6
5VkziT+lljT3DzqXpQlDOHErhHKgFeebJYOcE9FfX/uECge08SvHuvG8/kGue8F0
of9ZLlinJ5XAqJ7XkNu1q7iq43/XVc45PvMJRCZHjKi7dLNoXtPnsRY2tU6o/3V+
p+sZ4xIaJz6qPDfs/teLjc/3vhYPepIv4D+T/XwR6W9vPftnkpLpfCI+zv+83fp4
aqXJnA0aMP03R+32l75Foob2w6Zb4LpA+Zpxy4bKdyitInVO9Q0oSC0/F5vtDKOi
EvUnPi+k5UNFqWMr1WlVVLIlIOh8cSAtoa+pYk8uWR/7BkXuDyHBncTr4PPMrQ5l
hV1PNdmpxv2YwrJGUQTYVPSNBzsW8b4I9BXcz4qgoOGhJHiqkV+oxzKGDq+rz1Y9
a4BZCElvjnRdbIDsPaNPR/G35rw9JmkiIzuLkQa2nfJPzniDP2CGPsH3jOE6weJR
wDz8yc2WYf/IYl1nnmwAQEWsWrvgIIvwotEhCOgK6M4CvvbUT7HLv3F/Qh+C3Sa3
JELU5E8NDGRzIgnia47FKSDj8GU6+6T6u6TgVYtgvwUPBrrCVOna6Z8DcM1OpS77
N/fZmEvTSt3Og/AzKXVK1xtiX8DvbpY1tEOiEbduHSp/N+d4cwDAIhGKAtJmYAzF
hhBDv8HCRRk4VMT9WGZoe6vDKLCoVi0LqZrXP7U8W2YFbbAOJesst2eddgObMgZF
1RkILBMLeYb8y3h+ReyyyxMi+sExCY+izfuTNkg3Do2BDcyIJiF3v5BUQhpEIcD9
nMmGWDir+xDm0f29EXmNXQH+gLxVtMcgtZ0SStRFOLh7aPjbalgRvR4gkaBr5w+X
fJ/8cY1AnCSW/GpNSyHtJ6fzrZQs7Ad8Br/HVxf1lqNs6xi7HkjcgPdzUoGlrxhS
2GlRKYdQAnVzgRfyj41o+qOYR5ZiqomMIhfUIWTerh+s0EXjTsZ5XaPgKzFqVCgh
aJlfppSGO6CDmtTeS0dBNpNMWqD3FJI25Z48s/ULtbZtLVhvc4Ch0pk56N2ByqlO
d9QnwxMIJgkGa1QhA6x3S4rS8F1I6fxF5XpxVTziistZ+M5G1iCRnej7iQXwGY/X
25GICCD0qFCWNwU7FG6rjzDPUtT7P5z1C1+Zof8Pi7Qd9FBpEqEXElLaqD5pnx0g
LtZ8zr3s4eYokvLKvuLswBmFOowppE9dwYkgMN+u1iD5TTj+LfWicus2ggd40oHF
pM7bfmLiwK4tgnSrj1d9y/45c0fuIBLfG+I6RZVCk1B6OCNIvXpwdaqyjpuQDtCs
xFMliNeAgqUEZkYYksSGMI9vP3wIh0P1peL9M8oe+BSGT36pBmqq/4QHAbzXfVF1
rWpEv0WVi62e2vOEJ1xj9jYc8S9nbN5vbj5Z0dw3dpiEyGT6itWVN5rJJu3ct6I/
B2gqVWuJ5+AK+5RWMAQd5P7KBUjnCbYZX153eNNpWOVPBGX5FUU+ohP4WHNiBw5u
E+XP5YBdRxrsVm/QbbuSy14N0LROpy78r/DpxHbpuEXV7rl+GuiujLnKOht0w5RH
zPkNcq2XY4QA7poLiQAHLKNFp3DIy14nZDNzWD7LTWmw0Erb/oOGoRSAnMK9lfq5
WYVtLnEzuFiZrlKJr+7GCZYLNvMeE9YlPDkjm7M2+zs0EDI/AyMt4cpm9nMdJ3ZL
OlXQ6wB1ln+DO9Zdhx35vSHs+eum9Nj4UQ3zHzrIgEOif8GG2vjncLLA2wJOpSVD
6C7NIg5dPc+pZ+Cfvz9nAyiT62AksluXGlEFf2yRIhkvmjeQIRtHlbvUpOqxQviF
76r64heOjoaGtHrgeYBBVsfzeiLbIL5UKu0Owfo7h4gvX7LEMgXURqcS/tjGmL4i
Ivi9H3qiTOtCNUCSjkroiJBL8wVDV3I+R1X+n97lnj8hCGJF7XXowt3XoWzrlXAH
cRZyDsjww7lKb4QBqwtFZyUcLsrej8OYyKvDMspiD836bJeXOmDtG+sQAuOb+TRK
bDLBFiRG7ZAOaOg/JjlP9Aw8fuPzC6jeDjN23QCBIVqUX9A06T29EfRFmW/yOgeS
NHFANVVUGrWQTfNYIfc77btSHeBDOg6jmbqs8v4SRydu0ejy8NVcceuLzO61HENl
+leSSavTbKC2Z131tfS8Pi9UoDX41oxMJxBu9+DGJQy6e1o0nTeyxZynbVZCQPcH
Ue74E/7Q3CtGNZx6skQN3QtFQtbPr7q0nRfg9iTgnWOhdXYS9EZNg5wJ1CxnXhGc
rHA+uv0+xvzQkOyWy3oZMoECoZjqRi64CEwdGrOO3TKF4ek1kcnm7G/Ak4G5ksUv
1jSKirqUbIWooq7MyXq6xhiBRa6fIL273NL+e+5EvSMUFHv2uzKOfk8zO0nb7y6B
s32PQAn0LSlvppa6f74iSo/lmzfU5B6+GdA19bKWaeHkV7lGDP9TcMop+HOFlzO1
DgCJcUbzH0/LBWUZdCaQTi+p1L9/PG/NL3wCX/pTitiuIvlPKmnjn/fTraeC9HVp
mR4d/XW/er30z+9fHuZEJS9d3LiW05/g0hJdD3gzTPUUvakXVxar7bwDFzrS67ce
MLNkr+gBSa+4JBIh+UBRswn40zADvmqXhcZeOsLcTqdDRm/R5lecB85VIY5LzTLo
HleTwCR/K8wIhgF4XvZvisAf2/+wnZLMpxCmq/51rL3+d9MzZk9yiRRNKXTea655
FP+/lHH5+hyr7NzzAyjBTDgbhtUieKGyWAFcCCjRMgzZsxAHqru1LXCiQaJnm5tg
FER9REs8HNCB+ixaduNCHZ5xl7A3J9YMG2c4GB2pL8WdNdDRulOYVN33ktC36vtv
g+IUet//HGHIrweL9CIm79Db9cRItTsaWZs5NcOVdTA3j3DcARV2Ov7nW20QTf4h
+dE+c/Qsw0vQcy8GSOTJLaBswT1HnY3hpqfRe+Hu/nS5IFlTnxgO6bDd9oEqOOGa
DJqPfC3PRKYdpe+7di9aFkvOtui6sTTudlmEQq3T/7HPedggQ1ZMxp0T61hkmbx5
zj0M8Fv1cvLwYb51hqrQoj17GuXWjzj8c86DzUslJncSLaHQxmNd3DBjKcgeldPt
6kQNtUDzcrX1C9wN1OdBegrB/Z/+Ll+Fc85bHan6VP1i4ZZh2KXKuFC3OlnWkx4F
8Hcgnzy6YnnvoKzfyBXs8QJ574r+rxDPOteDTXGeWJuj0AT0EPfDQBvc1SCtmPO/
eDFAat6G+BhKMIN9cMyt4KEBFiFz5g74VNpnSGDbJ4O2asoIGtQgneGcs7KqcxvZ
oWY1yLRYkjbk3f19X3qfHf0wNqAFiNF/t5RH+Wacu5QVFF/822JgDTRdkTi16JqJ
xThK3KaCXbYsz65Dy4IFGpNs2NUgsuSQYDdRVJAB49fhgUnE0zkKTlbXgHDMPivq
R9H2iDivtrTj1jjFm52/o3bKFUcGnLdu67UM43YAR3aUr4qZ0CQQ48Qfa50OfLcR
oTDTHnEybklOawwJ6W5FJImsSmSk+2ksJltBxIW1CLxi7DCHfZdHzkeo2FcYHwvw
7DwU5nhPk/ueoNbloOIcl2ge0nHI/4Hw8avxGiBSsThjqCnlW9Wr9dVA3xFPpwF4
H4zTbsUdl0ch59HULGjzcKkqz0/+sWUoBe8nfL82iySoypxiiPuM279Lpgj0oP5t
AP9umlg+ef33lmR/WbFWYoEiqJWFEyliw2eJBNMPRS082aoalpuo6Eve+DK5OxFt
LfOUsBSxX8/MYoUEcUtT+am+vLSIRWZmlPKLfQ9dSi+BOcxAxZlTsRXhoKMCuvzu
+OIU0xkA/MxFkA0LgYkISJiPETSFWGPQ5P/yDfCccI+nRcngB0w22UhenmVxL2A6
BdjmKoL+0LejtV0XjWVH4JF/ZDyEOYWUAQtQdsOwJtrUNoNAXdxPP2FvYIAfWu8E
znWJ9y049SMHhS1bgcqXDLd0/UwdAIigcpwBTkxcNFxjbr2dQByIrXxdiq3VT4Po
bOc5faV0NQ7IJGKtEolL0I+C3C04ytQZ4aOywJf8CLMPnIqQFmsi5fz5VMLsy/FU
QTAzRCo/klPvUG5sh2TCJ+z6mXFsRE5ujVFy93VMulZsqcq0K9iZPVANNEpYwbH7
VnZJUjvwoRCSW1DTDueAPFcUM4oZIS1520F2HP1+ogfmaecGorlvAcJ4RwflB/PP
lEVfUetk3+oymlL+RwNoZ1wMnRpbG/wtTkUCOUf6ZubXGghvDeFAgmqxeA6JTChd
28uTSQL6RyPyVh1aU9SvMkZvN0N+2yz2zXtg+4L5crvIJG+kDJspBLgoexGurbf/
H+lTNzB0jeVcF7iw0+qJvAm+6B5AH+KQ/3oKiml3uf/6kZvNuFMAVnDtfp8iREmh
Th0s0cMJQqsqg7LHbRNc67eB9Hw+U4kbzJpcKIIVGot5uG9NubsRZPbcREd/2imR
/uLGm7TuF6902BPxd2KiVtci5xWq0FTTJdLwLRnPrVe+yMepxF2uNTLok73kUjpu
R++J0/y6/nR2PMOMYmbXpYoutoIhV9J0LSiefLTW2RAXYkrNVs5ttT6eNTXMo4+j
2jrS8OpdHCAthmaf6HzTOuSK0B2+WTDSqBEKZznah/dt7pimVitGh5shAT382PDt
8fqreUvHNj0ihBqSb1FiEXHz/1EtxqO0OfkCy7VWEl2KyWg6IEQZpsijn3qEEKcK
LBNxBjRn5fqKNDP8fTQE2R+OGOxS8JREp/gHf9KygJRphs0jXSviP4XL/kg6x9g6
8X+fljX8x6HaExS7/CylaWf8avTa6ym+xFGOLSAL4aNaiEQwNDrd1RCGkfNlL0QS
UnOYSrm94v9THHt9FmOUlZsF4vSmAxjs/tPlNPt78VCuMSHWlUUB73GOJCIgh6c/
9A2duqKHaxYdxBhS59+hxFUxsHhJYuPC4e0SzSjl8KwnKhLzGsxDIXiUUbPbIJQJ
Oame+sbj39qKEJSzrXKUd3LfHH08kx/LDQ76L29+qHJR1ldi94OBzky1W1YBux1C
qOf/U/61yC8Z/YdTelLKt1Z6VjFyvJoN/1l31M3MbcryCGmbcC6dDtfGMhgIZMcr
G67z2pju2c0u6L7Ly4nLCzpI+rq+b4XVu5ucd3tBDVDsFNGufs012LXBRpnw/dOx
U7nOi0t3VB39U3V1qAci82DrTZpFK4CqCU2L+v8LPfE0wtVsfcrY8YkhAxoS+mlT
s/VB+uDIwd7S8l91K8PwbRRyJy847GSAEQ3EJkA83vmneemOcG14UR7dWLeap1Un
rCTgs84mhxvhQXKeM1UB04xcSCAAx1mKUarIZgGo/yucvUNztuhq16LMtBGPop1w
rAvpRA9lV3tj8WuWphnJ4oR/zZhT8NI4Ev4CVFSCbIfPujw1cwvn8GIoA2sJIsJf
wtOb56IJnFCDWdaNeNNN+zdiLAtT1YDTSz9y72qJotuwy//KONgoEVEe+/G6aqfR
GDBmwHsp2hNpYD9klBBj8xP83ANwoxQ2mYUI0682l4114d0RP8mCemDhol7BHK7R
27YPewCQ4ZuVatFp4lkCKFgyaQtghUvkBq9WWcGdc6PlMh36vVHCeEznHzJB9amz
1YqTwPZ3OHj5StiwDIDbwjDy5AZw/KcIRpXtOQK3XOFjE7qd1KqPm82lIwA1Favg
3mBvT17DzJP9ONQfcHtIPLzKNikr+133mK43uujsRI5eOq1jI2X82oqjA0SWf1fm
RwKbDFTXjcrEg8BCgoVndidp/DzhuBf4tQFWEVhLuhuQ3POowiY4jpmvDq2QaHLz
Lpum1jS9cJxAyQJS7lUbbqbaM7V2ACmsFbVNzDzmqgESdEHYgfue+isLxAMUcu0Q
to/OLcI4J4LyE1M2Azw9d7jEWrJK9YG50QKSiXQrN3oO+Zpd5voV9kw5jaInnX77
63ZjcMkcRBkJJARq/2hd6hztqdnRUXUI/W2WVWr9jmWwK27/v/Kjf4VVuAKljTp4
Kd8TEFYVwOVR+mO7wRLCOspHqL0LhqvZn3OPBb0r5znpoW/A0OOa4EDA+T8/1Oyy
d28GdtbfkC0JpgAWgsWh2LKX/4eWv6+OT3mhufG2IXk+lWZC7FGwgew9Z+QpfsBv
b0htm495VZKBPGJPmo7cqKAY4GOPCij14NgZyw9VYQZpBPh5NHJNWHmR7XOeXpb7
QA1vxzHz5xJ0DGBPUDw3IW9UDxlTWsgA+LooyUWdtL3mzpnmfR4cGohOn910ZiX6
JW9iEEAmst/SBDDazs7Z6VYBIiTEPsvHMee/mzv8IiYfo0tMWpbqltGBNei+/cLM
3UpRyFIdxIJxodPLWwvIy5q/50bFcs59JJrDnCYS0B/MaKPqG46XOywBBQ9CmLRS
DH8+YAYu5t/RwY4yKXVI/G2AQiIDejPdfAU3UBmd9G2dcqWDEni/4gtuqxwdoKxP
/I4gHIzVTH6A08JMD3oqKzIK3qSVjH5ZCIcgQo0I8idFcvm1Fn+/5mkye10EI7Xl
iQfbvjOj9Bc4/K9JL8S/phSmNpQvAA4QRrzTD3nAZuxcuBnmugF+CFQCLyyaNyYt
gQ2Rxp663pxwsc9g+hFHUydku247ibNllBG0rryMboNG+KPfaPJInPGfkt29r/VR
Jl7F3iB4i/+kklzoyidWOVzPeUDPLECDPnPdDr86BvU0rDt8oFeE8fLcVWjy27Gd
vnHCOxwU8P8rUp2SYviwDysgssHk06gYX3cFxcSTzdq7xgU4hPCx4PVpDKQo1P03
VwN4oiaqabweyrvCBjqdpblyujQzAKGOeemqcEeUWPiAXnRF+rD5pnx5a7Oq9Vyw
0YF3xnfF8Vxf1CCM5l81xlQ50f8HmhOQ2tsIF3jpeSjZ3RNpovb7JdsbOEroV8ky
J+ytCu9t03IAyCAAFp90g+qFMgF3Zfh0TOeaOVIl3HQeZm975e8f5DrsU8VaIewp
6GquVUDVTMumAzn9a0hFADy6bQM8vgAWXqwr0Oo7H49OnbOfERmaJvX2rGJfnvsx
dIzsiym6m2dntz/EUD+N3/WaQo5O1tZrqZgcvt+jSSNpyIDpBLNJsVOIde3/q76s
e+52OFH14Osh+DFZFN5x5D0QjJQGMUrIJjlL6XflMydnH5QEmR/MTSQCYrKOxxXn
cQ3CI7x3IvAyVbtz7sdgq4BZBJudLy1z4Migr3pRn6RnxuUd4A+DUVW7h28wf6Wb
1GZtMJ7OESlK0fM9ffTdIwPZtKmw18AwU9gMM37ZRZTISaKl62TTRiAsw0bIpR9Q
3G6JmsN4pxqOjlTBb4tw7Q6cbnu7ajRDzUI3KycJDm7WSsMv/aHA/2nH0gk1ljOL
Qas4KBpQ78NCF+3FHmjWlCZriwoPaTFtamROxs0FZgWIQ3eyIU92h8wCJrmmIqjJ
igg+87dbwhulgaq81QNfJxFmoGt4apV9U7G9fDrupezVuXvv17qMYvXdABaXNfZN
sK7QBNwokEAOD1eUcI3kXZLPJICCZduigMp3BqdUFTuxO7xImhlRPx6EA1NZAHHR
5KK73waDmnytQC/GFSbFSg2cB8Ks6oKFyLSxVEY2WeWIWQ6KLJcUOe2X9fez4+7k
SMQbuiZ7xDA4PUv3DsHXQvqzeFH7R2g9hmggTUvYSFoqdCy09LGBmUWdb/MSLb6Z
7OT34qZzue57FfzpCSFDFrQhpGZYULhJlJHF55jH2Eq59nYYtIORhZG3AEg5AAf3
upeRqskNYCnNfg6DN7jcatgrZIhCr4ipiiIEXP7L1NmC6ii7+Ro7tyZ7r+eyGM/W
PvTu7opOkIRlt+t/OepntGK59ILvPkMp4yg7DOAuil5HLxf+tGnHyqZeCgXv+X5p
Bq+aVaOhiluqai1tRnC/esjdQLZTs92pLuv5ic2QiQP9K7vm6Hx4QqTABnOB6h1b
dKMXhGYQfKitZnZO8GVT40c/kiJdIF82tHiJ6Rr3GvBLyGn8z8BD4BxuLRVfnOyL
RBl7m52X3n+Y6GGCG9UdyQcdiJEM1TGXjSCjpawKlW4GSlVvFfQiNmD+Hy7hB4Y4
+PdI1z7UXN+BmgoMCbFvlrNuDWFht7Jj5TRef6QYwyGMcKasSin4E82DfDXE8HD6
vK1yyNgcP3DtptQzB+v3z9E2/+miez6u+8s0MSuWpU/8O9ittOfDoHuwbPlFu6Qj
SXUt63T1imATMQqGcyhB8v7vLPQgFlIm50VJClA6Jol/tEYOzVvEFfpnhz5kRuGD
2tEUOiKW08r7MLup3oFoZXy71YlNPBVyghURJdGU+y+JZtmWLJNAGXxRXnL2xoOY
TlkfKmrqpGWYuBzgTyNaiFgW+W7CCcRYXMp8IyXAtGlE6HWtRaHAGjzi/Z4BcrsR
sIyphNEim5C3wJG0U6NuxDaFhZKOZYbNVPm7IEPU+9GBEe5twK1NFocHaMrN5Feo
nMbCGVSH0JC/gMdzmIU67sQrmZnM5Fv9imfTQg+oplYUyZvFm8tCdwxYDwHwdafs
CNMchmnVq9rBnxFTT3g+lpUVfs+JJsQRNYVdl/dJ9UVuJNS2nytxB31ib3kTLKri
6FTF6qV+Sb+BJioOT8mzKF9g8SSOEbEUB11Os7pejMv5a7kunt4SX/vCFnq6Z0kQ
XY9V/UFHpT//nMG85pbsHFwyn/fH50vP64165oYo6bRS64X8WeTUMTH7eJ8Jask1
C31joUi09FPld6rOFNVjPSaoYrBGS8/Rfds67PuJDFsorifFGnwJvRsAHUhrl5ar
EcAk0sLdqkHHnMKFb5lt03CGovcjT+tZ63BX63iJ2nv7MM8IgNIv7FdYCw9rfIGK
MygMubBTajkPYTWe5Okbke6GXRiPqUPTX1EIPYsEwBXcGr+IMP9OeoBzFMFx67mU
w0yQGSFta5ZU7PqOJNw6yqtT2wPW3wTXSuDTNgLO2N3MyskTJg5BhyJ1Ly1qqvhg
+ZFM+HTJM7x5xqgTtiOC1uBIrQICRXNGcsLkZs0/vGBfdi81TKmgLoF/iLlfGmlp
fmpKOe+y9jMzjC2jAAKIBFY4XjmYB+rjAFpdJww+tUABb6QpV7eYBO04pCy0ryRE
s5ZjQ0wt2r9bnimB7iZhbWJ7jmwImd/wgUA6DDB617YyNwCeUr6GrkEgwRoQugHP
p1SV39CqSNN2q17UP37plsPtC15p8DwN8UQHhybBl2bmhZKHPUs+OEgI4YlOAWrL
/5y1B4tcRibMCsT9XPdNlxEWngvtan7tvohuxyA+sor1J8v88hrc872ZxgTqAwfZ
tHeJBfZ+4Ns7Lfue+TxpBeIkbrWLqSYSVjSiVwKojr8Rj/y5HrPf+WUQR00iJxjx
KK+2L9w9hDDgf9+FvcXdZ3nd9Zj9l40z7oQzzrUNJeH5xGlQdANdgNMQpD3Iotd6
3rdZgo4+JewTRQu5bK8kaWEtypdfdcTN/VT9mJCuUQ5ZVbfzDfFujZGcP49s6uzw
7lujVf76M9mhNML5rhXAyVsDlAUjWuajAxvZUbPNgoKA+zXhzJG+91SuuxJAoAyu
PxzVmdj3p3lJ86VKde8R7z7iK/gbKWPbKcqjfXJ0jObA0jm/79D8RbpmZL4vOFPn
H+vsxPz9uz0UTuFNSmTt6MgtGdbX2BxzAVj/gEKmHwjFD+yqIEAILjmzfcBcaJXj
mHDwPyBw20ZVK4yP1W8ibhdUk1Lbg0o/1R/o+ltSxJvQ1g/xdE0pYNJW+JVMKZ1C
w61cTvR+Z9L+VJXJtWEBznJgrZ7mGATON6nL40Eq+Vl1gDmSesXSQEE01+UVBJJN
UJyRGHcLW2uo8rZbwNuXl+RyTZzmTFTFKDsAntJvVHYyvBtv9pPwPSy1PQWknMBs
eMIwew6eBV6URou6WU+2LwYS7mhnQ9iY+feBZe0IhhsKyOO3f/0UrSXve51nUsnh
JVkzmCvGlx4d05nmMNuZe5psVxuKtZDqPkUKdl7uayBxHmL1d+bnuZeQsMAMkD0m
G7JAv9D/Dbbk//VPQSDRfu4+jorQLL13rdP4ejrTx7+Gf6hRVV2cm3HxKw0TEu9y
uL88/2Ty5ZXb5ZvTo7frsg/5szXRMxflUuZ1ebh2AhP7s8jud1hpUYBO6KZzejLp
cRqXTY8IBVrnxo93r0IV28BgbrIRbJnVUu5BXHvvOJwZ1geONQgnpYcLGDjlf03k
jMg5zMye4a+gTVsXKpObdr1No1QapXsOvQTnuzcAagoqElhFlIZtceig5yNCKEqW
vbJYTF+GxbP7Jed68OsfNxYXgFELp0zjSk3EdGGJ7s206ILFeqSy+ihYR2gaApF/
pEuj0wGDFubj3nQxecWcRr2oDAI0VAe1vBUZZKGFGACzul/5OKHt25JUJGqsqIJ+
nqVy0nGJNndL5lPUZ1V0GRJdt9uzb7VkgztahQXXCj1NWn5knzAjeVyimRvO0Q2y
f4NBlwSUhYurhESQdyPX/xm+RYdahPWF8PDaksMliObgS6be3/84zl17hc71Wpkr
rt/macQf6WkOEgMv+Bqqc5Dlik54Zlr9hk971l6kM631z5A8myk5zV7T8IBfsaUy
5lXWB7S76sS3WGfjDW/LeJkHa0UF69jVOau5crYrKnCUWP2DoF9hSvSNoXYHeLVw
+sdnA4LLisHr8fzkqYsP6xXy9VhvHB3TUm1ymwPPNtvOEAQUkv02Qk0TkKeRBKRt
KQwKuKqe4Dh8Lo9As8ib0MiSvIz3+czQZksThswfiVWuvnQBWkHW4yrKrabW17rg
FDqjvehOGNzqlFwwYmMneyIbFEymXSieUmg3Q1vKkoZkNKOQzcWlTcRuydW8GG5A
pUtPYSOs/iA+Rt1gGiIgRjztwFyTIGkOs7pd/Ze5bASeW0Te5pQBWyrVuSlTn1Xi
BwDHZptbH4Cex0bwLFF7i8enL3kfyBpXP4Ucve+75mxEiYdn+PRw4KhAMM1Ibg5i
uVZ47syKa8Svho7BgDgaXPkTI3TDDdXukwwYoYYRV5Lyjw3DcJau1waoKKE7Dwko
YDeaCqWcrU5SQ2aAW/y5DntTtYN69i0svNx4OyOnaGFT9KlABbQSZ0Ir5H7nvXpm
AGdQTimii2k3Y1v2MTqjy6y/1i9LCOY7JG+UzfZNJxnkYFXzBAiwb0XzuAhNI058
yEiz8Dkp03Y7qP78av+aJPyWdTnHxR/fYFZM/7OuHFUBE3rf3ThoGo/37iW4e/Vp
Pi76xQT9+uxxZEa59H8k384MNmYHUJa5ydWRoXgfoXgxYdZfDd/Qsx5AVjESLo/Z
euCMWI0+EjkGdX+MaZ7/qKC8LblZbZucUNy8gPEABfljefWYhQ32eCc0j/duZ5M8
7xX+IO8B8WxHVqwCN1YKu71Wo4NenzV3TEcMrCNFywXaD6NmwBvbvuaV3JWtzV4R
uTwSWXkYDSmxJLOlP3BdvlCe5yb/WnnfPBiMXwoBF1z5CILfhNEoGS1Ak/2j00ll
Nd9DDXQhPcH8WRy9vM8WV6e98CiMVi5p/52ELDd6kQ7hPlYE8C1BhZlwsouVPFon
wEePFHTIkOk4jDIpewk8dK4zAYvAvT8X58V2E90cwYXnhLtiGVq0iM//jyDCZQof
FHWJ2z+nJ7n0KMoOo1CmvFV9KTsjnoWVQa2h3W8y2vNo/6n7mHpZlfiihOqcdzU6
PXBpnHf3RAIsTiiyPHd8IzjvyhHX8VOptdSv8AfOCFKtt81yfpdca5UwxcSjQC/i
8/FB+xmrJ3dbA5M8pClxFodFrykg4KvunqsUHpvM/BI98pH2ggmTOfEBAKso9nDj
s0djJrcR40YJUe/sIi9yzXTipmtSMdgtaFxylI7afTVNIDje873CkeI+SKHgTCuU
fY5QSUvWuMD77JpFjW4GEsc8h3Aaj7N151LOnTj7A5Gg90+a55NtELHTD+FELAHB
ozqkc8dQIl+5N89PSxacSi9Ih4wUdpNWEm/Z7tmyltVfn840CKyxdH2YS9Gnrsvu
bH2HhZPcbBDQ4gkEadzXqSlz0zZU1Rukywd6CI33X8uY40Sdp1nTN1WZqgiGitmy
9Rg+DN8eAupoQvW/KukkyhS3S7vE1OV39wJmDRKUf8wLmMuEsQaCVeFUUoRYSRvM
Upt1RztkNeNeCVUdQ/jTFO/ZBISyyDUt33e+mKZG2ccMq5ouxcTVooyqFgVmp2dr
OX5NEw55hpu1QCuN2K9Fq//mkbAEfrYq87t7FD4aJ9MfAwjA6pmPC5LnhKvFkSKi
DGmKeUM+TLunx4QbgdHPqSRWK28sDBnK4nXjke9yoplcE0eohMmj+PqOJ+S43Qyu
hucrOhCHCubFSchcahRvPMYa1OQjOCzWl4SV7KDr7jGOiAu4/2Z2cP/sSgeKLECH
52iw6320+p/G6/jj9sxHuL3nfB+eTukyJFsYAS00TvbBenTWVuLc8RBTkCZlwj5U
Lr2DemvxMQGdATBvkjSf9dTkqWjobv6iBvJ1QPK/ZGHViQzpXhNhxW2robbvkX3X
ias+0tRyPPhjK4w8NersuiyZMIhM8+GlUtGQWLDR6HSkmCg7Ap+p5QCROezmTjsh
7RuOU6E8ZSOvloOI40p/uIPwqcFsaW6kBIN+pizHwQ8u1cHZoQKmzcLH9bCqRw6/
yklz5GsQCCVzg0WF56D7RgtfZHs7v3XmxiJcozIfMFHmH2YoGfNfzS0Xis4rD6fb
yeF/UPlAnm2ePk98yzbhxCV8+uzu4d4SZHCqteQSwQdkSem86TOlJHzGta4EQ0UI
uEnRHceYsmwBlaCM/H4BGaLJO1miSn0zSV2OJqZM77wpD3TLzCDqc+qYPZaEYoXa
NlPIyL5kPqIVJ6c/9kqHZWMblfSQlMVUoORwP9Y760CJxXL4waM8tJDPYZGPf2RL
hU1BUGNq8XDLbK/dTlRnGePUf/TkKnKfH7Occ1bOMRH7Wk32QqK9GsIGv4wlLmM9
AcqLNl9vCplkvWo0Yp+wKMJFlUVNOhZmhkC3llLX5CDN3Bmdpdz173ERA9LP2YHO
X3jLKk8rLqAMVjQWF6BmOo1mWxSVQeC+qLdpFTqGUG2LNlzA25/+UeCO4Rbk40fe
e1j/G+fX28aO1IKNU0UU4is21N7UpQfSf6wjy2flym7CN9KenZhoCO0Tf9zxGNkz
tpZjjaAW9RgwO8MIprFGI6Qyeo9swQdlNwvbZU3dr9tC0BOCm1PbkbJmydRM3NU7
7pfrB5yz4k4iwVkFoUtBI07209Jsud+D+Yk99Xh2xZDj5Jq1jwZUU19rxtzxEKhg
hyc4Miim1g8GD44VnijjHfPoJk3ai7xAfbrD/6Ru1cZNafUSHOWjKsknGCeBOjF/
J2Ka/h6xWi4J43r9uADUSaMHYZSvsUgECD9F5C+DdOpgEBPNj6pAoEw+kbXw8a/b
s+dqk3SwGSAgaI9hnV1w3Xi8ov745vNqlsNU4BEb3sSyQ6Ero95FthN6VpvWHgPn
fK0AZJmq+6yH0RH0joDMSy3q9HR1QQGVOqwGriNXdWR0SHnL4//yrG/mD6Ko9JLJ
EJhoOvuzcqnpNH4MwHLO9QGjlYmYS3zOTLPonzNeFndw/40+m9kk3ZHvqv9ajX7L
+gK88xC8TBtZYBggjguujZR+kD8eaYfgG3un+6dl49pqMrpSR8wcuv5ItCAW7DOn
U845cuCs0bqDLqemthU3g5u//hHanmRrNdFVfbwDIXZUvGdnkyC5/UdMeQdWa6of
ieWFq7ZVoAiAv8yRibh4K6qZdfpkfu0V+noTHH02Npik22vdW3WFTveV1fGOkr8n
CEtRdWpMiE7zKH5hdEKNDXuJqJ/algSeqyAkxz2dRqxR8vskxGJDQ2K2d+8hhePW
lFgd/N5iuVPZLezHIrpBNi5XkpZGgIByNz4AdC4oOvg5uOpAiixv6X2TSQHfATPj
5v4JPM7VLaUOszTV9MjQsFS3gcKVU30XcSvx4QjPkMZQhOj5lFYlZ8c3cUPCrybU
b8PYX0rVJJ20v0Q1WlQ67qHkvm/1OgLNPKqU82Yi2tfPLjFRjjvVfVkh6bPSRRBQ
kWF005QvOsnuADthZrQXXSszA93OLXHC3BUAaM3X+QhUr8wE3/JdEs45PVDAe0Mc
eYndasUPSLQUd9/wZ2m5vT00RO0cJ93hi4RieQOhanTU+jpsMzRnfoCQeupYa/ei
eYCwzP/hhcvx4NgbwIMwTIPeT/U15GdIM2AhvoGArhbJgq/Qj//fbwwJ+1gErFST
UWPalqrEJX/l7krQb8NSQNkICHqGS/fLTACPf3qUMviGiB5E+ua/umQFDcdjO0+e
ahBdLMZrYCg7iZia7tekfVU0nRPHeFRwNJq+sJXLwDmmofqWdtwDLcdz8H+Aik7p
EcdrTVYOENW72Yyow41V5owBP4BE8EQcPbyOpZc9onNvM6stNAmhTtZnKxvmN+ny
+vRyBCNZvVGF2VNHOZNsoXJ7cIGKBUf/z6r29DhcvB0CcuxKAjAR0BSxWigvkXx8
aYCIaftIIItTZVTjXNdFk4LZGDtsdF7dpWzp0JH1iYgyGkSIQr1kRbFgfjy+mkBm
W9fPuJOFe6uO4OXcN4oCIZ0NRztYm1BhFNtJvrPadKipfX2A+NACyWdlrN9oFmhv
lXinjkQMNwfkohvGj7tlqeX7n7lS3p3DOCK+EzwAPkhZh6Uv++Wjt8tTxNuqgedI
wrRUk52pLkiuLqU3zKNTY+b/7fDGQATm9gqI1mPv3B5XBj9b2wZu7ygQX2n5GECX
3iPOZsKBHmG6pfhSJoLU+T5EEtW8xv9OJRnda9Hlbae+OCrHeqdofp4uDCtn6AIQ
8+iVTvSUe8hSMR2DrA4Q1MQ2LXZhS8gXcGiYNBP+DbFcZjEKUUfnxrA7p/GaS+aF
3QXExLfdR8oI2V93tsKhDdNxLkuEtPgPNy2UwQY0PTufl82Pmim8ahjU7MFiI7LV
wxbuNu7OHrD48V/RsZC/YVG73Wrn1tpqVUgF/NorAHgoiuUhMN94OR5aJdMhVAhk
eC0CbNZ0svWzy7L/4rTQKDxYc4XsLiHSWo9wprlojz2tK8M6lmpbjLfMDYDfTnXu
PILaQxZuVaFYH7UofGcNfdDJZz9I6ZGDaGAlxLGphG76RGjVz0qANalTta0GC8qs
m3Ve0XbMJURJ7BJu47JTh010kYrq16caJmnUk5r+ZoGe8BU/4xWKuDyXYPFQIeez
5N1krFE9znIzG64g1nTDvDNdS38w+6w+BCBtyf2LIKgYppbB4MWnsUT/S1AF63q5
+NYkpxY4ZWuonSEx0/7cVpk8RPxJc6DXgrocxP6iVriS5kihqSPXPyylwBYNftyN
AUNuztvN66fnBMLbEKM7Ex+HsTmBBKbd2nKpsHer1DGNU3FUDdTWws6PJpoRMqY4
b+LqVuAqSeOxbizQ8mnkP9xP3NHRDfw6tiVE9FCZ0W9vgGYOA9c+Cu8AcUkdP9Lo
71ieoXTqGGu1uN5wF2NioY9kp6tK/O8s+zvC5wAgLNisOIdxZag6wt/yQh4eGlzr
fYwAVEW6S9LT5wWzwsmipcAM7I9Z8nBfPPv9gBfjZxloJn0/jYTGFlj7c5cNROYA
ELiTh7SHcKTB2gavaRtkQMidafn7F/RMXPgekSN9BegkywsxeleENZgSN0c/DJvm
wtdGN1phKHZrJY3LY4U3tn94M7xl1YSbRIrimO4AGija/5UrIcTVQcX4S2k9mKNq
Z7JswmAgsV5TEujVf/2vGYzU02fms9hi35UJAn5hWkCZFqQU8ATfYPGr5E8cWxEk
c0P8pp0XwOSaaMsXbje97LJmRZ3iusLO7IIh+OhAmmroztUqfo0Qgk1p/CBQh5gb
Dc+V2cQIS4xhKMP6S1etokcPAlh0DEEJQwBo1iAEIQMNihrxB4SsNVuqMI1sFlg5
OZlThga5BKpcL1p6Xrah5mx9ZJtTFUfzCoOfdDqUCOMWd/o6dnJFvdEi4WWKrfYJ
ZMVptbgR7E/JkFtxvpppQ3lSKEDSA0AbbXoEeHYWnUjsBgsJyGc9PnoIlz1myngR
YapyNbY6Gt+x1FH8kwSzIr59SaMoOAoF4Eoi0Vos1CwdEuW9E2Nc5krHB079oqK/
EfynKEl1ybRW2l/fBT18FRMyVCtT0/WZw7q92RI+acQK3e+kHkb5bqLl6gnN7aO2
RPCufnfi+Q1U99Y6M6LRxaRrNSFDlM4bdyPMEEozXxEr3I3VdZsUsXNj4dObf6yM
EH2liHG1zU+GEQW2TqzJbdlL5fJmsHEMQ31CKLD9pQiks4kwQUPvSIX05SU5CH4/
FkeG3Q0jIx8ciiwQbWEwoUSWL33MlAWeINEP1KuRLkJwTu2d9J9jvVmUheGZTzso
R2RXdUpvFKNbCVyyimNprhdWRPSJt/Uv2GEnBx/nWevAIz4UaG741TIasIyKcJOc
w1w+KGeOPlPArzQN19WWByUDS3fbgHC/QZ6ZX3G8Up8Nou9pWTj1ISfUrT+y/cSa
MRymxz8sbNbDqpdrrLvVcjiYB4vo2p2/U4laeoxWn29wuGTuVo7hX4RhTCTtE8h7
S35OmVHGp3EilVW1bOP3TQhcuejasxDcpJ2DqGKT0gGF4RcpfxMmW1cJWQrWb+U2
wRpkDfEE47PYOlyN35TpmZ9amTn5omhi1Gt7YZn9zFBDMYWoOju9qBc5l+ct8X1E
EpzO6HjnZCUzpg7PVtdgLjufKR0IdBJ8iO7eYOEEDgwht1Y4Swqfi7dPTeEcmt6M
TlYkSmzCNXSaIeOyQqVxaakB+G2T7cdttKTwhFJ3CKYe58oWDAQhSWJqvi8G4Vkc
6ITlJH/q9mrLPFCJbGPThq+w8tRBikIlYlBWTSGMk+mms2zt98cvi3Y91l79U935
T7ht6xudjERXoeqOoO75fY/nQm+T2ijdtVuaiDuPplePA0wLABUW3YaALS3Mk/nS
ZCBZYhS30ppk1eHnhfRE4ZSodQUefzvm6BQyZxAr6/DOLxzuf2lgk00IrA6MnzF7
4i9CMhOtcZY+OzEaX9WWe1IaCutWzoatqZgo7LvyAjFhDrxM/7LMxYlCOxUOdhqV
6V92aCfkS81Ygv6J6iDntey8s2wBPo+d0hXrODuM9X1p7rop167qwP9WRzvLAwBK
Jf/A3VosH1O1o4+g1RvZZLOesvW0EDrbQ66BEkvtYbntShZHuU3XZ25l+eK1xoGF
oWBREOeNbjsifSZYqOBSZIKQiJIvl4/NqXA6ibTbGMtqb73q761R0Qkoxejcp7YX
OOTJF2+c7ZFcDkp30sRWvN+eJvk9V7cpvimeqD3XPDz59fmRglRIAdImeblyHlwc
RuKcJ1SEAw/xEc6o9SQoslVOJbfmetvJG4DrEl1N1TGOvHchRFgss4A90wENhA2P
sY3Tl8YxCIjVl6VZ6Hh7wbswNCCnGbZIqIXUWnh9vgpXzkHOZfU9br+LlfYB/4Z/
QwNqDbU2V8L7XMx2e8mIQuh+dW72ln6PA6AqwUBlsBqQDO5loNprqVs19qQwW8BI
HGv8W+ZVfrkSbHk3LxcLC3GR+yplwKJp1rAXiV7alKoUMrH2Bu0jhpYEZquuJpTB
Rgi3vtDpQvVk62IYWduJeAUkZ6MbGz1IPsczgrXUTSx5BWNfPsoDzVnWGXv+M931
7FrTPLl7ye1EhaVT1rE8hTaYzeMw8KxeITSDq9Wy58QLv/BvbUCrU4njhIhnNby2
Y4GScYGac5LpaOnNYGfACjVx+R96O511Uy9UpmbY2dAKVDUl5kOpLCeHljo2cKwn
LhJwfRN0lIRbloiPzug2JkFDSOgPNPt2W+9vFW9UR2sjmPqGkdoMFb9P2r/7WGEs
AQ77t3xjKyfJzWpWfRm3gF9wThG1yAMgTt0DTr7Z/JJ+bP5fsD4D0P4zsFRnzWLa
EV4K0Wn8h/Kc97IYa8KWaf2rmpIjCxIrn9z0IJuX4+7cWYjJpZ2VokLvxa77IrEK
/jhbc/1Ipg2pwZATNnAivMrblPBUc2vO2+i/ypqyRVsQY4nYxslCXqY6rEOAFHbs
/SU+ioZTvYl9tp3I5dyIsC3fzECUegNYlbU5TJQyhWa3KBGi+NVXx2d8pHVsYFzH
CzKr09HldLiXjOgEmsTWcwCgoF1bpl1Y377delhmhvFAE/lhweuXx904PSEk4QMP
aaZQtcvvwfXqFipT91PJEGLSUTF9fFjsylYhX2jgV9J0AXEqlDd4IR+WsE6UPEDp
Zd2/0AiFmcDdwjqYRL+0RlhC+AW6ypC623nGi8wTIa0bTaaCXpKS+od5zjuM3rlS
b6eOeVDKI4zku1sytLDwHfYaIC/RhPsfodAA4CJI4aJTO3Vm9k388Djed9RviPqJ
rKnXVZSOEQGyl6VEcQrMAZgLxG8lxBU7QKdKzgCOkHhW12hJ3WQ1JDSmnlkp+sqd
UZy0TGyMGyUgaV6AEcB4v/AKFvLIx52XWu4vOl5BugUiHdkF/MRSFGo+jFA7koaf
66qxXV87tPML/kN8Lv56lr6L7YUXASwlCmeVXMVEu+jjpUBes67oFh3v4X+vk6tV
5jb4JP0l7y6h6MjO8rTt0Zicxa8/SP2BY5SjHnSqatE+36liAlakos0B3mFhgoid
4pRJ197Qi/TA6fHVRHoO8khMHk2x6QteOoQmfbLM9yOD523+ixw+IrelHehuziR6
HVuqzWP8ID/Y1mwfAmcWYKrUVBTh9Z+3fUaAt7u208jhcQthonOb/5hhE2RIKjtR
I2Ci39QV+ziuI3uLyjVV69sN5Pw0dyOtGGgJzgIyfUI/c30JgxyF4PaOQq7O7IxA
F0EAN8JOsH/lDbyFu8YKlO6E+gUKfeaLXyaLD8us0hHMaoOpJGSmFMzqvcDxJXH1
/YGZzBkLMQC2D+QlOoahalO+tu/FhorG9dtJoo29Jv7VXKwABa3LWYSFzNaiKJOR
VAKMNMdCbswDblyUKZGkhgCYrSS0vgUEgaaaDXELgDI2pJVhnQ5kFwkRjR+49icz
BkQwdodyiHHnsGf1F4ewpSiVkgP/WX81XEC+pxPIXvd/6w6bLb7YwykCPx/RN3ls
VKQgJcea4w40A29Jxvq1IHtS2YS/seNhyd1IO5O88PAF5Uq764l0JEYWGgah37Ro
ydN16yV/zuNUwprJN1Uh5Kyx1v2wqcRG2NXuMH3RRm2zFFtGbk1HvZ56LY8UAXSt
J8V7iVPWPihepW/mUF9YCjeqDQLJR02UJFH/8htolZLoarMcWfZ/9X1TFUMJKpuq
p9iOOQNJ8lgZC7XBIFvmcd7FI/8/dEhZhnwhok9Lx7f9HG/GZ+o7grzZ6I1dUdWp
8w6qa3Q41pCB3zqHP9lBscUKd5lX+AL6PasQE+fjyit/AlF0FsOW/GMdsbtNyxoR
Z4KWwtpkfiJThYo7OZJKoIOqzb+BybJ/z9NhWw2qa2ZbNASGQ8gQUvuOxduMDGTb
kSVHblaBGKlPWpxyQD0qEvKKpm6Ben4fKKZJFjv1kDj1pjjGFpzYiNqb68cZZQT2
Wu9SPXGGVwB82HD844l96MmiSOsfZ3S/MHtVjLbi+sYHt//efn0iNYv3oaQIBHOM
XcqcQ2zNuNmsYVJQWKZnAAnjGs1y0KTy0+SnOKmvbLi9YHh/s8LSL1u8AdYyJkJ8
GreTZQKbqTiUcTOdW/LM7ejAATuh8DPQhqBM9bXNlmYDQBsqwqhyo91b7sGFSFyw
pIuBC/c5svd+4Q082fmk7hA2cY9iA+telyORCOZh28VAEpvHv7kwL+jsSQmLGeLH
8l/Rcux+oXgZN3x24F390nj1bC4hYFQuAqUGYHZgoqu9UXXv1dSDEBuiPu41Ktac
1jE8CV5H2WV9BTmqB/ts7zQull3L8QEbDIeek7Nb8xPLVgs5UMOQmbgTrPPaB51b
fE+MRqOuAB9Mu3wvnPMukpqJcdQoB77OeZQ6OYqWY1OySncgCSKK/bavUcjw1eFQ
o5dcqAUg/c6FWLIt1j0PM9wz8dZHUZ4dOYyzb8v75vtZtTaYt93HqpMOUGabRQs1
WKwFmp2d8Z+1ObKHmt5dNts6t6GGTMgCn7W9d4i4O3oEeRgbjgpsqUyycFjKDZGK
N+Nvc6MU6MLRS5Eo38psEwjBi0CYkLVdDpGnjgOIp9eancwvH6BSgLU7Tz9rYOvW
UUAOxzoYhFkjEPZNNSu77VH7sjokmIxeMuKgRSX8DHLUICZzsmkspbkiyz8H1nX3
rkF9PqZ91hwwcLZ090/bdTY0vpEiLzoZFkUK/fA8Qy2bNkRBKY1hBxNExXLWSiXl
4NV+x0ZLflyZplPFio8P/tnRBK9KjKkWYAMhoh83vAYHLj2NQA5C03mZGuZjEfUQ
SXnRX6wkqgvhljltaGfnIQbAnaAg+07njhC1wcFdIjB4XgBd3HCcnZpiXgf0QD8U
8tEkmeyT0a2yQPy93hjj6dKgC7ftZryGoQjBMq3tdOnPMNgDQjLZ6+LxTrCRnBlg
vmzqS+E1w3feXIzuFEySe90VMMAky8K0IiehrzkPj5JtWF1PQTcbUdbYa149kfbc
lpskdTJ9QbatJgwbgKPVPSkzvKxE5gai5vgYnoGskbIKXR9KBsKbYE0RSXEt/i25
lux34Qy1hnMOuPRLI7m7PIjz9C7T+z5DPRwMoGCLBlrXgcHlNX1eFWPDHnlX1xiJ
g1PbTf5WLdHqFEQi2vzEcXPTTlFjUm4gPlw2/qKZDZf507sYtzxFkptiX98qdA/b
fGrAG8FSIluQE6bv0Lvk+UFvZfMRRqld7BY1mJPEVN3tQK1TO/6MiMDyA2GoLdwx
s26T5ZEaFWk+177mc761SKW5tmAlkiKIsMB9n3mJglX9dYXORXoaQ41/Z+jcKEn9
FsPh9RkU4wxboS8csz4j2hPtnSVHKd3q9/D1mEaNG5dYTh8AtaUGMSpSdLPZAkuw
scNZ6EDHZKLheU6pTPFXr7oP81P7I0sd46o0DkrYRFIi0kDMXajgXaXFuNQtvpeh
L8bFpfeiYomxwmuQcXbrnZp1eZH9Mqg1qQa5HMPaeidkn2Bj43URx7MYEtZWwUDc
q/K+jEmzknSKfxd53V8Jka4J+rbBVem4DbJwpI173ov8nHhUjs+nGjX2zC1SsI4l
P/wOEdo0HVBkEj6rTfk0paEuR8kHoJhXV00rJo5GOiRWK6SrcvVxsEKfYWD3/yAm
rkVWOJddFOW6PqOK5k9pvuSbzcokOd7202clGdg2VF2JOiJJBY/90vn0/eHO2WVJ
dkhrapbVa507qpXjRMVMoK2DbLTYLg5Q8ux0s485gT5Qp9/nvp5bMtdCYQSuzLbg
+IdhcsPt8Q/RHZ2R3KMIaIUBdEHsO5zhRN48vJhBJv1pAhXS6WznJ2bW/s6nOL9l
q0ywMJSjRq4b9CetNzJgQbOUAxY3fO0sYytB6QYI4qp/OfdVD/ervWPTYJ4SdNU/
1HVB6NjwfXsd8MWKSTaDQBR8UtctXB9ThjP1IKC/6/pvce2UCCeWWmj+J0qIX/b1
KqWbj4jOWFwu+aai5MDI8VbWL8JZU3lAA4XrPJPcYxQucU54r5LMnC1uSYPBn6mK
0RQU5b/wNwMcMP/Sows8aeC8CCLAC+Lz/oNbsLX0OY4mDQOhwqP4AeOszwqkusjN
1rMx+VA2pSVRrTwAsOYcTViE2XTRX/y/W8J4ySOMbyqBdzqGXXMFsh4oLuU5ghX0
OE21YUeBhNZ2+OmR3fCtMoO+kY38JHnfzE6qizb86t9USpAsHITQzdIZ19VvlUcA
pvku4cugVKUhrk+oyxiXDub0Cm02P5mctX0m29YGeShpFJ77S9+EZPDji5jpN+xc
nWph147gpzBmslkhrsURptTEmlUm7VvFgFuZvAae2pHnjZT21mCSdZgH+KKhIf+x
7UW7EU7i/KirI1sAHHD0kVBQWWqsFaNpm325kLXzLNi9e+fTKSk5omQpnFPvnnlk
vvQ0B5ZWcCMmsET0V41CWiTwOL1oXooxVAeFWHagrVrVt6ig+Fy36tO14S8J+LCp
EEtvh7YzOIWGAjBiAUajiAqB1Tngo+ClHYKIlPNxb7brxH4FR2CbbEKdOdZtqEHp
KXIp0dUiMYZkf3IBGej/JcCm9ZxNpUOZiQPlU29zl6ud6PLalQ+lQoDs3VSuF/Ba
535WQd0qoS+YGWU1CaQqBIpYqQUdlFAaEJz9vvoFwPypdmqc7NXPUpt2k1+z3v76
sme0lfYi6ZMh7nslW2Y+puPhrXWA3psWRCPXTXdealHLMjVxuKw0RtYvY1HkoLxl
AEhQNfIpWZsOVCF7YSTM0kYkeC9V1B05bhYdNJNSU3KzkV8pHPOMlFsuf2IKpQj4
00Y7jFWxqtMmxsGXWnSIdcY3OIvuZSwhhyGIEdb9lsSvb4AofO1J3GNXtFMcgLnI
WyVnOvdMhP6kvKMNX3+PftdjEUhneDoDeTGTQVvyklPGLYlRIFjrr0eEqpvyQdDc
SOFo0MxcFvzWskgTXiNw2Yf4SlXgL3bYyO4B1naydYPp/sSKFEuL4uCWP8ur7ZDN
OqvyVG9qe4iYuXZAvpUrdK1O2weYrcDXIAN3ucn02OHhsZxAXUKutPVRxRtfe9D2
TfyfeYmiC1tv1mQBUh8TRZSJbOez3VlCQzaSMzdo32waXbqUxI5QcSt5cZTCubwZ
03ycFF1n61y0QoBDBDwL9ffoLFS4h8M4gvAh+PFyB0g1fVsZ6U76xol/ngNOjybM
rrilkpnGwUq2Yo5PAL6+V0Hh2Al9chGw+ndDWXj4UneZ2KcO1WsMWcRjjcd4GpSj
deUdU136RnYxjE5PQTffKpHPu3icwDdk9dAwXtFpTLKiz+b0uWFzIPSPlIDA9ECe
9ripQlhaHL5VDP3SqeNsQQJ0zwEo5/SoZpRh9ZNSVg0QZoZaJ2mfBCKECYwlR0rh
BX5lElpYt/4kEuRmW9CxbknD2NpKe2uQ1P5N33u6RTtbraSseLTofENwa2G8Dxg3
26dx3e3qM7BpSmttlNYQfIO8EDXZX3noHcFaP1LVYChKUWlsPPFAiBQ1nfTG6012
uxuUf9do4CJUwJvDOlwqrCU8ADrq327RYUAj6ZRLj3cWTZwVFTUSgcDYDObol/Hx
H6PpksqC63veQynoPqpP+MzOeWRkaKC1lQdsubs0WpCBD+gIPvJiBz1UIIBtF4Dd
CoPtBSAIBEz18TI0YcPMs9dz/UoZ0l80uYUMhEnZxqCXwsiWeFak+rtL7lhVybs0
aw929ov+ZuaQ6nC7k1k5hXadw03rrQdwEKC4RRUqWXt+EZIiqJUO2ehWW/6QueSx
ADR5KpSJKCD+SwQAFlbzmemBEmK/DgFVAT48h7DKfe45iUOGhupYe6BSGe+yCEH6
mD1LTynFJfSOUMlymoHCVo6Jj7Mm0Igzf27vzFNR3uNKQcK6VwA42wgvZ4HXjjt5
RHBx46UBKmeqEF6Qq4yH0bWoipp+pm11nLG2CR60eOEgFM/uIbfXiN9NhuyFdIN1
M/zQwundfj6CTXZqlgIoKPk20LEi2uyahPo/oiuynrGjeUmVEl3x3hKpIjhbqQKd
B2GtMazwNxFby+GcCaaF9/qewxkJH3HJvZZ68Qo+XnzZ2kcWP3m/B6y0FIkjEoaM
G0gSRIVeLdFWR4Rrl5bPgbK1k6axEvsjZiZl3BfMelh151hiFHtlMCj7QViTDeH+
33+efrz+I+X3PdRxG+ZpTbl0pGhSn9nkAq18riBh4wqEMmOmJBGLmPu5F0/Dupnn
RKkc0nfRuUcjdSYabI/EEspeDwRAs04jT5Nuqg4HsWfA1TMGMFKGaqvSnDzfBsIn
u2pmOQQkxy9KQv/VV7cD8+d4OjZF8P8Tlxs9+1GnvcBvYSMIFN9v3jpV4NDlWgV9
9t5tn25JoefQqQ4DC1DOIa+6GDICBZ3S/mJfovLVKnlWg2fPn6hqtkybOJmzcQlA
62T++cXN+W1qpeoK5MCZ8nWm0+TO7IPi7Q9OPo8jUv37G4C0B/KS6KeU/lJKuW54
C/IuZXRkekR6yqPV3kJMxXjNt6qDAvXs/5w+baZuS14zS31tHFoE9BQRHUKFtNEg
dvVsabp6l++U6QyXQN4XRZDP9yHYEdNMdeoOV6Did4WX+mi5ehsXrIIm0bQvi2lJ
zur3Mcl/yIEQRRD07NlYelw7pBlGEQdm14EOInBufJK3JV59mMt9nLwG0CJV29Nj
357ZnW9YKbcu2CRM/BoooUcdIfc3XhptSoP41i2+8KKRp2TnZ5nmaVivLK+5YVNE
Qzk0TK2+0KXV5E9ff8LwGoFpLGnlzoifstCD+/0BfbGHUt54oN6vupUx5wAD5boc
x/RJV8QM8LoFH7jpml4hgjJStStziMMcgSxSRPnR5mfNiS6k71OV+OhhgakESqlW
NckLIXw90bPkGjX6OOoh1RGHGzNmIoIeyk0WXroKP+Dq9YU/7pvyISs4IWUMdIPW
WJMhl3370Bii+0LOd4rNxe79LMA4OwSVuBx5eAssXycA95E2r6IPO7phN0KDxsTf
0o/jry9Z+Ub4d+eJNZMDReaPvO9+UkzrRg6/Adov8bF1teGVmCSpIhXqqZen9DXt
Cest8cfVZPJTbrTP2TNLA9UWswx4hCGoCHWHM6t+xTyTW6peYl2XtTyWMY/SatoO
r/pIbK+rKuhOnTmeaWFdw0qi2oLHR2hxlfOsRznwaBiGQjNUyt9a7iju6ge9XJN5
0EZ87XDohP3sCjpS6evnG70WAfETrJ7Px1/rOW676sUKWex/I1GyewKBgrOYm7jD
3f54hvFrgYaGyKBHAd3HjJ1IMm8mIT0nxEHKKIgckb9mcFyqR8CausFuABB0I9cH
QFOedhDlrfupIOuFZgLFSGPcFJ9iKoUTF5BGosH+45vuUoB9oA1Z9Vle+RRup0Bj
okrkaBigvnRMTcgFwWiuScL6rcq81z+pHRy8WXhIWl5W7hCPncWexlTpNy6z3hAf
eCnAvYup35dKEbBFuDbTtrpGyEBETVJDcuB463ILOZG5/s2b73xsDO7mddGwzmJQ
D84c0zZlQXDvWbS5AgHdO2i/RByzdzMFosK9QK4m8pz8MPzavpwN9DhfvzY/2K+J
Z8XnakO8FitZFyoI/X2PDA8s9F7G/aiB98XJvn1a4kkras9+ar8LQW/o3oPbM41O
l5h9dxgSyjwSOD+mr0Oz6lO+tZlrN2donS14pzMTNyIzz8/Tzj3a3DtoEhhwA/FP
xoWS6CCzroaCO05KY85uUrrj4eQ9V35mbPr7uUZKXAlya9T42vk8JLOEKgxZpkzE
la8/XcKnBVxVEg8ZWJR/sjns4m6S5iQPK8n8SNRlFxUM5JmwHPeOusiWGNB3V7kQ
1u2j2aWgQ4wAuU3sA5E4syqmfa7lNLh+B5PdjOOBcZsvI6VsRWTTTVIdhjMQZvXb
WxRgsuGhva3bEDD64aSV3/fc7LH77r6HX6bH722w7FlI79KEUS/RhAPxwPYLeC9W
XiaN6sJ6Avawp3SAjTzIEbeuDIlbmu995LNk3xfvn4IRv90GAkQlULP9FErjRzEI
58baebtshic3aYkxKSyD8nOE3JyJF2cut39WZYoyjA/WIhV1rYDucDmwCWHCXneG
DaTUjafYSP20awzwi73somIhC2cWcRB9JSFwnm5U+cDYk/KLlgXcvngztGsGVjZ0
f+IJPYx/l0sYlK3n5eOgDt/m3xF0pG4Hpe33axRKxuzY9bi5wl1K2Ai0Gxv1CPnn
1TzhwZ8RuFygbkIY/8KTcFWdHAYCrqON4XvlaQ9XbMcDYyZX9cTmoJRTdz+iTZQk
ERNnPi10j+15OC3zKbU9cl8r3qhzLGlSPKz8hfDhGZoSGx7mXoRrCbjlhpGJ7BME
n/CmDtHs8YS0k0EjG/IPO60bsYhdxHSxB5eJ8RNpJ8bhb04r47wEZdilHOl7ohHM
PRfYDYg5BNisg2p6MgEFjom/tcTmJrnXmW6qXbiPjomkNll1LI6G3b+X+xyOLGIk
vF9TObNYrXqMnPw2qgUjutVSt2oN+1Jy8JUpPHuFcFfSMmLCOWIKtZyRlnLc4/J5
H81OL1EUS9+PkxEIbG3cVTLfjIOve4Wimbg74+hhiMhCgieMr0Jn7J3ZEvmWtfiG
iDhop6w9DIUsFRtTsPpv3juGq3BkayJFCohtkhe8sKVpiIESj03Ps4qNU+vyl0t3
GrRmRbfj6iEa92T980HcvG5vmXzZ3jPXLMFqABp54YTeAGVqlxROiUU3Xjx3d+QO
Wh1j9bc1NOkzvDd9CdSUtIEU/A1q9F3KvmvvgSNuT5D/lMa4xW+tVlQc1mcqCeMj
PsQ7pUN/JtVpjO2+z+srghkrsNtQ+EHoyGwckG+lwo7mlHCDYfVEKtpN4Pbn9juI
tnXFpdOPL3zkStDHT+lkC9EzmkfS9zqnUJ77EYINlZ17HFuwvb+K8hMlV1gmuKSC
cIVAVrN/rz2BNuDEfIZWWuzyNCo7A+9AyjYevIJu3wLtrLhJjO6uUW6Et9FNzYXz
X3n7dMdsNriIH6U/ln5xrTjJTblQ4+3wmESOKl2gYmqN8DBJqUmmcoLwhBoWUq+D
KVfdJuENRaTS0fTcGg1TShWCw7ufe2EjC6MosoyCar3KleWgdeHZFP3+0wyGLckD
2RIhOx+6ECSDvDxmNs+o9OQMPqYPOp1TTDArBJkDOx8EUSMXUY5IdbR+Ls8xCsSR
tv8yeod17tcnLy8bpSQo+gyjRF7HDBaPVIsNdLpMb6x11tBfpxWkgRdSxmFGyPaM
GqTZEunpVPn4LWxQTCe+1bEx9UYGEnNWaQ6wCdxhDHGVoQApYnJ7MchCBSAhFIL/
HP7qxADxJEu0TX6TdheNHdEVSBJ0dw4p+C7FdRvgkrTQMXvGlfLsTzNdsgq6EadF
x0S+jm3dfDplUu3cnAexnw6rNZCMvJB9PVh2Zchk0kpbRu5FebBMrwUwPzYjtM/D
VuUW2AEq/HIRMEw6+rU3ONMQbrOLSyuTpsLI+NLaghTbn7wz0BhCVdcyXEyzMtgJ
jY6rk3uDj5VxOudE1TrpC2O/PO9VbSCqol1EpXOFAaCnEXOuoHJDD3/gXGKIueYQ
VacmcPptu3o2M/LyfbcGlud+ZFZe9xD6bx4DFgLAOAGgWBnYZEmMW7AKyg8tMuYD
aEwStWHPIeydvFB/5RjBijBZpNNFEWssliutDbn42hyi4YxIm+cwVz/0tqxWIliW
80tcOJ6eRHfY38SR5/GjWfAQItnTPlca/CciDeg0MhMXPO4m8R9gKAu3l+Oy1sYh
iEFltith7X73W4bUaoyd8jrNKN53i4TcViWgk1Ln8fy3wcQNC2dMr89LweqLih19
6YN8JBYzNt7MW6mi+O8hqrDbKQlA0mrV64yALVezwv5uTotjvf43Qb8Z6h4wUr0R
K0nAEXy6EDmVtPFJEqy2u4nPm65sxAt0PzHxb4pIq65sRgVJYUZKjjvsQuO4hRug
y572+cdMBHRa2T0xO1rCPM3EUD4it+oPvTZO8xsI6R2I8Je0F5RFVRg/+HDPrPKY
V1zyZEOJjqFfWXilb07STsbIWN1SfJc1OeZweOehRx0qGxZTCWl5gmWmE/jkrVNn
7os7dfmfUrvbViL+u/6eqzRUhGBF+wmHXkIx/BFTcLChJ3BBHAFbXTuLALQQ+qBO
DMnnJAjcSaeCxJGElmJ1iXOmpIc+wvy2SF07hqj4md22T1IZum89WwAWqOaHoXR6
/Mk+ruUvkTPrWg6JiGxI3ndDjQmO5TZzr31xKYJ+N4LmmeNTEKhULchl8KYXAB/t
3Aqog65gQvEZFpAu4Qc3YGidi6wm/vS+/9nfRMkYolod8OAl1W7EPCC1AHX21qtP
9fTaJOSC2sRVqUaqn/RPWw1ISZqS4DFtfeCIuc3dmTKec56mEfeaGyrNToMIyko3
uNqrdLARVe5AIPP+lKjjz3eg8stjsaZ9g+DjKyRxkvQ5xat3t3ezIqeygwOvCVbQ
rAu1pfMENw9CoaXPhRpVA6m/JImzivLnVRmSEyp7t71Ze4R2/V5cIAs6AWTL9Bi2
BLzarL5Iv7s08s9R9/VOG+VaEISKUtw2sVO6UkXcUeVni0d6QtXOrAKOkyZqOUe/
gLJRsk22xj+PF7c9+zj3xBWuNEvPEr8iZDt577QwuqIhDFA65EGYv4w7ODy3DzS8
BkyGk5KVdJvJ9y5qOY2rW/ld6A4hI9U9H+9u81NZPjosBOeE3KdHVz34FGjoOoQh
i/oOPmO4gXt53j9qC2o9+NNxhLwNEJrX/kOwfJzQRCswiuz+vSPEE3mM6zAsAW79
kIF5/vR2DF4gjhdRG0vbMcV5Kov/qJVUpHoK7jVmDJ+0TfSxKH06cwXzSTx0snL1
ZZwlMdhD+T31rGK0/JRBCKm/85SwsTPADqEZpeTQ2hqMOkgczrvd/IGwe0+mBO0T
4YL6yENxekpJbDFBJUF/yHfCBFS0QqeeQH6674twR4RnWJ7EsrS04QY1BcRIqDFM
PUCnDdy7+QDmX5yUNFgSVg8qcK+8cW46CIzS1vjFMs9q8Kwro92R+DXpI1PifwID
aNwcqz7iIcF1iXlpuY4HLXy6alfu1/IbURBEm4qEiMzKpvzaR+u/x8rdXae5jXB2
Kw/pNZ+rVsC2d4r2HiSPpcpeFck71tBXx7H5ROGz0iRYmbT5YDBfFvN6/taNk8Ln
JMh7MOHZEjjTYucnaEEyBZUSTUpmxROqarbGYglR6KfX02jwjDOZ65l3p0+9m7Ya
kM7cXH1OxqC0rk6KhIIi4A0+kiiyVu1thOCIvylSIrgVl9cP4WYApU5DxwH98Q59
BZhnsFueiJbb3PpeeTmq4ZGO88y1tRhLplhD0aCKPBti1qJCMMtsbENat+puMlu8
xDhIL3uHdQRM2MgU+W0BFxnKLxIFTn0a+o4axSpewIwUHa8+a7tEK7+5cjKR2UK6
LVTsVB3JF9diKzelcPCU4g7/uF1mec9ZMWiLiRVPAkjS8rNxCnL3fOszbD61Vu+0
5uWnwCrtQ0xH353e86GgJA10NYuP8Iw6+fCqMtuLJRPqf9Bw8z5+qYzngrXSM5Bx
tqwIzt2Yr679JlmEVDrCz+U/zOsoNZ5uoHIgcQ/+JvlOn0OwnZG9Ox16bYqXglb3
MJOoiWH/OLi96pCrlgKlG22xIgx18q3a+fwIK1AqNJkZUDs4ANAOVggLZHdN7+34
8mknxf8s08VeszrYWVRYeD56jKyxrJ72cjDkQIHddtvHroLWdHexN6SWeyfiexEj
Om03nOtZLndvydvjAlBAi5n80b2H6fF1WIHFyBsPx1O7g3wJPYBzhJ70pRSgHhVA
VgBdxTruZhhRgby/A1wpVEi8YnFcMqg+yuvqiwgOGmEfOOftoWbZo7iS7r8SLUfj
n/Tsg1z+r4nYoCzHWRKEqTX5Olcb8rhAxHO6EXRxOvLp5nAJQuZ5cnnKYjXHMDKX
3G3BRsxrTk0a3boSoSFOtyh8umP9Vg0FUSH/dQ45Q13RqzOMkB11ibjDvVvgPrgQ
NKIORdhaC6arviFoOgQR/z5IgFhpIw0PWE1Flou8ElahT1JjHHQUqPQ6LZ67cydi
AqtM5L7FbFAo2UBvH1uG2M3EAWV1tX8vtc1ZumMs0aZtEM05RMP5TACzp3LqjJm9
vPTJVzAdhlWv1YVRSId2oGfM970a9Nv20u04Tfb+EAzII/0gPsXgvgxClbYwY0NX
bqU3RDNF89fovpOSKf2KIagS/sNLRiE0KPRX1qmDnG0IMNvszdV9Mk23u6cF2GLG
EmzLhg/gDtnuL9uIavjr1etZnAczGsyqiUeVVZxaL+6lP1GIcbTZi7AV07kgQdRg
m6A1HEueD1N5N6LtFONwCxch70/73xgbTmqMMCQEqUITC2y2blWNHiPCpcn4mDeV
DFe9HYYof0Ct1NRsaB7A8pd6HWG0xg0JI+C3NSWbO94MRnNoRAv5oeOLDEfFTaQV
8EWbRnbCFQ/0wgpZ25McuvVhlwXnaqaxqJ+RhF3q3HicbBPfa4N/JE+rtmGnoq1y
TOjJPUCSYutkX79cV+wPkjg6/g0CqPsseXbnm0HmFyiHbpMbBHcFcpGPBkjIpW1Z
3arnaH8hHmx51JnSCrp6zrzGV7nkc9klY4HSTRhitEDMHB18v8he1Do/EFd9BKdQ
Z+C3FLerunr7gslQV2N4Agh7X/zhwWYs804gvuuxeAC3aPBBhlHsweiNBcB0G6yM
8vKdsWHA66ikdcB4mPKIgr+IWjH+fFDPm7eH9feU+1mna57swQ+JI299Daqhgxy2
yck/eOfCa44eQ6OXgjWyeTSHBiXMirbX6tB7qlG6vXTaWBbPratKlIazT0zuf+m+
QmfeVyt1mVcYMFWXykZ8kpWdnCWW8jmSWUXG80Y5J5+4N7mNddCCrQ5ECy8V7b8r
FYB3cAtAGx5TEDKsphgxB9bMToQ6hrjA78zy566/QqlBDKD99b2iS+ad3UgPEWZn
5eukfyOn9mhc+9PHkMT2tyvyDNr5GHvEF47NNm5uSsb+0q2HA2mUxPzh6mu4v83y
kkH3I845a/ignGfxt+w/dz8wrWhSxnICrmJr+oVGqRNFw7GMxLgeocDEOQW7ashJ
PP7r8DRV9D+6/+aKFRxXOHAbnjuwQOD/CHatzYUS0gstJJwO55ntJGr3zCVB14ul
AUQd5iQrwu6UcWJrHDpOl9pHyK3O8LSwUxlMMiNTRYD+xKkAcaUEsNqDlehvXZNm
NDK0DHvaTrMp8a0bFpHGHc5zPOnL8MGKDJoJkxQwBU73BX7+5JSP3DlYDJJfrP34
0HQVpF4HBadWMndvBf9xlz6g4IdW62Hr3BkFLPwJgUdAeodQHCl36ONLifWfe7G1
uyGpnWhNH2TS147HfZeQZf9+r8J86dsD2flA93G+nB1sBRQXAW28RQe3hRnaa2l0
rN6CQ8sofAx2z2CyKuNtGElq/G+EU3N5BMCkSgRFBwwgxi1IVkWzmisaylEjNpJh
0qfybyII/PXOunEZH5Y0d/BJQ9siyWkaDveMoY6IqyPNy6xbtRxfEAH8lyuxqvGZ
LusOQC9PFuoZk/EWDj18Q5G4N9mXvs3hgG8syCJogtJkJU+Jb+S4QbtQlo4oGMhT
VYY/vIdi7W/k5sZIuNFsHFhoV/LRU+kGw4u009L4HHnCJxGoLuRFcckP00tRKUKj
6fDHnv4R+2+201DyTR6ELbG0tZJcFHT2zgu46cNZhZNvXiUqFQ1HXwd/gw1KNtx/
hbYEmiaxya54CrG95JnWxJVdFmeW53x1CBmkmWmiYXJqGhpa1wLCwr6O/+msH/CL
0JxhGM59Y8ndfScuuCp9vseYd2ciuhf+d35I/Dgz5pK4WMu4W8l2L5UXFtuQTPpr
AfobG3IeEQ8xR+FCIeB4qHV+KVyDMSYiZrQq2AG1p9sFEYRgBzbAHJNWpL9U5Rkv
E1KgoxMmLEJaj5gVc1HJk7vI2lM+gS/HpwFbbt0IofuCSajNO99Ptf6j9HLHSqiT
cAIBWvLrk8xvgiFNGp3S5ICmgyo0yjCiVEuUnFXJMxyUJe6no0dlrx09ImCP+uKp
cS0A9ALOB5COzSJ6t8x8f6VtAG4EVcVuhnPbKyV6FQib9Z1+iJreikxPEohWly39
4pC3U3k6Oxp6aDFYMW6WuQHTUipQz0nGyn2GQBJNeJ9aC9vYlon/Yv765NVV8qpX
OL3XVv0D96YRhrapRdYfi8af3NlXmIQ4CE5nkqIIRXndtaZ7cjd5UYcdHq6u5pd+
AsxfHPYStyQvxHYSqpAPFN44irysUX9re0J+Ms7t+ZzPiMKQELp+GHhOA/518vpr
++HGOlfCb+KZHb611ZW3WwbCBion6g35iFfG4CbMSlN+iJi97DRP4sKaJw72KB2m
ZVrk0dccuY4y0xvl3cvbvfRc//8hyM4S15RiDLuDCgw1h5WReYszBt3zb6mFsprj
O55TMKoEzuP2a6ipZWyf10TV2Pe4CmyEFYK5F4v3+FNCG+4aetvJm78DFJU/VvOB
ociUP8rMUWgYJXgkLZFHPf/CUYcm+NAkzI5VQ0hvdDyHka8lXRQrcjK+69/+2QJi
eREivolxj5D9u/FxeAWQ6Y3Wrc7IOFiji80P3FGx5mqqmWm3HoM6W/M150d55fBr
xNGXFruMQTR7UhHUF28rfhQFF5WBgszGyuhHtiG+DHr/m/38y55ZxzCGE0TpmSf4
qr2SqlH38SqzlosmvYtlpLvdf2/ZzGi0KX6wk6fAgQDhYZ8DgV6QTc8WBZ2Miaa4
kWQbBj69YCQ67aKJssurWuBmEq0pJlQcAmzmS9ykPhzQiLJMAuOZc8YfMYTlALEQ
QqNspP4m5e6lT3BQCe8oP5YjvdGsVLaDhNsV7E8IWLPJ3AbG2j4gnIb91DxfmA1R
+LohARzbP5ZedT+0tugGDcGr/bMnCy63WRe7QMpdLstjOHtPnNXOJ+pZXoH140W4
wJhJepCT2axgiRpQ7rYU/edCUGs3wmJprAi1pcsF50n1r7cUiCrdHrXJ3c1uFFtw
yDaQ1BJfzPZxe6OzUSuvMKzVgKSrXDDAFTNBnC+ttiNJE8olmlQUmzSEnYd8NR45
EFW0UE2oMR0wEUOQCRKl5rUVyNarNZUOvkbyH7xykiYGX/4tR0CGCf7VFgEiNcBk
XdRHA9UzWr+g31XlJnoaLAZKbyul1eN/0NTyI9upxtlKfP+NNsfw9intIQD9Q2ea
EFTSIntpzoihgh8O37q5L9RSKVUGmblO6PYGTvIrUIlHIIVfxC4plz/YqrDMxi4E
9Y51CTNCpj5n0lMwYwLgcKCh0mNG78wQ3/MUiwJo7dtmXGEejQpzyf5BNuehp+I0
ln1y1pNLLYHjvYhsMZHiJovxC6+JgtJ6n7rmDbUWUsKEiHQIBRntfg5cY5TxgDv5
MF2iD13c54v0RpBpsJYox76AvcO5765qvsGsgwk8UGanQFtvfosFjNw5APW7OAM0
xixY9YSbBF4yqWuscdkbuyeJl/2SOfSxCL9IDB7qCotmnAuynUSHsnwBH14uak7E
gIWQqY09x+AidQAbTeg8PwMP8XXqCkrEYH9OaKKoPskzyVipT8XhJT1bd37L322f
PC1HgLy2+HzwE0ozNVnZN4/lsk4tabNQGHkzOssFhOCIbD3lRPkV6egzXjzUERNU
6bPhfbDQ2dMvcm4tcYBuRZIzdM6F68X73XV1jEhA5hWM2N2blJUUGJETqyqzzCx5
SGleLuXsb8SDFE6DirOwEvsVraShpMBk5unN//TWMxKbBVuLQKB+sxAMiIakbg1l
NNF6VJkp4PHU9DOGr0sFaXKVLtkzFV2QPMQZ+K5pJTi5tFK7ClAKczzFSPZi00Jj
C8vufeAzxtSvMT4EXL5LaWEtmT5y33KLAAmfS1ootUNXdOiYLkI0VcvQypaEFxNl
uJnTpcwVNQl1u9zvodSvsJOgKCDxEmFLa8m7Fpe1OgF5Fhqv0TTZqnxnpMGCicqe
9B2/MXe6nJmn2vjWptFnkd5HlKSJRV91XjQxIXD9z0WGWSnJQt7QYYUty8Enyo+B
w6Vw+L9zMr4lLh66bIMleLH8M3eItVeamOxIu52tznRqUKFJMKh49NItEONdsi0O
zPelAr6PsVe6zCQw5r+qRUfZxhTLNVXPAezhBTmpinRxGlm1iwA4uRCDEF5NzzqW
TycL3fs1tGpEE9YjJH44SakIRZJ1HVfxqTHe7FuPeV1UXYSXKpPWLC76dRWrlpJg
sPiW4Ll4UHU9M3+bTSeDI245SxAagmbWgHLiYFPAYvRIcfZTYTcI4j81O1ZercYx
/Cemq40hMqeBGKC1GPrS30lV4SrZ33d67IPm/uL6sbf2AS4LowpczsN+WHoq4js7
iBSm9KNCkd7FzP6X+wje9epdqCK3tunYnMkNlvpM1i/ujBTkZ3vBoqimyZPLhgJ+
2+NzQfRqqaChakdrKiCImIlMQRAbkD8c5HmBJlmrFh98pO1x7dLa78fRjGX6h4rr
rNf/h3E+XPGJK6W9frssFDEHpx26QAd3fxpKXdPpTxHOLWQTWeApBHYJRg+qfg7Z
OA11GKrU02uUOnuxdtc70PPnqw7c1CsZjN9M1X6ZZlZMKypympflsxTdv+nUw/wd
CdHvhKmJ7KcONPo0HWhZjiBv0t3KeN1qrTk1rU7qm6Ut6QdMUXnoK6wWhMMuvMXQ
x9vMPVxclE2qSbCB5Bi891VLsgEzNxg6pRsGP9HtUyKOzgtcCTWC8p/Yc4ad4lW+
sD9tRaDZQF7AUr/pdNd2eh+KXIDZ7SdGMr00HBjfc8qIl8nJ65+IUZbSw7fviIt5
kWQEzSGhjxQf8pX1d4rA8S4O9y1ItwjJS+KSGj6xH+nwlTRMKa2WnV1viKV+vzp3
wfixa9+kd/GAxCdbkzjgR5KaDSt9wVIRDUsrv8BprBYi5/W2OBwBY6H1D71horNX
cJBKQgS3Mcyc4UmGmZUPiTXxZJGzADycc/0hshbls7wTTNsop9I34SUXGUs4Wyw2
nBfEYKdjJ6YAHlGPuZQ6cluUY0p2FSU2ZFs//Cn2NzZsHpjjZFPt+Bj74/4QnijZ
lR/N6p0CJ71x5J1JLnh9+qco7dBw2NFvzIPYQrqjDJK7tgvAvgIy5cYqEwB7DBig
oMiD77gmKxmDgP42xmmspI1mrVeAod++ArRFehTem0k1tWQeoSkcbni6z74nNMZX
cljnVeOeEVoapY1jxr4DBKfx/UqczgCDIWyuK6iewLzuRLqjOpVtlGgYKZos4a1P
iLbsqKwfbPsgHMS9NHNoND3HA8Gb69OZWClrqk05wxz93fwr4SxmroQyzhHEF9lx
IKaZ4XKkjSXCNfX3+jwprQBmUIg2RMGlvHPhSobE1fflqPoTaCFgcGGtOAjVu71d
8omnD2LUw3Zp1wwQq89tyMlJh3g6hpVibUNEK0trerclxUL9RL/xQFQPzP3cWFYO
DhSTQo1a/72bmyWOV8714RrTe9SKmNrxZVAkfOZdEuNtoiku9TBEemOAYwxH8rpC
YLSJB1HyrsXTS4JtWQl1mDr9pLKOTdRjKiPDUQtr8iuTzUtKsS4dw2bpOyRnOX3L
8tYwCIyXdGR2en3/1dTq4mp+rPAxMCCJa+NZJxmgVSM0o73wj3wWzbhpV7p7swvL
1g95+rIdbkAjNXF73fondr4P2UIAhffaG6qDr5zQbQ79RC7P5Ynki23re6Xr4XIq
m4EUFCY02F0klRhpaeTdkUdNmdLz2Df6D833Zi1cGrFLp9hcxyIO45HrGFj0txqW
DvswqtpDoDxz8t2SpGO22vLL8uUlk7kANWN0Ka94TygpFF0No/YRX+cbxFCIjasz
S05cgT3RhMc97/zbNLCZHoDrZCsviS7CPoidujqRSt2+e98lkFRvhR+0XGWuTPHv
4FieIxmKC7UwfZgDT2ydaX3JD+e5qzsnBeSuZorUX4kk/1ETfpWikRfTjsQ7JVf9
AwRRDnCtv966ReYdwCOQK2vwLmjrGwrCFJSMwdiE913c/4ufJ9tChgWpXYxnPDn7
EKv44kXBnvmKQWlbQPhqs6NmFKlj+ideK+fiKCGuv/Rsp+N7hvc6G9I1nWk3wUid
E7ltOUSaKjCntH1bGvPhuu94tAFI88JJ7axodBeUxRAyzqGe1Y5KapO5q4wS+oDT
d0r2Y+6oiRwgRocvPvEdXuJrWX5PUkLFso8Eqxk+KZ0lRhFvvfrUy21DOOjYs22M
XoucmfS0KWZyBpmBUayFP0RefqTE9yqhUP12V6P28shhyq0UMAwhCD4MS3lQc+D4
TMeLcBGDWMx/8UHs+zxvrx5TzqWoxbrnuYO8dxpTxQ/6R9QE6sH/AiCnkvFDn987
j6aJ0DNf9mYaFI444NF2OQm3e1zqxh8cMGAi5elzri4SVsb1JtlyEpPBVnJ3xfsb
CXPaKdz/cm3DCVUbqDWLL5z7rO/KtKyDR1EsiU7OP5pEp+bFYugYWmOZrDPlOlFX
Vp5tll/MWzWGT+t7M/1KmP/nLlNtSV7LFVZABkEgI0H4mH5appHVj51FGJ9ChRPB
OEzO5A71BXOFhSESf9mE/0c51KIZLQDgOp18aJx3Gg8FOzYPT1sORJqlsvqoLX/v
oJ2OCxIM6M7l26jT1rS9QTW9yYce03wpmmXWrijf3ENVasAXmmG1M5nxdzPKVoAP
Lo4P5z6BeJ5S1v2nX7gL2EEr/E3XSQKjLfS7mUaZhQHcaanwnixnqIl7voBRb9wu
0lp2xiNWIj+UIv1jsHesW7UGu+AFcWQiA4QJfJXJUxk/SY8i9potcdPAzHUaY2sC
9ee8ikpaqZJoeEwWfr5NY7oy00lazHvHScL/ibfMFORSwVMukVX84CtjsrMeXbdH
JSWLqOXPJ1hkHCeHb3myKimEGqr0pHV5h1R38LOQmk4ETeSV8vA3EW4xj9j+jCqA
zamSpE4Tl07WIaKc7eQsVyCY0nrIGPGOLdMkriwRgMkC9gznmCE3XzIpfpxrbokN
rA9HKuamK9doP0+P3OlOlRvvTu262p2uKIbfuqbYnQ4UzqZ7rLZVMbm5RulBEKBu
rvzcYIO36auLplZgmP0ump57UYh5RFKtGvsolJasQtEi8+Vcv6gqt91W0nlqU2Gw
AxHJm3PRRx53iTAvNdpq32W+t70gR0SZsI85o8x8do/x+7hMikl06VKWM+76piuv
ZNPLepqAm5cAJ0NsyGN+WyPfsvwCgxK/7GAWY6YpwM/UrRQb9+mcT5duPR2UOx+C
hQcaGHlj+ovgIgM33VGI4nWHGNdckJ21+7DlVCE+7YAuKxeIoP1y6CnOLDnjegtp
CRpln54ot8S3ihcZus7AgLrZUyvWzah2A0wMpZS3cwQYN2CGPSGAZyvnStK/tVuP
M+BQbBgmfPeTJM7B57KGtdPS3zq0VcOugj8WgMstBs7xh/Lg75dR0wT/V/kDHVhR
JnD2tFEjci6F12VolxzcgkdBO36u5IZs5CgAt1c+a8/AL990HH7fLc8ILq7wLVwo
wq5ET9H7/GNe4pxocRP57PUP0kc+W+bOss9RB9AXPBOrGSDMJusrHtWquncKxzuD
u2OIj6HCZqvN0Gk3A9KMzg6Jp9e4AGnc86H9ZrEnZd5hfziIFhzpAQnCZ7EoRscx
dcxhFVhvyWQ81LZIgD94I4ITjx1oIyIgR3LQgfvBfP5Wg2AEmwsI2ALJbI2oyCAt
ZSJkMAjca5o0IpuTEjHuydtNbbKb99epUfc8+DTp6BQLveRlXd6s5C9dU5r3Mowj
Fvm2i45RyGbo+TjdnnBooVBxnjN1/S/XhLqQmxR+lGO9pvL1eGx15KlaNPG9gHxf
I25UNLZq5CxYSOD1LoXixMBVnbn/ZiEx126476SXq2iZs0BIUTrQ7KOgoWEbjx+R
7PpNebkHT5oLTFJz80j9SV2cPSKhNAqTjd/dEvXS6L5CQpP067g0eZ4djoLf9Yug
6ollKGQ9JzBmr2LFK4dZKOO772b83yVYxL8HNbUv8KLdniugzWY5XBQ8gNl6QSY3
pWL5ZzXaZt65hBgTiAMg9+CKo4BiSxVPwBKw1IKkZNwvyJ9kdRRXQI2pqmAxB1ce
aKySo4uk1ORghZTfl+Jd9u5x3l/g9VysBvBBPEnf5XMLM6Ga6XdIU6qW97dlPlGM
g/MyWJryJlQMd2gOakAL5jaYwVOpEXLHhniqDcXI6mFHpdlJ9nLCGLzwS82ZGBo2
3hUVbw7MpvvN53B6JNKt8Kc3rHlmMKE3xXWJJ+Of6i1sx7hPcmKla74LPjN8B5f5
FI1AZ2VuWgphSYVRdr8rYQRyCf/g0i6g0ateczcTiCY6hpta9HcUCO7pPxVgb+1K
+LNCAbaTqc0APac6x3r5F05IQ9os+iUvw5wQVj7iXRoB+vK5wNRa4Vx9QidT9U4D
Seat0vQ+hL0pnnRu4KNzes2Ud+4wsnU0hw1x8zxpzdQslmPd3ro/VA9quviDKGRV
gfI5xZA11RcEl2SKQ4EfMYmFVcYBPO1HgFmRcT8g4Uld96Z4zS8YNWqRRYJrCpvM
B8QvL03BPBZiCBhBbTrRAFxdI2kwTCAkzYaNJiXBOyHIp59V3rrhI8hmi2b6Na1s
V3RgISCBhpC194T7W7+P2VqCULKgDdOA4RsigpQIhvqCCnfwwReE8B4bhZAvykCt
kaNHoVc+fH3QZs432RjaWl5wUj259QxBeGAsPLjgrFI1YcPjfh8EPrTQ2EMm8K7v
TEAoTSqnQVWc0ilC8PiwLUjJy1w4CY+Q/wW0ctw8oxyYNmdcsNhGx0xpycKT3aaO
2005OpvCaaqoqheiQsLLyhaEmgJoaTxifvVvZz95INiY2DlLGKcYQSENJP88paS3
LfrUwmqxeXLvJx2g1mTWeFcaDKqrZE2+KryXYlmMzzwssuGAZLE1G3cg7sXrSdZQ
x+dEFfO9hBduK3oxeFL8sT+Kzr+pET396XTI7j9PvxdbpAvCoPbXIhQjv+HA/N+8
TRVgFcxayfzSbGN+1oBP/OXVKtmeAfW9nMGBksl2RCaxS/GNHLu2k1QdNbRa2iYW
KGQB+POCXzib1INxWcwhRZ6YfATfcaTeP27m6QlHvQN3rOiDn6iH5SFTr12mf5u0
vkngIAf3iM7iJF/LPRkaxqb/NYv0zk1dk68bvxKnUU6YqWEJomdgAyqmFlT5dcnQ
QQ3yv2RAUkWOgBAD+4KHX1Is5u2TZkmNi5UMfcEvSCbcFFJVym7+75lk2xQ5nz+4
08eegwnutFhASVNPZgVHLzl2dcmFNpzyXoXWGAP3KyjBA5QQ6qlSiNPIEq3j60BJ
qO+LkLLNNc5je3uHhIhPznxqyGzTNTPPDRnPqqlOzRKs6MeZ+X+b4R63Z5s5xj3/
PMLH/EGzLOdGWzSocB4LVWB8uJJOz0uDahB85bKvnrOLSFLEerMcn7Wp4SSWTQMX
fKaG+XD5rOU0mhodk91Qhh+HJ/yjCjnIo0BkR6CK/Ge4eoEzG+hz37MtV2V+5LUF
n81fzGkH14j6whmfzSX1LIIqRDi8oooP1gnmW1Q0IX2TiABb8t55I5Z3qbVgR4hW
r48hsxWnC8ecDD8IR4JpPPVkfyZVcNwn8ZChHFOdFfMXhMzjFo9w4Tt1c+ZAVsNE
kds+y03jd0Jz9HGROuPjIy9iyKJcRmxDcB8qyO7btZW/SypN5flkS4aIKjXtSuqO
tVL4FunO29QCscSwsjZd8F9yw+vdKFSv+Yf66u1XFIqZoWZXWuco1tQvpdUEDMew
iOKdCJFwI250hqrdtsqjVAEGyb0oNEEjD1nqZ0CA1RF6m4F26tyILqH5qnKBQL2V
UsFp8YBggvLyHH0zUGF1nhxgewPdbGvSQBgjvOn1mlqJy4o3mclnFaE3bXlitvaj
fsP7VrR8Q2YKSGZftrfznXTtkvIjxcgfjuieZTEwbVTUmKBzkmDKRAe+Mlxc+kZW
+V4v6musSfyq++m5T6oM/DXZPZ8N3U9a4WN2L3ClXwiEjJr1q/i7JgBfjyzE+MX6
dKmhS09ggKAABU5oSpIX5fnmzuaQKq+GcWsID5dp2yalBkFUBHbcwfbclTrMyJ07
T9dGd0rhCtEQuTA9ukR4shd49npkGq4iX/UsVb/HYzgWMdsVIcNAprvP4YV9jx83
5W88VrKbgUrCV+4NQVMlEYb2HMnSxNNoX+RN+zL6352q+RlRj9KyEU/dEPSiXb9U
HsYED8eHbrSNcGWE3MM/gJVOD+lT9y/bii9Zt5C8jOe1ppiSuUUv9aQRyxneAliy
ke6zu0srQx/1EOR0jIdJPzXQOxYfVkBkxYOBQwOmg43mrb2vSmVNgD14qNpgibOz
jThkuEQQoxKXnYnDx/flojccq1pt19hlbxQtpngU8Qh3IY5lCQHy0u4ECT6/n05W
B8LGIFqVwrtSbvPLWCNIndQGFiYotbWf+zklO++D7nLfzLX3tn1xLVBIhiMN5OW3
5PlMqlbtMgTi2VqnInjBhy8jOEFtlsIgKtAowU8kOgWhaBsAW9BZ0Q5aMJS/F/Cf
ApQTsIFI80N5z1bD/5FJRdLikR/kj/hRe53s8VY5MVTokbC1QVykGZhGRWNaYQDM
8zHtkvkrYCTTlt+bdJmVLU1uN15s6DwfYyrSwFiu5ULopeVwdPxzNNvegA7xMM2A
m3Zcj6qA29UQFB9YEqQaikpeBXWU1i8agYEq1Mk7zio1Z13CcXHRvBQfvVU9VYsw
/3nbVJyA/4PwRZG6SyRf8AkYxKvAEJRXrTktXRNwSbwK/BQih4WEfTv7FKER0oDG
PtlLfEitPtdg3/CUux8oy13C/BGiJeKdf2YA3TXi+S8JqsGbQldd/cztzMSFCNkH
eVVR+i2h9qGcwQ4GSBKNAVB9B3CLMu/c58zz9Tm0VVZV8ElrR4Rf+mnK5jmQY+Vv
+YvyIsBZ8sV44/JSftz4pxdSRs14ljwELAVTZvftRqgxWjJa29Pj8GwfSpW2FCOX
MNuUsKoMZxTon/OobjqOxpiRIy5q0HfEknz86uj+3HopUlSBClg9yqcrze0+nGI7
SZv9/k3NBsmOsROKGwDUtuAI2UaZlm1ZCZc9RXCe/Z2K6CkBIrRuGwOKp2OJAt3I
J1YhZtLN44w4VI0Yv3ymQQSJimKeQVPKtRWGDVeeRLJayErSyL9SDy8Hp7Uyqebd
LOZySIF8asCEYkdo08qkQPo2f4mB6zaUTdQG8xEwhDx5jiJKId0+5VZUHI/iWurj
KZJc0mE/nYpLT0HREaNW2WYeRrsVReVRnicEbM8FZbg8ZM7NY6OwK5c7lvx+qgXb
2LBh5A45LafsoVVOO5k55NrYX10csoyzObYdMvAXtOjInDqPlGhwcRZjAm4njNYz
6dyxtSsV1Fb5HlvJBdukOplVf4EEtZXby+tQoUQXMIYcETUuygL7jyiIDPskwaBn
DHFZcWf8nGMXkZYq70lrFSMLcDY9QpyM0SvaM6C+UzsEjWL2TYWUrCwmBebGUEHd
3BtTh3x7uAuKfsFUf4WC+ZZnpLWY2pkuRkHTrNtBt0xXasCXntqayHix07/mmD8C
I/Es7Ru6/E6pGkEjBODj4jldoGqZGUgWgbbEo2GjUDfZPClwzeI8cMKkwzq7lALo
8HQykTpTjfmnpNDKgzi8uMg51PuBXZ5nASt32t3soj1qtkCno7doSnSor8+n4Jau
pQ1WTMqGox2iJR6LfDcazAq9Mybgv5ZRJICoA3kSQju3J0MRWOnBWdIfj9aza+7y
ItCtlbdx7JJWG5Ip0sipFJBhV8kiRo8clK7s3U+14uQQp0II5IRoeXB70YIn7N6v
x45XBeFHmARm039cpIvh+mw7qyi8g4D/jj89mu9tEnkysTX65K/x6jQE5kKJuSwt
CdxqBB+HBTLL+bdd4c+X7B/4iGcQRcLQIhGHXOkW1rssR6XpSOr4rQO1Oxg7u+lp
//gc3eF9uvGDs0NHGCPWJHQBxlb1kOsm/S+wEpZkPkYw92kJqu/WK3E4sHaP388Q
z5WNuOP//mhsJOVKbI27US1AkMPBgucVB1qTmbk9RzpU0WSzHUc+LuDj4GWV8ppu
Y3FCYkEiiFZ0y7b2w4JUYdDcnITV3JDv1Ig7+3d410QWtFdi+3fMM/bdkqZHIcsK
dKscIyli4VRij2yqoL7dpQGMZKdCSTpxA8EO3vWNJjS/DMrOhF9mkDaUbK4n0LS7
wtCo1MfVQu7w4qhpLvD3Hwk2ir5iJajXx3yxdo50HW04lBlkjH6T0Y5uKlrFBteB
fkPy5B5jUKEOFlShSP7mivkxGKCxFlFmmtJDVU3kBgJExBcpJeOmr+231A/pmU7R
RFafq0V7qP/d0IRVDI2drwiSWmGNZxm2OW1uoLf09BTEACwVeR6RUM6BrSwHMGRA
cxrXm1tTCk3bgmmJJFgmOzM6l9t7Z3PQqV8sRt/kUOgogNqMnfbJ10XpVSdRoVea
pahE0yu7nPOvvIIgCICx1yTqUkFOWF+p7tZIJ3HrQqPXoHOLJYgxXS9eznDF4jyg
yx7GD+g18TwAnU6NDcXNHN8HF1zs0FLCYK+YcS2rnkSrGdtdlkeHdJenWmrlDM93
4MvSE0WblCVO/fKWr+vHB1DqUZqMC11nu45liXq0oXi7JaKwQRZdQyz8xC3exvTX
/cuHMLyK1VgTHcXjyxfm+7oZiLX5RAvkBi7bc4vpTZ9dodH1twmLksl2mr+OpI4d
nemUqSGhQNqbY2ZXjaWlVyb3NjGsDBSE6xfWMfk9u6yYFKaSKNvdMTlOLOnl+bxN
4LQMCupz7rbVHnyyTYc6IpYp0nAPEhgYrmRkxc9BOmABFmqFmm/4Y6zhNL5BCkUk
OOHVFbSvzPc3Zz2+VgZmVctjIHM1LYl+IVn2toG3j7dFT2+EOwFuAxfv9XP1MRLc
uHtT65isC0ZH49lL0LrItBG3ECMf54uOqVNzMp0sf67Q96ier/lHRPmjg8SQcDeB
ES3UDeMZluUWsw+Q6+tYr7R545tGbzEEWB/tkFlrQocGgjBFHH4+kViwmMQqLX6x
7KdFdlhyy3cjDFIIb+zEuDJhJfGBqZGGVWhMun/fubFPeVSAv+OO2MeDkMiV7BmP
wMagK5pQ2umO83vtO7kuWcykDhJletF4Q/TVzn/60kIK+AmMRmMmOKwusqV8sEyb
N4yNuXVQ0jmRkgaPUBqXZozFRrI7+9/uYvmFi/EwyAF1NVjQ7gjHbjOCmz1iHIxc
+kltg4rJ/HKWl0W2E6EUVJisfDrtQgpHNeSIL/A3gezMMsy55q7nD8VFctF5Fa6X
6VK0orjqXeayuvIphJ7VDsW3urgSaoHoUfU4dtUFubqSukjjGvGqEjCkHkwl8mLZ
kJIF4L4i7uEVdPj1pQ4+jSUJQsKXVTZ1Cs8IdgpGj7UVSXFbhk8V6GJhxzBPNsHS
2AD1nzjtMPuK9l+Fk/0Urry6WImVLRifrDVdOzSAzo9jk1zpG6wGIeQbO3uatvql
Le7O5tPv+fz0jycKuWccN3uXObeq8K+L4DhNfTaw1zgTDwQB5AJoIdZbD1ScA1R3
89zXsJZtrP8r4SDiwDEaFFQWGXilBwS4lpHxRe8rXOBuoCDSU+MNYSWeZjtlqPyQ
xggyial/J7WgKkaYRgeSyNJrzyPW4rBJlUqaolgGbml5mF1bTxthG6Wftc4MuezX
/KF9iIcJRDZ7SHIT/xYlv3MH7/6vCtPd4H5MKIc43vp4cJ+P1w83zpaUmuEfDc9T
qbxDRWYg7YPL5BbjSxzFixAxVvorGB9/HC4ouTtKsXdP0OtZI+tCJxtMeOpSyjXr
FaAg2q0/PxJjEVeXJ96MhVJm3k2gqTNh2k8SwIXIuZIghkNCDYlgW9gk3EpZ7i53
V1yKyotwAjrmiVdiN//Ag4YIV4xtC3kHfextbTI0IsF+bJHtv5aUlnIxxaK1s+UD
8qAXXkcO+DHdagvOlLEC8BoVcrJG72q8DR2o1Em5qJrmoZk+AlFKPJ1TLPMc3VRZ
ZfkaayVMRMBm8G22ToJTR5JujEXLZ7KNLVXgTzFffeIxhqJAQ/WeqgCEU/lx5Cmp
Q5NoHH74M+ZnvmvvVv4ajMXQLAHvk+HKGcPw3mMN+0oh2WOBosFO43hEy60W3WGB
Dujnuzz+Xh7iWKJ9bdey6aULCu1jotjcGxAdhql2XlMzR9B++w1+GBllGnbnLS+6
AR05jNrWdy7zLzHD30QXITNvOV/UrwGOk9Jfbrt+MyndnrPbsoAmEBcg7omVytJa
0i9JSv6cFYAY2f2G0vb58fiWqk4nseT7VW2x3Nx7NJadSIZ7206HiEf+OqQ1/M/E
1ufIAyi7xrvaD4umpuINdpcQw5P0nbZ1bkckHRr27/A1MVStflbYDtsCHwqVP71v
9M3BqZRogC97mh1WGfMOe3qtakT6ATUuznKh8iwVqJxqx6H3Lt+wJ+vDP90Bny7B
/xnUfDf3a1kG8m3Frj5wd3LUG7A8jUv0QPMyKwpigeyvixGyjjj/eY5l+ebwW8/y
RUrZhpR7Jez/2LROhcwxJ0XlCrY0f1Nc4s+ik5A2MFYYstyZYSyaZfWijH5ZvCxu
JcsyvJx1u3WFFSRLlG5gBLEX/PQBIi7/hMQpQc/npCKZhLO3Y/iWyqVdNQPbPtBA
zw/WbpxGLtV6LfPV8NTybjb+rSMgN4Yy2dXv2cI+evKImzIS9H5RgPX69k86qISB
AgkXHNjVMEH1bZqUQwlCU6E3G0R5lhUkBMmZp6M83hPJRC6MRVNvrufruPNjBvOO
SXTqHrpE95Sz8qjIDOKndkRqqIu7qyZl+H6XgLcDXm4zYsnYlNbnOoaba4nVakTs
mCjFhwf4DdFbxxGecbrYvZvXkOxR8PGj3szFuBdrUh2G2yBuxAyvumIX+nRqYA8a
IVlaRRNPNzVKYMjrG2DJ2fdqEW8TCD6UCCPwqlRgGMWx6cAGZXgh1PxI9YFlsAJQ
npSrgwv3/+uMshrknrN6mKWvUFc53D9mzgftkn0N57UbHMQkydVbPdbhpfqPqfTn
xzXf+Eu/kCEIMSQXjRUnzmZVagdaNfhf2Jbt1HZ6kEcL86HiovXk6e2ceVe74x81
wW8oP/SFp4H8YgRkAcCdiAGo5MHLdHjqkxc7vmur1IjXgV0eafXdscI+LeGfvDBF
ZcvRF2izRW4Mnzoso21/DpS7xR7Jvjo3/VFkDTzZvhJisqIF0a53H48hsOkA1RB8
6IpaBwOHExtobEfXykOv8okq06Rywo+XAea1nAATEavzJF5HCvEV0pNChRLVtnmj
F4fqzEHtPrAQt+Z3RM9BMlwk+zSo3icVm6Gf2cbmS4xv2w7Hm7+UvpnRi8LbaZeE
UdRZI/OIY1jqVl8VLckMNjLRZ1btMtHqOSLqbWq13hp93ATMtIOlMkMCSZteE28H
5IKO2Do5gHDqxwhXDGrv0AM1KJipoztwrZVgspPY8byG0KdraT/4SBqcfWIjRel0
tyLwAJFytDBv5zrpSN5OzenqpqxndL14TeEVcGTmFe66VoPcl+tsJH0/xFdVbMUr
yzZoYAXevK8LFMw4Vzbuv5oCgim5G/8m+gETX7LGxHkZ0vAYnMJRJh6QRHv/GWH1
X1Vk8M1+qrruQTVIiVba3Xk8HFKpiwJbK+vCPjfReOBR/WADUrorxRb9KqsmjUL6
F4GT590bE58Tzs6XdPVX4q9dXboNbfvgeZK9TehlncewB0viu0RjgpuwyG7JiwWO
G+yy0apCQCSsmZPtdOtUnuG75vYEMnDfiqnlA4LEsK0uZ81H5Q6i0LlEOx5DPtXf
51DH9D5/q4FstY/8UE2GGD8c6Lh3xSFVIcpZTNVo8tEl6kwYeQDtueqY/ImeIKS+
d3Tw8SasO6NTYwv+XiXMTDNivSGWVdjp7GkJPOtyRZeO99aUolMprVlvhaj9uTeQ
Q5h4Z7pKB7YCdfudczInQbG65KWHhlltG4Q3rp9Qk0LLl9eWDBElX4+oF3+aVKA4
Be3N937PFOzlHwYxOUbkG5ubrY664E1x+vLQEHN7DReSBDuM+R3Yf0g55NH1VTfT
rzFq3ILi5WYET50ry/zFPaFimYSf0YWiaZtzDBvbWWS4FOmkv0b9JE7Gsii3QoXA
hOOLBQWRRhD06WWWhPgvqiWe9NhIYAqrs5i+sxieltLdYd76kH/U9C3MeKaM9ZGA
EDfbysUZI+k23en/eWu0jgtt3ijyf8WIo5qZvE83uyZhM3Nvqfd3xdONv3FjiBdc
qxR+WzHfq17mXmASNzUFLroAs6+9ktfNGc5/fqUETscRqrdldzIG/sc7ZxGiJv8P
DX6jhLXYWPisULD9cOVOx1Zbl4x5j0uKe9yhJz2nG7dMJfP8/qs8SKTHKt9lL3fW
BhRoFKC45G+6PZDeuYI5aH1ja+9pzNHJc2CWqwwMim65aWHPYSTt9VM1D8HKXX4m
d3PR2h1fsgCZltUh9AKf9vWmNIV/589xLuJjV2IzQQ2t51+Q6yTWGRNvZRtVJSOc
aFTgSJWhP3poKUqUh0sH4Ej2qcjw8axOZYdJz6bsU4Q9Fc6DevTYS6ymPc8o7Vie
dILl+AKBGrM9lrOJNlL7UalMxvuF1kq9Bo+oaXw1aGdPqZ4t5p0VMEjiIdFpcVT7
dkcvpzb0c+VDaK4jHqHnGf0L88GmnUsmMq1cL5P+n13YsXG91EFhPSJvkVZhB1Xq
Wm4IiR49KqOnR/WDM3+5aJKdmo2NT3wyqlNVN+OOe7ox96ap17UGknyYqIJjxVBA
ROuQlmeCzYHtzXQrFkQJtq79aqDC4WzNfQ7lPaTcaDa7M4OBrxSDLFmtDI9jVu8i
7DrylE9sVg1ByBgzJiaNOs6gECYMZDpd+0fuehEThkOUCqPNKuehGzGPBAuzPWMU
NZGGpFJfCg8LWaHdRa/LS3wPO8sM2aqi53ATqp3r9hyneIx8oB7vDT3/d4jRuViG
wpweIcDqnWhhsPoprwcJ8N0L2BM/A7k4Nhn13pvJ4kOSerU27prXOC3zV+1+Xecm
G0AztPDeEWsIBY56BMMyZtjcJQdN6bdd9rURTyRSKmC53O6U5+R24pHqjjyvDJ0E
OrAhH5QAdBDVlerM5vfZulMrrDc2PsHU1zyT5dP467BHsyYzDKT+y0knYKSReuE1
kQBjl+z7ptzaz8RQf/9C06uoIIXYlgF6L8VifWitG7Taco2aaDSsHCiypjjZcfoV
RILYFt74bYRpCW+wfSqALaMo2ieBVXB44bshcyJjKIysRc6CNGnv1F3wcuMFNnR1
koU44Axrj3GCIHvHTHPpyNVcSbO4SG9eah+KEFBRbsuNVmD9ahSoxG7e7Rs6JDMV
/tjavAbKxCgsESs5MBYzWvVtvaEZfSOE6ynommkD7kqXOqC1R3i/jJ5deMPOf02f
YA3OiQbBLxbM0R2lxVy8579C+wVeO7mWT+3cyeEc3kNRXGmwgIoR4ON3R1npydQG
hOUC9+/psdRfO0hZIrhYPEXIkeuw+MXMZGSYVm/feQ6VOLEgEsYDm62oMAfEhY6o
0T1q1d7WsMEZwRAmdSU1pGGdXqkx6wQtKV3wHuhs0kiZrTEZ/whe8c4khJbuJ+OJ
sjfTOaI/ha23TEZYr/oRz097UcvtxQhs3jbshM4lsw1SF2CRsVKUGVyv8emPCCYi
z79WNLth92ksvN1ye0gq6pDD1qllPSWjK6Ohg61m5nx8ojsLy6rSZSt8ZSYDj4el
K+zLUrY1w2pD0DpNR3Ynw+HJdhnZrI926sZuQOnBQE5wRsxvyEh0KZO2a+WJ6xfy
bhbUowOKVvzI5ceR5Kxye2MGJ60KlXlgs8/KPRSd3WhjjMheZBW8bzomnZtfSITf
ut4uSDBt7+IikgWbnR4yx+z7YB/1uR0hY2uO9DOm23NkkToH17sj1oalnz6JaFs6
2SG7o161A3dZclmskctu3eksmX97G7pdJHvCBpeOucf2Tg2LExhZa0z4BZuF2oUD
3oYPtusmftwTzhjeLDR3RbFhrV18Mwsa4Yz8un1mXSdTvIRq2V/PPDi2QIxVUxjN
N3sgoS3r5ySzsprJi/P/XZznSv0izCzuybYQY3IH5ii0xCuJ7CwotZWq6jF1gOsk
mV1oM+tcATySpDV2dO0q6gkUfcdEUFJ7lQiNNJ/ZBpeybM3rX8Gk/Kr1UCclEqSM
6bbSayJZJzp01fO5G5HWvvznEFcb6pHM0HuYN8HAypbhdEr8FGbHQO92rq0+0qn7
3f7nsabJzGsxWwzEYEZ96iZzHrp+tG3JIt82sO283ss0XEx60zylykzAplN0gjjK
JoOeeEhU98u3dkCL6PybUfrWZJsDHZfwVCExJg4adtdbDePMPkxZpNKPRWRM8EsN
mZPydVvc4knfnNgEYfPo6W4lLZEbiR6fw7bOAXdaoYndGchB2q4WiFpGiroFkNkl
FoqEUcdsJ4UZsoJQI7OEAZt7a2FDDErC6+f38SlDZmSfAhuoY9ld7q/E9bYZBwL+
S6zeQSV084TB6qym7kOdn/MpztSxfBbIlVgt6n/BWxZduQ+W7FxfAi5wSUTEBVa7
1jDOrjIS20zZU0vAb3/Xhmg1ORFeFjamFklBchkJx3Gu0F4hisJLg7MvLoZC3b56
ZqLgurfxGcz5jAUjX2tZHV/EMGsJmP8LdIASU+q1vfVLzQWztgsgmhHz+z4evIt5
XVy0jxhbweMa1j2HjwfVq/PZCDsIif/8kNrk0OfNuIsjy+7yKslkuTZ//eRnmjFu
C8rMeg7AwFWqKvcJM4+vYsHfNnvzyyxUrNKWRItFmsGI8SgdemMkIhgCgwfY/ylH
Vn565VK4vtdfc8FbegRiJQ7e3/nXuGgTzhKm3DQ3bNCZmXUxx+iIgbEEScFesqTx
WpwnwltseDjbKjy+FCutupM/6IB4B28rrEWyKjcmZSsShQtq9EjlNGrhBjKQF/8U
DR8uTifyxraD9ZzqtCwHYHyaPsHJ3JSX7WCp1Xahopn9+vkggzi0HctRRZoCAp27
OVcqPwtMiIOKprfPNAGfFBc66chKXL2BtiKrvGYUL2jQC+l/KVJyXK0M9LKsxsDb
+6UTa0dLVoQIFDqtYD0q92TniA0jNlYg8IA4TiEvIVkijvxYWl0rDpU7du3Ya5jQ
o8PDOEF04myVPY9RZzDaJfHMfLTtWDTfDYzx5IMDa97blfpT9GrDaW/xYaDxGRh0
ddDa8dhOErYMPANnLJfW9WVZCN0k9xCPUvBWVT1MnQJgH7aKUbq1djZMweT+Gc1k
Cnqka1+pJArdipfcvyU7EMFLic1Gq3PvXs71a9y1S+s2G3pnuns9LVCvU241smXS
EWaaM5QijOhFkGUe5q6rki3uTqI/7WO5oAntOGj3eXv2IwXVqr1tribIBCxfeboC
XDP2scbwx7Sy01MzFAo+hwyl35gpfApjO3sSM7aQavFGEcBtzw7biKVEweMbsSIc
w0HZ5g/O/oHl/jZG0do8h4hkc18PG29tGuf5lyBvjDTo93rc8Up5j5QyweQdW7HS
oXahNier9OtZz2tkkfeW3f9I94BDSf363l6hoZqcPQNEl+wGSaOCxYoX3+8N8rqO
3Kih9xHcTtTb/y5XpJrJ01IH3vJ5QCGRRIUO11hSHe4oGuIAoyCkIyV2bpgewey4
h9T0e9giBzEdCssb6epTb33cwavVTGFRVns7QB4PC4DXNfRD1IBNXdGqiYT1WHTv
srwgJXuWmsIu9BXn0WdTgqrVuAYK3OFBeQ/AJxhHsjbaWNUEBPL6yIuOz5d0SE6K
JETaeKw8QZRH4vinovgSxpjf1UlR3oUnCA/AdtReOXqhb9mLDxjZ3aUE44WCoibl
QshfyB+plzK4FsVLn9wmg+cOSWOUzT2yMTgJ+v6/6hILPGCMhsfM15OV9eq9kFP4
e8+HgPIsHtbYyCt5UHCshCyEgib+K69WdS7KqYs+jPCf6CJEh4NGAxhSOp24+/JU
hXpVtsxylnf/K78tucfC3phuKKJ0PKzOKiWdC0MxTjvOPn5OzR6Xp2rCmy8VXZGc
UByU/QuZau3MCdU3HD9hrIgOxm3r3v/p6j4XmnnkrXttiaAgaMIenI0sghKAun6X
OkRGWHDNFY7H4xuWNfrWGctflwxVsJ6lMzTWIwfdy5w3+vdmeeo6SfOWvZS2654b
BsEIXHsvQz+sxagXU7jdFPFgNbw264bq5r2JoZf3+Ox+jhYwCCoJA5c5aojse38V
nra0iCDO8MXCrX8jv7anbPTYM8pxc71/QLtFMYZQooe9YuU8lr8KP/c5Wfh6uk87
Xy7eC6OvKaZf2p3FfCQfExJNYZ7UZfBXKC2vp943DPsEp1zg/MSp5Xqe39DkYcfB
fnPlDKxm7onSt617oc1BTWQ8VeBN3p6JBZo8bms/xAhSCcftOM2AJ1m16GZJulXj
1Wq6vzE4x3LH+cHF34c7pMtfhmkv+cydrUOWDt9YoZjqSNfut6B/NflyeIKdWcQv
/SEVyVKyLMv/AL9MrzzSXOG0frQkgX/5sGov8OxPg85Ux1vPaTgxvJcWbNOjbp0L
QUnW5iNUY4wKJDiGeU1NoGgZiaA3rK3Iwz8PIQPB9Sh6DvJ3igbjgmXSJC3Oewe+
hHQ0hnkKTYxYFMYgHAadBYLcSinKJmwuNufxPBBWEkigBIz2pilFEilwWq7prA9N
vyetbTb10Z6Khbeyhz1cLVrEbnXNn+BrHQ5PXevcQRHw2ay8M406BcLQWMb3V0/A
3MaZxdldBzUh8UJRavbB1Ld8XagZFpRIYbVSgGsA1AISAbBC+wN4dRzTWIZAucSq
dvJnrDALp8/R07+F3rtxpemfUPT50O+4b3HcTJ48LMUNBarXtfs5kSvW0mHaZ4Lq
QR69a/wiOuRGdFomd6dnP/p+KFhLTqPbOqVUR7WSRnC5O6C4DM5V5/Oz4xGg7nrW
kqBbL9OJbPw2KoxcgvdURHJeAfxlDUPbZ9JLhbmbkf0IAdUDeeDi7hEbH3ZgXYkT
VtTJRA6UyBT+I47XdzHEAxouHRRb/BpYhc7oWa58S2k79QtLly9U54QQl9l4ikmJ
LGPGq21buoZ/G8ck7ywWjUHnOSnBg2nFAge0kGm+lw6yVMEAvV5smk055P42nfAp
EcTGfoG3dAJ4+GQYM13uW+o0mAdjbH3Lh58PJom3A8Sb2zVnrNrmSwOk64aRXeGo
TtNxeIT4z7a28Gg0tv9UNFZXYNnmqvZa6Aee6wYjAAIhNBrFGcOXwzv+Mgb58E2v
I8Hti+3LWCWvbq/BrHG7ANt+Tt9lHRRwY7ctFdgkhcvey+ut8trP+3H89NBngtaa
fBlZsNnMg9O7Vimue60zAk5zNu5JkGUcxPMIXoSDB4zBv1sT9oc6UHBNhCRKAt3K
8rD6Xb7aenKbpgFc4720zscbmJ8elKkJXkJrL4+rYr9VR/L73mHNVu6nUsoyUj7c
Tz+iRXx4nFaEJ6hUZpqq/pOL4GlpQRmIf0NNousNm7BvU7vC3ihnWYGCYDkjQCqW
iF3w+5iRHgGoCRf4O4FG8zZ6Xax86XzfJkwDdAURWKvRBIc6TuZQ8J1Mgn5q+phT
Lwjz/lQAJB2hN7iuP9disApQuXXyAJXuR0EWTuEpV5e0eAL3YmY2Kd2H7PQz638J
vqo7BTROdlQ5I/DfwTbLSnWzjTfFzPffBFBblITW4q1+CMLjd3+r16oLxidJAKh+
UhJZrtPhbaVx0IHtduEWx6dmuLeGYh8ZRFf2DXhr5uPdrJT8Lg5vgEmEWtX8KHdZ
2cZg9f1LbPVjNjqZwH92LCu9mxSHkqbHD0UNZTVILV+umKkRSI0Mg3QlAr9kGzMx
ewbRcYMjeQhQio3a9eRlRjgL09iknAsAqZrEdVYDV15FgRvuzBLU6pRLQE8Edv5n
0jIvq8JyG/P2i1vcp31RwFX38hBdA3NiCBXkTvIBeTjiZ3GqrfOTY8IhCBAsBC+7
hfeiog8CsL25jQguGMI+f4UE/mSOQWsYYBK1EtpgIb8e7gMmpsW/Zt5Gn51LRK7C
U72OjMZlsXhM7+gkZDJ+y35vpQ9bT+ITusGhBNdlsAJYgjIvSRNIycGcblX7m2ug
SWOLo9UcL66tDrKoNfHYX91zPeSkAeivInN0y9LZTOIKXf6xR/oGhPJ9KTlQZtzw
5rLYuDYaTcvUvANBrpYC/V1kXdiydbO7JD/qHMwQbnQ/OvEDfrpNFVM3uNlHGN8l
EMraC+1SLYpxB9KZVsF4QTiYXL0waDqsycY61Pi818yrImHu9hxBKCsMgq3groSy
/bVTUM6S59tNQ/xZ30N1jIHKE+7Z+Yh0bKSA5dW8TTd0/6ZL4ObpoQnVJdbIP4eL
bBy3aeEDW/AtGi452nPNRAzU/rFrFZeKaqAMNhSGD5OkJVoi8FFRxo5BWv6NVyP6
4dJTKBBcW8pAeZCPjje3BP4MHOQNn2eWYZxa+GEtdmtx/HC/4ZpXlb8LCGwIVqxl
ULl4LkGX9xjB9mPw7SgmSmPSRi87WUtAb8DQzexkoMz0y5KrjStODIt0HWTLygdw
5nTs1jxFTuoXWNEevUtFLeuOFRsBTmAkxxjF9QqSKGMxH+MzwqFJEzIzp+Rv9TSl
OQzuH40jPYn0aHDIPVvEPBCTK/GaI7b6B8lvLICiFZk7/M3A48SI6mdth19LYIVD
JWGpwjMHqbPHnl8k7bcl4dNID1EEB9YU4GNXSp+C6ABMLhpReTyKtJxCT7zyOvpZ
aiGIIaEtpNtcqcjCsxpdDZmvYHzxRITBbAfTEfgP5Wx6rJQTNpGgR1Jg7fHmM/Lg
Uv4QfOdj6Dhx0rfQuStNSitiKRUHX8iwz8RrURdoe6jVOujbBNtBj+L8IO9qWNz1
Of2BiE0tait1eZ9/pbnEZFgRc7mcCVTp7pA6btgmr8vKVjodyAp0/Mnjgqmu2P3B
J4lhhgcqFl/9v2zdZb1tnePdyaUIDqrztQnhS7BuCjEhC35s8q1nqlrjC5BPpgru
xyBz2XLhyLCAisvxt6lXANvtpZQ4U4lxDX9VbzsMpPoj2gwblcPIKnPafO/jZFL+
dE/xZXgRekqWK3ugM0Ezej2ylW0qytQXFQzJuOdiMthchsk+VJ+LOp0vYlldrbcQ
FAGLN2VCdEs5nx/8KLlR90LMZC1cOpgjB6Nmu8KVQk9Z4zXJWIudOGlPExkcXz0n
PQwkLer5dLXpq7qf0ZuHulVQEsN+1++XeeaEtGcMQPsebZLG+IBQEWTk7rjmsqno
gB7cb3B8ckngzIXYXU7UuPwnqXbbU1+oGRgOSqFmFA2TWkLTK/VcIa55eLfCXn75
yAiCJB8O+Ik31BMy/T2/U6sPT/tfT6MZ5auZEcpZ5dwdaxGZFosf3cUoteyeiJ3E
6+OyJlIy4efPA9W9vx/68zFp9+Uv7FC0lG+EfwVIvo8KEVTLPq1kumT1zRLE0xS3
2QwjHGUWKf8wbaNLBttcv8nlZF59RXuKHpdXJmdIaD+j+y/MY7XCSzNazpnK+UDa
sx3ha5KnWs9NaIWhFeqfTjGNzlSMu/0/kzFGHqpSoqu0O4AMu2Wm+mKdykYJ40Ye
lfJxIl+wZOi/Hi7DeAFexCNIBARRKUm2Pgyy6397qJrjzoPXlJJQrSuJxq9l531H
Bh/MT8EO4zmcPPgDUPlpKpp7VWZzou2CrswjQeDbl8nTlqhUUOZ9wau8TM/HdH6y
FKjD09jQ2TUHhKu8Vtq90uxH7gqMS+NMg6mY+/VEeK6Am90YxmgJOZXTwPMaiZiB
+TAkt46HINmBCFoffh5gbg4NiAC3OaHoLDOIlKh2eg9DnvAYs/TgsSxAdeg6R13g
EWa8ZW9TDIWorf7HsUfhDGkIsXYLND1k/BM7PgkZ87GQ/mdhmFkB5lun01jjdSgs
5XITE9Mt4ErzUipu4A/3Mx+OVsGLVYyM41Pry5hYiQp6AhM3OOtzwpwPyHGI++x+
gJPBZUg6WGpTNvyMUNey4ZyEwNnHq6N2qt3+sL6mAVIHNduIyIcL1pZGVORer0ZU
Fg4Bg9syHMKqfN22JZTFKH+kUItQdETRBuP65BrWyduVZMIhahZGWvf13i/IozMJ
aHrV7dHt610STIq3tPAFTF0d8XWMhQ0DquUdjdmD5LtzbFT+PhqYIAo9pa+I1HSD
o/AwDDx/ylB2jeRV3AXstDSkKYm7rF27RAD1becwJ/yyRT9OCDO6SAtOld+tUgya
Pjq7oKzfbkycTxBchOL9a5f6YVYHmq7ddOtKAVpO9pq+3Sfd/DBh+utNZLNbp9Xs
KlQKoWoWcje3NphKPpVW7ngoZ5boHZGlA2pIFhN4EJ/xGLkv5TznUacqIjd/FxJS
Ac61o/dWhGi+5r6vxjcmFl0yFu3iEEkXK3LB7XUAeRmZm+xSrPHz/S0i5nN8S5zF
G9NMACf7sSMSpLuNnNwkwyWcomONgXRYWbg73DTAL+hEwEYQq/pbnbm7uKLfGHfj
w56E7dmfYSLSfBsOHWSh7x9nJiX1YL6WnZ28jpH5+4MIHGcv1okCLNEbkOPoMl7Q
ptKnbzIkSODf3WA9Qyv0uXumNpuysvV7TBUFtYZezDMbpVOcXV8AFp78AByaTeCI
B2VYd3v6Edn77RxVSB2e4lnO5kLqlJbpo1APwUS661R2ry6fS68B+7xDATHLqLEd
ef95vtpwcV6bxMumGh4DwE9ZmfGoHUUJ0mZ18ZwWaRC4S0bESBJHi6SbQPzHUNm7
PrUmmGZ0/M4pj/N3fs72SrhKeYuhtcQOIyJdU18W2m5vIID260oorwGu41ZyRbKp
uwf2/1SAIyGDi9hN512DDqFfe9da57vSeQ0pQ8nhxg2nSyadZ/Nsm3heSW+J52Ej
qlM+mINT/5LDYlhs+oDzBJz8F8HZz4ZrXaIdFexjfI3Xx8kIVeUOfnLcTrB0+V+j
uCETFegZWTFs6CCCHTCV33ZMH+4pj+ABop263mF5I8WrrIuy5+CJcs6iQeEljpwI
gFxfLiKqTKUJeawbFrckUeA9w/kNVWHduZ8Ed6ld7UIqkveP2YOPlOw8lsqx898k
D/K3N5d8Fc/J1JaXHnHATKery7QVBGzs+5IGj1Ewv+/kDA2lPaMU2Ug7ErlzJAOD
ZxkgeMcSX/IGIXGf9fS15H2M+LyIYBV5fnC3/W/PlKS5HAEUCpT0Nryg0MbfECAb
qnikN6kbw3ZCUJoGcWgKVJT1DdmvLweLKvkEpax/U1KYNagEPPw1rTvaY9bU5qud
+BfhMCGn0ltgr4Tq7bV4/71t0VIMvmt5lngHvWtEeLuFeuux0kGfdx5ZUA1yIKjP
pzdrUCMe7OKtkpLV7bQC3Odcu+Ilv/WGnT0Amqd0S0rDReiFQaKVsVj+C0z84Ino
CqEGJl0kQxU4bWJOuNNunKzVmVP6BVVPGpTPovRvEPKDgIit7BR7W66w15zZjbiC
8CpjpQyCJ+EmlVQslnApscRMFNtFizdMo0gtDwm06GAo4xUrnCodT4q8D/husQmZ
+KSmU8xnapHd9CjNnj9Do8iIDsa/bD0ivsRlxaMf1HhohcgiBH+T/GthmFyPYuTX
EAxu6irguKdAl/CqNtM4X7Cx4yyuAg0+0Qot40IopRCHtsyBG3N7ZLevsDwAziSO
M8FtF/xreXVAP+3UnMZ5vdzO7nZGZE+C+qQQOCBPsAfFpHX2MOfvahuv6cCk5fcc
506zoeRhzySt0VZJyryrUD0VwiUZ0swRTqM5zDLUmb+K1fryph14dCJDP5/PYAeu
Xs8Ys559brgOtxFDzDqhGbbt5M+RP9mfK0S+B2Yko3k2taXN5i8vyME7FNKEn3NF
Ofbe94NkZ6aWHk981BcTvWaxl7SyTkZXVR1g8lFm5Oip4+alCwBmpiuX960lHU/l
NuPPmEs6/CPu7DwssRXFC3Cp39j8SWfi4yMJmS7ZKrnqESCw+NMBSI5hNCljdYW1
DyEvFkbkGCyjTKu0LL/2WArFG8wRWmKKQE3iE3OCj4aoXXlDUij5l1RTilssGVWe
XlaTCy5AmhTrOKN+lg+X70MzsBdPd1muJmu7oKDVjU/zCmCXc7Wt0SWLoJww5uXp
EEak+IqiO4Df5YdJ7JTlMFxY85S0QtoD0tRtVgPpsMmcKGS0uDgrSVMHlbOWKn5k
a1hn3pKZeH7rNX+S62aGTixvixZei7MRwzrC1MrUUMlLTHXCxKUt7LSjUMzP8Wfi
GGDKsITp1g2T/6Tv30lQYObl8tBa4jaYZWfXGH2+rHmHyKVTFsvXAdHT7poIvrY8
WEeNlS04G10j0DSm4lyKepW6jB2Ftu8ATfiyygoWMw+KPimug0RqDpeLbXn+BtV0
2JEnvcOmN1owO8WDCgi8tre+QNpU/wNwP2s5Hkny8sqVLDoEoeP2Tfl4zpJgZnjX
l801g2RSZZwrOa0YBNyI4e22kgmoQmwVUm2OIcYitM/kZoILEZ60atXeiQDz5QLR
TBrSHMvJP+zVJageTD1YHpy6nXo62tG0rLZZ0pnTOjyO70mhiE0kCzLBN7d9M/x1
MECb/l7faZbfC4a4N5xSqczhFC5xXVL/sI1f103ExOE6NXVOaaVDpnKCmesQxIzD
KnLMxmkDtYuNsdJlyTbIOp7DPaMTWlC1hgoZJNRVtAFCwyPllJ/L4EKqrj3Nbo/s
HQUTNDPf1mrko1Y00nu7jiZHNpO9VYPrBOYye5YnRSVo4xsv0bSIH0R5+m1qsm0N
h3Q1e0jG7ksdIQH1kVWV3wS0k91pKR7Pd2m12GxoJzGED3hgJ4EH6quGIVscZXzy
XfLw+BQcn0+KzUXyucrwEXMAqqKXiwOSDNXO3kepYXJE8tRyOCgSrChl4rZTV8AF
7g5GciIg/fccpvHmIAFyk/EBETmdDoBxAeOUncFdckGLMvMpUChX9m4l9HIahHBU
S2rZJgBNRDhCdbT9dt8BfFu4NeFsHE8vvwQ46U72WF5SrJp1ryx/qdf7qp69L4rI
UeFI6eb1MgZ+vWTtSs0lUAjSDwMwslGcreqRbjFgiZCxlPZ5OnS0KjBmXXOkWEpF
MEE4Ra0X73r/IYfoMEOb5qspD3gZs/bxnTyvniiogZ8QMPb8a/H7xXq7kbSG6P+L
ayQp8oEclmuvfhToTPiswwd6yzMcQMfh2i9Bk/CfOAd4nF7kYWJlSFwHD0fJHe1h
rFYVWNkbD0pdpsQNTekEfVlWYiS04ANGgRzmuFpnzTiPidUdahZrJPJC7Bz05vjS
n0JX01I+P9w51xN7ylL8Kiot9Aoy/U6rwfhnZjuOP/A4Z8j2Cc1+K/DZK3adnHcW
y/ht6m2ctK+uwvMrgsx820Ws8cWxhMYGlDHN3qNAv3tAp+CWA/BPBe1ndeWhNke1
2v+y5MK6nvSZRDwipMB3jbwcgcFgDC1Tgvu+7z+3SBbio553/5Wt0ObiJPfpGMrB
RW3Tybk7DCFSf+mcqkpiHRBqO6LftZLMTyBdhOkIMTE7VdsqUZOQRHGzxROpSoSC
2FYzWxrpdauRzLmzGSCyjZi1abgILGCsmLjbVbaPCbKrUpBMOh9njajMHrOT9wZm
4UHbV1thYlEEsVswMqPR8+t8f78xuECmh2591KbYLwktBgR1NRaQb72V8Wt1ioea
fbAsEyXUKFAa31x0WaiqT5i6l19CUmh+YzLAvHj9I4JGP1wNwX84cVBgkbpsK12B
NzN7LtGVLOFyq/3eaivY+ADxuTGhcM/acnsezUiRFKRUyhx98ci2PCjRuF7UgHHF
5YyGEic/VnvVVxSOpnSx9pG0Q6A08kuK03mRcspnkUmc2e+sMgRzF4KOYxOhlM60
Pbg1gl4sQPwUM5lT32aTv9stdsdBsP55zNdwFRbP2oUNYI54AOWJSLEA3DCQmqnb
i07S8p14+VBYjMfRgiUTlF+G0jSsChCKaKm+zwWLuN5pDF40rkqIds4BusfmKF//
HG3Cx42Zu44VKu4QVBlgFel+N3j8WI342gOWbiib2urjjb270MyoRDk4QkZYB1gj
HZYwN0mlBaqy43t+yHIlT156lGTS2WC2DOlEkx+GG5pK8eu9iNxcNon5/2Xw+0C3
DOWmWIl5e2a5d9k/gXbkj4Zsj6sYF1J5FIVs1iki5DCEPItcHBaeDP5U7dXrWpiM
KzNpoGMH8TXwbURRGorKmwhIZwDwVn0CwrzypWNDkBCxPPr6fzTKNkwom+m13F3J
3VhdZwmTzuY5lXORgWySGI9O4Nljl4jtE6LS8dUmwirpssTS57IXP1N6/GezSV2F
rUGadEmU5SLYo64xOIbK6WuTKsNfcyl5IYsj9V4IinwnzVUlPqlrENljBBjSCL1m
S7PwmPYdrwmvGrXgs99u7gfSNjGPANMY0E54rt7nUabuVfGWg8r/NwHH1VGgHCDj
2wQdLinpZqE36DcnvlJP7sHIJSid52/VfD6CSYgC368EPjnzjPKXyezH0eIxCwLN
894J2zMLwyZlWvNh8AEtqJfBH1ak2TxjGawdPOFFVTnhF3wxy3q8yLn6B8pOQoh6
s9ugnrcX2oLtWD8l/kr48SYM1dlhRi6Gp2gTxSE2y0xjQnIyQa8M4Rvv0wP/9knE
yyxXHbA48sZj0Rj75uWgifdjuyeHEFv0zjK47czYtc+9951aLFWj3ZGDscynGq6X
F6x27p7RMz7OAhQJzrZS4XCLUd1ibfiRYR3koqnOO65rrvX2YzPbxwkfRwtGJzzI
9OaDW4omXGk4BEWP8T/ncNw8vNajPvhh9QxtaqqYz+7gaOHtzumfUI7bc4urSG1h
5qQeZiVhuGrPJZRxrDRLPSPa+cMQD50h3wpbenWdXCQSabTnH9ktyeph6Y7kmTQE
rHKbfVC1yRBVa0HMShgtKBxkd+LmnlRD4dg2AiYwGQbTHzqRyGBDfG2S3kQ1TXm5
gwoaV3YvWhMWTqoJ68NgobGGi/0gIAUfeBR15aR727i+MmMzMDk7oyehriStBM/g
R+E2prSinbnK4G+QNooML4vCdO2Qr8zntt5z8gGI2pcFhNc+9GPGYpIc+MSZ+7t/
gaRBYeqeIFZCNKk/5UkqpUdEJahrvIQVwBHHLikcStnqYXBTs2TEVQ8y9ghR5qjF
g3ZZVFq/6ZtwWJnvJS7CPcudqxFjC9nesdvmIA0DMaOXDjW6WLE37MfczGHnyVgG
uOAtP3khAYXAprkGlD8wm9fyJpHMl0vkD/QXD36P4FfT6hZF1BOtrGqZIoQJ97N6
YQfk7ngCgho6c1hWBtE4YY/Gidf8bPKRQj1FftGCUx/vr9DTPvEYRTPPQqVfM7nS
v2wrPV0DeqF82z582M+rMd5rlky1awaby8KU3rd3pwGRFJxCaIO/1jzqIagE6R7w
Yrj8GyRBeY75QKdivv+Ms8Nx8jKvp5gG5ZV3jyg7os0nM9CJJwAA7A8GvLt2xSAQ
Upb9OZ+aK0bWvmCX1c1MP/TUWowS9nige7iGerzxHKP2vKPdBzMBg8BanwcI17fI
ynO+ZUEC2x3Ajtjps4yOpI1MXCFs4pkdXA91PI3Z2AwGp7Is9kb4WfnChDTJZNn0
dRZwsWBZleWe4OqlcSoW4E87sMq+iTA1GRgFvlbMn9sT0EL9AUBr5u48Fs84/IjD
M67Gw2HkS5qmdYkHYkWSlwmIRtaMBFDY0oAYmm+gNh0GLllD/XHbIZ6TK9mO4E9z
KG29mHdHFrSIzuuwK2Wpw5aT4SwYxRU377BoDl/mgwhwEhTfhmra0bKTHVWR3IWc
aCkgPZHVQ700IQ8s/R+NdQieAF+WPIg3U5HKfLeZSghUWwYM9VJDiRCYFo9+z3rr
HiUwxXM0QkA+K5pz8LOOUe0ysYdeKm6C06nFTX/ft7GZWrIkXW4F8m1cyi7HUDID
Pq7gLAxnFAngPOTxySyKS6pRglG7b9XLNgETDe7eCkMFnScLTfY0VvvVvrXvgn+6
9t1t/XV7Teidz8NJ94DZ5ixpkGYlpetI2/rySwJZedODSD8UYwgactaZaauwF/0C
fDF/pFiv6ZsYri4c3AcaRFRT0uVncpJGlFrelHQQa2NWS5dcX0DMjGlR4VINq0Bd
BDQfihPHzdLWiA7PMHbNXeH+NJ5auFCoHnDYgpZtxAWrxUTm7OmFCCh2iNA8+J02
vGl49S9Ea4R4KUtVnWFw6InuTfsya7u0DZ7ehpb9SHO9lJHhFPbxV9VofrfQZT2Q
X7U5p64LlcyDCmc8EimSIByfnNgoTR5nycEKIQLiN2jdyvwQlfvofHhHmopFbV/K
i8U0QUn4BQsvCcgRYZ8yCwHYeKT+S+zJYZmW1HiG+qsXiG4CrLDQvlR6w4oGBPHY
bWa5lnbSB+/PXApsZtXfKl0J83z9QGZ4es0+gtYaKNrL3ZhvSyefpZCJqq5nNfDP
qyx1fAs427Nh6aNUnHjsUxQSZ5dLh3aVIPSilAW7qht2brhm3QRj1vUYSkJIVm+d
m9niKuhSkOIk50qfqtJiosOrwOJu2Kin7Ps1k6QClL6YKbGR7nYtqZDc+bLkFYW0
1N6XYWd+zRqEL4RRMHZ+M2sN73OusX2RG0SASjO8WLJz25cTjNua9ApxFCupGTyI
vcwIuFsfPqZbVXEhYMtb4oxXIV6s2alkI4vzheY2PWHq+thBo1yrFuwsyTfFI89M
hWFNqfXOrOMvqm4FUCNg7dbHBOPVXrT+OFTjU7w85BvdKfz5giz8NCAaLapm/Xyb
tD9tGZMV14iJhD7wm7Uvl+U13taKUdZHF/7M1nLdcmUm1s2IerIUXT1u7RMcmbBP
gnGXKI1zltwmvBTw3XHsjr+zH2HgWF8KQIL4iMSkW9tlLeIk2XXhy3S6zc4quMy6
pUyN4UgRiAX6hECA87t6C6Hl8aHToLUmrMBmw1Mz3HitB1/+VT4PUJLkF4pTY7CL
3GM4svNI/oi1pGuOfnbn2S/pQyP1Qh2T7bmvRSmptw3Z/WQuv/poqPIy1NKBfqjy
shm+fHx6XpobZ9ZeI9zaaRf6xJ5Ux4rFvsfZshufIqPHgpNqYpBHJb/rOi3eUiTx
l1XITlnOrwIA3rqB1ZuEGNpqCSlzlrbMPiQV89UDOeFOfxEbofWeOQtmXbEHxYij
DqVzNkNDZb2xGRRr4toaI4SZewdOlwGZ4VUDdg42JH5bm4kwJgPjvQpGXPkzz9DD
0zSJrmIZiRgk9WiFb+oTEWws9R38eDRo8jBuHa9sP/yNWjotdrOHtvrK7D6bXeAn
mQxIbo+qUaVaEwp2i1Q2cBO2SavG8go7dczQgHKLMqvSzszjiD1AeHSjm20GB7Io
SJaXjbPJk9diSjOu9QeE6YedPTjZ6/ZtLa4FQL9/5vsuALt0eU71qlYghRBHsXs0
JEvJaQsS6GRdUTdb1j3ly1DnldlfwkxTKHHMT77ImOqk3W71Kas03CTxXHaxqdRy
5H9XKerQr3PCITxoS80PKjGYiRbQaZLQFvrKJH1z2ZPhQ3a0ACIxZLNs19RzAnsd
Q78d7143i0guMq3dUpYLy3wfF9lsr8qi5riYfLv2zDKoS7yxklpoubY8exDtILCG
/JwRYVwFNMVU8fgpuSGpZJA6LSb5Cb9K5mpoJTufrKlXgZ8j2ctFIIykeGtaqcjJ
Fm3MWvMN1iAyIvVQR9lwHwbuXlZIIoOIu6OHj8ppzInbDhKWVNv4kSGph+svsjCn
Tdk0sAG+LOaYRiJU9if2EvbbLO0HwTtTqtCRoqlcBKpx8pyg4cM/R1hJ5URNQ29R
NcWyhkoKOoZoxyUda577wxo61Obpyg3EDJsIsk0PFuCmBYzG97r1VZcQB9veZoqF
vRbOx5a9rJp8UZACgp0l3eylyOCWuonM7EpYYOUf+Rcx49i3eTiVc4DHoxTpjBcx
EDJP8LEww7eclyliuawPmgUIdCxWGppWhVsj+vTHvwbP6qL7pwMwTblPpQBP+1Cg
rbHVrcAAtqFWZDQrCCmFE1RMzzcXuTytP1pdC2Gc3eisTOCNYdouUJQEStgn6B6E
DQksD6m1s4RDdxilDu7d5FEslbQ4oZfuhtUUgym2MC/430b3NK6htNFNcWI5k5X7
c0sGQB0H7zFS/YW9swhFrl7Oyf3dIRu2RA9VjFyoo5wfF7d012mXgorUJBiq1X3C
VLl/tTFIDwfVSKjT9MefhsOGyaPNEI/wyi72KvfJDWI8Qt5T9h/JJGTruVJQHxWU
KHtFXz9umERHfnx7zU7f4h/HY5rO7xLilZcCIWMpE2A8zEQft/7Xi7hmZZq14vV6
9iyJJJ60YWTK75rWIqyuX0Nz3Fl+ZtPs8Nbj4dRbK54UZYMwfJ0OPMM3vc3Jej9S
eZrdT1YDE8yf7GQ1qXCoEMypKTLUlrOQbQWcjXMv6zwEVwSOUsTmWmKYNNDdc7rj
eaqQD8LDezsYQ7ibRdWMR9BgQYTgar2cnhEsqXlA84mZ7oozJeN/VHlW2esL7HBZ
QnQfo28xhAuLpa/RN7IPFh1pw+yPitTlga4udxIidimZxrDwLE5aVbNOzyH4Qac2
rjr6+IWAkUXTusgxyiuuKlK9cYlYBPu24COe+OkukgY7w0DV6XVKM2a7GTltiTo/
6mpqPqhAI/MJsgQT+emcrKKWmKtfYOj8R8lAA/J0AX5jRdNQ7e7izpEu1tXMA0+I
YdiOXc6dWnZQRzmL+/MTfYKtZS8iClZ7Z1j7VUCOtyCXig8G6sNUtj4UKs/nY2V3
6QI1SmWgvEpwuzDuLjzL2kHlXpYfz4zK6lcRMGlddiJF4eN6rGl+CMFwiF8sAyjS
mYcKEMMhJFY6daPXUsJDGtNwLSoaseCiNyayI9LnivbXWaEFcPnSFT/5LQUPcrlY
nmzmRwXKMtfP9aIN9YhecGH6595q4kdHbFCl6BHsXHDI4frlRCkhJzofxO04ehnL
AGHlX6mYMkTxDqIJ1zaWNmiycHMB4VUZUT2amLyljHQN+Yy/eMIRvW4Y3b/aTial
TmSaQkP4X3/srOSFfQ92uxuWl+W6GvR/GENXsrkCkNw/fjK6sOX9ZqXsz1mZ+F/j
bRpPVsu4hcKOsuJD6s519foDtYYP0NUyRpGBkaXBZsou/xAE5qQUh6Yd1vWmjFkW
V3NWibkcyltuoZk0Tqjs5PxWZlJr87m1Gy+KGp09Ug1TMuxkvinOE5RVN0wvVTaa
pztWKzHw2rUgHyVM1YUVfM+qi5qwE+E8T2pHJHEz37t9omp6XqB1/2Rz2eA1Bw2M
exqM0jsr/1uRPDF6lKimTBCbxiEaHUtJbFdkXfyWnpU0sTlpspL/8CEL4Uta+gI6
c2ZJVKYTgjbpC48beB4YOohldsQiHmyYQ1f/xQ1BdmAzLFH+MH1vsAd8XezAE9z3
elTuHmESqW3B1ssmKRgJ+k2/67AgdZU+PkL4xaGrunAAgd/Bb4AqPDc+vksbt4hK
wL5d+XBK0/jqqiwHW5bh1uG6DkVbuo3X5cobjRSLsss9cUj0H3Gt88GfiUo5JJEU
uYSplE+7wB2FMUA/lFgR6zNJBat4ut8+dvYZ90MJjPniAIY0iofBwTXl7gwfoSL0
u63s9kBi4Xa9omvmXq3RxFrbfs9SB5KGTVwF0YXJ16Y2a1t+2ACrXKy2nSTExbkc
dCNCTSMVuI7tGg0IecF3KaIgtpF8mRyTLrOXCYMkB88+HhwqxhZR1sLQ1vNDtIcY
MFDqccUZGEVD4NEhRsp7orjzs8P2tO94uGmUdDO9K3gdZFUXMXFbnvwqL/VkXrm9
8Ak2VeLEa8lNFYe879CuJQDfEkZ9nE0kFtyzGdUFiIpq2EShYuNu3A4umVUw+QnH
hA5Qsg+Q4btkoS2+uYuT2MLT/a3szKJzfUiKRa6soU/ush/rcmMYcrCCEwUcSzhm
YbGvzcbEdRoyGIfdOJM2NXTow7bqElHBGcCFDngTAScAiSWjLg7BKBhQSOBwNEE8
pfYXD3f+tZX+l9W3Y6pPNDCazU7j/0Sx9bzWKpk1UdEcn2IZUmPca86qofdC2MWF
o1v4wcqsjRHKNMD1J5nYmoA+HeI2MhhR7FZA0o4mtzTRU8H0myfi57jyTYvM/POC
FBIwzq9QPDraYiSPPHH08JWjMlMVSPhUWWJ+f/XuXGryz4LbecnH0KvCpDQxm+yj
Jcuwy1H+g2Nv8B9d3DgSDxOL4XGhTVRrkYoCblbdWuS0BjoxE6pk+qCxhwpw/tFV
WH7r6DQMRHZi22BoICUB3cP3x7+lNd4KD7OYyrDCWe6lDAtTBJ0mlrxhVEjJH7ag
VyjCDS4RY5N8YfIBpzuojXqRNuKMtTZMpUlUXfJo6zU5oU+fqB8Kj/WIW7PzYK0n
jbnG5pWdyULivajkik08HNLD9xRZQzSlJyBuEK5cJ2tQDP1eKvnoPY76nb2qF9N7
FjOGDpSYGJBV3gcLbtSCqNqGGo9uajXE9XUFITO3N3nZbiQQ/H2Xtek+BBJ52/FF
IdogNtCESwCi15QTpAANTxBKCqspnnG3JfMDU3XbgNC50vQmf0nK9Bw/Uspru2nT
XNKMMzfs2m9DqMi9ZmLr4666++L0S68Z432f6OXfcMLC7ZnwYjFhGVLMqtzBxyXW
KdqZDUNGYCRZ37G+uo/yxmpi/MM0unMKgLo2CGEa1tpE0lsqKxo/7LlrMUYtipxo
Dc8F5Hi39lrE9tzDuTyGecs808tDIajddeCS9tY5mR2bKf5uL0M34xKmbHolN/Ni
CVhxtZ1qD5V3fjIxMRxJCayYQEVF3QvYKwUKpq7tfD+DzjCYs8Vk7KqEfWI532pq
MZ1iy4hap9kHFajGhXakqpdVD/sIEm7csgUsOn8IqMefI88qkVueovSpODtl+UPh
xovQywETU/QYpxl80Bd4Nun0R17y/HaTmAJhV5PAveLVFJhb3fHJ2bfrKo5S6ECC
Fo+HUhr2PYvsRevMYMMpkmAavs+EWDOabwVCZDHLBuRKGDD8JL9GEOfuFsk+n5PD
ciyHE8hNN2d2JfvinJpd9tbEW31PDpy6Or6PSztNcsbdRyQxWLKEY+qGtqYc7ZJm
uITtllW/uOmIm40dCLUcR4W9KzHrxDOEmgVNdPNO5pPDf4OrnLgztQ6PyhgBbdQC
OJU0DdB+Yzde+FcJv7WTKHlqnfUbJHT6iarADEBm/w1PFQXn4QmJREW/6rELzutC
fN4V3lMvHKlUxE30omAzovpTd0cMaMGHz7XDtWCNx/f8/leMZ22+pvbgQKX9ox+/
IbetgKGjhZKUvyhHnA4i4uhLhfqINjpPV85FQEOVKvgDGK443YCzrH2Ew78kldPq
K6MF6mDVvwBs7QRPybkLM3WvSTrBjwGavjK60yhGHDuF2Hk+9lT033DNQM7OKonx
Y/g5bhJYjZaA/Cylma5oGfGklB7ikBwVk+QwuirLVJ0AaHB/DCzrvlOaHkeVva1a
t1TBdR01RSj7Dsvk29WTBP53n9e/5n69tIM5+vvmKQ5BIGXK5jjU8/j0hOj4yeze
yEXSarBLVXxnBi0SKlXI2Z9TdVU5fyd62o2oNbzoXnudhjiYT9zUY5ZeX/Mcy1c/
p8lOodyxuK1pseQNTn60nmR4DRplHP6YIXwnRzBRy/SiZWfmik2JIC2N+AI4k04e
DSzGhl6OOECjH433V72MGlZXJAuNHP0lq9Hjq+ofiltOuLMg0w9kY71im4GI7+59
dI6NO8im6CsYR/Ebh0bnUIx0uTzGBnvNYQGJUaiwWDvp0gkld4qu+wwiTabBFBcT
Iu9uOvgF17ga3Kyy+RKYzUyEbn79vb1xyQxljyqJ+rrZjuZNB4Pzl3OUdgm1f37X
l/KCBIpjktFBz0p0CC78LfMdK6P7N14qgS4cc9yQ/z1B8PK1qaAG2vJhmkbrCHTF
ocli37It0ksKJRxtN+LR5Oq6vMus/7Ru+waIhKzs097YkCxv/y28vAgePkS4cD3J
1AuxEAxrCxGiPY+XFls5jhjmW53AKLpegZ7vFw18ybqAdP6XqLrKyFPG4gbudsQR
hLx7nyMnZ5XjM5awFyWWSh54sRj8WFtPrwKGDYxdR83A6OOgKfqoD1tXAxJtEcOo
VN2j6jQ4pt0duF+hi+ww/qe1SwzctrnRJbkRatfJhFdJAebkzZrkMCevQvDiZjGx
OsI7luUzqnmPp60CZPjBRqu3hGo+CxjCoJ+tF8CjdMkyBDwJIXGeCbBN3uyTAagN
amcrT5PRSpk/IZ1HkOdZiNIOlDiVoCSpc7TdbT04FMVJ8Co4OKbZULcz7U+nMCLj
3gS9Ngt2ZqNNpVkuVCIANaTW8qxAItbpsTXWEKGJ4pVBqbZlfQXXLOAvW2W/8xoK
Kj/Zw2EW0XbyiyvprIm9MyzPSBaHUXi07kvqsZvn/iXh2BiZKDMNCP0sNBDCBHgy
A6+xFiSq9kFvCi74r2UWHb8TWrRg6ZMcgBdMEwTzICd2eEJT+FgRn2JJp6HDyp7G
LNnNfU/3SXBLnjIgibDVB1FR5SNSYCeag/tJrz+cxZUTws3sAqk34LC/zbDw+PlB
zHel3sn4QgSaHjpr6/6S5fcg5EOsOfU0bVl+U7lnH7LLwkVH6vkk9DlKJz7eXkB3
qVOwK64k4LzW0D6E7xq62wYuGskC27CJEqENrEmR7S0g+6XHWuUd5CMUO83DTJ4/
yc2ZfJi4WUyoD8fqzFd/wwh/tvI7mcE8TQwOOPLgbD1JO+kVOmvK5pxfCylXqUnn
7J3apAXe7dFzBdX6GmSZaydTEYRoSDtN0ZjtXvxiOx9XCTxQfZY5MmVVJjvf1s0Y
1HBFJ6M0yPxl8s1i106xBApu363x3HqB+ZhotcIrfd+6sgQ7U8qhZEfFMxtFGpEv
3NDH39hDPvODwSVH5trdVgOC4hLuWJuZITiyj9qgQfL5I9lKBn7CBW6efTEC/uZn
Bzrj7tzY1qxJfF5htfas0gZbnGxRzqFqzmb9pqdHGuMywzSv9gL0+uJJCUZTHQiC
rXcWZzY49r0+qIfNGecXmBntxnun2gj+OvFP2OBFmzypdyeEE+KwEJBtJmqGHzc+
d2pJk/qu2zBFF2EU85ox7PUmorb1m0nKQpVZIvAlzolg+7u/8KqXD4a1WSsibnND
SspvXk26NPc7pa6GHSoWG/L2IcuEVtVfAIge7NcLzJdPNo+FgXGK4RafQbmzmsvA
buSr8V3UNB8cxflu/ZH2nnQXKBKXyAU1Al+XeNtOpL38MCuPlhm0HLy87US+WEek
yaah0rZTefWIgZS7LS0JYvRjWqHfxS8tZBFNf7EjZHGRw3DZ7r4i3YqixiU6w3oJ
5F9Mxf9OlEgEq1HzmOBMAAYEvBVwelCwmiDXYhgh85eu6jHv3Nj8FVUt64WoA3xk
VO0Uw5vSNN1FYRpAEO2ofbqfCCopDExgWuY9XyTG7mjC+hwTI5H9Qus6H+qW7Tpo
t6UU7kN9SO6XfX6KYqOacJp+xqjMrfJZi/8aYTUehpX0PGAYXXHjvOJjuQCIvYtK
re55dI+2bd5cfz7XaePucb5NsWNSjGbC+q6itkku0o85uZUVAI+BS3h4kS4HgJvh
R0Xxdr1X9GUe3GlIW+Q0hbu1LzIfUVP0Xad4kDnH2KnXctKjLBCKvic/+HJwJoS0
F8nTzvtVkQPNqSGxGweYP+ZUhRlX7+QezyjjyJqZBVvTf179n0QilY4bikz+xjpY
wWvKdZPkuE0V5fkrIqsEpiCMMEMAFNRqCcYfV1BcXzPXiXi+x0gOncUaxZjYbRVs
BK/IFn9aaQSwdwZ7UcS1KNqfyATFX0wjCiZkQT7lWJ0csSalLhJr2gKhbn1kSetz
VaRo1ihRslG6saHrQSWNOA/4WDxNsuHovfrMn/2abLDxccoebtFIDAUU+M3ipSB5
1C+PjAVy3shRCmIDw+2IXOt9ZOQU0pkvYvhnxtPs8p5rc7s0839Swgt5dAZqX1ir
jORqSrS/jxCFX7zCGxbqoXuzJWfNcNZ6oGog5cwuD25Gnj906pP8qNF8JsnFAt74
pVzyejZFaWNG/w1CG3E04utazAx1F4wihwv8vMtRhd9QsOn4hKTP9eO1PlqMmXAP
8pnSBDOHn/u9mUg9SaN6AfRrMdW5k4GNNbYFLjJ5AaKiOqD5eVcqg6AAGztzfnwl
7O2sH0CgdT2NtIZzNvsLvjV5PjD0djYDHyW2J/nyAEDH4Feiu0y6i0EevI6pCR2w
aLeHijc3v/L5zu4+2D/7FANL8TKpYCvgfmu+jqJ9CjSi+6mkBeA4QdB/MWLyXRsU
YUQIYg4TRoDRBqcXoeH1tMPLb4WSFfiCu4w9Px51tq20SOQ+qTy77voYqLtxiqWa
D5lXj9+2VUFmFphDsRPIWp6j+1I6dRiNajNWEHzRarMp36oWe861rNTkKRXTGLMI
6HhPyk/Z0YG+tPddTWLFBWJ7ODtbyYLKaGqidlcU/CPyOMB9+GGu0VMED8qJZQog
lXSVjHF6mcY+cj83/Nt+trK/iMc16gI84nGc60S1ZEAbcV/aFiQKkxPlm44kXol8
xEBBI5jKezCa9KGAB3bnWHZcwptZglKCzlqkSNzz0lvLWnOz7yYvtztNO4o2oEBl
ZogQVE8UGoB5SYVH0+4Po9U86Z7WBww5T2MN41od4c45a0vBfIhp0frVkYVbUMPj
fnSVfeyhXcl0rbuXxqCxZlaUs7EgdZytjJD3Bi/8H+W3xoiizoX40peAmXzLbYsr
5dhNBQ+dkG/Kcr1qEMK1eTpOwbwP8eTn/nkJf61+Z53X8VT10QY+qf2K1Bg7wT/k
VH5HkbjHV7CKJ6c2QizcZ8zbFJw8JsHxU/0FYaIvS6TF8vsTOYq96AmPxu2OL3xE
QyWoBce6upi0WnHuNuwTY/59FP4Gz6JVBiGDDSeMdaj49SlxsnLc8UjeiJMPsolt
TVUueL+y5CM+vhPnBEe059H/+zrUp/o/CjjMi8BxN7MRBwgJghlCH04GDwGjKR+Z
e1z2oCG9uhXpqXtF5HPrWHVEoHAXtv5NV6OMSBN0dekirOJdNjDKG36ITWJBW4RK
wuCj5kxvZ2ZGcQOfEkTqwyEisWa6x+1t15pDU44TgUWh8LnUymkDQ9o4+nK2H5XP
8TAKrl4kVrsHp8+6xo5vjwIS/Ma2vqQeAvb3ivq1mpVih9iSilmAivvtNyikNuL3
uK/bi2NyzMiOOdvlGcnSfgxCaJQal8o3L2YqahXto5IYMLsrZcAATXCeuzBifuWG
uYhra6/eyi0s4NYxVp898uEjBwWvcfegnWZg39BgtU1fLecuRk9hSlasNiWZF9qa
nwZfwX8h88Nl9bt7i68VddnnHMb5L+Q5nm0rlWtn8t9fYTQYexYDiXKCts8HJzgF
pcdwsvmUebFQYBHZb4rvlQW0uxf/sxiv+Wa1CYFhHiSk/nuzw2tihvJc0Xkk5rMS
g0no5eFmvli8ffmrgrf322H7n8lNvkkmuN6tWlinPp4RKQSgpXsNJX2eVjblUZUb
J5o9ki3bUexAUiP4tFq3GO2mi1LbB0AAhKTGRHUkdyAcfR4mpEw9bwyQJ4AqqlWz
WGFd+uPqmSx2z4DraWd+iNYOCfRkbF1Du2osrgiCrnrAP/k2VwDbdjKHAjj/Juhi
pvyQaiU+YPVnPxOxGh1lApMo9Ct8LyHR82XY44scBsocbLv9DIvtvtG2rYnnuVb9
iZpdoZiemZQUMnq3OtDbYoqI/XzW49GHyCqXiRz9IKLknl0R5Z+qmhEux5x/9+TE
dD4fG7Dt3uAWpbIjT8moB3cNduqz0s9N4gPHp0e3hvI4YxUISSAQE0eo9HaHt/rX
7qGWxjgDjFkvdTeT+xPy0zo+Ew+wVAAKM6yC3J4QXtXoLehQSn2nFwHhzqUXEf9M
8DlwNQOJ1Fxq0/01ggh3L2h0OiI0WooqB8msX7fZZ9rh4WzsD+f/1jxWdJyNOnYn
UwVvRL3LoBad6b+ZU0NhGzsqHyngTb0y49QibUxjBxSfMA/WWIHEK8SglzkYNAH0
lpkey84nmW282TKPf8t3DmYphWZZLoLbklcXpbCAxztPGt3XEDkA7zJHw+I/7jdf
N6V1f3f59byStWaKUwYE96Ozdr5FWP0c5Id7amlsA0WsM5MtvxTU57hJOqiH7Uww
QTxSm+2XbTVfvTkw5cPzPVW1E/advgq6munkachTZ3Bmdg5IFpM+p4JkOI0nSz9l
NY74lY/fRlRsgCWynhNlJ9Q/TGPzX+7qz5sjuJBq+eYT/SD7ReIs1P2F0/ZAU+1x
Lvp8GY5GfXG4enXps5gcc7capzd7Dlf4kPfL15UT/hZ4Ix+pf28XoJJJu2bF1BAK
hzMUvIoVNvJBzdsnut8fbuzX5QqfCPmNxBRJ3O1LeEGgR8V2BTPLyVnudIYMhZrV
g9ur9ljzp/aDibGddV7jjkV+GN4w9Sxu+HlyKQSvOUvv1q70F/btU0BHSgHJSCXB
sk7tp4X5HWVO9QfGP0LMivXgBzxXnA4NombWmEFrwM1z5yY1Z4NvA6yXJFuUmE5L
qY68vpKvzLCqPUcWV9TadU4e0/5xWBEv9twWDMcxTRQ4ehdZVf9YVRfYGAT2eazQ
8nhICbPwhj0RGCIyD7VgVH6n9mCvr9UWK0elKrXLn9Bq18lpeC/xr1pyXhCPF1LR
WuDF/+gpmD0BiGwUmgDexPbwG+Bl33zc7IZJ+zQSNiiWe+I6ZlcvFwWudKX2fTum
ZEDbz9Rw6whD92FW8SxBWxoVrbkDd88LHXkw6Pks7phV1OzlHufRqXFghhJ1CJ2M
hGK1YquLmDFLKJN4FRJZWbE3fofUtKiuCuZGxNh8EEobsgfcrjsqQTeidapeeYGX
sacAj2Z2/w8ZIfV+Fg0h+zaObpIPifL9EanUQPhsrBcDSepPcMgO9ltgzsf9eQBM
IklNg75ZeuGVwenvr3mReWbVR56vfOmM6ojgl7CSUrZhCq0apxBKoaaUx7EPuwRb
hHSEh+HPFhd1mNNec0nUbdlaFLD8fDQx5p6/4Bfx5vIZbNHiow76hgS3yd7V6Frx
Uzzo+qexEanTsBXfTOsrCpuH1UTceCAjStf8FJ8LcButxkrWQPYlxRhoREaD1Usi
yR2lde8UupW/HPAmq4zZ0+9tVkMDv1SUDhYGUHLlKCnNSb1Qcq6oDAcVTgqkOHf2
yYLVdqdvS7w/xQ7xC6PFtCSOjDZI39yO4KY3OzYHXZhj6BTty+5qPcUFvsWavmhn
2J/Lh1ngFwfur96DNyjyh49GF86nvC8BRVEYwDgD9E/vN3SqBG1Lte7UxKn6teJI
IDLnBKWqK2rFxpSdnbKsmrNHi1K2wTjPdKZjeESyc40+oj/P1b/panwIfEzQIKd5
1F77HxZzP1rMmBmEx+PnVnPRuQlkoVSJiHdEYjsHTJnrq58y9yjKrS0XhB6ND/GH
ho8WOK2uFFkIL7KlXifZeJmJIOQ3JK/xLIfGu6qx9oxG7klcITX4230KAUbeWtVk
F+NQ7W7UmM+Ii2ZZ2k3MdYSCBouaJ+eWyyxtSQ2iFayfpOUzGnQzZgJ2jnNPEy5S
j8RZcWJFMqfS+QaHVKRqxEItJlPAJoCyVNkp5J2+3bCaMEeJ5JmGx9lcxe3da+0X
pdDbdNehbomosOBSVe6FIQHzYB6Mgf/QHCOCotY839HvzSqEalYOs1ih+O1yQGhU
EaW715LYl/EHnpgZrWyCWQER557nH4sHKYyjHSIl623oXkagc7pTMSCPrbYApwS8
vcWgnv8Le+zabzgjs93OjMvk5evjM2TABKJNW2gxaBJDf7r/Nci7l+qjEIrzIyC8
5f4kBZ/T4AT5Frt4maHg0dZMRwMgMvRPOTeOSsl8yYbYi0mA5BTU6wv1AIJANTIr
VAnRoVIf20fqdVENtNg9IDCLnjSfTpW2uiTMul7S84ZELaKQzjPrdOIUIWiWB789
rxbsKO9X3fwCC3AbvPjXuz7cqImZ5bezPo2gTrJ+B9DUMB0a7LhHizbmDgIuDj1k
slmb27Nl7PMv7kTiIqW7O26/5IQ7njVsAw9pkqjefC7iBR6Ps4zuwMORFafOxMfO
heha4w2/J6vkXK81xaHPEabGaB3Cb5oGK50d1ZjGh3+s3fipRFmxQuQWTtJgWS6Y
kCnhmYS0zrVp0mT9Ax9Xj4pnnvXXWb9C8v39osOfO+WmRqcriMH+njYNaJelao39
bQF/a6Y2ymZBREoyMFS0Qe9hP1R1eaeT2dJmSj1dQJqhT9bB6680FeE6r51CDGV4
DSjpkpvqNYJ2hmqhU9lZuRtOqHitY9fWh652h1GSioAPrEHUCmMaakaL6eCcyYOK
VXf85fQ2ZvRljAxcuUoUt430QFQ91Svx0MbJh4QYQoSkaQzuI85AzFDtga6aURlt
UAm9FZqzypkUyWj0r5dTZDlRNhFuCRQNncUMDX3QKhTAyxVICrQVpO3JiBIi0joB
kRBgxls+eCXBclEq8p+/eyU4hc/CpMSPLb7PAW0RZotSA9h6PCx+wVxP9L09IJYx
IBWk5x/GHavpuEsmgUVr1BDiPi/cFKvGk6hYH7R5BIXxQEbiDBYb/Cv3i4/mBj5R
J3x8maJXngpJ0+qpJv/kUfyfs0f7w88N7PZ/fetEIVjdfsabQSDgOK/eGnSOs9KJ
ypz5b2iY1QD0wENSau33vzxwt1TjmQTZ5+zpsACGqYk9s3TcIZbZZ4BAgrm9CKvC
+bkeJ1JomZ/J9CnW0oigfnJW7EN1bvhaGkTCsAM1nel8SnowFHoJ3gA8rLGQPKpX
3SiPGNqdCDgP3d5IZDcbIz1pUZqqZpXFye5ddY2LyIDHougawW2tTbw6nJhOpqRA
EG3M8iecB8woVck5THPCHTZJ+LaiwsFmmimezXAWyfg2cz0wI41+XDxBSrJkVaiQ
x2HvN+ZCWBX0UkNJ7RjeBCs/LEGqVkbHbFpqlkNevSyRe+ceJ/MM8G5aVwX8eTAc
Grej8KAy2nhv9AljIkxmywgEUtdRBQroeoZyR/H0elVn7GNvduInadFS895PXcax
CG14weHsnc/7/x5AqC+iB0b7J/L26uFzSxTybPpKsXQly4EBOjBAi2Yvx4p82A31
krZh3hibkJOUFPJb1UR79eMCORxgWqZv0ObvdDP7znDmz6mRFd1/VExuxXP3cmCq
kL3faQ9mbH6SGNr9mT8bJYLo37ESiAyOz+mJDGFJKrBGYBisAKaWkTc7mFW4sBp6
9fBJOD8JsdIGtMqZyZqat8HH2vg4BPGA39L2lQLWT1TWBabJBm7p7Hr/VKnhuRQi
eM/6jzJ6m6lIurjNIX4d9GoSxOdjZ+L9Ks8/Et/v86fAdmozXvqwqyl+Lz/dZ4s6
sAuswGVbkdOwN8mqtaxEbMynvjLXEleU++d5yxXJ47zjJJgpEULMc0qxgnVf0W5x
7dwichCRomgK5bbyKazK8ftjBqikSoXcH7ymOfnZbqrLAoRsFMYUGjmjC7510Kg0
pljhP12GvdQ70Xdfs0xc0hqB7ZgAZ1Hixxt3Ym2Ol1yURjTDhQgTOt+GeQY3YKj+
lXU+I+9mmBIHh4VYk6KQIbTURz4dLzq0FslIQ4qVV1cv/kxFBIkR4Lxj/4e3DkT9
jW0sH7h3MAGqzmNrAE+x9tI0gGB5mzTewd8HAIQB5kRehp9bFxJSt+Igrns4bxW5
ibNgEg0vtJ1NnlRpsqbLaMWan11DBLcjwDhben0QHaHiaU7qOUab4SRwxRAQFUHt
zL+8pdnl8ppT2tLBTp2cNgp3k9j08QUlobpwEj3x18ZaIYn6nTU8eA6bLc7beF9g
8HH/YvjK6yhXT3FRBmi6HzJ46hVHHnFutya2/8LeGXjGBANQudLI+iF4t53YPX3/
G54I7XDHOnCTKL+Z4KXf8CrhONQhW5yxyfMhf5D4vQie34zdTzd2umfB118LGDKw
oBOIhohiLo2zyz7A63A/vEqitN8iKSNxVdR1/UARFyRxqvC84kKPCqjJwhj5pxT0
v9tRrrMNf1U1TfewS2srG5F2d/eYOhYXehouWOqPNk8sAAn4J57fwlV3Yx/uY2cq
iCzbNFzYo0AOLQK4+yvoVLIQhozINv3lFirJcy9YNdH0Zt8J/fn9cCqIKXjK16v9
S6DIN/4epRvCPf9CBLvTTCS9/opRtYlaXX5z5VyyOr/ZttEwY37/bqib7+6hZTeA
oQ6NcDudzFDUVbAXc/0Tp6AIHAlTsUEQK3AiH0i+gnJML6pbRqEdwhd8abqw2tD8
FYras3cEaLT3/gbpo3yCIlrBQqA5iPeEXywpxDNPWCFB86h8uWFoN1o7lyf7+f5h
VdcmkT6LpfuhZm2tZ9oEUqd0a4EgljmYj5B3AgIL5fJDhf32VOLj9YRIUH3Cq0X3
wG5TysUflIHd3toLPZm2lQDQ8Fa7/R/4s09IpXNsPnAHqW2/2mnRAuH6aR+O7Ad2
30QoEhuxf/TsymFoScKFzFYfBdP8zIvlVk4uDGIGDaCD2j2QyulFE3j7vRgLHkAp
FxZR8GWB1+3BcFS5kUyOPra2BT42tGqOhNaxe2aUfZwMSqSBXXsAdcGD5s9lzWfv
2gcvWdeVJpGSBqbys+KvU3dyW7MlcTZN4dSOmEG3PBsb4GTDo7r4i33QaFGzXUxx
OxcsJVVxR2fZ4D+JDUj2WSMx1Di+5krLxXA41GnR/WM1AMjcvSbbYx7kXH8jMFSW
YHpHFlOLxG66m7ygMRhlYnM0UdmS+dVU+9cMJoUqfXYWf8nVU0Zsj5YuWk0xshII
s4B//BuPnOCeqA2EKikw6nGtA4CG/5dBBcP9tRGvtlGxatOA1hiU2g//0zXFVuA6
L6Rk55/KYOUHoqRPNijVXPDEMwkzUg4dvBLdoY0Tnk9wiKMmZ3KRQh/nk48tIrX4
8SBxV4pzQ//3TxAewqEAw/uT57Q4dvD+T8OiDL2zA8JbIfKO6pUZpoqiDSOqNdH+
PKzCjQS2kiNVlNzbefuwG9+ebjYQHwur/c4Bg7jF5RcPY1tQjIUVPNdASpJVavvm
GUGRTECr2sEXFyL3L285oZLbiYMTYHleqZuPo3dYqOpx+xrk1aoXtGAabBtY+Iui
PFi58MeFKn2Aa7Do5QCAcdfbrMonuaRF7SsmeTFHJ1IaE9sD0tSdc3d0tt9IGI/3
p67YrSUyTYgJdivSSf8xkYa5vcG/ISYOKmTGH1Xpq5Gmd8vSyv/r298OGpOIdpkJ
8xaFHID4JamK7aCBCeQR5wYH1WCyFg2CkpfvErr5FUOJ3L2DAQRCy3Ac7bA0OHhQ
xCaCnJWur8qJoykrGdcitJX+ipF/Pc5qni89hLJUjBEjSMOz5ABtnz4m7H18mO3H
ToPW0bgtLxSYkejC6n2BFXB6B31PkD6tiBGd0Um89aXEf6nCfCUiWf0IU+h2mEFJ
Ot1RzOGc32h6vfJdc89y074eEo8m0q/3bBhY8mZppYOxQJbBBH1GkLJiDuWRK+LB
ytIt5zSdYMTsgVtyD2AiV4gE27hBHB4ZBX6/HNoT/QvzSNuo+3o3eVlMEkMxgTT3
gcC/AjGFU8qWV2e6C25yh1sK2Q26RSOewhBf9GgP4+CPmax7onj38SYZoihYrjin
ojd1GRo288OEE0zCbjfVC1BQIAsLNA2sshOYEGC/XB0QJm633bMegwlAsu9vaQJh
0b95DdO4ItdMGZ3Y1agjjmB+ilrGmBdQY3HvNdaFjPVpjLJhiMZk6h99nYpljNsX
B6uXx9NXaeO0FlbTJflJZvHkDduOZAn4PXTEKnxB+HgxTqKLhmlX2NCgP+rq3eJd
MxVx+otw+zh7BJb8QYk6CJ2efO554jAqoOWo6fA3xcKYCBUPFVuY+aYdPh4G0XPf
bxUAddOZuCfwI/OBdToOIE0YXazuNaHuhI6YqrJO+M/3SwuOKZIjdm7UdyW7WB1+
lA1N2l+zL7BaSMkQn29SYhem0SVgPujoA3xcABFg4frikruPsmg6quL0u9cvfYOQ
5whvCrPSkRVieLxlyTIqmK0Vcfsjx7/BoxVMQBz7CssYuUXeeZZCCUKO4zO42aeG
NriNbtsrLp6Ox//nOxsKohfklCb+h7r8+WYm1JvRPV8zw/DwTfmIlPq5d2UV10ER
mo+bri+KjP3jqYwksLBfZirpYZoAXk4kulHGzFK0n3eI9z896TobdmNvEdjtx+hX
qwmQzbnFtWC5zdi9aTwUIT/yAr0rJu4zygakqUFBJvUScJPUc/M8fQv9ybCUepO3
1z7+h+P4B+dfoys6EgAWLYYhlWhAgyXu5RXYiE9iUSg8hvdpIA2BdpxvjoAIL94z
vD5FhZoex2d/hgp2lJ4/8HDh3CSW/6Lpg9K4XqOxk7PVfyw7HRvwCDlXBfHUj+3L
z/q6o9ACTUvudi0Skx0NahlF7/F02D2wSSszGAxfPeANgzhS7E+03NF0/RHqNGwp
ui+dNfmS5OLZI+oGm8NNvxlySGSARlMGBuTXNW5WXesH7iMxb9DQDWJ2cqXR2SQo
+ElMa6ohf49Eawbo80NFC1/WwoCA0Vm/Sph3YLBxajCfwbYIkkU9Nd++qQmRnfMV
VibDm4eCrNzVKh1QT1czo3bv6r4rdjZyDNu/dRlZ+bSuexrUbwG0Em4mYWKrxAnB
FeQnlrKBNUzyoy6fPRiJT3mow+yrZDKhCsuFKvnMsHWtCYGkViqomte9cG2Lthhq
bJOH0BuV1oIS7mz3LJY+DT/naB4De+heofpomDfwrjP43MeBJtDJJBYD9sGiRNYi
SIxSXtwD7F6S/p2Vb25o9qalR2Y4gEYNIvg1EHdccCZcbS6YVEdMibQUV6Iuo4Er
yTpF2PAdF5W9OugXA3W7Mv/TvVb+5XCYpdV7tu+wYZru4Hn8Reg4WwXhUh7xt8jA
Hv8qJssIx6hARXEWNsFOC6EgXgvVC4HSYz9+HQMvTodbNR5uCrklIY1Fxpt+nGYq
GU7yLM0+kn2zGaPu3j8sK17rwUfYO6txht0aUzFahzhvC8glwF0ROIG2Uw2a5kdE
a0iJ47I6WJJpIpmH1Odl3JDmJrWv7SnS1PPvwABeI0TeLjaFyJuVproQ4AwgHc10
9hga43QyN4cfGr4jPWijKEA8BzpTaUVnAm6EOydD13NB3RXM91azI4ugRTNI9kVE
0OdT0BvW/Ckko97zSxtJ0jzDjzbZ4xHdEGxTUzUg8EMuOOj32yQESlq61IiFT+2U
pM6eXa71CrwedT4Bew8/ulZ1lFmQX3rrNK0emZLBMaGsNKQKxc4BPq6gRezL8/pC
iMX1t+HWDAAhM4E5YWKwrGr7VHfZ8RQgZVMWlt+vYI20/42pOfzlBm1ln8FCFdlM
fw2M/tHUTb0Crz4H8J/0kkhjLeY07rSNVmdyBV26ohmZp1piLYWl3IOa4QBcAo3C
40OTA778VolHr52e4TyLGwTHCjmL3xJ06LvfC8QiU8GtkH2iG48uzp5JpsAqlcwV
NnzZcJqnAlG7SACjc5JXanMMCvDKnR/NlP5ZnB4dAWtaQJYenCh7bLpca9zdoCfH
lLHdKrs+BYRwhHX0BHijmYwdIrlyEWcv2OGJtVUMjLRFLiQDx7d6esJrV+PjMuT6
k3s5h3SR9wbo9es7fzcBnGKAVS8bRwdJOlEyZsdjaevVR5Q4upJ+zCzXNxUbmR3U
SJiLNDmsIC0ygS8Q2uCE92YvSa5pAY0F0DWIQSXFO7iIKnUQ+9Q7ocjidOInYnjr
qwJ1tBElCMNCunjUvIF7MSMWGsJEsse5Bn8OvxG1JmojHNyG8BAgL6IQAQGvgdDg
vMKC+izngQU9BsUUenSn8xSk1hxHOmGdJOMN7w3W29t22crTsYYg7JpapSRzmIrn
PwIyj49o21xWXvqsD2HoO05BEZPLr4tW4tm2OmitS2T6Njw67PZ95viR/aEfy9nE
+x4+ClY6a8jdc6/pftAcN4gvRq8bQs4nOtsuw5LjjtaPvw97g+RIQOiSyzmQlSlC
mbW/j8NNgbz5po0Y3n+GdRRmSpgY+iJuQMkMd015/P413bRHYbHVh/TDLc3BI+V8
h9XIp+iCZg83ES/A+vgk5SyGt8a/vyhA63NDP9gwfJ7aoAMojUcmpI4kpmjzLg96
V1eoIhmbR5WTv6fF2HnuLlFKRXvPHnY1MOKQiIBAr+ptzyAjTZbyZBQ07v5Fb0Pw
YNENic6Y8G2101uRsWxjPJppanalE7sfaMOPMJToIhp/TRb44gaMcOrTKH4XtFwz
wyJhb1riTTO9Yqre1H8D8qpm/Yi5VBV4bUi4DE7t2ncxLSCFNKVG8bn4VqggEARN
8nU9rv1etQ6R3so/Fz7TNtoDSyUB/Z3/tIbVPXJ1AcuAdWcZaY6i9t+VEg0nVkvU
qzrHHYB5BH5wo5z4exFsysqnN+OWu84KdMDmdt7BLXTW8DDVnnbUpMe/0Y6G+LWn
cnsN8EyPUkqUgggAeXldE2QgdfQx6mQFmCLthBoH0eNQv7/UxXBKONW3/fMJu6mL
K5TC/OBQTfuAPRPZDE3Eq7WnhgJ5ums47HtLJGLjiKWN0Kstw1uyQk/6cZ0EGAxm
JCUDK/YpVjxMun5IZ+WexvRX4BSXTsKiPtPUnmoKHA2Pjy+2CdJ9nuPIBgRz7mFY
QoDjgrDrVkNDoJXcoe3dyCeIGYmvYcdaDIPRaesA+3bF8iRz7aeXxAkHGd/vhFbI
4tFHuj3RbJ5A0/0TrJhEXwXRW+mWtCohVf6gWOxGEPz6cPFvOsfIeAWndJI0CK65
ulJc4Nk0RiwjkYQLX2nTc6jNsp5xkJN6qn7HcSCbvHAzuutvMQqgda0k/9EPT2/H
KxqHV1wfE5ZEFxsUsbZSR3hJUUIFTwELqgfmp7SB82Hnh3Sh5iLEuWLLrao98gTi
MH0AohmclcAJYvaYVU0UREVXqblSiib/Xf5ujEtdyk8umZ8Ci6buI8q4qoFMFnBu
YgRC8MqeU+24sqnxJMeT6hGI7bB+2K9vP+ozm0MdxWcc0emS/QX+w52rJerdZvdh
k6xk3iDlZQPTfzhy2aVjGNJM02hHT3tGRKVkBZQ0ZeGEsQnlNbLBC/1HM3QsQlyR
Ou0HSk+6Dq6wYbN1sD5yc6G91xEwfGTtHEyA+5HcAI/11lXaZjw54+XsuKfpVteL
klqUuq+ACvFlKu9mlJH7aVMTt82ZaDcsx0FJ+7YWCG5UQ7E+1yt9jbKJSx1fe2bb
G1GfhudWSn11XyaguuvX6GUv2+hzC8F133izEbj8RAz8H0kLK4ddu7FRTwPQIhot
X4fl2aZiy9ci8pcQQXIfXVILCWcZ8ay++fmRh5u8ef2gf9t8oTDOcvGOYIHfn+G3
qLdzI9m5JcL7Qvh6xViM0E7QQBCmuhtz6/Bwb9hDzD5ZTUSC6rx3+XzgjKwDruNe
YIM4CAzhf3N6uymt73Gv1jSragkyXRfZljSBjnGkYpU+CzcgScI/UmdoT3U/J6Ub
ffmltb3dFqA52ntnjm0/DywEv/7YawA+7geuCREpDrqM3vBOQ3giQsZ0R5qoYPXK
9jCkI7zbbaOYy7etChMkY2g/4bNA2oFuot8Z9Sv4PVhsm2zRYVwvnKhbSt4KGwPD
5H1FFbG0dCAWZJqxawVuQPbfoeCBFFVMbHBpvCRY3dn3iNh/t047zBuzll8DEFRE
oUC4Vhwh1fYy8fqQ7FxsD4LaNJeAjBpRu4rtAfiYI7QdALVv7n8y3NWDcWTJc0Z8
ZwcRIl/t765rrL2QT+cTCbgBCfbEmIlG8fy2RALiMRRJTBwhXSJ2Bk+zCYvLH7RB
xPPBw9ONufFV2Ekq8GDeYQ8vcPOND1YKHAYrrt1BkNYLQvwbpACIbe9YxLtQnPJG
lmkqbwxspjNLyMdr1i5szfNBzfPtOXT2ss5ExgJ95TJL3/Dd93A/uciZizJnDrV+
0YV9e8dCt8gDaualLlcJLjRXdWp0J5hmxRblxVIz/an1U1SeAti/jznLby4MN6vo
y9UstkE1g6ROGh6DXwfvOWL758ehq8IUzjDtIP7Q5/tZopOcibiY1iGYcOc10yim
Og1ilxSPkaGGLAhlGvx66u53AMp0CPG7gnAbn7bPSKPlZcoCb7gzH1dOYJof+olc
RvSKGe2nVWWTmy2BNwQ7eAbUz0L1KkvX4FMGA8gdvERL2QAP9xxImOXoFUGmdfMR
yJ42zgyWhWbq8U+28dLA8YrTa80H+u/DW/zh0URftPCOE5RdNC5CFqKBXDy6vEWZ
sZijU6f8xuM97UKVS0R5MZtzSymxLXQRsai+Cuhz1+ppsTGBcvDg2Ielh1PeM0Qa
iPN5nqJT8xzjgwoWa/GE8bMx4eRco6B6GfV2hC6TulagkS5UphVLxF0R8qb+b3QZ
qR+vpzOTUn9lodkWn7Lq+XIFsg/vbqiBA6gipzHRt0SkgJMfQQy6dUHHTlb2xSlg
9PgJwIHjx1IpcUyMSQWKk2dzR8yPOxdbIjZ1jctPS2M+wPMr1TYZFnymW1TK1awJ
gfbpzJG86uheV1bHJU8sVgFbG9Ot7zrOM9IAr+iWqhCEzyBgKuv8kfyTrVbMChnZ
YaSqYr1+GzNQHf3r2uqQKUEMNfT+K+wkSa0ay90QA0s4Z1f7pdCsAuHNtBEolYsm
QvOHgfnfvtdK/lWHwSZfUANq90cgyJPnj5eKlNq/0vxW8WnBChlChvA2pn3uuayB
kwbbBpnZKt4mV2y+eCGzpoyGBy7lXXN8+FMoxYJ2ZP36vI8vBGFZMMsKnpzvDbO/
jR4y6CNeVNB5GdBjZuxp3DEh9beBYzAEdm++8qv4ysFusTENVqtm+xV26J149EU+
B6XPjEbll4m84wUNsJKQ4d7YS0rJ4P+lDoMWJe1a0aflpdJ8FfpivrybsYfEonxJ
L1XeZKz7vJ5Il6ee3vf9xl1osVclft00IZNtGyspFcm+GbZmC2vjGld5XToOMSVD
5JspN0AnaZTtcRJpREFKyZ3WUQ7SlMZgoiuYlbOTS4eZMUrgmQr4F5tejLbFWZMj
qm/ga4cRCeZ3OnB7cQ/v5IGKUZR8Rtk5NCTDiEe7eg14nA3Wt1ceHTaYfOJhtors
vtweGhmxjhc9mwPnBD0g1jPP0dsByz/8u9Ws4Bz75VZjufvnJSeo4f2I+Ms0nMat
fqf4eO33vnZBIxkRukI8UOvKZdf+TQev1/leIPKNMK6UClfxXyFLEcRm/cwusc4t
5omr4qIoUOHyxeLsRdHoNlRoQgsMvfSsAGuYz5btB8AfZWJuLnlHxFGPpnxULnzW
PdVv5MSLYmKNjPbkMVtVyUCz7Y9+UL/DkpkaxBPmwkkBaPzTN78xnwhispOc1nyr
HQ9+7acYmVyc7F/gISc6u64corwTkJ7AF3JOqv8x0vxWlGLGJAYagDgR3O2k2eIE
qg5qtC2k58l7hrVbgGzvYnKwNzEjsDJuZic25t/nieADwXdseqTc1p31OGVurvtw
4jmiJKmVXKBqO9j3ahAnM6cIYwUOmOoFasldnKFjRC7/InOAjHxtv/cj1n+n2Guk
A8ZdcTFWiQls/LbyugCbtfvoxmjFd6F3vwM9uKONGfrXvx2iTshgceA6fYemVt6U
zhFYvT6vPdhiHBN8W1Luy2+c9xyIwcdDm4bobihzp4RzlD55G/eWF+QQaFUI31Zy
mfUvBZVGS0Z+l4ck68N4DKcGNFpTlzk9b/Sm0I+f5fTYAEW2y9qUBKvNpFUTdF0L
cMAP+hvxCHP7WreQibcS5vR/sdzniCRgwvrgrB/zW1YpsQjhlfYTYOOOGm6cLTRk
CZEydc5QZ/H10olkuoCu9hhtEXtCwDnyW69923cJeYD0m65TTGTnFM3wtvCvtPJD
COztweDKKfHaplAtHx7kUD5QOq4eVFpTArWXeWdQwRaRDAbs2U+ezegfZuEZ5ZIB
M8Y05oav34j5gUSTYsGU4zgHwEWI1kLe4XgvJy+YX27rT2uvqhwswWccP9gMKcm/
I8IT67c2H5xcjEreLid204vqzEE4KSWJ7lcC2tQzKxBQFjYfmBqtLsBeB/Az3nR6
hAc45OuZ/v4Ybfv0Mlf8zlxdVbh3tlXq4NmRfkkpnw8bsh3w2GCGXSaCfOl0HGMC
qnKszt92SHwxm1QUQv3+h786FpI11sKKIUyf94DNJMZlHC4Ze/0n7lllfY6xZl1r
sMBm15EaXOiGDFOcqBl+WXmZYW9pxnbGlbXCPJcjOJ2KJaeFJ0Ver3inM4ZkrdOm
mvHhUpRJLKtbiTUFBaAKWsLNEMeUTIPW489+zCzDqgXZB4MOlKuJosnxDYo87xGC
PbNHLen3+Bj3tJ1HYBRDvws95F8HnHTAwDmBn5munlpQeg2q4X9RPe7rqKhOTOa+
f62BC0TijsaU3ov1whfWkU2JcF7yRGpldMYl6srSra9uy+9gjpicTNjxKyFYbbrV
LtYWINhGszVSB3YjpepK7UWOh3J3JsUE0+RoDxviaXPBlKzxGh18L3kgRuWOglPS
GD5WiiMysFTfuO1S5vWcVWC+KtPsY0oAhqhrHdBpBS9Dv4F8VxrBJyrnGEjCXQzw
Xt5nYLdhCCzHGo1sGTS6dLPmUrn1nA2G25svVNuAazKHqautCgzPi7O7k5wo6NVp
GCFCvl3XQQbtX+15y+oocd1/BoBKRlngj2WcPP9mA1q0Zt4Q91zVYWohEI9qtn6O
c0hqn5cQQ87hiFZRpzv0h+vdVyCmdDscUu6gMVlnV7oS5FgaNtZMU9hNf0V1TV3V
43ADvv4C1DeK8SUF5Qd3UlnWllDsQNxj+KWghbiTb9CKR2/cGy6Y6DWwnj2jQ3De
Jb9Ek9rouWsWmj3eHjP3TCTNGlc206ccnkYTN/iBeiYwaf8ASgTcFLr+cxxJPn38
5qQB7UmVa+wRaSOK4Jvry37+T7uwIsHtyxI6vzTcleTfY7u17YkOD5hnJMtEvHOg
f8MhNMotDBEucOb9Qzsq2hYEPGOt1x9HRbQYuel+LL7EV7ughmUAkhEcAS9PC+op
ERDwfZO7ZrVa8bwYTTGE+msjGURunFG/SorFwLB8CuPB/PfrRYOyCFTs98BQrg39
NWyYURODxYacXVC7hddb4m4oNLaGO3T9qYlWZVQlB8I/kTNhARdMcbucaLD0URCY
Kbt9iAytdZbmRkR5r9KefotaMSg2oWkBbQgcBPswR7x9KQOvv073/UkfVuAm0rbB
J5AOpbdpqFpJYoeo9g/eMguHEIHgD8Hv5zcjRJzwGR0hf/DN4Pz+V2W/p1ybeJFw
xIqhCdY5brF0lpefIfku+Rth4kwLTXv0gTSQsgoMWDVGdp3dKeaVC36O7UXmdZYb
FTjzaLNJZ9W17EKDgN7BVBxNNlbgkUlzpk1kS3xQX6qBLl0vDDPbmMqqeZlGLJ67
vASo62xGnNcybQFKrCH77hY9r97D3b/RdO2OPOUSB+9TEYfqf7Lhxq6ba25laJU9
HkbJXK8+PPt4AIzcQVev9BeXYSykIDe+Rmgpj/11Sb8Hu5gHw60v0geeDk5RVHbU
6Paj2OZ9lrHcMtc5kwChmo8IjimRiCTQH/H7DBAFRVJzUwyqTF8WMO+7jUrtjx4q
woYyVk2YB0qlbgJ/WeR2WzbbX5hZ6T5bdOdbQpZ+f9K60xrObtZmjcdMuaXTxcxU
eFA/QCMhye1JoOfDW/Xc5rf5T7H8Sx4KKyCUcM7brwBkiUpfY7OKF1BAFBRx82pE
+v5Y2Mli+gjxwyNDud3M2J12IYBuDAIaVewbOeJv8orwF1ewKpwpjC8vTBYGx6o2
lRnMARmyxk/vplXQZtK7dpsFFQwTxrCuojB4TfYMz3MSl3cUmSbrNFNnH7o1UfD/
jaxnSmy6ldVw4zk1TLvjo0vBtIuMRI9Uon1P6MboBmzauks0e6xlqT8VM0WoxG9F
8fMcnK9xF8RhaI9/TELzNGnKZJshEguVMYQQSD5pr+k2WJfGyP4m10FmNwemUQfF
BEsuxMf0DRZWfEL/WshkJa8WYigjaGd8OElYj7nhATCgA2T7Kkb9pmLeMGVDA+me
o6EsUs5m/XZsCealkASPIKdOXHmRYY388Mm3l5wsEwLEzYOykiLg/0EaIlKx1y9w
aQVV50dTLqvWwrRtnzI0gyTftFM+gadR6yqx17x0+ht+e5f7obqv2baaFh3TQBOS
L70Meh/P4v5hOSkJ+IJK2AnyrHX5wH1R541uuLBCfxenZKApFB7YR+qUHQzSQFL0
GlheTMc+6utciVGZfrmtfVNy6O5S008qSiLx35lOaob1+F7gBnlOD82YxcUyKZui
3je6DarNKyGb3/Gmm2ICRiv8vXI44FYCYkQ19tFEa59KHM0f1UnDft6al6KMEIeR
QUvA0Yld+QF0tpDWShV6TyCiiECfln1jGIBHqrfV9K5cou/M2LNNJyujEL5vv2nm
2U2rUtq/S8X/oL32Yyt7zfJzLEZnzh8N8ZfzJgF/xG0au4FNxDZAQ1CqRyFHzUeE
qDd8JD9ICD4+5muHqxVEyjijP/JZBpGM7CF8bLcrbDyR7tk2qngevpQFVmdNwFdo
Wu8aLg2vlZaUbBGXDzajIfmA8RImlj//yr8udNq702E/V00qvhjY1k1zXcYPBkP3
uLQGzF4ax7b5Vv/saepR8qpFtIiSYklKqrBFc8kh6fzOGaEiX03v85nIv07/RlCz
M0wwMpaXIZGVu2x76onC8J864Va0r0xg8AVU3dOzNz4ADEWC+JRm1oktKj5TynOM
2OfG/na3tuFcMohc0E4yWHW6Z4syc1AWGD9a3Qiph+oAyaz8EhZXRor0gFjV9K9r
O5YSRChwOwt8APsNqDd6ZGkHMJpAOe/AgBHznpUSSJFxjpq8aOpl/PIzM1ugqP3b
xvj8oNU7lxgXQ1dr5U91cE35TZk7+L7n1XH2xdglBVZo2j/6pp79cXMYSzytCg5h
iAcdlmPsYAd7G6Ixg2PmJlxjqxO5DjnypMzxRGxHbcZPLGnDmVZ+6anhn31thMht
ak2QPrBmiCBuHQF/4TAyfcztb9RLemsVD3JpbMSO6D35tLMwl37Eb7tOrZME/pVq
VDbMS3YXEKOZyI/ZYrp/tr+DAtovlYh1QMwlpVKlR2Me+MP7qz+oLeKbHKrPNLnW
aGt0Wz8XdLJl9RwT4gjoIcfgJXJ4eLsjhLvF8BMJp42zg/WpGi9RuNyyux9EZyAI
Bsmin5gmyhaZ2qjGgjA3GvyrksaFLywngENabC6IJr5bvKQUfQzNK8aG/3pLJYxF
/CZ39fd1GjigDLroIfJEI7TCTORc9vq/8hru3JEe8K/JzE1xu3A5cNhvje9BFDnq
wuDqMBbz0+v35sChXIDeOY6UYDOrmAuK4kq9+WrMlX9usV8NK3FXEK9QiDzGIuCQ
Iv19K61JTHu9N5Ee5a5VWk56QF6iAc9c4LQ3lFvYmL/YRTJHIyO3anfrw8DDhoc6
WIesVW823gzQs02//Q5guTqTd4YeQLVXlhwPe2rvy465a3nO1pkZGoRewUqV79CT
feNLT1RqZj+DeUXcJP3czw9S2dkOxf+L+jqadZGb/D+tZo9APb/li88dbt3XK5O+
nlEvsPl3Sk2aBENwQbxrorGdNmxFhJu8LeHiXfLEEN4BuTJddhmKr+KhMMZpKYN2
qYQlq0LEPOWC+0irIJnG10qCHnOZFXahNza8eHhIPkgE5XgijV2Dc5sayBE97NGQ
bt7ZLbCmkfLc0VvBJflywZv4DQYy9MIjgCxJRRZOkW3q7fllGz8akWTcnb3qGoKB
ucNimwvcrZx8bfL/KzTsAVNZi4IO2F8tkUTqSRXSUZb80j7jhbwNlkOZKHCGED3W
1qQOY1OnMS1QBqOlrj47jhzNTNyutMx+r7gqCdMmbULIp/4TBEa1yOSPQ0UvE9cy
yiFaUTMVUyaQ+HHNZznihAgzfxnzrE+qJboc/h1eNB1pRKX37SrRZKtPu9ja4dN/
dRlhu2zQaCqlShuU3J2a7dHP0eREqM8eYMV58yBT44F0ETaNpvqjm7m0EklMAY/y
PWq/R5cnXHIqGMvRyNG66o18TIxslHq56FnZUPJBwJa6ztSVqRVfbBvgfhNdSs3u
852DIuNJNMpGZ5nTu4yMKDG9Nntcihs7KxF7spKBadqoNIXuoYBGmnSQeu84PxSx
R2rWpcx76MxAbAeH/+nlMl5tkr3hm7ZmsEPrXJZu7XYHLwW94TTr0scpLeQql4Oi
+diun1OsF8iVYo4fLiXg7AvbceyZep6QSSPiaUMbxzre5pTc3h8lhlQ3vqllsJ6H
54rVDUH7gPM8IrjETKa6zfnwlu5zblpPYUGdY0iiUEUoRduXN0WzPNGOiaA3h8tM
56ROqEHM7G7E9IRAAZtra6Eaw33LvouUPRW0RhsYmlXVSxHAey9mZWWKlxJtalyM
NJ1VsXswWIC+hJiY5wfXY+78jeiqQ0RCosgwxKjdqLAy0FHW+htEOQN1S+ufTCpp
narITp0k1s814gkXUxEO1RjhvEPInpPQF1NX9FCqGSemtAWYj9isz60dRnrS/hfU
xnRwwafkCfAFTtB6P3+aN/7fWQ2xyi7nt9LBcTGM843LQ1GZj6tj/expD/1SZ6Bc
VUEZPslE0ENsvAUoysfywr5X5x9SW4Zoka5dkNexPa/bWFyKiBp91bpLjE2GcDIg
ovt0hxqcMb68Ul3h85w0GbKN9HWjLiXDsNQj0IqnfvhBf/y/Wz1QAegLjMAITmQ/
jAI53hLqQdptjQzJua+xF3YCzkErpUdodz327lTVwd5Em4ymRkL1bl6Y6pgO+Ifw
0QL1LiRtGnPA+t8mkQ3VLvT51NjsGTUfOP2bxCaPbjlSpvus+ImKL7UNgMlmgWfJ
ek+Bj7BIntQpmUWUW6MfbUt1pjWXTdlKi4znLRWI6GtTOmEOlPBM4Z9aSgZhfEBU
07p7t/toE5Jz+0A4Lb1EC+PwqnS3c7ed31FqvnfVyWz7wE4+a8INU67Is92BSSsX
gMyvSC7S3wHwOM4VdRlO5m2FLIepvH7IJs66GThpiBe57JW69AtLvx4GtJLPrS7f
x1MFhgL5fL7MPNniN3v0C+KwJC7HZ3ivUu1A49TcVw4D+3nMMdryo4yNN8J+T3K4
3EzN1/t+bs/m8jjdK6uHeYGzI8ZK9TSVtkt9pHHKV7f1jpE4OPpPP+tMy5iwlnRd
qM+w5FdrWs4Xjv5RCLragj/FsmH22fEyHQY6/W2OAh3mJtRLH0b1s8T5KGwiojVg
JqtEbwhWpPEuD4gzsHFSymXW4JC6ZjhLGUAhSkr4fTHbwrlufCiyGB0X8vG3nV/n
bh4Oi5VKQeHQqBIDH0ph1Wgj5+E29to4zoOdSUtFfqw7XXncUGvrHQpLFEwsgRAR
t88RyxVN1u7slV90fu3C5aEkg61ThJ86TcMFvkCLaw0+rFGkZvoYcU4DmG49pxpY
wYgLOHJFmDAKrtoclXLXqJIEp5ML8IrRw2gzZ00vrrL6XUuvO8PRxYKLtxGX3VeM
Hcf0/N7L8Keae6brLfoImyIEb1pgut0xraFDPEKFmwW8l0mPHtO0tdKJv/vSta8g
46NQmOg0lJetob/FLtGgYBtJUPEcymE17S48w2FCiwsEc5mlgetOh21+H6i3I11C
QggsAv93pMjCNoZv/NfaSE9I9A5xS+rqbu3nNuH8ombYw1oObJtREReldVZLhm9w
X37/VaGRT1BbI3iYnRvhctnK0CNhRu1Pjbc2Ukeq4p9PFipEPNFPimhEZM8XWvxH
k1AhqujfatOunuFBvSwGohGy7lAdDH015DTDYqLkasWBx8wi5KeQX1gsOOB2My95
Ud/2y5dZrEMrsrAKuDnvaFh39P5CoY4dXOZWTi9TATylhV3e0L7SPwBQfQl27MjP
70+6ph7u55bKguEx2dEcLcu6tUd6jd4gbKU9jBZNHsmX8yOKLQd5RgTaNw1/qGLS
U30CQr6iFPnDXZCVxKPMbnvl+WUJSJ92jBnqA1n/hs1Vh0klv4rscOB70yve5EJa
FE0glIrwVwF0pMj/PNhwl2UoA7tXBU/lMX8vXdnnsRPhIQGx2/yEwmAOiIbVg8V0
mq3Ht9//12yrhTx+rDEUAfJJL6UHeCrPVcwS6cfRKHEE9Mby6GICOeT7q9VHid1Y
VBAALrejHGJsmfhzdY12XQ2W2DUjzpc5xluWgLKu7cJfKBRM0dgxLgkQPI0xUcMa
fhnVdt7ot03Ov7nQIrjS1pLREEcZveEMwnQ1LuwCWOfibQ/2IAclADEp3NPeqlwP
zDbwcfc34twT3fw5tDlr7E4dWBwV4QxeXyH5RVcT4pnJxaeiJR7BiQG6yaWHFWE1
nqPwhkIbKBh3VUp1GXIwMYlSpjQZ+sTtTfWyF5g741rMyFfmVuO3Nworxkd64iXS
N2GEsRmVZcWHpUS/iyC8ygctBu4rqYZt2c11V6vafKS7GRtNrzBEdFt8QA/NIhIU
WDoYVLclBgokcy6cOyeLnxtygM/LMnlKROeCV8Q817f9xP6PT9RcxcQLjLthijVq
8Iw7tEbq1kNwqn/VIWCR6O8Oy/WGQ23vhyDVfBiI6OAan41CvSzU30w7ZNI1Dnq3
mlMtrb7+/bH1OPF2rq5PhesE7hgC6dYn2TORpHhYvrTXZrxd7mdzg2pUiLdI5VgG
oWFqa9hAFfleUXD7ycLDsTIJlHj2nPaEXm2u3GoNiKzLFV4fRsRWjxP7AC/sTxCl
InaKYd6GJFHYkgWaUO2qv33WvxqfxzOaw1KKKLy7/eQzm/6qDeIeGxaR2gvMrXNQ
Q12r5LPvd0xuBA8ZVCF+tjigf529oAHwBvuiKbfXhxlM8lY2OeumT9EJwyMGBC07
ySeSX6MuzfAZ0fkZtKGsdQsNOrfnBOIYHZLP8N2faMDA33H1CzukPgwfaw2rP5e/
mXhjdM88QghsnyiKeMVL2z5wQ0KxR4E6ot9WbTClXh3hWQRBTSY34jec/IqnOyQi
xUZESk7cGC/Fc2M9WEBfapFxsW7aoRuT6Zfx9a1t7caaIm795tcf5LTvkEYXvf4l
klsupQe+NAzpUz7pkANI7e2AuPn0W5weJQ4dyBnmReCz1NLYVCETrv5t7x9tpekk
ETJP6ah0ZlACvtY2psSPNdNbTHbHNIAEa2KdeqDyPaPd1165gAx0D1cpyqOUj/v9
vSSuKyMy8KjYFg6ndqYjlzKyOvY879lcUII94zxSOyRHkXPS3VzCfglTFaS0qNVh
hHztmXFhs7tcK3zY3VtUaZ+c5yY0uSfECwhdZnqU9hO+CbYmWUkk+K27U5eHRrgD
eg6hyRiki/+Up6TOqGz1NqpkV1qdY6JPbCyY54D3oQb3DfklofrPYEq74kQHVhee
oSmysfMvmjj4uR5La+vnU5ZoX7QwF2EBRqpiOCQRDObl0k8VZq6zqsSUXLDUmKBi
5OXmQPyjla9VXhDvSVme80Gllg7itljk68jdRyyMgfQEEXwabJFAiNn2BXgOBcfx
6WHN+114FuNkULSU4t4jLZCFHqCMJBAn2UNNQQDLq6GpNr1wmxEpEX6/zOxveja3
V/HraGhD+TmdJdRgzRyxmN3Zor/E7wWV9GwXmrP3hNfbO1gHshEY57q7p2x50RFR
uJVKFjru/zZWv8cYQd9T3C63FqjdfIFle89SJxBIF71/S+9HNZ3EjXYtriWk+L3h
2yYnjjyeciZ+E3Cw5iNXIH9rsMckS00P2CqvO2XbZ2H8KqFIQgL2/sF+oaXw3aId
At6JolL78plFJuqzVMh7iZ9dA5/Ez6QJxwA/AtVz5+vZVpYXPfVh1lgg81PLmn5A
RAeP60LvfsecesXBdMfCrdzvNJgpIUIxuw87zUB/kBhDp2OA57nkbFQreQMB6fS0
yEHXH4CSjUBK7ra3p/Ddr53asNHfeA8wIx40WaCsG4B0NpVPRJwfqbBgTbS+cvt0
aLzresjqXfuAWlTn95JJ+bBGPhs9WHhv7GoFhn7T2rhYrkl4hYW7+IXOvLwgfEgz
UOmbdG5NZGPdwuym5lS26tmtnjTQb+mBsXAHTaqNLO5AYM6zCWvaLl57AsoOin5b
WyqsCWtCpBjjnFo6gQACHmrjBZWOm7uXCQL38kC/u9N7CVr6BVpqcaUdswqL1mGG
Xz8dFGOKFn+RsRjUF5ul1jfk7APU83xZApr6jPLHRw4sZV2UeUxUQjhhSg0ROvGH
4DW3GMdqFySxTB3frwVd9h/On//X3Aic9t7ILSL7/DQFPdhRSi0i5h4lH+03TKmW
RhDfy0KKCQ1y0qIvbubeLBY/hMQtKcMZQiPIlAMxJP4zouuBcp7pefuKVbcEeMnP
1cVFwuepXQ12SW+9GGxlmAMEPoZLHzDP7X7IQpkzjIsbwRY8Sa69u8rLQ+Fkkqkb
9YGlKo94Tot+6OTDQttKhW3B5r1OUym4OzCUJ7lKgKSashZtAYrkunkdy4/jqoIk
MCaN9dCWoixPdLRd7T6hnKm33FuSzOe/7U8licciYuZ2VmYcoxllndeVwQGemYD7
BGXbDp+CrKXhnSRArFXYdLKs6+WyGd6gYA4JSYa4tI3Hvyyg17y6iffB3j0foPTQ
OYQzHCRZdYUb6hKods4X3+UloFwql216bB7cYx1+Gasr7Du/J/0Qyiv90HZkiVUe
lHwaPEuikeKp5xKzcBCHTmESIJ2JI2b1mph/WpXyAtpiTnU0TYKt3BejgSnuODOd
KxISELhZ+351d+UN7BpHcUh0YoegulpVOXDUD+8FnpqKrk3nvoqthesIpvZwAy8b
nwX27xfoHIvuc/AtHtyZki4yMC7n/Blb4JS/BKS4P+lNrnBTT9mfQLVZXq1MxqBq
E/R8Ohvhe32PGqaVPegJb06lq0gB3zTyA2HQ6VJ3O2g9tszANfYJvSpRY6FWPMx5
So3SrQmoaME76GeCG2KykFCQXszHRHWNZur0ZDcXSAq1SmPxGy/RITwtgbc5PfLw
+5CxpfFFLcm+R8ETROR1aSS2VUXITYn/3I3j0H0HAgnqXnBZEPuBqWT5CDfaQe4M
joOLwPAaeQv3Du5xSEomuqW7YCBrvT8DXuWzfYAqfQ0bE27dzwu3W7XByGkPFWcN
iYef0hnP5OTcfNjkXhWTIvTcUG5yQQlnscvKqJ3MR0XdQhQoLB6HmUstBxgdr0Rn
h4jB8nSJXBlf3/1DNlJw43+jHsMZsVf1QKiKML/+Rn6R0+NxaLhTeXlIh69z/VQH
iiPt/xOpFBJV4e/0xH4YKcebaliJoDaZg6Z52yt9ePcglCX0X2lzhTt3iO1WQVby
Ge8jUVyeHeFHc1zLEwpTqNQRr2CsoRvDp429oWLSAjBzREg6r4b53bnWBCulev1Q
RCi0rKD6u0JYq7lLzOVeVD0VEM1kGdJbT3ear9HE0IBpa0iIZR7rcH3JVyCHVkmF
XizibJZCov0u1yyHzgpnhUg8qIOnWJ9Mj7drtyI57uE1GnyVjexFSdCnj9uLM0Nz
1juuczoAizlH7uUkcJiIEzu09apkbiFTB2S5nrobMEUDHLISGQ+NK9ltt2VbO+Ji
V5E1nS2XXvNqIgYBNJXau8hlPzblPG9kfwWv1olV+9NMDTN7LEkwHy9+0QiocrIz
KFgsQ95L5aryon+xxpuy1JosTjQXhxCoq6bF5MAzCsC69gvcSrPoWxw3MO0oYvjz
FbS07GPJeJvLsUvWoU8aA7s27IF9pxAcSkuxM7nIFDNV2he1fmSNfLBTRqZGzDmZ
wc2NkMf9TMFnTjKiDaf5+A7jKwo0vjPjFiwvfvUnSrweP5W4J3hkSvGMPPkLmF8m
vl4XGR/bi72z3Np5BY9A1VlUnmeCw095EP4QbcD50n0Qcqg0+vcLy/SiFrpkLLdQ
ZpG8wrpepWhS8yn3/ukelxfArwmN9j1O2TVkFqI3kqkf8TosNh3uCKwOnad1Qlfs
HMTimhMVCQR1cI6up6zX6GJyKIyJtvcgplHlziCycMlfGFFTZleascoNwa2OeVSI
mI+ET6jixTtLcTkNbN3C/DPrnJgkIB6ctbbA0nF2OfFrbFesFFxpx6SadZyf6AUu
0HufU8h4EYe6Dz/rVf9peKNYQRNfpWQgOy2fhh48P9s0QX28a1agE1Li10OCy/eQ
8wIaNPacyxBUdP2kHbPYmwIOxnHqBwGh4X9mFycOrgBam/cf1HKzhnkPaeeYgINo
JXe1H2Zv3bH3nkEuB6Tfyv4kJGzn6Z7CqHmc1muYXQnYxEA3KbXV/unVDnp5ufNK
uIMnu/zXPhgHVD7X3VpWMqtCDNe1pYyPlhOZSXJa6OJi0nedorHoKuJRlyhEs5gW
YOmGDUK+FKv6iqVb1ejlmFg87j3mf/xzOF6qbVmY+7b0Vgl9iwMmZTaBkS3ql4kE
59bhI11MDKJpt30MvQOX0Y1IQpbrNw4Rn0cNXK7Fph0D+eWDwmcvU0PikftYth2Y
7z3WBQJboZfzdx3f8W8i51i4f1s6dUu83Mz8AlBohSF/9YoguG6zjc/aRPxeby9+
NCsG8DUsIafO5O9ENmHbHyJ7PZWW6RrOj0wLavk1dt0rChbKZHgVeKBVkl6yx04q
5cwhwzO083kMsvo74K8dIVz8QRkR9LY254VA8ZAMrvtkpP+X7NaTvh2PcnyJh3tN
iPzXBXJoeGgT/Qc1oASzt/OYchzoWKO1KEX1BV/dfPii1NoZwX8xJeyBGYf5hyR3
+hqq8ELRAgW/iMXRWjNYXnQanhTO+/+fWCZzycbA3QDzisrM5QiD44K4q1iXYj8A
hZiSbLQIcJWR4XB+VAV5pRlFm4tgTk+Jz4fC2KpFs7oTc/HTUzwONhVcQQRWzCbW
DvUUoyob9GSnp+2rU6d8+kXMc8jkXGRcXeZmXFynfeZiDeY/Yj4/3TlGqv4bE8Gn
sF3IJl13kroixQsUXQTAJt6OxkG9m9TfnY+7vOMfce9auNJXWha8bqtiolxRfPVB
QK4wBODb/zkq6391j2/tQk7oOHKdT6tiNjjHBivQB5Gyys4fGKiYwVrE3Gaq8ZSn
2KP+vQvW6vJOK4MGSknA5JWN+kLwJjs3kcRK8gk5cf4xrwSB26tAbqjha4fAhRNE
vX22YFk/Xb4InMP+UNVs8QtOac7QQoue2T8uXOx6/JSUeStFprKhykgDskOic3zE
D44tRCXZajBVKf5OQbzgREpiDsUPJZB3Qe64Zq2BuZN9g3cnXXkMWbl+K/KWTn12
UdjAiWOIegnlOxUTrFnz732G7IHoX6l6IS69RarvgNajG+dwHIRJ+ft8ad8QaUuI
jRipq9CwmORDGS5HwLNO/3Vvd4GDl4Z8Ln8AAysTFYQfXdioceUEpV+d1eZGjxui
2kSoahoUL1Ps2+48UY81BY0sgSx8h1GPfSMeZfqbuN8KBQTarjwJX8fi2JnXHyr5
xOueyDSUAtmQBc7bqwpJPkSXfe3Az+ocJfaFc8DuX1TYxIyCfDBmuGy6tnpneI6w
BD02CYXdhuRfUHrKgzuuh+uwdj8dOI8N1xyjpzl9mBghO+B5o9uNDQTPyRMrht32
vQgBOE/SOB5WRLI0UrRmU3Li9q0bKc7acIa0fDzoyb87CXNUnOzjFADrL/WbRc3m
pgYnFlApqEFMfq9vQMv0mIW1T5mhitYK/sjw+9DcQnsXKFx2O5Gue7waxDDjfBSV
dH0ba9atBy3gSyMD7R0gb9RgWs2g3NSmJemgwkejiV+tl7fCuDBIkDXGiMt+ovra
dD6s2vDJppWUrZ+69MeC7yfXq6vsPPR0I36sok4QRluWt7ifTtaTaTuHQVAa/i9i
RwweNrssi2ojXCiMfh86GKs8ZR8TwakQIKmxdwibwI8uyv81U4X+Y+O0CsQ6vAfJ
Sz2/uC/xR9BF8M7sRCXvJn/umSCZfYdf3NJzytYRaSr8g0ZDEoqPPVg2gigmABLI
crRcbRRL3000yw/0SAbzlcgCSkS047X03tk2B6+kmM8YPrlfEUA4axjnq4pERIbH
+N/BjiSk/DFLL9OR08KmEaZYYiyD81UoBzL9egKvNvOvcr14O/PkMSKhjfAHhZD1
yw6PIvdJWHsBMj0DZpw4VyBXb6Cw+C5lziVbXo/Pnw2X4rjxAKmLBAxAn6PHS3XW
IxoweHStCgRnh8rGFEJSMoIDLsuFFlGgG+LcJ2Uf4Np9tegoNtQPON1uWVFaLmkI
PAvATiTIhxOa6msVEVLWyQmcY2SlVr79I9Oc8rC8P99rqeICQYfzcm0d3JkEyLSD
4GHElFzccB8CqEL8pjzmo+LP6iej+ydR1MT2s2mwsYr/b367UchWfED/CY0N7ymR
B/BcaT5PkvmSg2idajxo0QXZlrAMp+9UMi1p5J3sTmeguxWn1Rmr1f1dPAELfPoU
w1GN+gOILSkY37McWXNMKPDJl1hKRVkgK2HxXc/F+KbDKHiHuDx0NV8N0YGFKWOf
XUXfd3GN4roKmaidY5lyXFCQllNzqiQds1dEo1ydw96IPAbyDQuLZnTyVdQ/BazI
D4mob4XzeTHpWw8Ie6tAlG+/+wkr7RKNT78gNyIuYBq4VoD11KCrPeX1sf7dSNjC
+Ls99Onn3adD3jHWbr00c1jyeRuXdV6409P5I8y3XOQBhDGyX2c2IxkMqqMksxoa
JtDHYftDFzFgG/x+UgyyPbzpwK6C8exSYxCrEqOLr6Px+RE3Ye/JkZnJL5aAttzP
A+37FuwAcsnX+U7QH2MKPEPt9pppsxOFxBzrq/Lp1wqDnyXvEZ8SPus4UnNlOJgO
s2hInhtHCkCHvRY6luScgSKThWGFaMZdpMtZ3DU0bPu4btj+7Ek0R3KC4O+TUjpb
n2zk5BQFt4HQAeQtd9eLSrSjSHgjh9eigRIjCtdRGc6fSc4a34kOfzYaQMBCbYbG
/nWouP66oa2EK1IhiHIN9VHtl0c4xndNjgiXlnW1ZUdkMdZu8raqP5IvkmlrKkxC
Tk3uRWOcnRHQxO5tmVbxmLDBtr5AB1nLMl/r+pnDWdFlEHiVyo7EJ+uaNy5yzwxF
4GJKwg14SYceC7fIzkW2/G3cc1RjwwC9Tr8DeFJTDFH70xEW/e4PStgdHS2jbdbC
SfnnR+ezXY3fFRSOCTavgigaG+WFjgqilkEGRxOsVvbnqGDK0OCHs437qcmXugs9
duRyT1rZ9lnIbvw8VCe+JokG4wGxiKQpMPZvytYnXkTeuHC9wc9v5q8LncZc7bTE
dZ4pvhMlosURIqx4ThMm9a5IsFXhkXo0dJ5ivq9clwcuU4DTUTU9UlRM0Bf41C5u
vqoP1hQM5iQkU0y0ywuR9/G2aCPAx1kFztWMTRqu8mr7lANxhAM5ScapECDLCPi7
HXHfk+cYvjx0FkRKWGhPtnlsYtXznz4VIH7BtSvPYSatnN83ZlHBbD1ABiJLS1Dr
6dYv13e+LrFtgfe7Wbjf8YgBbfnnOUhZdXAD626mPlTySqSuHh+xllrWGvsoWrP+
4LAyfR0E2j953GZUm53YrwwtAK4igsvTHhBK4e7uvY7g8w7KPdIEzDknDN5QuWNb
W3Em/WwcGas5JpilAAI0xfUAo66ivvSqyN7WL8WZBIXHFFQFNB6QdJ3P+LsmxnWo
+J+RPPNvP6MfY8CViTJ+rfctGZHPJ3EOYjiq/z0jaF63H/EWg/sYYZ630tYNBC76
VsFbWIz4E2CXSbPZTgpNG0iViIcsPpDH9XFCt3VshakNsra5DSk20bCYps6FJe2u
52Q5WOTKscFiH3cBFPcYvhA5CqtZtmYVGvR7wFrYdAbRchoLUDRv8IlSnxhCgqnH
jXMHhgn06dHr5ssLdw9zDi8OTV1PLYHR1mfx8u3xQt/ieFka4GeqDau69U59tEZ1
IREOnHaTrlG64NQ+Mt4+IDVfjKn3LtJjCuZejzV/XV+6C41wx7mQZD7NhD8EOdw+
NVurILj2QWKXG2TzVYtNjzUtopYSFMBz3djQV09Zz2XxOQjgry+2DnqubwZJV9jh
tC2dkEY0tlrxBqp0TyolmG+8BkU9BaRWJTMd8OLFtzHOQclTio34TvYM0o9xRIQk
Jyv/LGCosEX5+1/pxvjh6VYH0XDsQm1VQ9rq30ploYJDj6LXBrOSkS48kydNXv0j
Q6HLyNgNNaYvHm+i/l0L2WnYK2tngMKHOLculd52VJe0mL5yVRCB7jWllAx8TvjW
HLIXH4NDZPUHDbvsn9pNqyakVdoyL+3OhiBSX79E7Pch8scBAoXcM6SvrC18q7SZ
bD4+VWLk1rgNIFqufG/Y9LOLtJeaAWwopCJ3Ji0U5mqZrG3ZvFfty0R1chiA2z7X
sBlTfww3AszXW7QwZxNsnb4u4HR+DZ+qhq5WBfqCHjVEuernXCdU2YqlhnI1vLZh
DCYIIr36W9stSms/bkLFtMwzuWSealxjjFdO13rebnnbgNaRN8ooAgVooB8reGBQ
OY0ZEhsla9i5wwqzSEqJLSlaoIkGmYKNMAuTwrVTRDZkrxm/WLJAFR33ludY8Z+a
b6Wfbtx+O6xX0KsVuJhG6rVa2ZmmL/sYDzq3qY7KpKi04BlW4+4PHvRTRjvqHnv6
7N0qjSd4W1vda4pg2eCkPfiQLOLykI4yJDjD0JKLCtLcvT5UyaHHpaW78thWz4Cz
Vrh9TRD26/N159aBfAaomfFqPT2ZfhwtYtiBaQyY79LwTtUZm1fCgCMsyNxAurRE
Pf/aeG7bp45vuppC2OaveaT3TczkJPgIGCW0KJZphtOoNaWyh/LU7odoASYnk1eQ
bJIHaU3jEAmWtDnIJlaHGYTZZcdkwQ1ortw4qf6ODWwfdYK2bbSOzfoIdzHzexkg
egPYdbHDPSZlpUevZxii+pWxdTPHND/Ot3cqJbABGuemEcMlPayjHHBPnlzOGT2p
7TvdAg9B7wFGHWxqUBxC2qHI0JZyGMadpGi+ww9OhDzflAKFEPZBW40O03ryhwr9
4fW15gjfz2MmDpBAW6/IVH9wQtYfVl+xtVWpn9u9d3LGUmStioR49Q61WOK9o3TY
qoL0aYhDIPglESiSwzCKnIZpM/Kefbxp87ZrjhnVOLy3lfMduzvco705Hcg6pQZ9
nQshbgOyLNVZwnWE+9lb6DbJjHG/aLI+/1LEwk5xe5GK0lP0cH2aQOunOhb8hKnF
ESDPHS1w+ZOTkO1TWMAvXDI175eSYJw4ZVqtPVVpos3BeWUuS/uVz+D3/mXmteRr
B8XKlpjlk5D3iWI3n0kj7BBXHsws/aviRKE9LY97Q/7CtvWSpMa4XFQUrlIKSP/R
CDStseqTmrJLmjXEO3AFj7qODVAJxLoACyII8A7i8WS//qy6U4KktuWyB+Q9ZQr3
FzoSaGN9dwf1n86PgkP41JfiFz948ia32wyB56uJGQdEqU1vqFweC207+JI/pqdh
V21/P1SuUoQ8JfV9q1sgRtJfI4vlQEe6y2ZmF7MkMt0kv/UN3cV8ARRg+ljHwV64
TLbfcGpyzv+wJlnqeYpzfbL5rIuLEg+0/y/yxxwHRD0ykWRezVl1u+7yYQXCJ+EV
kd0gPHeD3HBuTh7MO9Dp6w5jxS7LNgCDzSwnCi784hui3kKH3dJkjoE1vOTT/hE6
Xge9ZU1IyhtaKi5LeFpkcXPm89a4np2dHFgE3G+fSra/HBdkDeheO2T1+88oVAR4
yW3locu5sEj6F3G6dnMB/a/c2vCg2NHzyT0D0vGTgnb4dTTNo/OLEk9Hm/RNqzm7
Mw3pKGCIxG1sa8Hbbz6BPOnIw3Z8qPhBK4WIUoiBHLWLQX3k0JK+Fx4yYAtmLnIM
zk+p2YbP61pfvQeK/yjpLrxl01bSova2Oga+BClU1UkzoD+jJJDS3grz0YpGy9yY
7CWF/q2yMlF4/6LYRWE4wxgJd2TPASEsVnBM/MTQ6aLZnHA5abdTSwmJdroCkeXc
HPIFZhoGgRw3pqNlPwsKQC1josWTh8h0HBfrs3oinp9IjzRU0mbjS7XQvSCZ+S/w
ukOZma948ktaVnlwcRkgvuETtPclX1hNeIrZjkLsrTx2Q0jX09PcsMXj6qwdEwbD
+XK60cVzHnduh1HcOSEP0QWXefQfcCdgIm388glv8pBXgz1ipf2oGwqdoOuus/KE
0cp0h0UAR8CycCzR2rKUnf59coYDYDJUSmH5DhkUIwQfosYHifvEL4hymfQJ27S2
kVLMF0XuOjydX2NDNC5KZBnSpDe7M/NQHG3f1rMP8DF/qMbrsW4dGTq5er6/ffWd
yQs2QtVa6N5vfLCk3/PtAZ9nro+OXakKhMcm5ZmVzLqt5rE1gER0RQV5N0nVqzOy
rImDM2sOkS1A2jXbG2ChqF818d/3pwSTJmVEFQmAWNyGzxf7NPjXd7FhCNJkS8nm
9vB6OfiQ9ghKyPF4mq7ixez0fz4BOTjE5eKA61zasW7ntBPKrnv6ABvUi1bT7qNg
vDQJ3F+rUxY9ARVG7/okwi5UqSWP7Z+pMwQ5/DtqSCZlhPDbVdoUwXyfev50uxA6
+iIXhciPRpaigFcSWrfs0fbv2soj7wugpims/wSdluKhCcqKoOITd7wcXwI2NXOa
9UrNPRMiW65irSTydx+gOf1kBcSsaelcOIvEG5eSVqcw8F4cTdf2mqj8m+LUxEi1
uR+/arD6gs+DOHjRUapL1t0tLDceFHi96mCKBJSng4M8RMpkxl6uxGNCjijRLwop
TI8S1S2wjJ0AJ6C6LpoAQwqZm/mUSEX3UKZE2UIQvxqfda5Z+LjS8M0Jh6R8aRZA
kUyzTCprr7tk4DvA3WScVtAEKJlYn/YZqXKsDJl2gFYaq0oCPgfhkFokQhfuzuME
+03hQJ+qe1GxiH5t02AaorAgVCwtH7d+s9Sfzi85r3Wk2sWLnWI4jn4ZcdlIl8oB
kpZPoHnIGy6a0uOGgF6XF6CvQyArOLwy5sHriFEmOglh04s7z9l4VCT2+i6CqviE
l9slJiRCgX6nXmbLS+PlawPka8BA86ZFn4T3WALPMS+kCTNCmdQ+qIsKGi416CL1
jTa6MQJa8ks14Ee1a964Rth1jtk8vxhAauuwwDfncI0IWgb1XrbvojmDTUta6uRT
ePxy6pTKyWq+604rurqwtInqRLYwFNTMSSS2SOWjczX2ABbRxJTDxF+svnAaOYlT
vdDM38g6f6XvsNpXgbCMOlFCNQg+0R9iJJDGYes/UsFjaqIBKTUc1h980/30xmfB
2SW9VHBUkl2ehM1vvD8ooavlA47D0ojL/fiDqL8ycFfdkBeed9LaPy9xLOn6y7uP
oQuScHRrqqRETqOZ8D/2yIEu9SOfkFoSRfIIMAdam70HrK8Y44nyEvQdzDFrvV7R
fvXkGli6YrG/1qJEU6M++Y9nTZtpvwtWmTLiKPi5xGmF5mSFtVVjJtpdpwLQ8V7n
Ls6EIRXqrvLml0Y2VO3aqvbHGyWzhOoti1LyJg0KhM0z11YwJOG/UV3F2/EcgeMq
K92xd+a7WPNcY6gyP0RelbNvGHTuQ9+Dfj8/0KnVEBQqQa6/ktDXd0XzxVvl4gjb
Xl+Ofd96EEtYJuFvxMGgG92Scku+7BPlWvsXrQ9DnjRRbSnKhL+mLIR09afgzOB5
CIIBesUA5w1M61F0DRlz1sck1xTSyyD/hjk/Qs5/MeZmvrxetJMjiqdQmQQvq0Sd
+ORrUf4QyP7K7B32lqmwCOpN1/syZbRq/FqGGfG1Ymobid82Z72FOeBi2dx6ouVQ
9gtDkOI3+kDqbi5WbZXfuLV3O9CxSWgX3f9+YVcLxpd5UZ4VO3AltshO+gIga9x6
qEFW8x2RH8LfmpgUTzVQf2YSmetojKduqysDSI+ObkzaOnouuXutAwRBsI8dnvLi
lLWvBOA559tYIDQZCRTd7LTxqVFLPGSOc3hoTz4yY1QFUqbHaUs7ApweWC0+z/Yq
NIZgwm9Auj8RGsJpH6UybBV/PcTpKiyLxMsZeciEcT34I+PJ7YRHlZJkZ/Q5nErD
AB/elMoj0OniUSi410c5t9vq3rgqy6vNViAKgeH0r1zdnPc8TBIwFqhBAEphkYx6
Z4n+7iXQFEvivMAq0Ophuz4ojYq7DYQuU44Xc5pATgcAlR5UIhmvQugV1h7pPG+o
RUlXk6W84cto9LQKdSeDEVeIZX/s7p3hFWQbIa7/s7sIZ0JaTE0diW59Sx0f+haz
WgqLPobAIhyUy9x9dvwSXDErkW12cWyqOeAgT0rYFKvbiDUncIAxVpi9IFQcErJj
O1E1csRV08gMCfTcSd5jQvgJ7d4mGLNo8o71r0FSryvcaO06sbjwWW3SvbqAroYw
StqZdnxhN38HOJ3EBndSw2PTul+3iecvGehBF3wvtaI3xtDy6+UJ/7FJD3nZMjho
p7ESZXbb5yvtJTC1MGQ4pAC7OBgrkxsuvsO6f+LbkyZ4d5C1uJLk3PVqvY1xuKYg
Cmd335QkWWO7Ory5B/s4R+a4Y9N1rQk7pufY1phZZKPESlJJ+ZxiYPQB8gQuKYug
+Mb4jHcXOQeFokk0CMNyGpgLWxgDYqVC0DxQnckxQQg5BKPcsxZzb2w1sB+ZzQOV
KKMmqbQFOjuVRSfgCpSEG9EHc+fjn75m4sjcW5VXsis/KFuWdD7xf6tXPGt0kK1K
0ZKUU98Zso+ME1GcQXIZuqKdRQqr+3Cq8ahVjtsoFe/46aCFeLpmOApcMmQaPRdi
Fd1Y4NKDVxln/R2nP5oF7m9k1FXUNAKYE0MY1dVd/0gN5vRNLQ7zg6y4qZHYdMkf
XyopUoawkIUJsVds7s2+gdctmUYaX3N347QDKGWZ9amgCpetF6jGMY8OJ9vz8LDB
KikP3hOxkzoC2pF2QymxZgAbBwVh/q40fuj01rNZEerrdPIHJ+rRr+9sy6JEV0nd
0raaQ/Ql4OUO5FWzaKalhTT1Zp8PpxjbD8u155mhZXLO0I8Vz4PDNkrTC6fYFCe4
Qw2uAuRD7hvBzY35F82VEIDz2qe7UNBWdNMACsRanbWNDZnvXcTGRr3eD0It4wkx
2chhj1Hfx3ZNQ6O4v0wcucU38EWVdOI7kyoSbV2errKDmwDXzPUsmCMLRxYkpxJK
Nf07SmQci8PcpMj5BGPBV2tFBTjvQl9b47A/eI8mq+va34tJU5zukm8e1h+SsqVw
G7OzsXXVYQ3gSndDKoRpJueGgpz5g+Op0P55+fIzxzxWiTIPerkgbQCOoiXmMqOm
ygwfV5T0mHZKW5aybcFp1f9zKQZUn7PSX9IqsnPjlgN5HRSsX0Vb1E/8oTLilKxC
LM2TG7NUCM6FMvQ2G9jMvl7Dc4RnHRgADa6fbu+Lhk7aXsE5KfwO4maaZea0AvH2
ue4zp1a1PETFDTPOGfLvSjCGwz9JR56S1XF/KEvBDEh1224XqQGFhjkz9m6Em991
pClSuiQsssHgPEHvAmUBe0uAeyR1wq5h1qOj6rxPpIIjtIFgVk4v+LULRSzAsyya
wIbz2yixuy4eZwFJns/xFTNMuVg5Rh72fZEIBfGN0RgTDuIcWxm9szh1cFT9y6O3
dP5CPEOPlSbZboqJGT0HN4feyyaXRDouSPv4Tv3TU86MkszrayOy2JbkCOhSYq5/
8mHqnEq41/gT698sQDvFDMOj0Y4P2+kkq/d0ak3cX6rlMMx7ajpYnaHs7i6ZR3ZT
3m5EQ1uFtwCYayGmbfDiJxO5BuZKzBWcQRVdH7XHl3HgzO/Si3c6zhbQC/IVzIg3
1aB2NmrAVuoxcvXoNNkiodmpgM+rwKouiQMi5ryNMfqmXdR6+i0HZF7A126ajqAb
dBC4ua5LNAWrLd5aJ3Tg9hR3wLjt+fG+NiuU1Gjf8/qL9Dq9KcMJAHzIt/nogc4k
/llIVtUests9Tk4G7Yb2B+xvRhA3muE+rw1jm4e0caAvRXkVDOFXMWxwULFuBfq3
oAR0oNZOBTdj1sh2xBLVQwtZqpQPb1oHud8Kk3kn5BIQeHsh8dtO7pKUPj5l3uSG
cPiRJa9Y3s4M/Dj0d5+Z8KyW4kmd0AVtWJSLGm8BIu88zTyj2vLUSWQ/T2PdSX1h
RtF0mcQLtrYCRKqpkuGra0Cnq6mjTA2TFyVKFtIVBXow3Qt0SMu2iAkOEmaQKoRN
Yqei4pOFoHb2PJZJ0n0tlquUliDK4PMCTGOvTsjhTd9xeBO75ozRiUhVCPXk4FW0
boB4rp0a+0y4+PiY61beq1y4VOS6AdiKtbZt6vIpwqUn/XEFMKJaPYuj4t3jftBk
i3g9gD7bOg654qvRGcv9TtFJRBgA06bW8MxS1BW/1mZmZDCdRtJc2mDZWYvNVFkX
NWishs28wFGBMhDvryGXLYe4XZI+RTD2xzp857Mrd9OmXofT6IsNZlDM48auzcn1
l03PmreUyz3h54rZQJGItrU+ILzHKv6wu/eHXInXUgKD4BP7TiEGsRYmpoya41Uz
Ay8viH9FlTyemyWLmg3FKur7o0bW+ktFlIEuhqhx268fpNU3aYh+E8OJLE9lDHyv
rcU9Su7sVVoCIZ6dnGDyAHimY0WO9peysgz8COkGgjUja8d7KEt0E7N/KDMCP+YI
wcKrNACyR9gPcPNU4HUdKt48ZaVqfxbYhNO3JmotB4gx0KX5hagd3V1/b+UYwWW3
xaLLsKBVpd+LHFITHER4Y5vPStdN24L8AuyZlta0f7mU41UzKNfNvn+eegTdTZVG
S+YFjG+88+oM+zSmmEOVegVGsXmUQL6NgtQPF/7y2o36zO/MG9Vsn3YpYLdWfXVS
ZEmLwsKoiy1ulqz9M58/tnAL1PF4WPMluGuKnfeB+KjzNBn6KGxnXYeX8dVoU/S5
bTgDJ/kpQRQ3O9hcdSwqRyqJ7qtpiCO4N8yHAjJpuJ/5wLl3KxiPEWwAlWrS1Jg4
Rr3l6YRmLLt7RxiiJLJq8T/YVdOLZUzkYTQ+OPIoW+2PWaVfIvKLw1GRC3LXHS7C
NjwakJ8nFfWuvdguWfkGZRdkKxVZVJEA/ucbAXxijdER4L8MWuRZBUJ+/XIvvD/o
z//+adZxqUDpA/gytNftUBu/zJPpAKNgChO2+avTfxsCNSjN6akbsuseiuF0RVhu
FRyALqazRqV+zdjG6DYEaIg3fy3A2kREqFdA9yfn0O+dTUc/jIhe3A67OYTskZjr
L+nmvnrqYBvdguoHlcgJbGzINCHs4EFF0xqLVXTHdOK9B7r4HGwW8Bt9v640oVuu
oCXcQHpSk9U1ukaclaGqPHgO+hFfd/5AcC2u1NVWAPWAN3plgEEHDuD48AjQNXvj
GQYrJitn5Q65i3SXrGv+sJ/pKMlVQe9acURxAIdF+W14YsEfSS2NayZT3Ch6hhxw
7YiMn7fLtJEh0tQmeOyJ/q5vFS5McwpK3xuO7jOuMpmFff7kE8rIiK62ZQOSArcC
jWLlDU2FfVrC1/JlW9Uu2GSfKsXAE32p2784cUyAeumBdba1ZRu5ZHzsNeSz5YD1
XDM1wLbBFjpMmXBniW31h+eqKAnoEECEtu0TwJs8XK6TaWCcmLq1PwSeK19KqFl/
k9bwWEWzwXJE1wnzYdE7ADj1PMCxG3SsguCxbFsTh1JktHGulWBkvnBi1Fgvhn2f
JzRgSBY0s6OjJUp31GF7Qv3wBgTME6NgoBg8zNRp2u06GfRHPABIU4oduuYAGQUD
jQch0u5EjgusjhWSC9tz3BICgAvNUmjaQrk/ItCMGf9VTJaVwABQ7eAbXoZHyDLC
PEPRw9Mq4GjPgyimjBsBulzDkgVqHZzgH75mXUiXQzzfpkA0o7RajTohF3Vv5PQJ
q/AcWCNavGGywapMRcQNW948XToSahKpcguPwCBT8SJNb65lxit9CqKU/TghSDj/
CznFSSl+HqFPzMBJ0byyTVZprjoYl46/UbOX7FQE7+ozhk5A2TD4B9RUTPzSxUJ2
RaXUA8LYIWDyZVw9jG3bCBUiOnSK3oB6Swuc11kycy7zcbKCVfAcWzTwE7sqefze
bAhSTnSSwPKEpYJoe6se/YaQjDbY5C6i1KQBc+G/d6yAdWZSrN23QBh7GL4EWJWK
gMfN0T4FQaRtI+Ada1eUYW8MkHTSZa+IyR4AtBWL9Q6vFQUsBzVam7k9Id6tsfsq
QCTfRO9LkbcfVejTQLNDF6eVI/wpn1aT1QkcBGOMQWbGegUV3qZk3G9Qsqh0jLRj
u4lC4KiNCRplf2/6ZL6gnp5MA+UelO19+xiW0k9TeapMcahw+z0UckDQ7JEeN3r2
tJgreMWPlUzGb6ggj5lnfwqK5KCgg17uO2woBO7X8ddlXQ90rteikGZLlpxI9YD7
ILKFwQjqLhtQeLY5Ec/jziJqUUpDPt1s25ZZbI2A4gKrAHvswttYKVa/w+SqOBbh
S1ZLzJ81Jn5ZzRArpkH24jXd+YtuO3GCE3hPw0+0AjWZ9dKf26+E1GHxMYoEmkgV
Qf5AzMLEvznBnptMusHkYQyjrCniWbNDubi8+O5HpOQxJbksvjrqA4olpsYiCGBh
kheHodhagJ0PqdRryQxurZj0+k3DuAOL5pXIazJzkXes1gBHKfmKXRH/bqEscRsv
5KgHd0CyQad2iWpfYKW7xfI6K394wApz1X1Au4Vy0AwqC1fpJctmBOmI4QTIIz7c
rmdp8CuGvrqyJS3o/ViLHJh78qfPnknXMOmMaasQ5qjbeUb6ncx//YtoF/KxE045
IADdM4Fdhjs1yDBHetYpbHYJx+nSNaUPaIm8FHAfJdRgO7YSZV6XIQT99B4t5QZ3
3XgEC9upIPtzAOmLduBh34TJH5U0FqN/b7Nagcz3oySFOIQBhYR8R7b2tKZoqH1k
RUifGt2xTZq1xSzfpeh59u8HRr8c/Ul4eXrLLETD71f5uuHPU3FRDPaG++HnQ62+
meYv77bppbtqu6JrF2u9YVE1wXRwZuJzWbLarqKUoDHMota1PDovqCmt05AKsQSj
hkO4zGLnUMysvopQqh4E2XDcPEfY/sF59SoK9CxZRfmDFcu1wUf0kaE/wJlxCWEH
tD+AZYIMXhLOhKTxLo09YBtjhi0CpN+VUmBERJGe1TAAOXb4E8QxY1BAqPVV0ev1
rcG6ydRIB87LtEz1mD4f9SvG4QP/Rhz0wcMKaJOT91s7VGUgI87VSz8JQVtB4SKN
MTT7q7CaDUP7aUBNOOOiOtnheGI21i9q8QR9ECSs04wL367HBbnmU4H1X2q5/LK0
q/D5jME67cTYTeej4GEPvlPCj57IX2iJjrN9QgYeDIr1fYZU1HTiwyZkMXGk8OWd
oULH88UVlotT46QTISEBGmltUgXUsxrLxlLad9hEGLt6qWCDoDx4tj3I7+imxpq4
mo7dQAZ5FqO869D0c421A6/zEkpbK8OknXGF66lmEOHMVTMgLrCbr8iQ00P+qvLf
ZC4ypqIjJ9OfTMMWVS2h2AIDwUCvLkfHYR2pSKtAogzHVoSpRhJTWLCbPt//Mj8e
x8GaEq8DsOF5qOlqAUPWJgwIjE3hIFC+lLnAkNZawM7TVuftWJ233f04Xon5D7ue
zVuTLOvA9ksXY0+ugn3lDrSKVxDXEA7zzI0ew6QlpqM3rpTCS8M5aFriN573qn73
stp34Dcjcc5sFkpg4/kYW0rbHCpIrNg/s2z0V9l2r5bvKkAQ8+7wNhA1HhNfNbK3
Hk8eEOyFi0ngAU96OwvK9PVPdwz2v9CG2PNZIn9grwtsQiakWLxL9uID+d0y0r9t
iVpdGDLCOR6CuHxfm3rqMCFF/m7Nd/c8fXNVEhxEaltX/4u7VNW80gmYaKjqh7h9
YOxYzhnaNeQiMucXdVnTWHDn04c5eD3llIGFRqhnBXwGR57fGRXxoiM+bfIDPxBq
MEzv+DfQdRceKHyQGCHjfdBfj0gfikEi7snL4tCTVsV3rE0ajqIWSzvqIdO9l1XW
Xvmah9QaI0JIkmDw/s8H5NuAL2YIQctxsbuGdCtObs5GOH0VJ3bGU7XtUuTqlmR3
wvEO3bNRtYqSqg9M4ZgEaXqdM9UaOMSDqdRei1weYMCGNo6X+QWgsnBTwHmHj7+o
/X+T9jieV+a7HI7RCCsWKtw6Luj9lmboKJAoDv1cF5tgK9e7oPeBPVOGsUL/ufr8
K6bErGHJhncPf+PO6Rcjxj/lKQOFcmIf5Nx/VzUViISL7xKq7579nUEYVbR24LHI
aYop+p419K/7lL7rlEyrhNsdFQ6p41/Wvl5mbr2uOtybKr42q335yhK9S6U44zOo
/1EH5Fw4+Gw2D4aIY+lEI0acjEMwKfKAMvc9+8EIA4DTJBEhWrLgQUsD7nsDcidj
qDeTqEaxnCy3exC5aLtBpiprtNqno7wrbTsCxJ1jHvqKQPFmok1p/jixyw+Qe9kL
YSG15SejvG983hdiS27Wl6GeQL5HPndLdvr761SNWm1n9DyOQ2To5oiG7cqF+gM/
1okce49j1Lx63EcSR1GtKQFWNjES05DbywtmkBVFXxJ2anXiXP2iyLe3gZMVA4Ro
eKbq6Ssg5bdJZtf4RgXt2RwPkFGh4JIVyM5hiO8XqDa92SWA3XEZHW+ct0LPorEP
5pbwcrphuDrkHXyzQc/wKwLFd8EN7UDNs9ccDvWnqaPh164/zl6qH4xMINV+/oep
MliEBn1kZ2t9GQcHEyPl0qjJ78cUFM6QkDvGhSmwzYZAxWI3wrsKklcXBcFs0Wva
ZOcXwJWVcmV4VQxwO+0BKX8ZQwQ/46FVBYW4t8u3rmfhWehCV+2RXAn15UilZvEg
S9W+vWAvlnCfhxTWFl64jCjb9n6E/++g6sEwaD89ACgjAEc8lxSEd6Vf+Bva0zQw
dOCfPYafFEOoKlgyNWWLsRJhpSCTQp5iLcgB//1ZmJOgyVLl/KDI0xAipnxefBjg
T9boLe840OLzjlYH3+65lY9x20zXIQriZg+RdaUOGHplDVg0u8YV86TSXrinVy48
51ThXp0qzvgzLU4qtpe59e4mi5/A/53XjtMI+YT127K2nk0YoSXpCr1T/A6x2Aan
6RpRDf7O2eJjuPComZPEQKLUlrEB+JeFdzgh0unoqoBDkc7Km3sAjJ4bDrpHGc9K
wyrqyRWCAj2SD9GhwlIsVDxPaMSpU5H7KzZtCHX+SFRmdoazbw55wKLovh1j2Nv2
nR7ZJFV5+aCdrv3VXRyk4tw/DXURlS6+Nq/pd8I41O46Z1aJ3BmNgfDV4bhD6Esd
xT13v4Bm6V0e8hProO6GwGORs3z1hVxxR5+uOxslF5f7rOWKaLPGB+ll+aZQuIp+
uRlwdHpJy2yq78kXA5QCs9+w7i1+A65qsC4q4OrsSwus2wpvHAxpu3igUV760Vbg
uHGbIOf6W+bUit5es1vHADGYu+HUTPP8xaSDfcIMIn2djr+EfNGXtnNFpYjKweP/
cWE7xt8lmoAXJ2i0ldWHTKmHeZag8efZr8b4ZxNCcCOUaCnuIl0K6KYlOUQcJMDs
LiKjUq+S7WGvgE7TRqAHT4scrAoxCobfsALxGZncsA5f1nwwrk8jMMTaYstpSiXb
Cmzupe1d3EHADITUzzaef3SBAWKnT04yq34LVRiXDSrpzWbL4urfla7/Ba7wA38k
AlI3RQm78I9zApIrH/2hoMTWTDtUNBo7VcICusS0d0zcCN48cOsHkNZHwelk059d
GQw4jtUxhzslVtRZKkKGBqgJHwdIWSmeYHBWvmcNCmY4abo8ybfAVXcBEanuHTla
Ixe/9I2Eei6xPINpP9zXJwfa7AdliSAXdQfpiwVInxkqH7vbVRyWp0UBFdhdeDhQ
IVm4kLyp0u3PuTYolnFYQAI2lLxbsEov1z7vmvJglrJ2lqZMY5Zxej1bpCQb2xs7
VUiJ4GGrtrWzXPIJcnz8cz9dh+595BLuB8c7FULsXEdPhIRlkc4JDtVW8wfloDuC
XJjYNQiz+v2HS/GO2SJclIGpApbFObMJvIrWNrSbuMtxhqgHKJMMWHpDrE5WIPpl
JCuzO4XKK2RfWvCyEbEDKcLZm+J6GQis207Q8AxroMjZX9q45lglKCTitcULpxJk
/0QcBQbjrBCUKA+J3icTiEZe/D9gIzvbXHamE249rydq9KxlkLu5hw+Np866dBlg
KRuSIO36yICscavdMd+NwGq+XGbV/CLQmYdDXPIroTzrzhz9jljtsIh8W2Dea51p
GfgVE03ZpypnHuAY6ubzOvxY2LNDxcKaR+zF/XV77CMiD5wkraCG5hhLY+LeYWgy
xXD0ljuRBT3Wp3rSGOJjfw7qD7p9f6ai+j71RPsyUirD1WnPG3gLskHHdDlTDr1X
0pUS9NwaPW0RNfj1zZzxDp0shcHdLPt5GI5nHCKzvGLMxZXnR+sbWXVE5b2ajuOp
pyJMHSXF3mScE/CtMqqN6n7k7g+g4FgR1vOu6TjlYWO86iZUex07uSG1x6iMUOpa
VAjADfprbS1+bMX5x4AU+qcq+TRIc9B63XjwGM3Tu/ji8v7mopAACOX1EKee9sga
oBtOIli9y61bLcSDnpdaYre/1AOLHox8YP5qlPsUbkne5nV1++iq+/nJdcf0EBQj
iOkMM2UbR/nG7mrxSmThs3gwtEib7cqyIEmr3MpmkL96ZuXJDPoVcVg+UO8w2mbX
6nYm3eo75aVSIbN/Yi2/LPXx4wxOyYDTNU3ZKDxb1W6D+JHy7A4aLGeh6iDq8Xco
361/osROdYXOK4VKCnMiI+2fLIzUd30sWn97jM/NUwWBwz6jqVzhA/5MqNYvNV39
0cMNOgITjHTL4QRr3QzXN1pEY1jHw81x6EyqjGf7HC4/WhfMEd/6FmUTUW31ZQRj
0Qd1q5O6oQJD4g0/rdDjo3X3ruzTYloVxL/irlv6GyevaPWCV8b0iErfOQNz/Bcf
9EK0uFpw0mHK9Zw1wWVk6C1UAmhu0YfHJ2LRcN78WM7qfpMdQG+PLmK5BS+yWZ42
3LirvxvFGoSkkicde56r570IZxGH8EU9R3tO8bov+2PKPdOnDXLvHZy7VYJjWE9h
VnlsVWgi1AvKE9oQZw49NOaleUeUgwNkQdM/e8xJedkd1lsql70Vb2H9OYN3Vqr7
F/E//gOee2TOhie1RLPFMF5WjJF3mlg0L3psE/TtSAPiCbByo7y5sArr5MjrCR5Q
ku+uOHLdIa7RLHZCC7aAFBWYNqz20yp3kKMA/6S+muZ2Va9SPatv8+x+R7If3aOd
x50fHvLovtZpeXNoRDWmXxuVXXlrlrF8N+3jsnZ4lxSRyOPVmSAm0XGTz25Csy4h
v6c1quJF1oyPOvRCuAnz06nVLFtz73KvDqRAA8Pqj9S0xoVQYglBfpn3DVSjIHc4
9xrwxe1q+FPF4hDgiRtoMOx6ds99AH0VdaLPboUno8wMspaGQkIAy3hFIvzW4929
wceUYfGnCoLY8B8zKHvYUWBeayflPm5q2vX+TC9KWQ5qkGis7oZPdMIonc5ln6gX
dJzlIm6T3bzQuoDUIPkALMZUf6nPRbitcCrAVG/FW5Nef7YKKwdkAbuWLyoRxsrx
j4SXjWiy9Hs2sq8PNpbmFWKelp+V+XMtPsVNXZQ3UALn5EnExjwbWnPr7Jr96BcL
YSBt08aHmTKY6Gp7sEX8t2w+AJnaCRWSyf7mrSOk1MX6fFsaXXUfWXDO5h1coJr+
P5SMgTxcfaoihZfXs7FQDcPhM/rFpG2KaXfsjF5eERbSoj4r+670ZUEhCof4nui5
RL/HJYpRh4NbnDFNJkdV/kA4VSbNWPnocOygp9zKwqMP+u/VNhWbQ7ko/egjcJQh
aavqEZyK3BN7S21CNZhgsj31y4+saYch7nW7iDrHiYuR6q2RJxhURyOeBoz3FMqg
ukb+Bcg5zXy2STIwiQTYss4APg1wnC7oVpVnAO+bzP9uNn7eloe/HeJhBanKTa6a
NJ4l09ed+/M4OAHxkStHmR8bpznqktsdxtINDbnfp/HBvvyQEeyLpT4+NrS2ZmfT
WDN42I523Yn2okzE27kt+ol6q7M8+gi0MbaMr5HXKv9G/TzIFIAfhtw4HG/5ER8u
GD8bngcJS8Tz8oaLX95SMmwsidPhqJyNYx6XT5Jyx6ZP1XRvzUF8icTA4elTw7gi
BqbMKye9bfc9sCSOMetJ17S0uTgJL8CetZmIdsn3fHgCwwImGSzWnbRw9aj4n5XV
oWgVgNEP/xL5cnHWDbv9r2SPqUz2DoplYB5X1jyPmE9Xcc5t9Eerss63RjtK4sVU
GbAAzz5V8voNG6a5UTe51Apk5/dAZxRBnmU25NRgIevKH6yxIErp8HXGykBYW2Dr
jvc9RJpEHcWKHfSnCSHJEOlkdR5a5Ffp3oogEizox9YwP/oeTU7gpS0iFiVgBely
7mlooee/2qkbrJY+kh4H4FaD3ti5g2Psoz1H8aVTusv5I62M+2OmV1f7mGkxP+Ch
Q5hQcuaQ7VWCMMq3KGl2hi9NGX4uJR/vx//HAmcF3rlBlz8QKjnSW8pIGRqwo0Fb
Wj+x1D7jC2wCa8XbjtAjpzxLO1tULrkeLhmS7rfDfOCC6cP+QRNTfQmN8E5Qxa3c
txWEu2XdglYe3JvCNWh8RO969ufla5pT84Cw4UpLVw7VQzGaFzCmOOjqRe9AGGd1
eHX344q7AHmxDq5PFu69zN/cF3fRGe3wYXS9r1BjPNFbXG2m4fVt45e1GO6kSJlC
CVZJ2v93ZCHh57SvvLlmb9SfogiPPGtMpCyHI6y7V/LKJlVntgNKoccd5AXfG1ok
A9srDYgn4V15HuA12LAnTQJ4Auk3Dha3Jtp1a7EMYXx8nuVmT+y8FCSIZvWIOx1X
7h11DGDg95uRSkCbBStvea5CYPFjSjAeCuaorOCYJh6OQWtfUf542YTopWQZ0pS7
KbbxtIWQb54EPI59XGPauLQPH+zeSyqfCsRrl2uvjgDZj5okt4nOup7FkSj1DudD
jNWTBn/fTiEFzenKyTllpZ7bJBMy2xRq5RAs9SY1F5wvdguZKT1Uq//YZMXyJGJv
AMdCjogjsABmwe2iGtqB5iJCyZnGqn9T7Kc074okqRHZBoPg1dM93ifN2ZNuWzz0
QlNvPMy2N723W9fc4xPTBPABjnvMVTPjbf7Q0x4Q3FNNdHtbaWnB/Sq6m00Pt3wn
omFtKmSKANOu6WFNtDNsOyvvtMlvwZC+36/2CaAIXwfEQOD9Yno+WYvpfupP2P/W
b9cbuEI5V4/1bQ6VUu8rUjywWKoSlgSm5gMOfYEckczKa/oaWvCwkKHDQx4yneRf
tMb3nNUZ+D+pQ+SsVscLtI9OSxpTWg1DtAh9ownL2TKz8KdIUaGxucIIyEH2rL1i
+Zi7kPTt9vYSCT0evbNvVG35I96WnTsnXZEQ00Okc12ptav4eu3UyCbjHAinx4wz
SjO+Wf7hADiSZPlWCi0aDQMiFYKqh/jhrmAA4PIV4wZP6osTYmZ9qCbsl/3mDIXF
qVaHUcSrWEN3m/KcjY2y6qNwC1kkPTmBhx+Q6MeUUE+Ho6gpobA8RBTtF+L52vPq
CivDlzZQc7ZyuuTw53WI6bM7mt4hckNQ2Vnq/qulVC1Ir1loJ6pFvJ5l3JVAY59x
S1TGEVZffbLnumgQfPe7yamov4PSCIBtmbzWdsDVfBgL4vY4KaRPE2KZAsqGnu4O
emDv01iAzAjIQrVKTWwFsQkC712gLmC98st8u/1jdZKbYoYOU4XBza2qBMPsehNs
OCRHCqhkVB7nEl00zEYjwTp5ned7BHi2dRBSll3hOcBXGxvAxbVTpEO8zlN54xvZ
JxHwsS1PILRtRFlGw9hCMpRz7Q1eaZhuVmQlCllMVD5Wvh1vOavCWN3LAHSCK+SZ
Ttie83+mYi6ZnG6yECr5S4lLUFc1E5MgyJKeO1ZI+Etu+xuqEhE/DKBsXKO1X0pe
3S5ghqs5rcmVdDrz2HYan3S3+EverVAMsB/Zzj1lXY6ezhWCLSH37PMf4F124zo9
BrRI20EmP8/JfHovPqJUHUhNfxtHcTSxGqVFP0qri3oWKDuk/oZJNHl3zHjYPdti
s/SMWs2F0+FF3YsYh/GpLz/onloO9nMxeGsvMBUfraDxCWkSWZSB22KTzREAKBzj
BA1g1CYFFkMe62FoSBEB4q04FRB6/RymkeiALK2i0rvN5fMpytTRghTlaRcSoWck
+EqTVjsTWOwl0EYe4CeVxaFwZNQnqn7xHvN7VtDnb28mTPb3CIm9hLrl/aWEr3+t
mVhpvSnDhLUh784rwmtwbudclo3Vl/thk3e69iYv81Srfhe4bMfQsrH2h7eeqfF3
exUWp7d/T1pI1wZQYHPXht9JDjH7Xo9cRGNf+n0XU7Icg65mHSlqjwei5FnNSskv
2V2um8N7CLeJHlg8MLrqq+TYk5/NR5MkoFKa+X2n9fZoe37F7otMHJBq3ypxkDuq
o11fWtbKSn0swes6653BsfHiuEqATE4Jxs8wKxFLuSH4QpXIS8ktUafiTbaMgLJ2
oujj00PG7Ryr1pswAFWsC+f3+KGf/VNi0V+y9EzbVat5PxffMj9pYL4vcg0LymUp
sQKTZQV4QJcNr+SMcOFQVdoM9+MTaJO26nSJ+9IdNBkKhVMUf/1NDjYMaBknsl+S
A6JmbcvFcDZnRHeiwXAvg4RDAxi8s7za9hBuBbkjQHSGN+RA2a2OzovbX75TDMHV
T5CNlGO7zau74tSm0giL18xT/mvP3OwR633IV+UIq/HhU5aAZKyVPks4KmKLsbUq
Kt6lDoUTGmq12k/RHCw3XizoiKkgCSIYAkrcewHnNSPqRq2Rbg12UQoRrNpYmWAa
+qnje23H7IC+9+iY7/ot4LE1KUzH9hk3FhddBYZgIRxvYLKm5BcMYY35JzQ9cDRg
qOcrbjVlOtHc++JM7Xi/LbwZMDDZWg7Qu0eYlNZ8AlW0hIPrexkvWY/cyMxpKUxI
8zGtatH9jsdYA46Db1kbHVXFOqHzfGPCl316qRe/UHyf4MAfr9Tixwb9nliZjvSu
QvazuPrczCkhjDX3ox1kwLYfJA3f8Byy7X84Ew50dp9f9Z7BQKS1Rug/vMECQ2M0
U2I8rWAn3hxD+O4G4g2Jq0PKtrjoUC0ZKckB2ml69hx4rwoGXl4l5hibpC20vYMz
Eqs3RUgtbfNoGGivESrDwo4f7TQntATkiFrQ5woBlQo8Bl/46jbM1fx1VlSrUZZc
DWBybq729nkC4Y7cPk2fw8197AuyNEVZKpWqUonm5LXqjIZPfTOpT+/zEpNkq9eq
5yE7wVMluOs7Rc/8uyNsG4bxylJ5ABPIBFULnZ2+A/ipms3Pml76mo2j2WmExMLw
lh/xYiJ3UF2l+7+oOTKBzdDm3NxrJBvgLdDi1OqUsNG5V/J80Na0Oqdnsj1fXFJT
VCipyOhWvk5J7aS/w4ZBolsDpFY1cFhOtzFco7x+Yrf5oJBAeg1B2YTPxCEWgox+
fLt4jQKXBdztaQ+7HB467E6OyNZhUO1TTx+/D6VAwohIDhClEz9p9oqdP58PetL/
2CUcjiEkXSBiUr7iZfwJBRF4o5km2h6EDkbkoRPvNjg6YTl2nTKNSkZDivQkv/7h
5PpBnKx1wgCTiLdqp2pOLHvJd7/Fr+AK+AyzA6rqBHc0CUDv0kb+Uru7IVPTEsBL
7vbdiR5U/Fyu7etVTQZP+nO8hmSiKER55lPA+828Yc0Q5YtGOpslQB7wilQHeHf9
hCZL3ItVjgK7rKh3CxQ+9mjc0QjlGTzCh4Q963NYwx6wGKaCo93VsJtAlroD21C9
TBZcUxddS49zJ5C6phZglDhUA5eyeEWwVwkBoizMPBTFADVugp94iethgVXMfHD9
C7dqNwIbu9lR+PxXTgW+QODuwoS1tD/4eHplrm+wfyzGtcL3tEsEnMqolnbSxsWU
dxkWNgrxe3F+DOBni7+Xm6t4tkDFvD363OoWRLyqLx2h/EPRbJhAet3xjca40yFP
PKIPV807jOAeMSKC1zYgXsRCWhIHkcUHMkbnNKifZ3mJu8XS1uy0zPwPUBarp0w6
S7+UYf539OC94n4FzatSy+b8EPM0iw7BK6AEPte2cvCTTo/1sx4boNDVtSNHvUkO
6G28pXMODQoDcj8EAOsW2zLYiGFGbiC3dAQXcvF5sc8pruqe/d5qXN4E7QrRN44z
l4cIT0Qxw7MkHXoE8rOUOVhhresJHFbKMdzwqTR0SL/M2hkp64hUgxCIG7je59Ec
OI9wv8oGKIrgNdPK9NQoAXxcUzMA6+XBq+5ttI89OPkMqutgDj7u9vKB7f/B7+p5
uElgRyIudcYXDVkr+GyBlEGceMpCRLyQPIsvuPKLMRG2EXDZRlkA/VD+uvQrrmDz
jXv7Sz14R5spDxWsMPHe8Fha4lrbJgGjRpm1ADkNhSuefW4rhfaTKRM37VBHdBfM
hrJn/VrPYsGcYxtFKwGVISbl19BhWBDFZKfYzAALd/5whAlKkQVCEOnCQ4pRKFqY
JA/w5jYBcUcBk9e5ZEdhyhOgUgvjBQj8m2dvVFJ+MF7lhopM2WK41hECuPWfr4ny
ETiMjO9q2Sgy0x17cFnLurAz1eyOK9UsuSSPo6Y399xyRKS8rnzQHaEx5OwEX8Mc
oMJTLulesVLrv/S7d0q7eJbg3ai2MxOJ2FGvXa66NP+Ti0mICF5zdN99z/N4FkqJ
EJXNl9OY3HWDvow+/lqQKS3ryCoamzpIGEWJhTB1pKtDiiGqPQG9bUijOCJQm4Y7
b3UPE1rMY3YI24HpL3+aCBvrGjJsrcE+0DFE4yAIqP6atg7fD+E+ZSD3rk+vDRQn
UkY67lRtqpr76MBTJd6aQKTS/JIsmo58gFKvF2kybMMbHLt/CSyFnkXXaoKJQ3A1
3RkSAsAY4M26csWQ47QRRQVKYi6Btz7Tnu5OKFs/w28IwblfLAn3hBvcDYurRbuV
XKrKphGD7Yh10nhjOmcF5hvrP4bgNOSunbltBBBkTBHzg4vMyU48MuKEzPPikvzv
K0XXu1cBPNQsdC6h8PQevcMecm798TuYMqqzRC4OigFGfZV/t6LAlJNgW+LRedSz
IcCY/lkkrEJ43m054ebZWtcZtLy8jVVuExNy7oTteflXf5VemgNRcBRkIwFgOUWf
H36rfs4Z2zb2jb9YdeTEEMdjJReWSrq2Yf4rbqb6ULihaRPggbXqxC5ZAHOYQ5Jw
KuBuAXd+yWqIh43LAxiVMgK7+SlhRNZiHQFCsF/aY6lTp/EmpK+hTazEc3LkPSrs
AZ/xApUm5yLe2BVRJRHwIp0UQ/HulTvi8lJyY4C/yZaYtTrvFv8rq/bDuteYf9q7
+DQSHHqMdMQ3TeRKuw6QWUArJcxaHov0RAQB3l9ofncPdI22ob1of7Rh3LI90S/f
KgyLCQUvKzTa2mZ94AnzEwaGR16UN9u8+31pVHZF0EWSbJEwyaLoVgS0EGMC1Yb7
6ZeFRs09SXd+G7nRptIIgYr2pxsAvdBE4R8PQHNAUrXf4uCC4xoQhnu8ivpgiFdM
ptpKWzsEkEnBkF5dJBkRhNoMPzCKjCOGazoVdgNHf0VUDcPjpRLqv4V+e2QIb5RI
i34CFgaxsDQ3fyhTpDdgMuZd1gd/q8rkd7Sk8KSRGpDTJ1fZeNgJoP27ENz5KCEX
xGa0hEP+TnP06YA1cPZ2XQ0RUZTwOAY1BC0TStuQNLKWxhiNr22si+glzpQ/r8Te
YFtPpwWP+hRCkQ+/mc6Re4rPriZjsrZ5Oi4VN0aeCV5llFIKAvncxaJ0iyeNU9mf
kViFmwJN9mdF6w9lZ1IFJvlHqoE823mVJSHHoLKDWwRRU93b6/OstCVL7/ilzLi5
FgjjCyqPNsI0l/VlxIlyMPd6+ozLVAzUJbcrDB9v+vgVPdAecukz7QSFOZbuHhR2
0NdzzMK4vWLFTFcSujicfTXlUVIJkgdoDVjXDX76SWbq/mbE0p7wF32ikujY4OHZ
hgIC8Ibtd4qcXy57cnkaqU4qpcPkWfvVUjy9f1FuHnjGHil096AjIiegMj3aNZIo
bCjW+uMjvhLCgBxC/XhGgSaD/Chym5fV2I+vt4aWWKtEcZRDpKr1y85qtGsJJT1I
cdvfAGFVB9aaMSSyQw8Xe0juykzlC2L50jpOaXNJwi7xReSG0w1Ik46UxqUe2liL
XAPdj+PkoUWsRrvPCvsXKwRiM+m4NwLLZivtRHzK8flWw4FRdIYfhUDyqwqc6roS
TCtYva8FIdTxyVZ73ooiEr0VQp/ydYW5xG4DpzdgAG0AOAbB31ONrRyvoMB2ubeZ
oenC7SaE9PGwJnKlWcAFBGkAgPed2WvKGCpji42hyMm0a3usGeYEmiz+rAakvssc
fkf8H2P71RbEJCVB2yEfyToPEH0duAVZmCLfy/ux8IjRX9I6/3NXf1tiSaCqkwId
a6ju1yJkIlqhunXEXlJXkBmoLKcqxedxh+qOa37BPyOHMCrb4eGCOEw4fbxY840Z
aZOKR8j9+JSCoumPn6rA9vcYk0p113YcNt0IoLxRPD1lphEOe+rFHts/WkuY/dMy
wueaQFVN6X3ehyZDS6IgK1b5UzbinPcUTYYgvnCGezEs54GBwo3ZyLWtyi47Ac29
sX6q2SKU3T83o/pRJGOE8urkFms4Tuwc3qI6l02fTL/0a0/teq6UXZkzTvi/496G
1en6Y1X5BW6156oEv6oZZwImerfn6iyuV3AGYqQmHepChn3w34dtEN7P0yqmPhUl
WppjFeIHLqF2r9amDAqtiXEVMIYCWbL/dJozCjlGbrsLXSmLGXEkkanjwMCMHMx2
8K7s+HrBKn+N7CgX3gXqNjfhrx+hbgqrqwiL39PayM56nG5RjxxKUZdbeRKcjxKo
+d6Zd5O6HSNTmbU3BhOosbmJq02dDH6hRZBGBvulEk5j+LlbTwFHJ+wTa3frPOy4
NU0lKbU8z+8yz83lhgN+ziXF/CGKL/+6T5x3z9AU5kxjirHzX57p8EiM3VThaDBw
LHC0hYV30cKAy/Pz//pcfoWjPSLWpe+EGo800+cyN4HyGGnX7qxVwSFI6MRTU3Nw
71xZvIf8sFZVzjXZXCqQJyxSYL6kNChoIrlgYu3vLo4VBW2AOYA55U1EQovEayCx
y3Wlio/jfFQkGBPqhnPWGe7G6MZm8JpP1gkisv/AMbCHxsCAviEhMpqh+EfwtqaQ
BmZ1mbOqz+XrE17NNEErQqm4r5gRsBRlmAFN8XdKdNg8UMz5lJOCY7/aYWcLUTqb
xLdBTI+PWDWSC0wA/Hj+wBsc0jHdyfx61MrHMgwDcsoKEidixcgKa6AZqsuy6UM+
cgHq+rHu7owvs/9fxstGrjczRsEHKprNM5rGVK/DPyMYTtyB5MkdPrUEURMrFBos
HuMTpC6SerLdlzYcrLwC/DgxjA9Qnd6djtf/Gy9b64JY1Zy7wZnvWyX+x4BIf/SC
/YiUiKXQKZDUMR1wgrFyd3VNGdnnTOWZuOqwx8ol3htYKorZpCUAXW4A9VJQdson
UWf8AeJcCUnhz62l2jlR9LgvnWRcuyG6QTE0JX/BzVmmoVrdwWmqvhr85PYylAwR
Pc+g3Npw6/0+NzkroGJmjra5wwDHEaCT2CsaRxn9CQ7gaXv7NrGgHrxTSMf1N+mZ
zOrv5lkRBsJHV+ZgvpZCo0loIPREBNaWQ6gMW4cNgEnJrCCaX+z6J3+I1l6fwt3O
2gL2h+s9J6McZzBp6HL3Qbk0zIWi6alAAzLtnLIp+Pz0MzGJCOTZnFGxvOmq1Ql7
etiQkgrpQzPUBXtcmkMyVVgqVIWbfbOp9xL+e84kqWz0IEVnqTSBnmOmQyMzA7sL
oBbApuZvahoysjdMSN0EYjna+IoAzr0YAl0NMvbFL8LpE15wu3FUpn1QJ5bS8mYg
DiO0JY3KnTulwlz/QtXosjM/CxfZLo2aBuJ2zcJQ+Ns2TU3+pj0K/PlZRdK1n+qg
yOgGMJW0suGttCuHe48VGm/J1EOo4NbEdQZllRqk/OboTlcDlk/lcr8o0GMpLhcY
YfkpNIk+NzZByupPQ6waaGqYWSxEJs2jCmM1NQA8sMuTh3hSkDvT3lkxnWfvJYdj
8F4W9ijtoQf8d3yp/iaZpIN4U6z533fos995mmZgqimB5hw1HGf1xc9KJ60zb4av
XVmOiusxX/YFG2l0Hbg5Za4tHWKDFaaA8iCO2usak75NFco45ZjihB/6btWYS7oj
cB9oBs4dGy5dzJDCU9TAPXAKeykuHMjrs5qLSWWS9KK3S/Ro788UHTB3gqcUrS3T
AE7yOo2hGeMHBivK45LzO42If1yfOKrf3faPI42polfxHQaXKC/8S5xN5oU8XXvE
+DAmMFekmxgMRerRiQXlCfUIwhVlDAiJJ/3sZvS4BINTYXBkjtfMQCE55wMgIkiH
feV7uQ6YYtj7naysd9hu1nh607cjRhQsNdRoNfga1yga14P34OX2xvI4JFjB9Ebc
8K+DtmvptAOLlht7rBVQPzqE+5RCV9S7k1WA4LknAZiEKlDLhLxHTipSe8S6mY2t
YeHDIwowtgA7fZ3fW5gfwZTS7wiw7ya31BrKAzn7vrZs5MkL/8dLfh5cgWCODXXF
7K32urHnBgHhkAHIIfeAHh1nnFPjMy0qsguVFBPQs8FYxQMyi7ydj2VI/jsq1JvR
vni2ShmIP0h2lBm9bPu6U1lYH+wj9et0wdqxV0SZUqL5l16c9suWBTqIrhnJY2L4
IBSP3GsE5FAUO6pqQ9BLAKW9Gm1j8V/us6ycTkz1G9V+ye2F6Z4DaZVBIKAMKhap
IpapM/FcATYQ6v1hGRGNASvUrvXnNuCc1EHHfl4h3DP7D5f1da5f3LpytiHnoWuc
UjoYvgQZ8A4frsWaIr0CPrXlVGUNYUshmx8qhp/Znt25KEBbVGnMNblPhm5RHfGR
kivAOtMTw5Qpy/9TsYnB63hzmUuhNP1w0COIXwwFI52n1lhI7mHcvZ2cfAN+f/mL
oE6ZVhMi3P70ZIb70j3IBtdOMOsc7K3N2ST2BC8obx1HL4/knaBme7sNM+3ndbK1
15g3Vm5CDQZfLELgCel9DWySdS56kq9HQNZFOv+QYJMEO/0ZkVbUzdHNA3cte25j
l0WGgTzE7PqHLBxxALyQRwQuny55g3Vw7DngGvogV6+nBw+5ZMCne3VZ2bI+jR9o
1j67oMf8ywKJhfJDSM1fEoXhbuJ51vwn0Hs3ZudivOH03IdpJP+CK8a0btaEfiPi
Rw/jqgKUvwmbMggpuG6+9IJ7kOQ+X+b09t7OKcFciV6TmtLgdA3KYu0bbd9iXQoS
UulsEIjz/YrTUifIqLP39OHolEOBJkINIr1bBnRPDjssBZ3GmYSRS0Z2qNrG5dEJ
xgpomFsbGXUjMjugDcj3E1rQEv/8S4GT/YD5gK9Qlf5F6HQt2gC/WqrEoJOYKsjb
uKJLZ/A8mhH39beh3wO8bQ+GkcG1CMXYbGqvFjO8JoFRcBXg2eq0FTFlTyGm9xww
waN2NZale8Db87Ess5D9PUcj9TtD7uGAlW8b7sdC3QhxctJlXtHyn8U/+0Z1goCq
vm8uX3IObEMWs/3u7zyBUrSTQ9go+ASPA1QkVwKdP9dIJboHK53KnGvsyV/QBd5o
WPC5EIqEysBXDwv/fmY0FKa2TaMOSY/iLEv5T5mypcAYMqMd88s3r3Ts7p7fYEkF
nOPFEeNL2AMcPivGql/ZT8qoetciSiyzWAqcc2Tth/t0bmdUYGA7qdRTg/Qckm6U
mJ29L/LDlfqSOdwAhrs17eOAuZesyyRMAspM35kyFxQnnHjqH8wNGQ/Bv6VgPjTH
EU3yD3GZSc2354EvHOBuS4GSosBGVJAxd8HbPmPK/EBuhNS8oyDiEj0a2aFCna4n
woFgzRHFhTyxkSx/eyBw4vZAl89caxSbkwp5xDIYaQ2Vj5hIprOeON/IPM2wJYcg
pQJ2ZF7WkZGRKBWi6KPbGmUgxin89c1rkum7+Vkzo6D9htGxlc9+OTyfEnocVbP7
tjYgQp6iun9MjGih1mdiwRNZ+RXhS/SeWvBHxknoS+3MkBGc+HEdyqK92NE+xBqM
1RSHc3n+rKCBD2cGpVwhCl9YZLMkttEMgdzaRY+gvSBwmhi77orz+ApLhnFuHvRJ
OFj1PC9cEY5z58U4RYxmS9NtiN8iJoGUFgBZheTewekZ5hQ/8t9Mlk7waBTvyPhb
+IAgaJp2CHuDc6QJykeC2oQ3aWI8gD/LwGuJL/z89Wkm1PrtRcReEPtJ3thvIkUj
zIYLq7ed1wMJZnaIDSy4BPAx5vuzex2qm05Yu0H3Q86POj26JJeuWBfoyVjDcQ3u
xxsDpDDbjuDHAFB8jcc5S8EMg7tMYRKUsUV+Gap/Tk4jMKJiQif+iqE519/TMefy
VPwXjGD1IX+l4txMwKeL46KnhVqw7ryUxhLxIEurE9ePp839dFpZuXGs5AN5PJ6O
8oPSXex/avueu1Et91jtUYixj12Gn9pbP4iRGQEGlIfKnUjCSPf49cMOdldNdUja
Ze6+SyddGQxycnkO9gvpQTIGutoGc+DmG0LqkP9/8yvRTbsagMkyBarwV5Ud5psL
OTwpy/BZLPhYilFs+McItXfxKGkt7BQT1jYnrkgHi+DRCe0F7vbpi7Yos2impgul
NjqiK8yqGK8jgi5lFqO+bpl+5PFsusxYyhX3hCmqYlp84GUabm2yxr8O4bxH4EzK
xlhwliIAX9iZCddXUrq7I8NIazL1Sxh6ia7mM3aPj2JsRwXhWebXKwoHNpNw9vJE
ypA8omTAX2uNUI4SFrhE0sKsHdLdA7s37YNpomJKXa+PM7p9JT4lzI+qLQYaCIbj
p6EJNfVbaOxHKAAF/fPxonZ2BzSkjUCzcNqz85qBnjST8xLHexY6d5Mx35xLVKJY
TCQ/o8CA96qG6Wm+lJiTU7DouqZ+FLiO1jdoK1pd0Fz5qQ3lPr8hF8zMII6YbR4J
LUJODfpB7Zrhc53MKjQ3aFe1xnlWzwRZq8wLDN87DSfX0hGric1tYofC2Xx/+piK
2TuMqoVI2cEWeZ2p7k1pVB0+7OGqIRkM8JS+0ZM1i+kEzQCTFSwsYgbE7grnrYwA
2AZKZZ7pvPp/XGyKQiIzEaLGun+YYla9iwgZfSjaToc9vz4xme9sauAqqg/CflPh
K+WDoHv0QqfmBm9ayiIvPI+JyKKc3ATNhsoYKfQq7iFR25tZpsgyQ5NY8fbJpriR
aNWVdl6gmF+a9k3fbTY9T5hKNhE/BEpizZNZtDG8qf49z0sBx6oRSXyNiu3hgBw0
SVBdd6pGzvdtOWfkoKWaInSkK9CV9NAOnHGlaz/sRtvT6rUpj2RUm92kEI7f1c6l
BENvJRrOQqQ1VGrCt3p4dd1yT+WrRjLP7ELojmwu2fBW+pKveZNtwZSjadaETR8n
NMAdUiEq4M0djXD+iM4tLSxRI1n6V2qI32WxMN7MKC5m4Tn+e4NKLZS3ZQBbihz+
5OQGc9gyo0CgH7Y8SIeKeLvZir7QRlzjO1hWa7IhzQCxr+aAwKpm6TL6MR5lrxf9
v8sdfQ9PMzmbCp3EiUYnuIwT+z814kbeAjZXq6XbOuSTBeR/bkfxlpbQOGxrqypy
psZAO+2PBjHvwgL1C/nW7sCMr/irZ3/6kUxM/OLLnKJDsWfU8lG7PXdPAIamjukf
oiBS81bpvYmle8Y1n2Nk/3EvujVUa7hSJ87bX3v2mC3eICO31je1QCOSryLDbwUV
tsb7F2rIk9V3M54aa8nFF2lnzLDvR7rjYT55ZseTU4peofaZiTbyvPYWrIe4tKLO
AE29EYVzhb5XNFwrx4SGaFfmpWF2Hrm5LQmnHea0MUoMW2uvaB0TWLIxyHUZTcrZ
WwUmcjn/tWtytKITOQZYF/BIerpOm1wFgS2X1go/vXFle3hdNnrx9+8hTj3IHnjA
7RMU5EmC+AfjiME7kc+odMMvvb4RPoNn8FIqDb4wVp1G9k2FPgJc6yQ1YODb8Qf7
KrUcglrqSyktF+wnQYNzRZ+1vbi6pBVklezrrl/bTWetu36g+ekX0P4cCBi/xh+b
Bmvh3fztYbXAcWFrV23KQeLGbIayF7Xljrl2ey9jvvZE0A7Hikr3l1Z4bM3ckqZK
ivK1uoLOXDp+e0CjlJRt2L4ziojnpRflnhk+Of4uMzJ0HX3ZUidomdaf3jbIbZ+G
Uk/iMU66BadTD4ysiAVAT069Gh3xMCZiVgIX33Pq1czmzHvmfxXavh6D5Y50DKQW
/ZfmMG4ZXmyCRPBgdHvYpS0Vv9caJ1p0btyansdUa2AhD+qUbrOrtn1g9n+mljLj
RUQm8wfgCpjogTHddB+1JQ/yjLCu6t5drNZ/Epcw5GrKNtXEjK3kyy1rkztvzcrN
2ekj0JhtFyCNuCQxgxvB74mLP85JmUT9vzuK0pqwq2nHfhU+7joiVFjKXeJsrfZ0
xZyNCDC/f3TzNOleUuKo07zyGaGGE0PJroz4Nzo2EFDzzYyWcr0D2NS2s1yA+ATH
CrilubYcr01svIswEBIJzKMySU9avQC5QJ+22ugQWjIgXZvlUbTI5uRF8mlWRywq
sLjzKUv9lbaKwwNs3g8NGZW74fJ81uDmI3gfjd0fo7H29yVjvs8h3cqfeVjUUqGA
Zqb+ioJGZxD3oWu+IPB4o1sGh+2qbhiTklQB4q2d6ipjhun2KqA8PwCX5JjMqGuZ
c+V9cwnQC3GxpKYhqohHu01SSLDrdogA04uOZ20AC+3fyIdJgyIUcBLKqhhyLN+r
w0njI3StrRPRhgsgTPzGyvxXBKbUCzGDFbGFD3oy5kdhUSm2AEg72JOBOzWD6R4O
SgCp1t9Tsw4iXPgpaIAwKB7qF5EnLs5bzaYeZ1KYFw/0BFdCcxK3yB5xFG1HyfPP
5urjnIEkKKOTQNvJnCZJLuyfxj0ZPQwMuqzDQRucG0j8Qwud3DrUokc4L0KGgW7d
EZJTzqq0MOSTtShplQdqJkM97fTbpy4UlAdZ4rhhYu0UnCuwQ2wo0lNnzSPwiFOF
TZqzhn78aapzPoLrMwPgu8D2BMoHkhJQ5PFQGgP/9d4R76zDMrtQZyEg/PeFemoM
KNoytBxjZJxqMpbw1a84rQRW1Q/8+YnUu7ghumfGDhK9nZYx9XvF8STLQyvAUJsy
1D9qiRECjObE6yrBC7sPssdhJ900c8Ahn/mgjUWsvIxcBiqM6Lx/uO6qKz5Fom35
okO25PH2HWAb4mzNlhy3kHlM5Stum1cIZve5GtQjr01g0maVA7RrTUPmHQdx38nQ
u2/A7tzafEQ1VlW9yKoCcaBpg4OudNZJXfOnOE9Omh67nu5ilVCwKH90GFeE6I4L
9UzpNro4x+Hfo/VQqswzaGHQUGJgfkGnHc+JgHT2AU54pgm2u4RdNVhp6kk2WPsl
8thmcACfuBg04+UQchVmi8KoK5utPM8QM3Ammk6eSpJmBaCLimd8IId7QrgRK7Y5
P9IHZafAkW2H4umOfOM65X3X1H5Ly5jjcWip3NBSQHGIxOvjRQgQoQVUv/+Xl4dO
l8fIordQi/c5ojv/w6NuWdTXB8XNoK+L27Hc773ryvvHthvUajLIjFopWVg2KAEL
De+4ua2v5D3IV7bGC5Ip3gEbph8ZsFWEvYzqpfU9VpS+RYOI9hXYJSiMbsna8s9C
9KEq+IQ/AAmpChNVPCReIXLGE7isDaBW/lzgvor/ad7rfUhC6BF3Sy7cadJrbbY2
EkrAUYMhLDIZfWKmu2pts6ey4MXS4IzPjusvKz015ALPBmHtyU99fIu8eJx9zqys
iz3XNsoF0Vj4HiXkEXRacLEF10YMzdl9J1+zZetmhmxDpu56HrEXEE2a2WxQLTFQ
6+yKqJ4NQ+TrH1rGDxUmLk/9+YrxvN+PMOHp/aWJQ7lXeQPKvCKxJCrnPCXFkjLm
r0BUknqUcVEMYCCfijbPA6UZ1mA1u+owquaZCAoOn6fa5gOIzV7zSZmiGri7odAZ
+ZZ/aO4UrkNsFSMSuQSAAu2dDBUhcSUA48CH8fUzSf1tdaXsyMlpdes2wxBR15v9
lBAhnEcrRUEeLGD3dud7Z1MCfma6VlyB154PNx/dY/g15Vq14FfKNEgnGZZJ21cz
8ygj7RgkZM833Fsrg3RfbnH51TVePNWDxX3J6KUiijD913bhhvhJwhvbm/KY3f8i
sZC0s5DmFo74N+KXWAAGDzbyqM+Il/GMKbEtGfxzrbAUV8exXiXXrnBWWfmz7K2d
ed05uZgnKE94oPWOUUOS9sr7IgLeS3a/HHGVi+V01pSyDvNIAkAlYJzhYzZiwaCQ
5DE4mvsDUCG9sVdfkUM8CNhMt2KNTmoSb3TkXsvsHiWbgmPCM7oAlYkmwZjHWx6o
RK/cV14ftLyAlYMHdg3rHqBBzMxhqnthBbS7ttJRfsBGmbI4oWGD3SoW/ZO5A6/G
3VOVkAC/5BbsNFfF7WJeqDv3g3grRKyGKXxMPGzvQXt5KcCJK+/nWs9g6mvop+cr
DyKoRWNN4+x4tunEgf2T/2UCakGDBX0Ka78NwAGsrAIQvIdWYGc5v/Xxl6EhoAdP
yVyTcUbjPTMqxMf+ClgQ3FMWSeMc+MHj9nG9OJu8yoloaygd+yVgPYZZF7dmheJN
eKIX0O6XTZz0MOJfe++S5upuWy4osACUfNhhus1zGJ7psAs51CICEIi8kQw8Up/t
M27M2NkhNnJmVPtFKMBdETzdg1iBr4RVsxqpKROI+F1dXb5zay/tmzAb8zZ2VTbI
ahKvemB3WiSjKZJx4QmFMgcYAZpWoXx19B7TmplotObwiVnaziBYXf5X6KkbVctz
eSZYv7351biW1n3qUIkJVQP0JMYpLyecYeCQmXHd2Jw876Rib+Tz35LyCv0LsZt1
Q8+u647HfOMb/V+UrCQ6Eh0lF6vJt/2M3szVZRH/6KZ9sKIheLPa6VfLm5cdBXxm
82AwUK7GjYl2ahg2BGBm8GC5/7oFGGlbFZ8BV6c5/mW4qsWesQfVI0FJmWt5LK5p
CzeWqmmM/tByfxUHdUeMd12zBGDzjNJz4INQe1wkmz1DWiyIsSefhIdHYWij7wpe
xes7o0v+UlppY2BZpCoId3hHwJptHkfGukvhUE0vEWaqZcBmApBDWIs/I9lBrpCe
Pu338sbWiHYQbL1gs5vlsFB8BA0NiiMIWYBfhQw4rp5h9pTyNFMoFx8P9Jnez/U0
oHKwckJLI1ZRm5wYDCTz9DBw53+qSUXToWpXcOnGEwMkstyTu191NLcJyzFDWyTy
HmDXD2WewIEImbh6Fi25BrcyAz0RmffSlyuo85EAtlbpby2YZ8K0G/H1yL2QTYIT
u3MzegvV7s7y6sxffxzsSbeNkgL/udipNUvhcqHnkveDG8gZkVmC+QL1HHf4Imc7
uH4/AcIKJnjmihYSZd/ZYHnHddt4b0bdvV9to9WCquxaLFn+PqkHUtkokCCrcYtW
k2UH/Ywfy8a43t5gcRRIZigYLXlypWeNMxsyfnm0cH6HombiUZum9LGsEYCNXQbH
JDvMD+oXlkopLZRWq0IoGlGmaNqzyrSOv0U8p7N5zuvYgBa0bKB2VWjGP4zR+oWr
zcvXq5VwibkY1cENnELoSqGEedMYG2P/QPcrzNRW98AOFQ7Tas1g7oqN9v1jsDU+
R4MpHa1sHdZhCVNyDEelqTmI8Yt63sDMWD/9rx3Ii3dwGqVr7ZfjKAKz7KnURFiZ
b8Xfl3wkVu1bA3Cngh7S4UMSAZtFx6dfLUzBnRDD4RaTJcaEtU4f9njDD14PkHSA
6r0TwTByjmRIeLtKu81FNfn8uYka6KovgzqDHIPENx9pOwQnFnrZsDCF/WHBEj/K
buBqZ5QEsoT6whntOCsgnV0clep0hcjyRqlWSe/y9knSnIyY4RTXKoXV9uQKk6UR
1I8dg7LJSwd8zJhUO438+l41lJ0HhbfzebcaJGL4eNgcbvFgcfMqgljZ1lZuBw+d
p8TtPawZBZ6Jk1rTuA3owQilNa3uUYmrTuoUtMsHYgd9RoQsZHFAsz2Fpd34GAiL
FgTFboEPX2fqtqesFyjlMEpqvwnDY41xlPS1JfKnET/x25jT8qZUFjfJNpBWS2+T
fi3qB5kCmDwgQEU4FIIGS+EGpQWlbFadZpU5M8NwqkRUEtMlUzmy5h/8q+RxIWFi
rwkHlhYv+KU4MP2qdsEZNzIBXmrEbMra/Vbsr1KFDVYajXogWRvSAGEQQYILs7ez
MBlPRsOovyb7LjBJB8lObzeOiTxcv3kUNtOKcYzNdaA668fJxpwgGZTrg3iTm2WQ
OvGcFM8EU80n7qFp+2hP8mon+bOuc0tKtuZ3FMjyf68SpPGyn0k+hjtNjLNFoxnw
UIQtp0dy6C1wWO6yN10fbbZSFRKghfi+HeXsjQkQqQYBe40a/Wyq4KA9U7sYq+lm
l8ksTgrMRaOVFREiEIFC/qN+b9qkrAXcBV3IlTK8rpdiWt7Ga6rRvluGByNdBLc3
Gau1XHxA8qmidszSm6W6HcNUQHb2HQDPeljBvDRZ2pVu1pXOJAUf+065NgE+yAU8
I1ZLS+JV5HlVblJe5lEvQdhcY0gnoq6dwuRM83tSS2rI201pcYcfyjF11feDHKKN
QFF31nJj40K8Nm24BZIH8Xmv/P8zZmDQwsDqmf4WrUxt/HXUbdYa52zFgTCsktYE
8OtRsvPQ6zc+MODcB2fADDlmv9F7WwEQ8tURCz8v4JEzyyy5K9VoRaH1M6qkh3Tk
jyBOFihOM2v02veF6acmysfBrJ0OI+Sex9Av9PDUidcWP3L8OoYX+Tzo/6xrLLJW
znXnRQ2rARexUQN1LDVKP4zB0n698Buf3alerlmp3vqq37EtprIN8VVY3SR7itTy
JOETE8gPI9w82+Wi0bEF5esrAMzVFH/qNUHCi8kbYgR7NYk7VZGlfv3qIM0VagPO
IGm4AR0IDKVdpPm4r3LtKf/qipDNON/YOz/MV045s6b4im5kh3RkgUlEmg2u5l6o
K/6RBG9waTHiAOBCLHp4aDatR0jl/X3fLMTRFe5acYCAjK+XSYzcaQS/1cxlsqHY
zNAy0JqeMWMc1whb1krQbJwB6mk3+rIc3rVwHuwjg+hqpvYiVUSguZ+2QKXZbO/b
agRyU+Pw7soBTJ25DAPHkDt3UXETVTeyZBvrms8yvIKF5xOrP/odldEn+oTrzWXZ
elHteasV7BMyTIPzq7WpNqzZ01bLfaGoidB1nnuI9LdHl8S8z7RnGwU3kWvgFg1M
Iltbapbj0E93zKTEYPQoYLJPHwETcC6vUeAWQyaG6pJOqSdeqGQoYjhRvbsRo7aN
Ixbhx9JPwD6KCcNJQhcP77XBhCbd1PEeWvTBWeUnrDSBMG9Inv8CJL7PmB9C5zj8
srz/Wc8mVS64bGDB45BH6hOSs2y3mrWgNYJnxt/AcHLSPAkqPoSgBAVUTRpwbqUc
NC6nMYTxUwFFTbrk7i+Yz7/7zeRYgRcfgmamRU+EXffEuN1iuMSZsBd2mX2kFuKJ
6nHBU41KAEqgturTKxW0kfpffxg6bCN8+7RF7AUjv+dUPEB4Y5TxIhOan6X5rQQz
98ROkKQslA72LD1nm3x7CfuU4OaLptNEbZ4o0+CGH93Re/cm0xBeI7ueYRqbsoRQ
bYbY6XEzkOj6oqYWX0cPv8IWQzfrgIRtYMaj5yTTuSZ+a7yxpE3S5y6NXByjdzrM
qtzzqXhNRi5lKl6axtT87MVTespuwNWUrvagjv//Kn6IvqssurWEOf5ADzckPwJL
XKsNU5EakXn/mptHt4Wb7RauOOtwPQHkod/dUwYgXAFfhEFUI0U5RGyH2bcWVSrb
1lYsQmOeX+pmHdpIWpU8k5vIF7BDtpdTffdAJWG2qSJJo2+1X2Zh72BXIUaCrBti
wzitGy1yKyvQBk1PDWRm8ZDosPfp49ZOQT1UO1IfLvg6cA41gKqD5+FfTgSH8GGe
uSqM904iWyDR2Z4k5+v4seLNwQi1tWFHLxFyuXfZuBZLlcxokIYQ8QQtxgtb0C3i
owTUcv+JUmVhx7TWVC+LiLAKuSSuup3yYn5LKGUSKJhPlOk54S2cc+Uu4HmHNPhz
BJVYYTFh67Y8UXkkDJ5F70J/3RjnhoBjU2+C70Eas989CdLpuBeFQPoQ/uW449Hi
k5EOvBe2LRHH6rtd3xyUdvP88bUqEvBfLf7ovwqLa3rHDzV32H/BtxIXT4aSefbA
kEqiwpf8DzbHXd/u45UDXBTYEhUFS2t8cgWAYVNiPYHryDcNV853NtLo3IyvU2AC
HwbrTWNJ1DI5Vdoqc1nC8mLTB44FRyCEMPPsnQd23cnr/zVtAO5pznc1UfP0jaSa
j16Nc/T60FJK2QkliXbHwLYkbl1NhVbydxUIsq+6yklff6nxxjvCUx5mpX7qrZoH
peJG1Ard7XsOy1IUXtrmGw86mnR0M27aoFjAL3nvLb9t1pZToKDNX1V2Ngjg0zAI
GDX2m/y8cGMfup7zakiIxGD1gA7tlItsyBFf6LEo1muqJ4lqNcq+OGThx5ys5jEV
oAFr12cRSafiB8xdJ9JVKAm5CIuNphCANt/O2LJxjba+XPaJcJqQKJvojhZ0o7kD
iwsVhz/6bjP9zVBcQSnjRCVXwV/EvXXAgeFZtuad2gWESGhkFeccXFPOYYhD0+ZY
xeW/oXlCTCWJf9AF0OEiW/ekIAuC5EAUD3EXkz6d2ZWCcGBIuuuasYW2d0dS/2S5
/IQ6Neeuft6Yaqm+RbD939K1DMrzTUQgWmKXkTfG4h/8aXwD7eq3CzG/0RpY2g80
V6BteYiQix8t2v4Iu+BTDbDdT27hdoYz3gtzykti++Snyh8m6CK31XIPy9MeO7c2
sl45ZGkv5C4nsMzBiJiiKclZ8JQ8ziAcl/hSRdr4/glACq6dcI+uyx+gu/Bf73UZ
yFkykDoYLicCq/Ism4OSCQLDy8cVD1oorisj+CFUL0h8mqkPgeREUwUOQf/v0vw4
AcZltpFhjE1UwtBUfAZ2/8yti1AiKpHI3NO40sjCG70F7ZHSx877jesWELgo+PGH
CKTilPzyY07ph5zEGIu5lzENyePyHPI5m8YR/r3eplV4aZROK44TbHoO/JDFESoM
jIaUaKCkS2XNPR+D1sKAbbIY/p8bjJw9LMdnXIrJ1QZ/N2SAp44RW1qBRS/varWt
EpEx0j0qUX0oZka7sBS6rUZ/JCVb0csP1PzkvpoO4TB6U1aASgLMdMdkkVIqDN0Z
NHPVoihe5OYL3ahj8xt+5BiLs3cnc9kH1uZKoDRfMP5XUev7yYzOEBkiygIB7RPV
wrEC6E+PTwF3O2nzBCOnXd3reZc0LOiHMyNd4XaZY4pBrKfR1aMsNi11Tb5rALiJ
M1H8nO3TSMhgSCvoY4ZYwjWg0e3OTc41Yn1uwq0c+sr9wzqRoYwTQ/9HlAHng9D+
79bePu64L3DL18ooxB/Omn4DTirb34xQVmvHS9pydc9wcRZGkKll+2PU5yokm10J
dDeywciSMPs32EyxSQomPirePyxrZmYzs1pU3WhV7coZ8f7HcnRhXD9BD2qQW+xg
fxEvtLNWT3v3D4PrY6td1rpc4q3DSzuE0f2uxxS5XZw1TJYhg9KlxQYLZh8PXkzM
M0RJnZK/5vUm4dryj/17YgeZEkEvDyvMhM1DOcFekYtBfnN2XQFYHgDDbbkMa35O
BWPLPNuVZkM6detUx5up+L0I2b6DRHlxMKHh9GMW+qXgJ+NMd4fnGkfVj1pE3IHM
7ta6KW9RtWPo64sDQdq28Qo27gvk7ezTjGc8CNijDSbU5SRjfrlP0lvMQlE5C6Y4
SBoswg7MF883BQKo1erdChQGfgrVjddaFS9Z4H/a9Fkq2A6VY3WEcA4xd3mCZ4KG
yZQMaGGoOyHqnM04JofU5u3EBixeM/nmkrgKyu9ySAmuBuCF4Ox9OsKpzS4Ebuwc
JreDIIyjcaKhemSCPH/oyqc/WQRjSqsqeQ3TcXg19NQwLqrTHlRxh3H5WSqlhW9S
PljnRL6t5Lb63IdorwE1f7AILaqPegc9nS0o+aSG3MEcrpUyWJCaVruZkkmFn+V8
UigVbye6gzHC86BVwDt1aoJCD+YJjwPL0gIxdzTzzdLxbxTsVUZ2JA5zNMBxlb7s
U9cIgqkk060rSniSikF9UA==
`pragma protect end_protected
