// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:26 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UUAj5m9hyRUlMaKkwaBzGZMEUwg5r3Y1vok0RN1wFUyQkBVhf8VzB9PwuVdrlCu0
ZqHsBOCyqOFQS1Ym8uZbG9Kaz58EGyAUiPSsYFwcrx1JNfUIAP3GyoWERjXcIiuh
4KQr9Is9i0JXb2SND34a+8Wio6YaLDocSUSBydQj0II=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 93552)
rOSYwXklkdp/gAQOXJycEaLaQ5JdtUeQRhWsSkp4t3qu+RRE2Sl8CPrO1vHjC/Y6
zvdBXv6gcH6KSzlosZiS9jO28R6Vo+oIVASv9j9tvjfTYXbAZUtwoHZ32mUG1AZo
B7Pw8buCQ7Kf0Qag2taL/o8UfiYUViyMrB3gY7lPgw5zUs/Tp6OzaSmcFO8JNhu9
DpZAn7Pmf86p6ExBenz2yZourbIXvNbq4FImjbDahqoqZGO0K+2fk4zpc//LRyDj
du5frM7hHUfCZZSyzTQbg7RgXCcq9upwbGpu9B/h92EAJCULhIs05bYbdtBnOrnd
/sYaA2ZZCDJM1sR6m1hSeCZmuM40ZceBD1H7hKUPParhSJJDzyg8Xfx1vcwR1cpt
gl8YSN+5oUItoUAU0wDbou5CBnqJbHJ1JimqHqGDoy52A/sfIqI+g3mwjxlbvB3m
PoXRJ6WT7uJ4p9QduByDJ+mNhmptSdGyJK0SOrylyCSZ7XAV3PO1UioE5DnSGkUQ
G8ucsX9efzAbl0yxQ+4XLp2R5gCRkSlTIKotZ4YrQ7Yq1eKxarwo/U9oL/69GzDA
IwKRdqIahtueCC5M4eg3hn8GDt3vIeffnQT3XRFHUbFEsvtuupCueJ3Smc1XG+vZ
1SR6QlqzrVZNUKrozdIsCnBTND1UMklVvs0yw1UIS31rQuV/Vfe9OPdNfYv/cntj
AqYu3s9pjqWslFLB3yvMSGrfZsO3xHABhlLmj7gMmamm77DjPmUTtGApBeujpn0N
jexdHjb1bt3Ntt5X9yUtMn5W/tzpPUW5fi4oc/EaW13X+NJFRKXFJwuWkL1IT8n3
I9eGkdtau/ocrzbXLJeWrYEqr/R3+S37ktvjJfeCG3Ke0ydw3P8PZU3JsyA+SpqH
SLDrZfP5bFxuCjJ3UKSCcA6fn3yK8cEpqREI/pdPfgMwEqv+XGR1Yp0ZhBdwUBOL
NodWdsJFq5ZzxwrHiLW9ALlgmEWcV3TuXerC0tkRvmyUDldQwM1L/aEztQA1MfT/
428mSL1EXfAffH80Gud2pfc732ibrLxZqB25WcTDeI7jcFaYBvXh6rmyts2dM1i6
rDogno9nwC+ipM5ZkDQzHFekMmVYkZGDWjtiBqMM9zQd5EBB8QmtfSpPB57Ws+rT
NXvJmrKpIIc+1UR7j7EruwM1vGqL7x5ILvhj05MuyRCPcUGQZ4JMt4pLErFzcRWm
eTj5Eog6gl3INAYc3kajGp2RllpKXEjyPXcHaJbETP9tyKoCrFFieuuGCt8H5PfE
E3h9ElSLjwDkmsU/ZQet/CVC2YbzBq91RvKlkvX23GVXvs1+rrsBpejFSKRGiKU1
voRaTOfb/zaskOCOaWYUbJIn7K+O3/mftN1Qqx8jtcIDfv/V+/AZYfmPzjssAfFA
fB9/dxhYgRde91NMEiFQDCDdP0SvSWvNYNvKitegD/ZdiOr/mTIcDm+MeGi4X/2J
urQghklQCmhamTLlqe53UyPDm78Byucuau4myZq8XEIPkCoKHKv9hOSvrdZjw31F
hbfQcgO49XtSwEock9z8x0+NiyFA7zyPMv4iiAYwXWYTmKDoeVeK1psky02llmle
h/I0IblgwcF6TmC4yGLocozHE61lvceKoGgKbNwJG2vOKpt+am1sqqkbReHO8fTm
hOrzW6i5EvemXp2Ka+qpU5wRIWsSPjS253+XpsUIFJA707Vs5mfc3GTMwT0F1LX4
/bmtNubadeyzQD44mF3AuduZdx7nxuXEyBZvC18oU3cXK6SMQH8qe9g6i1AWhV8N
pNBSX3Wx7s+Hdaxb6rcMG/Ua0/OuggIgIvUJyQUHWYgSoOKM2FT8H+YDz7JNlVfc
27XqcKreMDv5AL0ThW4BtrhDFQViQgXpYTBP56gh/tF1vUkrc0+wMGM1UR+fZiA8
iEmo/g1uGJb7YY2DJvD/Doqrz61IrB/EpAkz081WLsvUaeIQKNdPpH8NbdMYQ/BN
jZsD9pOoYq9HyBZXiNnHvCWoR/xyr0f6lZqCbKxKPEaXo5r8goxG+jMRrcoFd27o
aEtKaSrKugkorChc3m2BTmj+aeV1tHBjy6oBT6dkl60nVHhm1O5aD0nkdIf5ELbh
2/VTNz1rIGmhTW8lmGXqOMiJLtO72yDv0e56d633qEHxm4pWCbG2hlRNAZjF6+2R
RtOK+uzd2Yn5B8COFzJ8HuPDsIDQylJ1d4lRd+dnf8U4arwGUu/0dtLgHBq2tLMk
Ik0h6fJMTsbs1IVA4AYhhXedk3VsP4jo8dJ4YTXmD7qufscXkyx5ehIf4WWRG6DU
V1EgXjLGZ7UC/GnjOG+tMYJY4Z540kArzv5bfjRi1KMwIeyLM4NyHk0Tx7nDVihD
swxB18ozxhCEkfx5Vquh5hdXWNH1CJL8gxaxe+SVyNCgYpBq6J483ACKE5T2Jblh
J3zclNIWKTuRYQZQiwYTCkx9uNSN4Kg97DJkckR9NtyWAU0gzDQajK8q4Gdg1rKb
q0YOPh+icQjGddegJ3MYmv2FZjswJSFD3qVN25yRLi0uyhNt5ihRpb8fntrPaZTc
VY9ZKmk/90ldf9t3RK1t+IyPtIXVurJE4QV9MeuTIEExJAyoEBuG0rJFeaPpnLaV
j4xMUjvo5xGYEXTINZ84rXoG49TtY0hp6EDcOhZGdKUufxbk4qcZ3VfDiEWgX9zE
RXwa1S/ni66CC9VKJ3DwtTrxtXlJ42UjYXcnaEWXb0pmBkCT340s4ONOhIZZQltG
/JeUPbJ0q2zkxKx1R215QpM1JsCaHTJ+IWs+faHYlAZcJ/sBGK2qOL/8zmFK2iQh
R5x+eFlWn5hVYd8VBOhEYS6NWG9HOFLSAnHXMyOC2pJPJQjj4RSKQpxjH/Kk3MX8
OCP3Jtv0Sh8nO1KGsYvQNksCtWfpYAnVglJHYhWYFJ6wOaCsCDYeHb3y61zkWjBB
y1eOJx9O/GBSvCVFgN7eCP9q3b9aIWDLVO6G0QqV6+aLoN5QKdqkftt+IC1l5oSS
VZpUrtyjXreMi2JKzVGxDgMEPIo8M0pscezQ/H1H5njQShTmq/Nvt+g62oQYHeBE
Ltcc6EwZJaVa/UeiYQ22zLfvPHphnAIORxXZvYrQe6SVWhPv2n7oTMoHLFhVx+Io
vl1Uha21VFwtArIqqDhoRzf8NJOf1exZ8DDylbU789OQQmPHED0sdkL0IPXeNC9R
/xOrVzIlC64II9N5CLtq4ncD88H+xSl/+RR8sSIGTVoEL54RGOPOdWP72OE82j6G
kfXR7mnV/dc25AMvSswDdC+UYMmP3T2UTtXVgrLI3xHvT8tBBvxPbJiQQKqdt4+Q
mCnpom2R0+HxLnMgqiSZlE+D49AWNGhLszlXfRMuMH+ZMlzdFfiCIWfIXJkcI+Er
5lQhOfCahmqt+sc03hgtzLiHy2ZLppnC2Csz3+th9vErGvl2Yi09tQ78ItbShHE8
U1vlWlA1Lpyw5fWfce5ymc3WoUnjTH65tsupZi5CDvXscmrEnVCqr8kPZDp+tm/9
eHxKnqnspB/zJdddqnG9rD02SxOGFgNVzwyghCLldqBjrDGzi/IUujZBHSrcwxA4
jLIYWPXBY3N87JuVXhF31scjrfAtb45ADsCqJ33PZF3nbVWkWdhOTSw5+nr46WUH
op6/EZKf8FyAj5YoxRUZusCYrXzfdC03luzwRyuR1tzzn7yfFyZpGsL/WWyWmmCT
oFvX8EAAJxGjT+joCurIVLvxzf+KeW22gc2PGJWUvYZqymHJIu8cT5ZDEEp9UWRb
7HChNxN+1LDrUv3jWebBh2uxGQ+yFGaewFt6o6ZEiqDRDUJgHmNyu1yspjeMb9ux
TFJhC1fQEx0oXWl8KDnF6lt1wQSHys+9Tb2mPpjz78cWtWsb/DVdpqpNVB04n80P
yMSIWLI5E8BBk1mzQIh0gnkdpFZkSwJGPTehIVzsvAeC/3AOVhTuxvnA/eGs3dS0
IWaQDS+jRyqny4pGdxbOY2Zz2/Q+q/6rDnwB71xqlQOvPJTNSzEeSc8+xm/GuvpT
/5gyZi8HH2F4tfsqeF0zkG2hRid+U9Sc05DaXh847dSKKK4MLpuZf8ZhLWRkwe6p
xY3mdRvEdx3TSYFDo+kBle6IdOwgOGFHw27l+HfP0gwFgP0CbiFSAw0TKAtmSf4H
VTVYQiI3w1kcT/e2FZp6NhrlDscCEUY9lJlrkH1sgepJaOX7mLYOfge3g809o6nP
lLKghPAEp+ZsUVLSMzR8bo3xou50J+fXLwcXzgckIQWlqP0VurezeI8yvm2yPB+c
DjcNthcZgT5tbByWlzxgfA5EMFGl8KFkhkeBGYOpFVAgCjhh71LWFaS9+ETzqulT
DTnRuDHbeboMmeG6fY5menghhoK72vlLWTgjT+kfgI1Ht4nZtYeLSD3r9v52kgN+
TOJnD6kgOjV3FkvhceWv4SUCK3uf5qpfHkGzRactfKyI9x9dCkAV8yPxy8glYq7u
lkm8uAbugf27O2V/mBkqnyUCR4XE7Hh49WBZAaUFh/VF0fWF+9W3NEDzyQAcZlth
O+wKuOIvDBjwBnvdQBZdXiWGyJrkUOwIus8MPBMHS39xrmR5Guxmd1v8tJ30ZAYf
tq3e1Uv/JKVC1sYPsPbp8N8fSJczHNHFQR+WDnjcEzDEtpoP2gLuIO2GfbqcQ/m7
ZssHCGjTo3tud+FqyPQ3CcRpZwWGzoiQOHzMGH0YlGvRMuGw7jyF1KojTSz+oi4v
D1B+i6odBF45rvCiCJFokXQWZU7p6jCojqKSzqyNyz3vM1d7r5WzVN9Ogwl/h5Tg
JLSDei2HWUQRnF23+I+buv+CbX5wlQyOofMCAUK4ltIfrYdSDfNi6z9hQD4gLTqg
JyFfpJmKWKZa+QUsopjNwHrSfI6+6kT4tFsxn2nAcN2z+IB0IgHiO6OMfuQyuqVY
Wr5nMCSUevxG8ooRihs0IB+DXlmF3YPk128jprNyuKXc3ze99T/wTyzEifZog5+G
SNCw6xzYVxXeVRHENX8UJ4+kDYSdoHNkSltzwdAxfYExAU8w3WSJWgQn5Ggk/Mlm
Onryn7opnNYVh46Jou+sJNmh0ug5XqUlefxVtktx6C67PBIWhkvuwcws4kQZpOeG
F8wSaz2I1JnOQjzqklc4zr8EQcoo0Z1oWp1gaHNyToUmhNoQc1jDMkdPwHPqfC8q
nw//pQsp53JyZZ6vATwVTjxG9QlN+DyJkBdFXvwXJcFdZ2cDk98Xf9SG0V9R2w4k
wPnvB3bDjAuorpN8tU6X0kieKPuvr8lO5R9ateWR48zfNfpHPGOM88jrL9Tu5yWb
t19F2SpnLKhT6I03qrHa8gkXHTzy147Vz027RxOrrZK7qJdyKeVAZrHlRomNpyEf
lAAkr4gdMrZGVxRZb9q2xGGkK9cZsz7CXd1GjqfjAAx8DqTdg/778qj6VFe+gbl1
r3t/FygA+teOVDTme6KSCggMsTaoUrAeeTJWomj7kRpczzxdrIwoIsAcaKL66HfW
CseLctjXTYgvc7R8nVqvoQOSkpZiTL2tf0kaJewkW6IlsZIzhznTHthNWaWH1e2c
lvnGtrvJsxrpe56RTKvS2sXsqJihPwhn/02bKEkyesnIqxfPi2A/AiXDPoTvxSuR
1kWAlKsa5hIL1NKKPa5Jl8pas3saXa/BQjIRd+zau8UYYbirciD7hKFuY4H2+iWl
jMjwFah4f5sWfyfsv2YDJG/cBhBDBXZzB5pb5A/zsG1DGRhBCoAzLbe74rTVxgxF
mZzSMd/O7l86j+QJ4JQKQnPducV5pNlSfpK4FG1PMP9n9iUQZ4vz69d+bPp9ajnX
BdGJRvyGpbUhIGm+pMvSq7nLep1uKg8l5/OHqJO8HXKqDwtGPXOmxTxChPz4ueeK
tNO6gAtsEPC3dl8baAb7ZGmIBSstiBxcxCtC6c43q8p6UDIpHaCoVf9sP0iwhyhn
WivDXc0RY/+fO239ZWMiD5EezpNVb5AF8Z3B/+zv+lENhWPs9o16nIQ3Tm1kd3x+
ZkCqXSirKM2szRtduM3z+RwIvTAiYJ7jCJnSsfiy3NExHO3xkksJqsVPSgBsHiz6
heHy+I+wxn7Rez7L5j/PIH54WpCVac3T1QvIpYzf72BEMXjI5TLPuvq1Nj3ISUA1
OIFQqmXbp2GqxxlpNJm1jnMEr9ptGeseFqUxT4jT+VowLdx9eG3ItlAfo8E0o+ou
OCpzl2eqd3Jy8qXa3uScOjB1eA0EiDnSnyGIwzUqKKZ5b5fDKDn1U7D4nX3WFu9t
fo5nS00FOM1Aso2QcHebkPfOVel9OGQ0wh4ocQ9laWeQUDcXlFLqx/cltOLj3Ukz
bfuMU/6UzddkFRRWp4Dux47dfNkLqe9dFJUI+XJ/t3s08Hlm9WyhsFP+x++DmPZU
lIYJB/WVEhealc4aSMU7huhl4JZQX8cL2qkn11zdNrYbaQ4JmHaF6h1b1hCCG6Rw
X9UlRs8pB9GE1B/OYD+GARWB7qmwaqfEIW0VCcmKfJeXZEEuhvugwj8bUs3eX+bj
T2aMPFy9SZx6PxFEd9x1r/qRkpDKagffeH4/e7tSe2HwlVgj8C39VG3xbbsSZBVb
2OgrP1BdGAS0atR2PEFfjzfZr02XgukhKyUPqup33zoz/3CTjR1vu7HdVEFrqDXC
BMUWAC/73SyE8jppCNnz4rlHTpohZeku1yWbYSztXdf/SKr/lNpKqR62upW2SU52
yjyIF9JlkV7D6Rf0Nrf75CpM+fO2usO0++zsXMcM0DUEa6dmx6jgD+x3HIMyRPaF
k+LNk+HHkzmh92dV06+06N37irFZaGzxCh0If9q61ExJ3b9QxFFPuK3XGtS4zL//
1uZN3OqfpGhFcWbsxcAJnD0SUxEPDarqQSMfS/kACyqAzZwbHhxNI9WmyEVort0T
o3Pf7+1aIF9j1kh+3F0LkVKfXWQUSzLNx4Yf3YKu9BgqjmbchAh/IdmsovjgM9Fw
PmKICXV70KBbBj13omTXDqSSFUFQB3WXq6xoSRVMDHIDbBnUtiAITm7S4Hxlm6Pa
OUZs6nekR4Tvlas0G/a0uXa6eKhS/1vlDt0BwPpZK9Tu0Q/oUyM30T4P2xHs6PCT
0wWlQDrY3Ek6AUT6U5Jtljyw9Vf9pJaEXiAeqraxu1Ce2b+V9HFJ/mbFgYV54sKf
1ILt73Sz0L7retI5zjs878L4Rx6LFyUWUkBtkKx75VOUFqwFLk2JzR8NYQHYORyc
rv0RJQ31YaCfbUiegtqTwJaRlTo6mINT2jd1zjNTXAWxBnMjeUZYig+iOiCTxeZO
5CzRqZBt3AN2Fiy+bmC/E8mhvLIL0XbIsGVfgJIJjX5mALJFL3KGI7LV7XuE+F/W
DiwXWOBc8zr+sH/vfMDzLhmnbejlYVar+jFZd2jNJsNJYzKkzc3UTzgu/ZFEetNp
VGwIl1+DOxvyqY1Lx9gJAVJg/W2saNkAm3qyy31TRRxkw+0OwASldBta16fMCFDE
qtiB4NV5e+W4dUn/ZixwC4rVBnQGEVraumtGkjs6Lsas2+LV0d/VaAvkn8Xe6qox
R7itb5PjO3eS1IkZGl2zPoBXZOFTUNTW1lZhouhcc1JqeMFHZwO12Y6d3xdVbLWS
c7s7B6pJh9+hXgif02jJ/kxf4Z+bozV2hTMYwKlp1ePjb4MIUQnIIVz0f/T81+4B
bAbMT+7GF5uD7uWFYPe3pAjnRqwT2uFZk/9RiWztm2guHFElSYbltqSGSiPxMsQl
SIJSl+JGrbAlwBrWuNNX/horrab0EllQHnl7L0gDUxt0Ln5Pt+zJSwavqjPS9OWk
SOOqWstT8NGw8LMCJ83HVtRCIy1zjpJ6/pNWhmAkcxApbop++VnsJRJLUp6EoTRv
7xvRTlSPrC7XpubtHOolSvKpu2JdQyT8tuIobSx8mvTCvI52O1roHZbQiucinsOk
bgxti5EXitj4vd6A9z6jCx11uhmusZGt2JbcafVrmVpwJk1fiHom6hGSVe4/6U2E
M3m5T/Di5vXel3fqgxF99xwf8l+gf52XkpdLJ2Rrmed6klm4KAmAdtA3PZ1B9XRw
wL9aPHAA/Xyg29D2VrksnJTITej0hRqlsFyp8WccIDxkIRMGsY3omQZjg3WVMf/M
jpWl5rPZkQAnxDClAQdZoLhV7oEXcqGypQvfiNFRCuQke1TmW+FxM+TulHX2ys2O
XqsnIklvm7H8E646N6c9NPLss+Wh7WdmOKetQVYgzrIf7wboMW/6neOFM1LGVipJ
YJdux0PEvFlD7E2tBQcFr1GJcWNzmbrtn1wreWVkMEWgBI8L5CJjwNoRmO7IB8CX
yRAY5Alb9k+LklHZVw6WJw2jpKHWtt33/zu3oScml562owoiVtS2o0uo8UL+uANt
32PxgEzNxJAiop5TUplp+a9q1HsOvFQt7xn0K7ZlggWm+srZoI9HlyCuI2VKqVOr
1x/tJekcbdD6AbN38rfQhtLiFdy/5K4LBTQgoHV9dyC4z4Na5aBTG16zBL46Kdg2
zZ/E2XitmczV6+733p5508XT6CJj1uNJkuVT6V0aGpV9TFo/ew8Hr5HhkGZhWTNA
pzUY/T/fLCp3C9HUCmz5Vn2hh3sKNEffhFH7RwOkVZntUBGWHx0AYZ3om63hnnM8
3VbfBIHCb2axA7IrQAFeyXGSM3hf5JMv060FgzFM4BeE4DcOViREgJzCiPYs9CUI
4rurKbABHHdFK5wqtuphndJWn5x299VVvDbowz59ttCYYMXAji8EkPnIpXLznyD9
RiQ0Mz3qVMI0oRBvXV/eXbjLlA9liEOyCqxGmozCiN3XfRICNUTIIXToD6cXkhct
jLOZ8c2K+OLkB4TpFJYBrjAOYraFaA6QymPkj+Qj3ENSvsiMZXibZWG67daDCjKh
VfWA7rG2SFyF9SnnXKzvO7YCSPc/K61xatbK+txEv0uWqOlKnoVb08i6bnirwsy8
KU8dPegq+nkz3Prpv1VhFy0d9CpDq/qu9I+ByYOd2OmOznLRb8A+VxDYPA097JXm
mDmE7kGKENj814WsKv5la3AARZyHMpjWlIMj+TlKzWHgcNlt+ks2xPFiJHrDcTgs
h8IRZ3j5/huU/ajbLbPbRlL+cikKsLA4+Xz9i86HbYHd+3p0NY3rEcxFxBD6nXbD
qUSBI/ee/9b9nQD2yxQEqsChsuV0dhDqp9tKN14vH/9GKC//gCLzvPUkbTMdHzUo
SVSB7bZv1RC1bFV6QWiuntKRjC48m2jz3/E0bkXxKhFqIecz7WPEZZU4bE6M/pnV
R2TrfMrkwBSClj0gA2GCHL1mrgUuK5T4ObgLpA9oGdk4t3bDOIu0KNrAY7OQW3Jq
F0wkmIYQX+/JaDqHxEqYKgQXozcUTCqQlA0QS2ppairbawKALhAvjBwFbvNi182k
SnYKEHWESxe20rs2FcBOTlt5Ugzt1xKnDgjnx2lVaYrXZejDRblbaExH+VzjlroK
qHxPEXzfelFI7Sw0dv7OaoPlnJFuaO25OFSEZD3Pqlgy15c4sBzn5tQdf8L0QMxB
0nxSgrXNVvRIQJi6szsZ7rqhwNc81GK97xgOTB62YZkg4NYgbq2szCAgxjr+DQz+
ETnK8LzA0AGFtApnbyDNbIqwRLcbXoYlRp+VZkGlyHFFR3YfQEMXBG23gz8Fal/l
jY7h4toJttsMCPMNZT3I8ZlUkdAn3DzJoLjzpH4hgEKNlOylozSiPYYohZw+txDI
AC14piUAF+f39/ZDo0eRNkpkn/VTinNVPSNlNaHtxS1mjFKe2CC8WwQk0Bw0cCG+
Y2Iq6xAMqZEvfTM88Fa2OlSaGJkhMWqM2FqRKQL9YDVPTnievuvta/ozqJ2QlWNq
X/He95reS6s/LkXmRYaC+nZcuQJO5y5YhFf64tetX20/o8UIkg/pAC71GwQQ/yVO
aeWIHbvT8E+4XmefP0q8Gk4FdD5So1boRL8EKF+J1Ky8Hly+o2qD7PAzISl2ayVc
kUPvL+zoAl4Q0lMxLW48VScI+tVuDTqfRV7xvnPMCT/3TnPyn8kc8H4T53FYtWJb
oPKX1uevpXMpnqzzNDLby4chtA+PRGxvEvb/ocqlVYbPi/xDAukDiVlzvE6LWr6R
JXrU2yu7OieSbnA/NWCkZh7NM1DpTKgPHQiEg7c4fEPdgIU1OGKmXvYHX9JLU6x9
5GRX6fpZ2LJcfPInxC5iGeN3EuCyp/6HO2YJkVdFo24I7ua+chHJKlzFbN+rA1je
HtlJJ12kMtMDoNTXIWmpAq1k4JeU6NIEJpZtMxpcZnpzeAqohl/04K05emkizqF2
dIfAhP85Gkf2IcxNZJPPXICiCrGVx9oWO/aIfzVX2u4z1eXTWW5FphrnPedsSQJJ
ZFFexenAJuVPCCwlqMZONZD0gsT2UaiHyLFl0sdfGg9VkqSL4ZZW/7xDTMD943y+
gLXMbVDxfZ4U1LNGPXBwMxIiO1WwsgkJBdFFRZxdfw52Zd8IpOw4YDJrGxYdVvJO
oHr+vd2sgXn8TOslgGOeSPEkTj7RuoShv5gXA4JESEEKkS23CYefWCMhlqCg6DWk
j3pgzEcvgrI5ex2d/BBGcRCy2XuQSpGvnMglEHnXGEATuXE3/hMNWMlUGKJU2tbU
PLj4morddbpIjsozNH5KGQHLhjUvQ+njw3RWb8YAUg9dSXN8TwdusfEnduDzzULK
EaC3xPpZOPfv5U37D3jzxSKWdeSd6p0DMuz8MAPHiXAUucWZ/FxWSIGdjxM36yZw
maWEjjGz0qBx1ThlDRTA2UGGvsZO4v4iOm5t00L7NjGEbalTeBJueF2aieMSfgGC
Bou5RBuFzTBOomfKbC0ZGnsNAIousEoaHNfUhLF0g36MYCIzdPFKPwuz1ibGYK5P
QO3nf3zWaVih1TQeUhjj2QCUhSY1Q77pOupBqq1C2HL+WKDXWVYhnPwgy99FJdhf
BEs4vplwLJdFKFKwHOQRUANgWgl9Awg3jnLmueuNd49n2+5LMfpTgxT0NlwDNg6P
Aj8XgCXfZefDBAV1c7g+cM07LUgZUwkLnUNhLHmNrC7TEDdOQZhniijixfrdONV+
qJ6Tj3QdfnV5dOMUOKu/lpWMbZlmfHX8EiHai/pjQP3VX8nlLXLM4Wy07D03S5XI
PWwuIAKnApiRAl1bJiD5LqEl0loR5McXaqrQDK1SBifmFqCJ/XAShKSV6M9UG1o3
QHhYseL6j06a1Wsmw2MINwJGIPrS7qC4DtpUmtmy+cScm1ywSDwz/nrlCPXkQk0j
Jv4cvsYdEg6LcEHmzeod3/XK+VhxCgzQX44oUm4jTXBv5KvtAQmWiVDcr442qBPI
pQak7SLy7TrdZQDeiumv8+De/VndZvV5ax+MQyLjJ26tooG5hTrA0YjUnwFkLFsY
Q2bOqCzGcVB+Ehsi0vxN59SGdm4f5a02EQaJ9KpNHq2cfkEjlTEMwwBTEHQb+5Uc
X/8HXsSzTjmgt3tpETJNHnLAoMuIvkwP8OfCxVxeSD/49Q8OQtQ6ad/0m4hEdtwl
PRssisyWG5upRicKB86ttr21dgKvQGfKmexAJd5NHkyTR4qvtXRYEzF7Q/y9zdyp
sJ/pYGnb/5yRcouZ3zF5DGTqDgkL9wqTcRmKL75u8ISQfEt6XczNG27aF5PeMoCT
kl0Et09Nvtheus4jIGom+zJVk6pMkKvpKcjyUWTHWUjy4cwlZ9br8IpzCdwqf9Bh
m41C16T6r9uoem96CjyI27fXcVkmgm2SjRDIjpJ+gXpYBHUcSzBJiOReqwOOLLTl
+OPVaFJFlN4CsOv88QX59fCMv7PXCTA9+js+zBnFrClzIxfmaD3lPQufVHFhpTgu
sBcsAhSU6cpBjoM2QBo6G67Us8VQEUQrj+tHAxit4ww5z/fE2e071CO/PVRjqwB2
TfilH8wMYsslbNRWiPqF9QIp81DtJxYn+O3NRVM3u1VMUlpjtCpRY6eLf9W+cBSw
nNbeaxMhd/d8rRwMez3k4iEO9F4MKzIoe5RWOd7L2F4TrOtCjc+g5/hxV0TMwCBo
l096dXypYouaRA+7u8l1w9cTGg7/Eo1kHl0ttEvzd5ED6REzgoHaNQOvWewM3Td+
T8ywzB9C/FBriokcc6E9mW6rxB8czPCbqhjvDbhYLa7R1R04ri5NHdwZDLNiUmVv
DV2O7H0QUsxK85KDFKpCIf9wGvYccu2+7obPN89xsA5EwEivO6USYQo8xdaudRrV
PCku+aO/Kwb9SigwkHOUsgrjAgEjIyafYOxiYEaikqqj2wsLHnmAUTYoCJl/cAED
Ra7N+Hs5yUpNYQElqU01B0lGJfy7sTLhzs9bwUeRI1M8mhlRT+x3y6hfxo5ImgAc
z+Oi82j5XAIDT7iorNzi5BsPzxFGoAnglnVE3yAsi9iA6MEiGBWZ6FCM9uH/qdEb
0wu65/29DLkPF87OsXzgXBWCljmi2a/D647onnK+YMkij/R59Llp0gb1Hc1c21C7
aPczKKXIDbj/6j1FqcdSnJ2ncEwABLmperHhBgO0ID65OU98dfKsz0vdVeLCH0Yp
/FvlXuIDDU/ZqWR024TTaPwUtv4C/n8yQUlXlG8OXZgbYwcqDK0bxP5Um116WGBK
L/OcYdZ1sYupucaOuzq4ctAKPg5+Hvu1HukvOgXBsaPghOomcoZLb34tuehWa4/2
6Ok3/TNY6PynXW/K27mJWV1SfZfWpQmdW+AVo+K/20vGaXQneVJTYYkM7qlyYUWr
cJsAfmop/xnvMYF/zX5fN6b379EB0eSLRMgjzNO+3i+mgDwNReYY9z1jytJc5abn
1OfnbhChuGvf1uuuu36gq057tLyTaS5x0ONKWsHpqEk4ItWvcb5+dO6km7tRbMEZ
AZWxYNdeFIzwSRTCnFdCXoM0EYzMwLraCMIzRgrCOT7Xq59rdFWfU+Ho8PwcsIy3
q3LYEq/gOJv8nYQOfU1BHdOoXHFDHPyYNaIYTx19WSKHo7aPQ4DTdzz3pXwTw9re
7yZ7rZmQvViR+BCwXYxLiE9Ds47KcCODUxBUYrGjKtrDnnl0eeCKetzojOtBVS33
7gObuxz1huOznlWRIUtP6WI74Qrd36Od7ey+8XtojAd30wkUeYJCefL3K7O8E5uI
DlV9Honq4FFAcPas1D0Wira3DIXjNflrnlH5KkF/B+8sq21dH/abCnA5vmBruBMd
PRV+bnaATMR8o4xFsi+34nbouaH77Zpj2pnV6o8/ZKUVQ/K9ZiM3wdgG/PqGkE/t
3rqb2IcKy8Tky3Z652JXirldCUfX7LHqCkjfMt5Bpq2Dg+eMvx6d8TLzHR+1n4ik
x8tjzJg+LvP3aN6k8QwTsLL6KMCeOJhjZ1JrH3WvuLk88EZmv9BGfXzn+J9JNXyT
bPdzihbb+aozIpB1Ir4n5dFlGCtNgE+oty/RGCkoxy5lWR7ggP1OgwsY7Uvjndx4
uR4PGNDL0vr/bJPCHXJ7+n2w6Zexp0xquCgtxY/+Iw71x3O5f2Lpc5uhzHOpRSZc
hGi4TwgBgfq6HzpJ3BrLBYq7qqmFi9wb3LGA0Lp2RA2FU+z7d4yjATuq0RUTpMfz
NFh5ZNszlOjn/mjK0ppbpg3dFf8nnS+tlcY9Yv5sTnHB2is4O/qtZFr1h//H+i65
4hMsFDmJwYYWDkpEJCEEb81RUojQ1Rx5NB9Whc1kKBYCcAhbUJS31p+ihliLaeq9
OAwNYmuAILwPDSeN6pKywmXo+XR+xvCfODY2k6iFMrJflKsIsfC6GBwmV4bH8M6+
TAihetfFG/+9ECi9wZhaxZjlh5N/1t//m0OwNzdMIp3wraXIYOXsIWLjsqggcKDJ
3TGGY64wJBf6n6Tpi198jcpBqQkvwlti7HSAn0va4adwisr/SZ7p5962r4d+ZXJm
o9hiNw2Uki90wLxU6d2qnqkPOsQPnqhFXX4T6+XJgZZePqUJfO9YSG+9WNJ2EgMP
OWlDJ0xgZY+fT8JqTSGKUzz4KY73cnakQYv1PYTsFb9MJEuBrvNQWo00l32KxrkP
sEDzyAGnY5i6mSVE9ZP5VuPRwJ0XxghfE9nGe5DkkzKeax1dmamu3b0+G5V/0mdv
covNQMTSK3xIMtDXseKAtA2W98VGZXF7vS1XZQbYGSxiGpO87TXuH+j+yJ55cOem
b1gsu+zeG54hjp2F+W+EivOpdbhiCUOMMynSQWdE/vZYdGsuPAJLGzf7R5I8lSvW
Ev+fSFrAPnxvs2N/2Yh1mU2tTjVF4ERyww8JvJY3A9xsqJcnHGawsJxyK6Pjhl+g
yBJyrMz52Bx9qftASsptVWyOQ9uZe06N2CHH7aGIIVQJpqnzdFVS7aX5CstIayI0
+e9/NxmKX7uKwd/WBmMW/wiZxpmoNR5js4iDT0jx5kX4BlNlRRR8uFlvLi9HoxNr
udIvtKb82lMITjH7Hf+YNO0F3uDZP9BJguMxjpBCXu8sSAhXw2m7YiJtuX1WdDsv
6e0pCbg/MxtjcXENp5/cIHxqDtyo9rzjFkvV10i9O9f26qFPEVOY9jBlRlSddfW7
zfyWEhC42KnJp1VvQT7A91tGmyRzct/IbvEHWRVnWP9YVqVoB7DuiM3Wfiuny8+I
K+l+wV3H2nZ9F8s2/NoINjy09EeFdQCWJ7PPYmXcdEg3aCRPmuxgurl+BYzrb9hd
+qqI9rVqUDTkm5dzgGf0UtI+GW0diZRJufn4XRG+5+4xDtsIpNOBB6zrdLLBtGNS
6B0bo+W79XUL6zt8WotrJoFaHM3aokysDcm3A3FzyjYZvmXMXYmu2BaWJvNDZZjp
JOvBn3yY+IjdHnmaj+H/o/huAItKHjzPCpba1lWjKxuvyol2aUrg8z0Sp4/M0ULx
1UniOvM8AlEjMjFS7GHRYE4GEQ82Oav3YNv52vtjrIhAe8Jmxin05+hq6C65yROE
IdylIf5P8F/hjHHDIAO9bLRYbvNnB2q/Yv3ADUgYbKFtAvr2vEfLSSZHYitHSFDL
1inhRenzDn6DAog8j+HtfkMm0ypJ84SUnS8Gb0ToaTA3gi5xuu+VxDNDg3zIubcJ
RBQNCWuIuNPpfF/acPvqWADfeClfC6LPZ+xhn06sD57JYBMsqrJdjny4IM1IH1s+
IzZrmYuPmo+ywDfqqLXMzBvNBvYbT7X92h+DkBqzYV/247kfxepdpYTrPDuAUfLC
V3Wntq6rXvys64RKxbwI1WmnX6Pt9C0MEPraS/Aywx2dDuW+eXHU4ORHftPfFr/p
FQHfitp895qrz3yjIYRfP0ydFcTxZCihEOgi8uZ77QlLat853CTkCAb0lh8BLcmG
6dA/eXWKcvWWxXHe+gbSMEBr6qKEUJqiBMfxcw+BTZprO4JFXtHKBYyMyI0afRmq
N5zYWCNPUlRxm6/dtbqntwhNoywvgWsFrbsNtvIi5FxTdzFbGlja1wVJ3qhiejCG
nvUCNjGDDLFyCzHG0WvREjrrsXkNlNny/5J8NRhC661nQvFhjWJscovRn2S/Kyx8
4mQ4SLAJICNrfYcxv0zMhZ+Eo1tMD3Z2/ZXgYhK4ChJw5Q85KRtKlJ1uacsQ32b6
+1niEPD1+xxCUCl0rDkiKIqviVmZFjJfa9RCrU8ryf7urhbDez7YKQTyWPhlycH9
Mi66EGyFk2+feqkqiQX6wmxXvl78l6sB03lTZteBySFtzdPYnFciGkeNG3JIzEcT
/TR3+Vu0dG4REpLsOOF0O4HAmZ7C9pxJViY3Lfv2XZOfyBn7gaEcPgbHR4ZvUDc6
K71KOEmRfGHmEo296Oxw5v4hnCI87QwZHgBwkMI9vtLeCHc/J+nbGljmpjczBftg
NPYrjJ9XTpF42bAAu0+Oy7E/ocrv7JtqAEQ0v6necFDxW0c+teWO4xKEUF4TnHBr
wuYLzgKT+I/2BD6+rkFkkRXMT3A+GrnHXfjafDEQyIsGIYvb3YfM5tJcvFXiZsoO
C3bHjYNJKgXgFNNiDFiY7ir9lhOdj590TO9yXLaOZvRAFNBZTi4zmAIFn4/PL/il
/Jf5hRH7Ya65Qw1vUUlWbfW45BdtZnV69iZE/+YvQX4oq33KTA53LBR7CbUCfCHk
neooBb7z1H8L778nwLeOcXIED3epRk7GhLbWCvWJxWyn3geSEB36h4AlvHMaIJTn
OfhxQfwwRbx1k5PQonxMwvqq1xXhPO6rQs0dGRaZ7xLD+pTl/UOwNWOmDSh7Oh5w
TVfzJXaZ1UIyPy8dDXhuyq1dw3xdyKZchiX+ZotI4SRZHXILafVW/YhlThx+ynbT
1hG4zNWxtBwezecD8lCoQKZUdU40RIAr6/Hfji7ThjhrPSRPFX7pRqi+n+rXAtQu
k2zxmZ+DHtpn0wyVXz7DS7bgSKisIJJ8R2xYpHUY2BKxH3c7mMQ2d566NVMgK2U5
tXObbtr7ajX++wSMDEUZSFx5k5Xpl1BpIjTSJmSAGIBSI/XJa06AI5pSzLqry5o5
rV5gq9OvhtrIctMbRk40b3yKzR3gOkOtolxeYOxgXLFxXO+UVaKBFvPcuLFBdjae
cMwce2ze5WhR4wtWwtF+53GXe1oOpcI9pz9GpE73Aw5FfmIeC+eQOJBLlDgp4KJW
H/DVUz+eM1Nw9+S+qWIOU9ECjY9BSAiYIEvH60nk/+ODI8aq8R5oR8akl70eVT8e
KQaQBNbVBpSGrJZ6QNAiU/lJrST4cWL8vlRFqE6d0Q2tRR0ct932RyZTZPa3V7yi
T/U6/wgOUYbLbfNEiAg0RH/4pKtcdtBUSibEcuiDsZYDZPrhbX+FH4fyA57YYfWq
7bRruf98xS93UCV51VXmkp7gqfM3t2WUZgVsvAzbAu6vUezSFQtuksTQJHXkttrw
Fhi1Mz+5L/JcFROGyZdoErcJEsbC+grPq83p+K0XAQG1SrQLnczzV70XRec0diKR
8qDQXNql7AvQVAtPpscMCPlUb6K9xNQ0QYzVLAiSB1x4EoFHoLLkwZ+YUpUNYS5Z
smK08HePpRAq7ijE3LBZYGO/WUraOIppZT3PA++hfsMK7M3uhsGtg+cB9h/gcMJa
vWp9dSGVN2enN6cgcyKnAC6+P/3wDgesgmlN0i+KHmutQspbtg7gj8K3JClV0Rcg
wFaZCIBa/dMQyJSx3A+M6BNKYocMLhJ3FX6PckQPOUaMeMfhOs+AeBmUY6f0n8u3
ZLHemfxA3Psvz7r+qyu45h7/fAa5N98JEp9Cihe053+ZwukHPYiilF/M5bbXK0zf
A+JRXT9ww5xXg8mZC7x0m1B3jFVQrCpAG1qVfAu32GJJwwxI6VjexDvMQx66uuhX
9THOD/UMBXhsaUROKo+HvlnF1YQtxhY7h/OrdoK41fAMA1R/CmH/FeLU+xrIxPJ9
9rBwkCR6DEpbs044TrltpMq6pmgXZhAAnJRNmPTmaiyH/2yhZqh4wxqsaTcfcc6T
KaQPSJCv7BBSqhg6xUm/U5NHEQO+FjjnmRyAazVt7CNLVDFxR8OmL0N09XVp2u1t
251aTu1OX5xmbmSmhhcgcNQ9Z6253cD06Mqi5htdE6/0Va3diBoysp3lSBjUSlkP
d+++b7/6Dkv2TqZj0Edtpb5Dv6FpunV8wBUI/0nrDza7eYev80X18NhEc3b4gCcM
qiq8S1SQdMmHnB0OlHCoSzLNoBFOuY8TrV6CoHyupX1mMEk4us4MNR7xJOSpgOHh
TmsFsNj1gzFqD09iAUIP1Jb+zbarOcBGRjo4HJte6wjyV1oKzCSnJS0fNP11aH86
OJBGHpMCUqHjuKQqMHUBf9Pn2Dgcgh6lWbq/BDp2b6Iy5yYuGMuiyPi7u3MvhBjF
GZFaeFFSpvBNe5nnZtn/XQugDFRoAYcKDxEmnSH1He9bTPp0Nr4hRZKjKwjXTNx/
H2Feyl+CzKRBzgfltkspvxNUsbGkSRk7V6dZyJ3L81L/7YBe2bBJMZoya4d8ojbE
IwpTybm8yz5reb9BohFD8NJm7uldEnQZWT3Uhvppryzcnjh3EbChYmbXqNWkoTBr
twqN0H2L0hZTwJ/P4VZdf0IdFV1rZ0TOxPe1j/ENSqxrXHnzYl4ONZgEfLlNDN3l
srf4RJB/xrntVNZmeeCqIH+frjKqJ/LkrjLp0gFCjTBGHSysrCuz5aRnB0oaEX/0
CxluUzqZ+RfToEg57M7OJAS1kV30rGSSm8uriM+MoZ+6O7WMSGrkrOS+QfY5wasQ
HjJwqzqeoP/FewtKVuI/5LiuqOYEIzKvWHnqmIenZdKxuGGK9HrRSar7zvucUbw+
PJFAPaXxbz+zwd90LjbhShXI7ECU3kJwPt6LzCVhFqmyoc1Hca5lm87cPQIVqJWz
VN7QUZVMQvYUec/IA65K8EfvHuPd66n0fElMAmVWXMM3qEGzbJT9qI+4WRMGeQY8
/PN/NPBuMXDCzx2kMUR8P9jYQwkWiwPmne81+e34OKK3gSnDuelv6qfuAmXJ9pd6
ko7hdhI6S4b4VplipT2r/ccG18AQap4OkZDot84jbAkBHXAqtzkmtRxGUjbZp3CX
gqNXEUwFR5nUqiMM/SLAZPvkN3+j26zoHKL/QKt9ap8NwFZPuPVFe2k3MgJo2oRg
8iJVhjO9K5jSW2C/m39HWYaNBcJVG7wAOU12w9kEWKJpo3cI/rzZgK5fahqN0Qsy
WVFdaNEPy+KquAa3joQEd3eUxXUEpwNSGsKYGvBrBrlS1MZi51QjpnIOnCjaydgK
5ndygxHZcEFRj4tc/QyhRHbUIObskzf3ii1g8R7MgjlJChEGqmFGcyPfWdq+9E+w
Vkj8KMEZmsG4E3Mmd0Klmw5k61nf5Awlnyh3+AN0/DosaRps3gVHST1On7rppbnc
40bJlaFnzu07zUQL7qSWAqkORCj4mkx6go1gHIPJE7tRieXMt9TuAwdLPBPTLLa3
j9/FztRZ6n5FDUpxg1+c/dB8cuWrpzK5PkhkULX+/b5swHzn2WWGu8XaIIO7OcHS
O5KrHS8GlrXguSZIcnAVLvvfhkeR15SOxr2fujFXPF+S7xE6JpynZo74dhBGiixj
YVsiyweNFRAvFgIWAZ3UyhzN4cxhrBfv6ByBYRju2Uw+cRgAV4+kxveCAt5eCGyr
T2ozk3u2NMTMIIjLgdPMHBiCrDxcD0Zj/jIkUzz85YGGsiuxGqrVkWZPcp0pWJKz
wH7wTTc+d/+u7j2bIZ72/F9fL1q9Tvso/gVisCq2OK/XwZR4nxr7PaMAa9c4ail/
gumeS3+q8DnFTToKMnEq+tP4XUC+bWSUgKEqv9nBtPEcO76rI5XQJLEAm6n5XMti
v+BIg/1tLRk3ijLprRuUnO7gamuuNbZrvwbudS0/vvmDFndN5ZCGnz9j9l1FyEtX
VQLL+QYmuItvUl3hk12+7R8wh/qLcSSGFtxmBtn66cTWA5lLGg8RZVS4CZ+asKgp
yaMxXFkhowtkitV2M5tJDd6KtPhLxVZiHpkRxgTJfa8Kss3G92wsu8dRaLjb2Bqb
kb/RRB6r8LPuVcL/CrT6e5YuCbbb31XQ028lVz0pXJFcv/Xj2WtZ/KOwOLtB59Vw
8ZeVNeWteht7pCI+Jg7r4GpM7bpMydXvE3Z+L29NRQCsaui6oMB7wjHatlKNYhPK
NYubNf6gVCUAtSBloWvqu5ITnI5olMJ/DKPSNUO3zU6QXeJJbGcbhvt+P9OSG9TD
U4Ewg3pOHmhJRue3mbeCROn4uCzK35nHecss2mWZWg1r7s6RCOW0Is6tTvTubD+p
cqOC0pg9jzFLY4q/i8f/b40yUJAI27LCY8yGXzxT6feUdNkN7qWfGxZJeQJpgRrd
fSe2GZxfjBEI0urW6TV+yeBOdqd/CfwNwpy7zPh7WbH8NWn/aMEFgOEdCJY32A6q
jzRsL/2k9AzFFub7r3+QW3D3NK7kd8x6tEZRI0noMms8Y+kIR/wp2WUOfCvlIubr
j9nixwDUNiMKuAeS9uxIOb0+M/89VsGI4elIuPQFfGeZx7axLEGJn7gXtP8HsnLT
JVHqpDjf0SbOD6Foprg92Cf8mSvgof82yIFqNeg5tKCIwIkEa1tjuJpDVCVTEDp5
0zCdOdr/8a3WVtEAv2hSs37z80Gr0sCHtAA9jkTHdJT1qipQivei+S376u7qBAWP
c+Nq4CFLuOLhnbsXXQ4aO4cHAj/evdnPO+vsVFHFxkSdoJniveBj3j3+uvVv5XH1
fOueU7s7/1Uzmr3HG/IvJh/1S3yB5hqTy+VPu003ftLSDK+xJdMIoMCth6HE4392
nTLl/jwMWDXxEzuSygmhU18p2C3t7eRvVSclRTAuLjBV60kBywG/F3RlestLr4SC
9QYQpUJfIG0D/FA4G48Nx5PsCT70wCCeeKfMVcSxfqHziEjBFTnmGyNfH/IA5wZ5
l79tcU1COTo4hZu5cLSRiPNsyRGsnu6LZ6SDGIQ/izbj2s+PxTLxAkNf9FfGXKx6
cKbbHRHfYmUVR8gQvjT99YWTNmhroAUJeu6qwm2Ddr8UlOXb9SDFn+OHtXk1Ka4n
hIZ5dN5mnr5f+T9SOBku3bRmZGUdekwzgzDQYa9+wlSI6vm8AsrR+CX0HEevt03p
h3h08AiqffX2gtwaLDDwDvkpbHfkmQfs1XdjSA8o5+Erh5HrQyti7Tb5jDH5UB5f
F/C9RiIj9p4VOOxCjAed0k9qY5N6n7nwatVmDl+6gpy0qX06qjVD9pgV3rNh6EhO
a0zXfe1cHY8zVnbfwoOyX1yx82Hp0xkz+GP931daL8NuiJ1SpTTkqjdSpW2kXgTn
Ao4FUbDn89tk+MgtnYJoyHuD4DOOxV5UbNRvxgLNnV541/Y+3WAZD0Z1klMmfQF9
ntcHrZ+pYDtWvzMIdZw58odbWZ2dgG/c+0WEZiAA94ZoAqOep3x63DlfEGqjsDs7
1ogMZh/urams+BfNGoIUN837qk3KgrxB3lgnVCBEaunVij57dilikIacmCNrfhXk
ieCXbBEMzh2JOK71tiVt5h4BMpG5PIuWLi/l4Sf0u96UMNmQzsFbc7vqih/lRnz9
kgBkLpsSCYXzWxN/y1he3wLuQdt59J6rLQ8MvwQdZFmGjT+YL60octIJhDAlcuT5
CAmqHDH5WmzCz05Cx1i5wfxHoEv5oqXguJgNIV5zvy/tEklgzLsXZpgXkKbQn7Mi
cBfXESwoyZjef5Ozemdf7pHlJ1W4E+7wlyA1AJR6BEsWXluI/2irokEcSpH1x4VY
uy5FNsBx6DNVp4Xi87+hb8BzwOaU1SIOEidkdmvXn7ufAhc6fWu+jLp79uQPlIqM
LlUOOGV36kIcdtqkeRfA5KkiljOmyLHRUTav3jcUdAx6iqMyYTbUG8o7QpIkG1D3
lflY6+Nwl2zrMeeaI/2SRwr4qgm0IzsN+muJeZvj/6kt5WMnUiWq6WQfJNB76RSA
N1WHulk+ugi3SY8x/iR0TUyjN/T0VGUDeXxemKIYyBsb7Ga25Bm9JOpsdCe0Csbf
t0nBnfEi+6rn3BoEnCWQ7jzG63pf7wE0nUUHD5vj0zaXa2KRTYup3baNEFfEwIdF
N2xEhnAZhWofeOkOiGbzq9jmQiW3ksK/yWasYGaEe9axtzltIsWuEmAgqb3fVMzm
IgdtPVRTBJTv4Fo++jj819oL9L1z5EqZ190N3Ms0sMx4h7nj1m6/MLRV/SLUaTwS
JjsyvJPu5KWSHPKoQ022gcuPY6s1NNoutRrUL+QMBA0/kQ8LYimcqu4uE6KO/run
TgwTpUQlj1fQb6QUUqIpqcN3usYY+Xp8ESIr+k2DE2+ybBwKWTDB6FWo2SIU35VL
z5lMZ74NwajovzN2W3VZaIOssgzeJus7TGhajNe11EMt2um9t46SccSyeRGJ72G3
S1lIJNbnrOzhMpy3AssOyNiJ1EkMeIGdiIEDPKlnwebmih12p+6LTip9Qr7evgLK
ehNjHpIMXTXBJ7/cjVnVBXkcnFRQX0uaAJtDARaxRiedem0f8nHJL3Sl5DW5jExv
9nCSkxazTs8bL5/k9//udFJBXl7i3tqgxGsEuf+qCsCTs045l62dQ/3KRQswZOm0
YRsNXR8R+m66MJ29A1EtURRoEAir0lbPsa4X6VRW+N7LJ8m5iAI3sde/vddIJHRu
iXNZBEJcetY9TzecLLdXi2Vl7iUM/fn84ri65N0IkvAqTbF00aSDwwKavl0bEVfg
a3e+G47MXCVEMneCKuyEIy7jVX9q75JJABW2asRCTuvgy+bJXX08jCuRyKiMhuQ8
PZWohjNkQI1M7VEeLmb40VEqPInp4Dhs//C4gcexvcOfeDbW+76W0Kxn58zC2xxJ
aed+2KPBVzuEtptNcVdYbNJcwbCw/xQJAqu6JkXsuO2INORpul5pwEP8C1W65FGO
d6lNPOGVA8+0kX1DSYySuYo4fWrOGEN9GJshiEOuCyWOrf1SKb4Dj7sDaC6D7dj+
4bz6rFjyu3AsW14K27LXsOykYDV28mBVNM/4uYT576ywNQ0S3o+eCdOB7ZCDkUY0
4QTqKG2KQKpTf5YEJHG2PI9wzvaJWlgAlDyCfqqByrsGRxAjdPcENDlS/+ig/UTz
dqpmk2YQ/Q+QDYZqJ0W7OFJS9tzhPKy7YMw/zm3ihZ2/LMR+kJcvjmtpwEx/O0iw
wZpcEwCpFOCiyczAfNzTls9W27O3DgdfnixWrJaPLcr+ZPGNIVewQI2nueYVj29Z
nhV8ckLYeCgpiFGnBhznbyqtl6ez67WXGz5+TY4L+wgredh96aoMA/P9l+3wHsDm
/Qw35sOl00trgJf9zvCobOsUWZ1/fA2BkpSkKOxWVn79L0ppggUWUyMs4JX8x50U
uSqy0Ws1z6r+VWvfKJZ9HoxOBQau0xsE4o0JXf6DpWhxeoeuvvSrO1I04USCRgHB
6T1PWolQlJxRLqbrUS4SYqAD7pJuPbZaR6j3S6mP8XmOc44NkhqBLBUo5gyQCnXZ
sZSTdz+cLo2iI7SAitBdLC1Ahe9eonhab2nKj/KkskSlE6xev/9wrCHzH4NYyYQ/
lkS8tV8FvG0UY+o4JWDU96s4pdsT/QzkaRFV22Bwog8mHZHllHzuAH7vyoobw20y
O8jiLa2ixldKJcvEDojPSafkI3LIeuHGAaqqANC40x+C1qMAiKIPu7OdX+org6yi
9IY/Gvv7zaeuqY4BEHBf5K3AmZUQgIiGQnYTGbG1X2RtW6oACZ6NhQe8kiT1PNfL
WbPE3rD8b3sWoh1XJTYKdNu7bPQwfXC2F15xly07uxdRJHUYzwdPNthiu5uUn/ev
ChTwyc8IFDC6n3w8JbLoCY+rivZXYJhVrMElg3MdzNKVrJRjmhUQ57I/ScN8F18r
CFmYxn7tlAeGZkltvVFBIlIskRzA8Myk9xLlxboDJbyHxvjPAFshLjCJD1dSzpZT
wKTnTuSVjlckYXf3s3BuXYFEiKr7WjOdCibPVe+tNe4Zga0fxw65RFdFimtxJJf9
muuiUdxkQi60f7lXU01z9Z7scoG8FbZKT4ls+FMtQuYPHs0rqy2ufWHg2eCDvK0c
yP00YqPMngxTEM3vHcl4yYhEr3bZ8KlWNf9kmTGlpe536S2227gXJEj/nUWr1qXt
+AOmYVy5KrYZYzohBm+CQp6BaoQtBiFIRhrHqrkZCj9uEphR22bTmGvEcndjKKME
Xuh8/6jkys6g9BWY4VCdBhiqWv6aJl9RS6Pz5onI1oECjp81roXEdP8XPPbG2SX4
6F1MdHzwBa2WvGZ8dCUpGqtTMwnexc6VgCUqQU7bcAWfl3z17ekxwkGZb5NiYxG8
K8+vmmEuUhH7PbM+Z1YtpRTvf+DV687dR2bBA6zOTiAvUCKxoOcZfhqP8ZjeYgOt
MnlzNLAJQce1xcaqluT/FdZD0BEE2Xvm3/jknk9CFkGCSSf0sPBqTZEI8VCseFtm
bWsY5ik3gN93mHzKu8lXRr8JG/v3H56bCmY943FvEwA2Yr1w5qlsJdYNTUTXqd5u
s7W+GXlV9bIv3wnk568PWHqcLrVn69PPznqvCEvF7rOm3aECOYpjLUMobje4SaiC
ODVieVHRDlNohmV9GqT6chj3uzzW82Ys5fq3v7QVny/P3LWgIc4SmLG7J5u7E/dI
rIs16c24x8LJR3kncBUcA1IjgOQgXZWGW2tQEdoPpzsVUazmvQzlpFipHc9CElG/
oR/oI3pjxuk5rmNk+h4Gm0E1+kz1UyZniLLxmYKDavMPSmFHWncpu9zkcr+IbKL9
bKmvVf7Ne+LM3OKhB/6nWRm50GWHBVk2kLm4U6AiMiCCydxBd/LV4bzGWTDe0ncu
7AReTJCGkvCpgG6BlHgV9HIZGIyT6P2qc0/Wmj4NceFPDBWfqsDPf+UfPByB2Hh0
M+qN5cZqjwkrL3qVbiF2mNf8tE0MSJBgspScpY9A6Z5nv6Oyrit7Qy+OOXaSuhVE
CfK868fVla89E8Cm91hz8tI7lehe2BGvmzXd6rMXlcfD3r0oCsf/0XjDD1CgMFSC
jPy99MuqjTw7gnyzBuzye5t+ZaYIlEDmX3l4Ca3xIFJy2dAgsL9L6oFeUIdpJ7A6
2S1JAmyLpMZ7XicmiOX8HAlsNSeF0kzGXTiMMHNxyhu5GUIueWLjtJYKtjMHRGMc
7J/d6IuRaoDGaeIdOfqi09RPDeceoLeUQAucqEbw3rVt0frsz1KMXe1D5JTKGXDp
18w0hHx/rk+Jh8OIjEkJX8mmyw0rCLtKJktSGNPj7yfeHWXPSWAsMDpUBLJbaX89
4pb4gM1VxET2gBY7WYqVDPCYUhhm5pC96kFwLNU1hFnNoKLe3b6WxrmoYVf/gdK6
Zk/jjA8nfsr2GtW3Tr/1Xs81BzSqpSQ/jAikyVVGyJr/VFwZBtI4Wbov56nlIrAo
FUhjDeoeJbuzrImBeJj6OxeZrqYrwyolR3cADwkJM7Q8FApsObQoFDd0jj04XH+v
2vnxy+9i2CDbhRnptW2QOH6yMdBmT8kvUfpnSIFee4ALxOJk4LMm24Uv8lDYt9i/
fYH1MEobc/YHWaxEd8i/okyoaXpjcuyATlzzwLpRmyU4PLJU81Kzj82R4fZJCDFJ
JtvO/bZpH3V+HDC0ao61YQxQ6M3VmP1ZvAnLgB8TndRqG0+NQQihSG7taaFlA8UN
8sbbM58FyTpL6qB2ar4jxp/BNu8wqpBnCNXXv+9wQosFrRuj8GX0uFEwvcaMr8Gi
CDL8cLWA3wx4lUDTcKC2kaPoVVgj6doc6RCg7jXl3Whk9sx9Eqh4UjxcPn+5V13y
rQFQ0/eUHCqeKY0EMAZouHbtaQeiodV7BKo8TFGeavEjkR4dMMCFLr0JiwpdZqrb
Mw/occYQ8HRFo087KIY1+ArhO6SJufzPwhaROiTcvCtd0OYjCyk6+E+BgZUuqPYc
A8Lgi4NXTBM/9u6ZxkQkwxdNVkxxqS/sCXDQqvEVYXDfwDLdyJFSX5wcGccgzY7Q
HS7xI59XjcT7B/MoIV5S0SXNwxYJvnA8+02aFW1JJLTBFlrD2l5IBGaQdEJyW5OG
2suU6qJWjDrLLTXHlSduer1caAMzGQrUe8lJcyicvg35kBeme6ziAHwOlT0ZiZaW
wwbw3IJMOSoSFnR6n/KxdflPuoMHJD+rEvIsApRazuAhkrJo9k9SWgMkRQfMl7M5
xYsWYSb44BdnQdMw7CC6r4Wgn2o6JBiPWNXJkrxtMKcnr/OLG1q1yOGe0Lvxx7Fl
WfK1dYmZ4cHGXgs8Yy7Vfbd8dWz6PteXZ0rokZGYA8mu3aR/sFph1SWJGpviD9PY
FeMwwROFhkXoggkwmPgfkffWOmn9EF7M4CFyJS0OMa08qE4CPheAn0gF0nAecFzn
1IMmOEbq3g7HY1839XKvek/KUaRWPYmbPourkzsW+acNmtsFozAam4fyD6H1LoNi
6nsdjP/chivPIoBf4EZWWIhnhHmynE0MsboH9t3VuNN/AkEXKAW8zoe+A49Hzx2t
CY+aWkL3JitbQxzSAsy2AR1wEpDAVJ6V5i2zyd3YlFP2JQ8L/i9GYv4FaGW7VnXZ
ZwOU+/Dt2rg99zZxwEr9B13M2/2BtTEPt9NulM91tjf//CucdfDo6J8nmFvygWCO
vF3OsyE8gyIWH7ClOGGjbPMbZBLjEguZxntjr0fUXPq47jYJRAGSn+xEwm4mfHrK
XSlxnkM39WC6MNEbE2fRPu/7JlsRF1ZHsFQOUQbaZuMuESwcufD4qHGySFzVhPd+
PTN5TiecTtrV/ETmpIHHbersXORG3B8ENmadyCG46C6SvVn4t/PzGJ+CKSsf44ib
MQJPguHFzTmh1hWO+iX9pjSutcEyBixEjqtQKsayeu0nhjqDJOKl0A7audFE4D0A
FIpbcwca0HLALuIpp/dvzz9R9u90msqrRFZ5XTZdAhNapWM9rYRjQC8RgQLEuMXZ
v4+dfaagFXeGhOTeRI251orx0M12oH7X6RpfTACkPGgQ8JV0AnJ/7mBXUS3awMOj
NeT6Q+Iiy+OTc+7VmNeXnh6alPL1DF8xgEoEb+tqyfUz15Qr0ddy4ZpatwOF9li+
Vz8cmOKwQm8dGpj6zSqt70t7d5lPZsjjcUslqoHM7d/8Jl1gsnu52fNanLZM5i+Y
irwmL6xitjrAXeEHWyFrlcKqEN65Ma7qw/isKzrQnYw1cedxQR7AM/hBW7P2XeN8
Uv4vr6KLrSISOnl7u3cNNM/gOGgLFtY1fwZpE/7ZWN4xP/lMNnqlhpuAo0npgH7w
lsDSRyEaEXXAFNdQHzghFBd3SQbg7Y32tYJ5X2F8srLPwEknq0n1uLhNH4zVQJjT
GuSYQdjdXnjECngJTslaBh6GqzlwL6ywlgj4qfrpjPiioHz2KkcLAilfOyzzqSez
s9/hnrtC2EkpLiexiE0xILoJrELJIcs3O26TAp9ki8fddBXnv0FCQ53gZ8vym6KJ
yjBMLCoO2ycL++pU6BXlRY6cG+jaYP3ua651GA6LHMxGROqW+O1WiLgMsBWq+nX9
qqrjM/rHIdiu8Kg4BDSZsKv2f12KU/qtZzbFdKlusZIc6foLcE2zrwRMlFZ6N/FN
85B3D/0y1496JyhNuzLL+aTCXDsgk1W+xiu1WjgudDsihkz4eYkAGkN/6gAiw6SR
uBdQWQZTxflqkKrax7zQVfCifGHEwSJmKwupSMZ58RFYH9xN/6x3ImgxQgHfU6Y3
+ClYcxMY21FgBMykMW0ISeW0+OlQtcNbWFXevBHQSJ22epNXw4InFCyHyhglvroN
aFBT0r9i8e8zG8mD57Qve4Sl4m1Tqj2u538UpUkTz6Tz4px+wjr/DPRpItt/PhjB
OxL9y5TKJ18IfzGMrXBd/o/1Pc46QEVe8aP8rNVsjFwxTuQW7lV0POGFCOmLhafY
jbF0PXL5E2R+fUP4hyF+dKiqwoH2eIEQ19mNPbBzNVXwwCMy6ENP5W9rDL2PbOOJ
p2+JCpoJvg26bxgN+4o1IHnIcTbj3xtizKbGECq0QPr0mXW6SnZT18EC4egnw1/h
vI6WRUs3XCGNV5GC85iogt84a+BeDJevijiSXverjVose4QPo/4OwTMVzEK8hFna
Nm7fGTPPfocDF7K6PPMZ13P2v6EF39gfx2Fs0MYBHRXIntYzWheH7+hzNIlCjAWF
lHN73+Dugp6B+aPDHjpKYqiwL9BnmEqfdeVf776RijogdYfBCArpExUr4D4rounz
NPNkfGC4vhI/deN57KlpwQ64ishal86gzfYPCXkFPTSRjwvw+K77R2qi1r/+lFd2
Zc2Ebh3R0MlCU3BfzJ4L2TJkB7Zv3Sbb3yynNL9YEKYoJ4MSo4UFUG9tKUjXdCTt
OSoJ32fKjyPj5s7yh9eT2wAMrbqYm6uWZ8wHsYkNbveOsmOraQxy2WTBtgGcnsNV
rST7bMLYfu8VJuh9dO+r4hKT9SX3MGaIu8T/97zk0+QVClDBF3WPo2Zdh65ponW9
FZgTEAuzpxlWnixIE8XSd71O07mPSwD40qPTYyG/AWd24ejOaWOARSZCMyMBa/LD
PKuHbSfQSNrmoH0UdkyLWRLGypvq9TRmzDG6p9cfMa6XTfFVLgQjBUYmJ3R2CZLd
Vq8tJgzhTAwwPl6ZBr55xSY4LFpD6l+LQgAzfKdhQCAhl3j5fACuL+4HDBP71OFe
WtI8DZXARD/LMTNThsgYWIiwY8/M0dWzLNzW1YucaJ/4tBsxdQUHG0uymZu58vG6
iFOXRVUvS3SaAoc9qqLCRdLp1zcS6pnxHHNRWoDJ1r/TChsNtDlSFoAo1s8LHuvS
Al3mjWVTPIWLe+c/EsFtRQySAIi9yQmtMmThYSQD6m2WB1QTrZl90AmZHt3y9fzS
1Nn8SPn8wZdLNLlBjLMXOI5q+btRDQII8ReOVq3SvbSto9n5fIVw44SoScV8pMza
UuW0+H5YsueusW/2Q4ncJoa3vtbwdYMycGnvBLpF8IAfnAQ52LaMbBetsk8SFSEz
+xFp3jqQdpNER0sdsMfMoAy1Uw25arhVWfdhER6KvSGOcnsiexvrt6iTJp8XR39T
PHlel7rAjDSQdOxUHrdKGF2YgwEmQa3k5k2uDRGhhYqo/pG4yJpJdCUB4jHl+cSe
IiIFzcFbElBhQj6I5boSBec5YuntBAz2k60YeGJk/yKH7W6sXHNX0tj7VSftiU2z
m07KcAOUsyBB3dltgpL0ck/+v2KxPNXiyhOAjI7f/F2j+qM497iU917s+moEUzMC
9vfnW9IbOmcnnwZ/vH807KFNziNcGyAB37vO5AHxCND/hd1mEEta8OkUm5SzzQ2y
Cljx4ECjqpLPVdLbpJv88D3BgogTQoDNOaJrKAfWb8nuNsqT+3NQuzmptl3Fwhn2
g9f5/rSZGcqnYEGjGH4U8Le2I0jdENWUQlcVXKEc4Imldi0/EP6S+vd/sgYlOpTW
ufG2t31bbL65aEqH+Ao3WVMJHQ4PPr3GthVypu5+hAhsxfrI6U+cZ8zQK52vYHlN
lKU5VRoBVRkLkqNXJVd29qWwAAXyCpZYvgK71FdzlbkcUfPY0056HnTMMyvwXJo4
IRZReQ4/PKEey0G8bFqXbcoCEcMvrPcJesXkL8yHGeyIeIPLGcS3Ksmqg2psbBUl
Tg/lc2yVtRT1MLEOivKNm9Bul90o5HF6Uq8BlVQOI8ynvkaQDS7mG3OMDJlg8cJM
orZYbnHUKwZnebcJRXfT//LZxjUkcVY4TA2KyUxpjf6y2s9pS39IklJyxYjK5Gg0
T+I8n9Auu2DH6EHlpRUTHzbuEUwcjGDZcnTvwS9/t14dtruBxJSKmUJp2F1aUcX1
469qb/n8pfPu1s8P0YhoDmMZn+Rn+pGRrfVLJkdqQ6RzwMomvDREXfsxn6ZUIXf4
Bj64DOWTE7AcBWrjGZ5aTg8l/mJlFnVdw1AZ/Y9C56duFyLb/uih0kP3ezLUEsvE
JCS2VitArdOViYWW4hwgvVeVv1JF0yIT73K0Mxu8Uofs1vS0KFUDW8R642Ki87Xa
n6jwZU/mkSo6zFyDSN0/hMuc1yT+6ZaA8/3lWFvBvoc/uLJSeFP8HHAvp/7NRefr
CWf6ZTH7llkc70KO6Rptt7SUQ7ZwPPFO2HCiOv9EABfHQZxCmxIMD/uk9YstaGXF
lNjV7tra05C9uKksIPnPFA/DuGHJmhvG8/+cc6FHfe6omw3OVOUhJvYS4AIX1f2V
Vo91mr2VOp4NIHUS7SRyDYj0+Q5/pHH1EgOIVFBczXtuh8F9+i7E5fM4mlDXKXtv
1MJhwHrpOY+khwtvA63eHDnyyBsF+byIEhA6wD0lHW86hharibA5LnaRaYmNjLtG
Ez4joaY727oCCrnZhQKO0dmKa3N8mi/VB7BAoNnXXI28A16ts+kMdCjMadUYwd8h
Vxi8Qes2KnXdhmCOK66bz06aUzOHbU5R/YaPMbyN+Ysp6kG3AoAz0paEsAUK+++F
yrw32uYIWewp4uUKbyDVMmwOZ3IJ4vZLPiMTSV6Sxe8makjm7YzP9ZP4d3mrd9hR
rHuV3dtYaNbw9DiQGMoanHSWFvlWRsxOru/oLlU4DhJIYlCBWK8AO+pcwtA5HQfj
YwYAOs7jx1QwhP+dHuPL3bmq9AFjih9m3s/w4uW/HxXZlQ0o3XQ72dfUhcU/DJrM
5eu0DdwbzJQ2EL+whC/oJHEmFXaP4bU9wtj8HD7LUvnTl971gtFZCZI3/2pYAYkB
CkGO63wCnJNi2q0DiltOf1I8cEPmhd/1lBuGabCfzyQwigk8IefUKWuD5tZqVj6Z
pVphMXj0DPOEIV8tdzYQwePBWGzzPOVOuPKHv4wFamKvwvk/djREWINSzFuuPPfi
NO21Mw7p7gb7qjmtmdUP7L8hr6TWlf1eixYqRkCyj8rUkgbQYMZxUJdOMXONnbI3
EwdGhlOyxSOUqKaBO5QxD4pl2+zbGMUiHfaNXc9gEb0dJgGzAaKWMQmIe5dIEadt
Wz5aO1xaCDvDfQv0SVSAo2w5cHoi/sGXUYLOxyyIKEX6fjYGstx56+PbdBVkX0yz
pWGrl1XHk0jLg2Z9DoMUQOcgWNWPIkCiEk2XGU4LW0VfAbfv4ZqgoUpTFju27EGp
sxPGetvU99925ojGTcQVfF+vkErdsbq3F5d/PkEI616hJaZgd0X2hUF2I9ahcUAY
ogNPsfko5C5n+qeb7j4lKCEWMgX0rcDDTxdy408LQuOISjiWxaQQqPkzYx0AGC0o
bNEEZudQgcw/z+JNRQJE4ebbK3Eigv6vDa4nW/xchVIVrPoxupj/AuP4lboXCrTd
QXV/tLzDuhVymU4jSRhqFiBblGpS1KhSXrp9QJ90iUgRk2M/JEut2tRPkHxjJXN3
+PHtStTXykjB1hEcM2k8ELbLUFNBKyzUrxomxPeLlbg6IXSbPAICkL2VBHyORKRx
hk2R2Xivg+KG1IP237Cc2Z/Pv7S1U0FgoHk3jMrpaBQprbIU3hYvlZCYy3RPpMKW
3APlcHnHCbucaqUDrTp2pEPRoxxckW4LunKOeqRsdjJuhgVPZQkZaApHEtKOPLKE
NhRoboP45VYlXwTtiYnXeB9WNzybGp6pJi8dgi2gYI4lyB17itBalIU30EvKV2Sr
PuYtiAwVp8zi8G9Y5FFCf/36tW81/b4VcXFFqCX1z/zavA0cmwwDD5D62uXxKnkA
kv63OdLe7GWki/e1SbmLYyPCYSBhhFgwZTayOD1VVlrnlNIUzjHiLUHiqRyy4ect
O/rraRh3t41XHMVKmS+OseeVciVWJMJHG6XkF6/PQjm0tOvCe8Zu9+FRJgM8sWjR
0VPFQheqc8+Ooxnjz0oF4aewkAGkxiaISKnCahhYG4PNW7Xmyz6+clHhhav4OF2Y
iS6wiPJFRfF29DRpZnptuyKJzU5kIryZW5BmjF4QBNPoreTnKG9za0JCKJ+wTKyv
YYQN9aDZkLbYVUqvMRhCVfUIUuXhDlgS+w7n76NAu6pB0U+Sc5f57KxJl8RWE5Wl
CDdG9z/QhPGBZEA/cckZQFhlWY5rhHIZO/yBZAnig03EqZ5PMwpH6K17Dl/NF/Zi
r03FR+QfRKGb/suns+t8kkJMsKtUOO175vcYTbE66gw19jBIf9/I6mjst4vnZDRj
tRDLyw9assjTglLQ5En0RUwd+7OvfFMZqytzp2Qrs51xz95GXk03POpwrit9Fwkj
NOmf2kEGCTZyE1y9mdRmjmeVR2zUHmJb10LU/tYWByKlxFy3TzqLKhbo2xjtz4uu
yB7Y8AFQn2QP545PEKAxp9t6/+VpSv3tSEpw1VrxPKUyKrctIjoj/rEAGDICu2fU
KGJtXZ2Ij1IozXw3+mUBcLUv7/1jOZt1VDhLgeHYdT1gamlQfAWvVqTwLUzgypG6
Sp7MWxzde5mpdu6P4mWBeDxy91JsDJ4L/vpJv+GfTjhsZ+ZV92CZIJdKo4cBk5Xf
YL9D1kUz3LDAQN2LrnXGYIKdSto4QBSwREOsA+kvnvP+RcgYE5nPEhbidG+0ltDz
SW8P+JJUUDdMtou318v2x/u7dOhaepm9vfqC6CtVeOzv1TWPPlEQgPXWk6TpwYmo
85efj53iG7hkt0MVzxyV0jovsOikT0yCBAO1eLPJ1IZz9aKoTyIKQijIKXtYikoP
xHn/9Ac1qfHjanMugUrap0gE8D2XyZh3N7IUtKMcBHzBojnj9cvbDIGEmXwye8PO
Wxia3H5+WOzB7mpvxcROEubr/57QiBVTTlguIJZ/GqFw0Y474GnqO35c/UL4eI58
Y/FZIhPqoUIRzZ++mSJfU45RRsJ9CXPD+w49zDX3ZG7DvCu6qjFNzqaZVwhYuMzM
fuKIZPziOzjP4DrPZAW+4bB+0V2p2VoTz7XgtErKFHKlFqcW9Moh7gY+R+OE/dcl
zE4WGTIKKp/CAeDMNnmBKn8TctbzA9i+HF/QupxKWEtInMQ0aeMr0vAifeVWWcjn
Xwg4LxzQ2M7YkPls4wjXtzFMvPOZj/QJNK8G0VqB7O3CV/e74aK8dMI6c0Fs/6u6
THglZemS54FV6uvRmsJlzLaEeGEnlzRn9CSeGhBYGSrdANIM9NMYIDoc+o+wohDu
FVB6TGMVoUilW2t3Uo0ZLj7uBMYw61MQMyV11ju3QIWxo0kTAkiTXLDEkomQ4hZM
QVXGykM6TBYrzW9FakLXjMxL3Dd68IfEc+sUvISLV9ZIg7dvr9hrnh6MNj+oOSVj
CWF9qKBerfS4dHWpaY4AKtxZcBkEE7ZXYWhCKfO5MEJ7kIKzqjWzAEb1gumImhFT
6in/trgGOWpAK56z14e8tF5ICVW2LbjfpxVU529LmfrZ2MnDK6gDhj8zbdrSgqbK
hsI+4SPdod1YUpq1F95LM3xqFJ14sdOJZU6Kc3cEd+FBCXFb9D1aWfPxP455GNio
isAmoJb6kpbsdq5RmAwP7eWPFyyfX2yd265RyDbO2pjGYWJqO/gfsh8LQVnQAiOy
4OAyuNQZhNiRXvQnVkvtnPi2gyG4dNfgUGjjjSdJDnkTi4nkX1wv71tWV13ah2ZA
XR6MJBN94iNp5QYLIA9FkbNZsrXbJtbZqk+BrVAR4NgnfGpX4HAWOt230SwoRHT9
cRAdZen9pCLalDQODCZt/l/kRoUxRSZsWxMdB0A2f9l9vZ+UwVC4jruaKWXo8fkO
x8NdZsZ7rilNM3/CH9ZCiWJgjp1ccrNend+73YGfnejAn99VZluM70SpDjGZIHpB
P/o2sNwLVDIIGEGgn69VaScWN6v2PZQPy+DX8xwJOfORr/IWLSE64dytPfDGiqSO
3w0YG/+u6JSMlG7wWbGKPd0CD2Sd0qQO8b+TU3SdZJOdx7G/IOLr4dvLvdG5kiPC
F8tmKdU4nHp+dofscsmFhk2rBqzAIVL6l/z6j9Lonf2Sfq913a66PFYAeJ0H44DV
R44xx5N3G33ZpxQ8boclkvVnoS+mgbKh1Z5CVPMqJgPUNKGVdeF81PFzENqjUwYa
D5QklpkAn9ZykAgmdZPtCnyTXszmumejGy2CFZEmsX/5hTXA7xrMjvFu1ebt8jcl
uG5hV9pdRyFV/g15kJ8pYxj2pCi9smUr88VZUr5vgr+4b0xjrDxcy1/C/ASu4Zsq
+gvddwSGMrEc8BIZKrdXR4nemzYGeKIcxU6nR+DW/B9lmK7dq5dJifKYu+c+bVcQ
20tA7yWJplg3XkzWXtJUujYoX8jGp2/xCOd7lac3v3F50ImUONXpQAXRWKQEwjUE
2Dm6r5jSwZBQDqG274hAkWDg/gTkdeXddTlWaxW737yfVAlPucbWHP23z8eIqNh9
9gdWhvjWeLwetJ7sybtHHR1Phzu52TVaxVfvJzGyAPjzJOX2AL1mW86RpktNQyJe
zk9SABEfzFiZe8lnV8otFA5dWKnYCZaTpzzB/6d5V2uBQxzs3yXj28Fstn7rQC3l
rJVifF57XKdbAvDKE5AYrwZnCqrN6VewS/eGKSerB9Evuy2zfl6vT/qlp6MJqLFV
69MI/rBeFAmt3YwbVVaxbPdQZuEqPbsNpGwve9+8DkSJxOzR7m7BNpFaFdXy3xhf
RZ/NkBMRBol/eKIS0aR8NbGfqdONVCvW62HfTAaTdzy42d6IjVTZ1pBz70qw3+eb
IQlYqGTNc1E6buG2Wr8NSanlSkR/dU4VDVxI1Xf8IZW9A3AADrnK3610ntIBl31g
rkhZIvA8NzHoB2S7OEpiYCydbj+E1oed2vyBQDnJCNxJ5SArbqQudblzfEbbtFYF
Gnj+BighNRW9Msz2LmcbcwaicFzzdnWnyH1PWvprVk+af/h9CTenrpdf/2tVhnmE
fwnHzT1pvlMdJ5v709Pdq2GFNQl4qWWp2dHGy65opnKGVOxkESjnyAEraAb2a72c
rYs/VPCBtMPGtlWJwcuzPVhNZhZJZQhLiHBM2FgqqWbqfy73NDyemIz8TTGJbNEg
hv1mq589pkKxtxk5HDZ0q5iBOApfV/y1iBoYfpZOnM23rHmzX0o1H4op0mjFFt4L
ibwbKVSpEtTR+0o7nkwqzHaKRX/aQBCmovF6l4Adv8hrusRtdz6OqYxZewkP+0ky
IoiRZASiuyE2dFS1CAG5f2TwzgWGkY0tpKGB3y1wBl7xjgrzx1XkLLQhInjuK6BE
pDKC6asJhtZ6TcFQeWu0U3qnBC7fzTawCm4ajUkX9hv+Rvc+tejmeALjLJWQ+KUl
BgJynhXWNlTlGmPwVxyj4vB13AmCY36pvgNzL1qOryT3kM5WtoJ9i92wcbniNiqa
WxRH2P+NDtVsAY+GAUAWKUHBaZkROjGhUp9z0iTCduv4UUyIm9JRQv5HR/rHCIwj
uqVqOgTQ997NSku/ItQJ3Y+AiuIbskQKEUb+7P4HT0X2bchshDB0UXCB2qWTO1Tt
CDjHqa7gLXgj/S78ja+T/jQPahh/0bbTEyvbTqCh5Tb1tF8Dsja7dafksrrSM332
k9xu+3ZmGF4QrN3mBvRY8/4aat+ou/wzRrkWRyVGyM14Wlh2IyvFtAOrP+tpCzi8
hToeinDGCfTu9+l19CAVp1OTrH0lWtzN6xizitOhSYuXCeaK6Hk1vdnqipRHI5xl
5sJSwjBaOY+r1ciTOtV+QzT55I8aXf/3zqYEqG+IeoPnUaVxRVFl9Q8MqmVjJO8u
eqAmrpvdIYglAju+Mww0Lr6hUpoH7mKki6O/qpfTnaC6N4B7PKLRa9DDcs3R3+s6
T+F4E/2dmURG8ANZloATKcj2cGeVkMgv+IniqEFACeZXLul6Cg6rsI7tnwH5W+DR
nv5408W2m1TyBiNs0Yd5LB0DaoHGjooOeOQkaavXaNc/QwsZ/XsSNNJFJvaPk8qa
WPV1NefOARBLPKBa1e9SvJjV7pyc1LB1Amt1tNQPrzbsIBEL8m4BL6ZOjt4+fPhL
spYQc68WDzWw595dL0bvAFT8wtAb6bswVzOUiDPkbd/FpC5x5QV4UJshmFo+2XAi
PbUgfjLvzoAFdFBqStpX1VELaSSKKMOy5vHPBQkai1d31VT6JSLQxvBtd0bxaj40
oc77u0x+AvqHToRtBPDWgKk1ofUsFCckVWSfKGPeAy7LSmXCGPPlR2NC9mizDUPz
9n7cqPwioa/SUrAHAs3U24I+7F1aoe9KIyfBBauxTIsMwtowEME4uDUa2Bzkeqeh
p5GiWFQIS22U3/QPmOqtmx8kzvylMoqLY7MsuOFqginKLYmcG2KBTU2jNMubRkry
ymW+CggU2UQ2iKsVeo2/CyuErC3U54C7FgGxmhx2GFGeGLHp9qHrvTiu5XwB66XB
jSRFtZFykO1JPbP/Z2Ng9OYwML+vk4vm72k2P9Db+38Hzumfw/SA+RgHcBbZK1oA
o3ZfkO3Z0NJc0aUpThwUBTcmgX66a28OlxFr6WlQ3xtF/eoGQ0CcgB1oEPrVSjBO
GRMS+7TlpJizRw+xh8syCQADfdp4wr++fUhDOyTMKVOfbETC2fYJXq+Eif0aQZuC
j6b/0/CTA6dmIgFGpLLI5kWzvppMHoPxyl+MV91Z6qDWJrkl4DP0sx0D8un856bc
9r+y9llTOEyxn4oLUhZAzV0D9ugVtygrtWhsYy9ZH8UmCCirw+Jy4TUTmZK9QTbs
JUSXXUN5kyMjXLqo0nfnC0j/tn9U4Qb8605Z17Ck2yFcU6pB6o9So6RUNwEyalpx
piKu9YEK6UO5oEXt2+eKtkoecDR7uOYrMwiN++/AsoJ2stO1nluJgYxz1/CP4/+u
92EFi0ljX+hzL3azx2aLCrc7djusyDfwNISExh2nHK5geRmdUt3z9sZevP0lXAIw
br+/0eTzDcT0vAfSXGfPmY+ZJuqRAyvdA/Ie8VNxMTZfqQbkD2uy0XdkQS6N9W4o
GxxSrdx6Z3zcXzfPX2gv2qoAC+BDkabdV+QASDIkr4lPHQTbIpxA4ws6EkxS99Ig
tpKjcVIVSyWcjl6E81S/7t4HFWwYmIcu7PZnSw0shko5dCbcmsaQzuSdbBf0V6mo
e7zTMVDBrjPifcknJMXhb4G0MDJak91vraizaZH/WRSt85BSkel5XAuirX9clu/2
CipMj+mavkvWE7qyg/HsMqYJoqpQwk1FWUlRmYFGOGDrDvJnR+FbO9dnBbVZf3Kb
fB/WDrQDqmGXpUv5o2nwlYJRPQ2/JJFw0PCt+bXiVuMFsbh3zuUejJulWXgLKu1H
+Vbimi69gYA7xScIGOU9bH7sOVOpSIHZL60seXj1A5AeuxdZfaEXOp9j8tBDBs/k
xqQ2+EXmjAG4RhaM4X/dAuQ6N35/PTPIc5fnNIxTjrBU6aIVgGhcF2WU7lhySFS3
s68zI8JjlNF2N++YwCfzyKudltVoeGx+xB6+ox3RlsPzXD/nHTesuI04Hc3bPDy2
d7I5YZB1U+CyZ+2z4pECJY4fKmJcDwYqMC5dtVqNcSJhqueB2RaGm3eK8HuinCW0
5lhaGiiupTK89KK28n+IDBiC22Y1+bJx602wfn6y6QywCI9X0TaA+mGlhvQLzgff
uS8LaWrny8NVLImdRieXNkt/tX7tmE5MfEGw5KbJ9WT0MwyaQCeaWGaMBL5hk8gK
bVr2u2XPTwvNRinHk4BFAG0cwrrIrnpsagB6o7ntqb20nDvYziWT3Thy/IjAPKIb
K7OgVUnZ2ggrmD0xRoQ0lxzX+xWRGho67/2Bzrr3MqHJPPrYHKociPBA96M1fmuo
yMJTDA7epPxazj7p++H5wvLKJjXPD3gfbcEgCJmkcdOJPrl0tQpwkEVy9ctwYl8Z
OduNOmubByeHII8GgNLL0mD/Y4ar48fNKeqnRbKpXPlC28WCSIpsJLA4p3BnToHc
YsCTfS5CaAToeTmtl02ntaZHL4YYWuakMTmhuWUfz18VYKCc4F/vcofVF5qhGokw
wRob8C1iX4AJUqboEHV19XNR/jSiTFr1+bbukpFDc/nQ3U9iPcpottuMT293Pn53
CRJS5X/wjOuY4exhIpU1fA7RdkCr9LpLGSX0nfLACSSHGAyl3fzaJlEWQzQuhlas
kbqbV5IvlCWlTy0cC1FAWCIkuMLvQO5jLBQaQimHgu3dfRpyoVoo+prjqIkPWoQQ
/EP99Tp6VtB2M8BCYU1SuJU0ubPsiqJfiUjtB6xMy1JDFXFJnYAn2gDfXNFsc2tG
cvJtgNoKgpt81vNX00wkFtPKcbOA4mo0CmFSSIbliuB566TsDGvH66fEHEixJHvz
JAIzGov7tn6r2+Zy5Ab33arBJdKx3Wn4nMAYvunHRyLfwx6cbgG/IWcCefZR18Oq
K4KKbffjbVNZ7Bg4mdA3yQ6D8UGK1kNQOC63Gs4prYsfOn+1XitL5I3ZzEROVQGE
yYePLbIvtQSmqpw+66m0P4hiD31HWkLiK7ZIX9Aek2YDgiAx0MU1WKfx5AwwqI/s
IaXILOJ9euI/99IMawHedMv3R8+kOYzqD46nnI6XOOAfibveTmTtXF9XT+H+Axns
s4TpGbgi3IHVU+k+WJQ8tTZyADizAU8jDKpg+FmBAWldQ2fAiO01PUI55mYth0Uv
t7B7+48bI0AJdlYYwFYOVed0lhFh3bi3o0g4dj40ZUNtxcrf+AfpgpZtyPSbampB
kzFh/eqidxkhr3xUojzUiEOWDUj5F0xAz5q7HU7aMtKDb+8ls2n3F24QPIwMqG8l
9yY+YWVqY6hKJAYDbgGPhNWUwJZTmXwgFXGu9WDb2Mc2vZTmrQWxqQ95WohvHuEV
fwNJ0l6ZlnlgpO+RSyXJ8JYI2UbswbqrutDKj+AfAB5sx7kvavCX1xfeuvJZlwYV
scUR7RnlM8Pta1hIoKyVWiOrndo+SSL01B3BHf6lhQ3CN+vFPxR13JUaWs0kQPNi
HX5/DZt6EVMS7D2cDXHyXmzOEa95b1xKoRuauwbl4khEiCYOFC0EF1TFTYEd44sg
eZdLEgOtdidIA464r+DeIYQ8QLUbaIisXwLF+77OVvh97KS3UN7ZvFA4LTB1N9+w
cAGgxX+rP6ViKgXAafT6Cm46byd2eoecrqB9Gxzs4VFaqwbAGq5qi1LNk2pRauY7
BbO4BpR25d+K67Rn8KAzWymC+087uSl4e6yt1HujNjf3kxShF4OV6cY2B1u9IAan
lGks0XBp2yRN2dU9FRYSUDPSpQ1MF2aQNP+qGi/kMQUgvpOA6gcDZxIFrzkRKPRo
K6tUBqcriiR5uUo0RkLrAL9IgDube4TeA+QtgX+S1DqeLsOxQwrUhPR4AjFxd9ri
4Z2HUpM4snKnDGrIS2kt2wgNES8d+n4f4/JaWC83DBOzLvtQcJh54LTs6pBdYvdM
F5tLSUULzdL1pcU8cn/84BrSemqqr13AuNsEsmPZ/1R1GHf2f/DjBLDRjYVZxKSo
i2/fNvat/bhNKSfGsW0DaakzqWN+FfiYXRSp1IH4ZFD5k0ah044woj3cxE8H5ta/
i+TTr59cqUThz8WplEkFRBE4qHsGbHgavtsAIlWC8erecL9wq39LlC+bsJ6rS4Iv
tn+dX6neJVO9JyD4uSG6JxmAT4ODHyTxHg1BhPmvFopFKEvYMQkEfmHh1TdRatgq
PxZK7Dtis9xorKHJBBKygw30DgMH9xm1VFOQPrc64Qe8m7Bwc9S95+aCqVnmE5Sl
+8q/Zul/kahDnugsJHdpCD4N5SWZ/fTWNsX9NfspgYunjdLKrzM5knc84fYJGdO1
Nce5I9FBWgqeXd5vMGapfPmGKPCwjwBlLik/KmpA0N7+cAbDUrWY5je4qbJX0C/b
pCfl6wfNmDvuOiUakRKYiSWcbv+ReUZiJ3ukXfUVCWKVWqIHU0Bwabju+0ditxcM
hU5yWvg+Jt+Gt+mO1a6euHfroxY5biUxzYukBxtBozFrPPmywcXnZYyop7QJ+w9S
2BIYwYa78DmXKo6Rzl15ObrgmWzmoTFAsVoj+8ziZB4Yr/0ZRk29Mza3gJdo7GWd
LdwisbPW4BeZz4n4gEJ8LPpw6R34fiHYvYX0xt8Z6DgvuuKVFCh98wb4Mhpft2nS
Yh5dCwUoTd+72jArm9ROgDa1oZuTIjCaTFc8dSVGn3E9cBneHHCcEoxgYDkdP2Cl
SHbBgXT9mC91q8t5U3UjfAkW9d/NbercujHLm+jfaH1x4cSsucufpatdRxVnPWy2
FwS7Y7LuffasU41jiz/3mViWyWyWnEYxOWvNzvIHJFUv4MoZerT2IH0DZQ2opfir
5xNMpusKIbxOniQCBwH18Da4qtz4+5Yac83taaUSoFe0kfWUxPwcMd4Ub/fnS0Bt
Ry1jhlDb0Y4tB7lpYoZPCsxcmGI588Z8R/jhyODBwcgFLV/8pftDYc1qrcZ8VDjo
LTG4CYJRBFeVOPUi3z8PndMoghroARNMp20gqzW9QHZ38+0Gx+pWUrIpPjTseHLM
SwllpLi8nyRel29xnNPAaVLSkLekPa6pT/BUqU0UYTNWdOuIA5iSm+nZPYEwWoVa
53sCXqGbDbXkl3wrFipE7NNEDHCSi/TSqfvwaGzvQuzy4wIkCOI0g/EwlN02Si1k
/J/MeyI9G0cCoWBi28eYkYreaevPY70+7XsaCc9GUsk7XVkQ071swzrQ+bTZp9ZC
Y94PJiatGM6ZDe2WPkadprl5aL4pr4bKdZqZZIguVMnhwmW54NRg7XXfMtEWV8XM
AeT+PRuDFbs/varF2L7wtHDK3+t2nfXTTMVGipHVO77axzSOEiuP1GKXpRITsPyX
/PvzxcMS35gzK5BC4jn80PsMRHdsjVrP3rS/Do7n1YdfDQJcgh/JKO0NDEk7i0ox
hwQB13BD8j0T8Jg3wbQnjAg89tVQsFFCac3SxkMnPobNOXxuVPy2t97Grs0SxuiL
iVb6Ier70UIDS1/sJqArpu86Xww6OZasMQtHHuNpGuw/6hIcc7hiCsUqhjRxXpBq
pZ2ufBMJFct/vHPTh2m00T2HmRbtlDGnrjlFSgMntQopzHpd0yE0OF2SXyGlhd2t
WP/m5QzsM+ka0yOGS7ICS/pnMnJXWxx2jf1rnbRG+rLxE4LhfcjIvgKLGVUwn/d+
dxtBQLJIyyyZBVMyVZmrVzAyZbflUS/JkYI9bpAkLNfl+844LymO+SilsdJvbSGO
9Y0LCRrfarUQvR6mpfEm49xGUjBOyTGvRjZM5xipShN+C/4jtqmVZ/lXGP8yWFj8
s5Ze3GlFkpRGZgDaNKVgykrJzwbxu0KS4oxxXGS1Hr/MbKdkfMp5XM+nwpaDqJyV
woHzocQSBw8riJ7uPVUs2RoB+cLA6pveQQEB7GHwlA+uIruf54Au1iZipSX8M06V
vaEd/SqFT0CujeU19KErt3bjDgFxyCV+Ey26rvvsF3huRZDIyj9tNKOEoBk0sK+v
//H4g66MZJAwpUFTOvd+Ue1rv7f6Y0F8peuc2drE4jq9gYBV0LLzYZg5Zev2TPnc
Xu2zHUrm8b7irSK4quXEe4Kf6/hx44reIiUWB/k6atdGkBwHSDGob0wDCYYbdLh4
xAwYOYtvuFOqZFhgvmezBVGkIUL+SlIMgu31j7KM/hA8gbx4pDr8Z28aAYwC7Duj
eUmnecdpJW45RSNdG57AiqxO2irSImA6/2PxHn5sdhKpba56wjhCJJTXlm8kodBI
t31M6qOCurup+dSwmWWTnA3jquLgoCnYDJg699RrSV24gtGoVqqhDkkN9VcYj2YR
1AFIYooOPyArYVnYuhiD74j2lP0FHz2lch3eAEobqBU48+pJqbNAIuQnDfPULUwQ
YBf/7MUhCAwlVPFurDM1JRg48aGilS/FKpuG3UFBEX7hc0vGBKqbrUCamdr0OoVP
ODAurbbJ9BoIdsmKYcuQD7CowgSJml33y7k9w08TX/ZGsi8drIk88aHfPGMnB95Y
XTg8CEmkBebQTWfzwk4O0t84xDcpH57z0np1sccYB6WVtlIgzGLCM0a7HoxYuAEQ
0PzxyVwPJ+irW/WzaSQZrA+k9OaF5OA2rn5/hpAjSZEZmzN+JnUee9k8OCS4WwXg
XU26venlD/LOUWs0DyYPZaJaEtQ92YR9GUNW4nekuOwyVq/9O8zfLFJSwU7NzNrs
w0q3P7K55Z+fGf+Ey/jnHGnF3puXZRIhrioPs/qvFdyiMsYtK1P4pn5p70aK0FiX
33QR5aTcmLm/D1Ks/3gfzqDLKHmnFYh/QnJdLfKUzZG5vr+CV/wXfXnGb012TNVK
leBD156Z8yUcz46jjg6g98S6//rL22B8cq9rw0cBCrz4Srslg4LRXuMK2RmldPw9
GWEghZ0Xr+RgYN9OrffDqYj0vFwY+y49ntPXPF4skdC0xHr5obfTaddfk4HPCEuu
qzz3BGUbv7DvEcnDyJWfM5ITdRLnGOW26uckc5dJLdyQ/hajZt3aygnE8A8EXXOP
uv5EUKbwGLfbsBgZwDxmqHG8U08HllZwfFXOShhTcR+N9R5DzS0QsJF/VG8Cm+V2
FDaGaMIzFip7M+uGQOkEIre6mI9tTrInbSwEVc3I4NsYpZJQr1JWMntgUC0Oebd0
E3UPkSAjpnfEDj3V/Hqa3rNujJQB8+aL9+lyiihLUkJ4KzA6GnMKXbfadOMFIUfW
Il+pC52Z+h/TRZD3oVaxAj1BCoOnPP6TiTzP+LCKUhyyC11z00FQsaoVnQagDSIj
Rs2MapdhePqCyKqyvqxJtktZl/EUjzvpRiZv/Sktrq6U1xUkkbwuTWbKNUcatS4a
h8ovDkO1N3UFv9hL2GREmEo37XPFunYh/CvVqxYIgjU2JMYY9P2qvzZtmCW2Okh1
fk9WfwfA7vo6PwYw2A3fn3NdVS/fLYts1fEWxN3RamnHVpQlyFC6ikTLuMbTXMhl
bJwXfnJQmgIFQgrBLnx3eSGdvltoX0V3q4onJrkfVBV9jZNg2RzYNLD4tsXruEVD
WWpaBwfByPmWxvGkG6Iou6Twwnx+B6bJHTmy8PaGNzp61vBke+ec1rymykfo/oEY
3Lil3OShrn0gAcKMzGjQw9u8OXh0dCeOenQ1T35Ke/6AybkT1xOiZogoD2O6d3dP
qRx3AFjHMjKX5wzyGKfrHau193HwbkbihoJtcVHeqgVUBmClJcq0Pv4S9S7ZEyqn
d8cRlzHH+HLs83vcl7jwPbF5/qRSeN1MjLyK+ATiVMeqdINom1SjC1+ye+2UliWj
88YgG23kxJo0xhgoGY0m3WiwISHi499olQvFeShHwsJ5ARN92QEkXmo+hrrjaBMC
8jGGP69kTVPBOpn1rRYL0u9aTXZT+MJFTYqCGAzhX1XGqObV3wF+UE5hslpnbA0p
3yZBMGF5zaunYCj8Uf+MsAOmY5GwchEjLO2etI2FDwRVO25CkVt7E41hkETuOHmo
M+FpocshERQBAa30ouIwwImKkwzTJGIF2Wb9xZKHSypMmzLLA2lK6EYzad51+PDK
uSj6tfQD/oz8DH9/J/4E5TkRqHrUUBvRCI5s0o2LRGaB1Q2c1VnHHGYV3ArMgRzQ
xSVLoC332VI7TaVPQwEcN5+6yXdTzLJhYKCb/WjOJUIOklEZ/ACraeiUK+Gjihdh
4DGqxKQPhUzfF1y6sDCiZYf1+Yh8Dl/5UyYq1w1GmpjpHspLBoRQEsOAHnDaS5Cq
ZflWvG+S/P7PJA+Tx4j0wuEL//uRv2237XqRr8hGCh6E6JusZqS+izIcV38G1zBW
Qu0ZCH4ZOsg3kkXClITRz2JZ/iD630wABmX6f3fWMWf0xppKHfZNIqvnpXjdZdRQ
O4whLtnUaiSyVPr08dDGGPjJdd7j9+5gsYhZqqXyJ4KHSBPfKW2xfjGRKNYwBZrN
62LV3bwUlBGwz7vKuGJTIzreklpjaGbjtUBF1ZStBD3yPkA3Zjj66ryXUiN0jhps
hZ48U5PbgQGe3X2aZHxsQYdZiT4ka0+zrKwXO4Ei6D9a/KcTabKjOa5S5R+Wq3M5
ziPhDzllE4oVb+kjLvi507+Gkj6Hrh+hSl/+hE/s7oDzzxliyyb24QO8bcvPxAAS
1x9xHxHoZj8vvxMk1E/lnZjPyydkd+SEMsQHUk9TyphCgren/HD0q/eRyvgIYMQt
MGB9j4MJOmSyman2c204mWawiINJbBXLv8OsNqjuZ1y0JAKKNK+e48iZFrEGcljF
5/ETUn+GYDgPGJFbISkSjd+y0noqJCvMXOP9ZhvFU7AArYphaGVPlDmcPnlYMRLj
Kd3ACzrXRNvm26c2KnxW5yQmq6pZchMekv6SEh8Nd396bXr/QS08VpLWaTSbwIJa
78+OypoY5WImaqEfN8FkjvKiW/uSvhVfWHJgujMnw4BqEa/3jf5mOOCM/0EmP3Sz
aoLMR+BrzNhODaBPEmSkmKDP63jmUt13LlP8hwVZ2+nCHLRbAuw8UbbIJ6sBpf8R
6ZMJdh1ecZcLx6izF/O6HO2Dyb9wZ7O0Ta6qPeXDO+36Z42DiCGsLi9wBKzbdq6l
WeRGILNNn8kb74c7oO+NrdGCE/O5taBKcstGXVz4mer7rp4V8r5GvqzeMj8k6hiO
drEqLEZZU7RvpgJRApqidWQ7cfYoxMHTs02pCIx5DwwyXIEyVz8pIJnD99igIAm5
P6jUbsFeXfwPep5iwpBnWULqy1s0uHICwP+VwXYqXpRx6unhFfGP5oLEtjVmHDor
TIJFEaPpZa/iynTPFXCyoi03f25aFJTMN2NAFw+Q5tnB933VtAbbyUVjWcOREkCC
SNku4Xww4yA0rEKk8zzXM2bin/VDLRyCHi4hhbgR+B2VlQb5r31DRsvIwIkSogE3
xlA+wIjFbwuOCs72H0c4j6dMD42lfafpm6x9AeHa5Aev5LSy+7P0pXFiWULwuNA7
f0UkqliGhtei6T3l/PBjtnbN8EwC8YM7QzEUBL9Hr11C4ZRyV3iH+bzKT8Sr5ESi
WOrBjTrmF3ztI4DwpFK2vcIYXun0mSN7uWCI4mdJtMvMhjANkwu5E9vnSSeSYW9M
VmRzqZ+Zz6DX1tz3lQJNVcy7W+JU83ZOP9duEayWCefAUCqAZAPWQMGkDI+t40XB
H3mn70iiOzjzJnXK1ufGyhpVPXZnnPPkR8kbHup7DS5iM/i8zzam55tZLF2b8avl
ZOS6TdcBp8G0z6emZGbsY/bSdKWHG9Nd+dygLUXQ6lSGnQ4SQOurQDSjg5xqn+2M
hp4T5HMohEf3bsE2VHlWVBqMZ6yNbraiMazPL2sR0ju9yye6abqJG2UXHjg0ygOH
R7KiEgjJdu84o0fxGZpWu3Ru4KK6diVrNuX8gaRGNuaHsREe1U7Wv3C/KZYzAMVq
pACQt+sv3Dub34xsHNompSPqo6jOwxCd0aHhfKOJOmUqJWjyppBDhaJp6HThLc72
E0TOLehGSwOZxqYFX7l0PgUCXa0uSbcqSGiXez0Tix+eXKdQmWgStZZdhpUSMNBA
W3J03U86rwfPDdhgaNgmtHPyqIK5oZBXUVrUw8SKaBMx3D7OlYD4V/wik2BAII3I
BBJ7yfJNbFUnm9kmY991+J1pfl/2p8+3oXWkrwzbCX/NSMzedqyhRmmkLmBbC1qU
t4KqkP5j7Mu9SmZYzKpNrMfNhszOyhqFCYkVnizu9qn3ZSaBFfzhxDgeBV2bKhMi
wu65y/XM2U4xkN5gvZl6FcQVSykYR7Icb9dMVB8CQALSjOoDUHvytz5GDgkWaTsG
UU58egvuY7zBaxfvJCQojAnZpKK7O23USeihNdFMYmk2uToqKkwsqLHnTMd8dpuB
UlYaZ5hD/K9hue/QY1UJZ5cVL8XSr23DCDZl7LbgAgKqn6dGN9QazHrQMV84OBHc
9njX6rG0dnyxZh+3tt6ZXjLjBSKvOnwbjbRpGIus5dnU5JZEJ/shPkeAoJ8reRKu
rK8hRq3SDIn/2JNDD5E1LRDYBoGuJpTGwId1NSnavdjNRjbLTK4jug7Pnb6A9E5K
I7cbU5XP5qt77bZiA9woZkKXNf2QCrlXvX0qWqGN0ItQvBetA5CmAuqHbqBEdftF
rl/ueZV4LBE2vzVZBOYLFYXV/fn4h/qU4k1dYp0rbJ+MRZ1ptuLBSkuXJpYPGdDs
dE0EfRa3JU1TnUxxOoQyrhdQlvw+xRIxJ/Gc23mooSmOf6QScb4EBDfNA3UNBurn
F48wDTf5TD6c5NBOBRGOOvOJJH8Tf9nYiUC0RVLyBZWciTIn+V+RuhnPJBzKaRYj
/U3zSpLZK+k37T+d1gniFcEmaMLOf/BaXeI0fswgpY3ZNv5zvNM1AlmYDAJbwLDY
xThmjHjVQpcdfYxsmD4ZbNLqETCpIDQWJic/+j8ihDfWHetJ1A5rHGJmnwZMSUW0
hQspXK0dxUk+RpQCyR+l2cYICNO8VRqMHayisEM8qS/d790zgwUhKKD6xfjpCSPQ
XekZJRCTLod9LYDk/t4cX+ZgHjCp1JnGgghcPA4ajwAYPV2ALfVe8xm9ANi54QZj
cXIHosszClbCP4VEjtYRB4gM+VPDbapo/ALABl5ciYi895mZMjW7XsRYQ8qk1Gcf
F37NRsORveYK51FPIeeVuUCnpm4bYyqF5hSQFzcMErgDhkGcdapHT58S6YQyi1X0
bR80EAB17Zotui6Y/nAjx3XANXvEkJWo+4jblnd/COPoxLUYGQzrvczM4o3vitnO
2A+U92NT2oz2VRuOm4KrmbHx5fGIrvibtiQvS7HrRmnENaDD9RgPxQ238sgvfJ3f
U/oRNuxUZJ43BA2V80vC4OLEbQSarfLrwUaEO8ejO+Gcn/p90Ga6YYjAhTxVRxf8
JAGZWpqfS0HYPfVuWWhH9AF5E+/99ZakGXRAR3mZ5fbDaCfvihQL6NvE8aX+FACn
mQOXgF1Iwleffvl2HKTkrvVATHvyBEuSRcc6ysmxBr0tpNpNi34yf0DqSCnamsbf
ny/FSt0AyM7OGhdhudTXtPIqVwjw0Gw+FvRCW+qAWaj6uRuP2dcWnHZiGbakycCs
9A6J4Yl0rzAjfLDPZitMN2hPMhGddSAeGQ17QdefQSqBoqVhrcwvL0/+gLkazZFk
k1iapj4YZ89Ttpdzjd6WRLWoEjbjZJpVbsL3ldadRrSXCq/dkxuZr/a4L6e3UInY
CSYnqjVe+eJfRjufiGIcMHr0J1w6fLBq4kzHX7JN/iwAi+avrRUyd5HIQyWpu9sO
PW82KifSK9e8h6/rwrxLxZUQGq7i6Ary80q0XLbX9dmqm3SiJ+Z5El6Pd776cOIl
/h3oCUqkv5YpJys33RUgBhtU1uI2xqx1Lcwm+2e3vzASwseb1k3qWGswVnUEj+zA
NgZFqmizod9LBIiViRZ8VvwPAaUThmjlN4JtNsYaWW79uqyGKZqQImVI7t8a8md2
PZrOpFhKg3pYUdHnzmQxyeDRngMMQ7uYtg8qBvSmvjMf3/RV2x0FHxkt6c/iVUNU
7GvslrFe9soGbVMrVkZPfHeI2/Pob6S8xumgXKRiw7Dvgdplz/7Qkfb7bS2+CnwJ
uFI0i2DICmCA3yHnNwwwnon4Zx1lllP/65vqgV+RZMmZov62LfKLoF5Dj7Q/ZRXD
IBasaSqFtrXUIZsjoQdtWVFP/NFven8LENniFI4scj+bgaEr65jrpq+p+kYdIzg0
ck4dUzD5dAHdvAB51Im+MWN9k8NhkdCkkN8ELXfdwPqtyYiyfQoSDE6E6MU+79Bp
gpaXHxNML2VGfy/UUQ8w/isnOO0JobLyL3yHLaHA0pWTWyDJ04tO64RGJP1wS+oa
+EBEgKqQuVYLfcOY0l8wvhrCCTwV5FCYotEhVyVClTeNxOGwpfxFP4RLX7XAl/i1
3t6O2cvagfxfvpsptxCxUF4Onk7HA1kW4lpNSi0lc8lSIQmdsf30mAm8GmL9nUmJ
oLZgp5uSM+V2nmYpQFajOhp5h7NuFuvT4ANccMA0tYGgCzJ7lkWFfIaJX/E6G3t8
6SfRriwuw2WZZNnYDMOcAUFvqd0/PTxjKIZZWU2GqPLFl/Ik5tA6Tvga+8+1Msk4
k/YnndKcMF7x5ZYkGEP4ELB9GyPpzuY/kkC+q3Qo2uGXPBGFHpdDbBTihtxEmLFk
M16I69a7P3GDgVxBmDxpIfeiWQj/zLC117acQPJG+TiS9qdJpWVXs6QVqmgCOI5l
0Dx6OvE90+M1BEKiXWBkEu/b50a3tdcJh0S/rzsIdhxraP0evYlICo7GIw5R62GY
WtF1prFsmk8FbV8pcR2uJdu4gEZp8xGgWKnEA5f98vLd9XIP/iWDYefYIKC3IS9Q
HhFXAkkChDGQ1BMuZf6WtJrU2XScXVEy9OwnM32r9JmOTTDOebbMT/tCMRPDowVV
GshXd6YQv/gSYUKAGMQfNxqvabQPfiTQo6JpILg4LknFvQWFIoOeVsULebOwsBAZ
xm+9g9eowmKAbgxncmXW7f7nrcJ/O7V3dnlcmueHfnQCwJkynUX6xuXwhAvOsN0G
C9r/7d1lOIPB2UMhrOCpzxJKYw9dD5H0y98OW/KTrjXh6KaLQKuXxocB0eB4XX5I
37J/mV2trsJoaHhE0bS3meqvOjLCrZRvtMGubS2w+35gXNLlzEYcYaaTq/065heO
PP3fZ9nlCXandAVO5IbxIrDt6/Rs+7w64vgucEzONgtVRSOWMUJA1r9LaoKq7+ea
KuBWpHaaC7knAKYoVWgYHk+66fjLYdn5gw0WgqIxEHgUb3hdatXn7Q3wsGwIa0Zy
R4rL8lUG8IQW+w8FbMA138JKPIvM4ixAPUpl2CS1RwXNmfDfiq3/rFqr7RTwIHc3
Oj8zq1J9VL3ot9GdyS6E67mW0lJOSv2MOZFB5ZMt7XFrzo9e5R7PmiPvoRlReUV+
zS02XPifK/DAA/V/J+Fj4UzD+I2R7Vz8uENePIdb6oVgOC/RQ5eDmcSX+mlGICwP
1qGcDaffl+fsLpTrsGU+JCygLf3KpZKq8RRCzfe1KGWyPFewjcEslPHAiz1SlFl4
dADp9AnTa0LNo8riGFDvS6dlzgtvHhC77baVmkvFuq4dRwMT55doDWuMaa9MHCgz
QWIqZNa6IuDMBEufkBUS/UWN81xo5H8VHmVUXRDiqA7+Tyq69XUvAskjlc6Bsk9F
bAfAOKjl5PYLk/fQiA67ELIkIQGsnHZNL/BdGd3IA0nM7RYwL8ZzHoreMKXMFevY
RT/A/IVWXwaJ+nVUCpu3wj8oExIhHmabRKolHh7aGJFNipVYlTIDB+QC9WSpc+F/
UmuHvMPAG7bLjwG2l8aXOcEYfYxjQ/sUsZaRt9fv4av997g6L+KKJxgTLYuihq+P
coHbtoUsDTAiXNQ6+wPP7jS6jn6dqu67TU+/off183K1/LXbSnmSCfzJtiiVFQJi
xnFBzIHkiw0UQtzh83+zNiiI9uec39/bFhmZmlGdbhiirQLxyttMiTiomNBbrSjg
UTtRx20P2S0izJo11wDdHHfbF7r8h35a5mppgzoMiZE0UYyUBihqEPzlSD1v/pdH
IBmUL6tgt1Ouf/sXUlJVtYl6VD9i9TagwlwFjARrkO3GxFJR2sgAFcbJcdkDkTRi
81VeQ0M0yFa1KCyGCNOHk3O8emyFyJ/UXgS1TP3OA20/JTvnUN0XNNPoowVODS0v
5hUDOKzZFuiDocwhoMfIN6Z4w5I7q8ORoBLo8/Vtyw7cxaTylwETV051OXYyfb8Q
62N0AuI68cS7Kh5aqy4GABagUoU2n8Sd6HvFQt6Kmsyh5/0aJzzMEznaOvrZMN//
o/Nbd0k6AHWZPyq3gvBsvOgFlqSbcBhyHPRb64gfa+k/7sQ0t8k3YS0qqAQzRovw
s8iQ0OBq6HTW54xjZGlAPrN/ZnozbUXZXu9hEtHmFwXgiY9rqVggEbG5nmnwQBh2
KoRlhUWoMMPQZaWveNobJDVg7AbVvld2gSxnTjHlDjtfkEyR17xZ7kVvL9Y8dUDr
t66JcrNlfBqBPNo4g5VwnQhsttji9QjEXkP4MejWhCsCaDHJdYdamScCxqyMVA+d
+BGCDk7TuXezohGOr3ku0mmt/9wdFPcxnYFS28wQCLuLpmVY/+SQz/SiJ4G2qt4B
2CSQuYGDeA/DOx6S/ZYdYpyPUy6xUkNRywIU5jKxVWIENfeqq9MEslIgDZTBb6Ub
IVfhVdupEMchIgglLz9e8bHCki/4epHkqsFqvefdQ17u8Bnow4hkqAkgmhjtwUFJ
+UOn1PKg3y1JLOqDZeoMgmdLlw/Tjhvv4MSdgKZmEc+R7LjztzR2HKCbkP9PHajH
walizoxYjjXFHFQYOsN/utK4/6H7TmZbDcXkjvkIT/YKwNKqiHNhMOuBUCWPL9Ma
zpaA1+XmrPDDPI7253FH/I0EOgOPnS6JR9ouRiaK7mjYHctQTe0KYp8Li333OofY
CNkB7Dj1Defmw+01YdBH8ENNMv1tCOpsWkKhskklK4bufLgzUwh5axe8HNOFSQx8
sWaTBrJRyLaLT1jHJ0yj/w6fHPdYNcU26CDGKlGPX0S1qvaZJ3kZzIC09nkPhY6u
56Nqh/CxM/EoVUXvWVZ0F8Zr7UJ1qWxv4bIbEOL6vHvmv1aFEUn6S+UCjqlValoC
5BT1oxhribRTaQ6UlJ3DYOnSXVls6LQqnmz9qG7KLcM0zgNjN/kaQFSHVWlp1J4S
I5lLNceL0hx8Gimk/R1fP4jtQFkOf9LA94sUcGzVIBvKTbkOUE5mqYwdyAZw6yV/
VY3xgC3m3M2EQyBuli336Lkqk3CL/+t7FSsJtrGiMV6lj9TtIKXCypnqOYY1trXe
pcFlW3v9uLoQY3cduVo7YXE7WEy2BixdzLETCEdAG90L4Gc+OEuCz4K60iYipHjg
GIXfOW8A64czj7M343q6v38iaisv52bs/ctibWp+noahdkLCbr6+MHQ4e0vnHEof
rF8UP1rHp3Hdv4Tg38scWRPRNCiM+dIuiVdBMPqvsWCkOlbCYNHdQZDT/zeS8TB9
Cx7BP+45PKYFttOVvExKsx/MWd7+HGjFX2WW4+pXzzYovp3KqYKy81LtZC3t2yhv
eZEk7aEdiy6CA5avyvMq+Kil2TOZ4C6jBVWLI5ajXsqDDUGufU95mnALa87byxk9
SeHjJMQx0CPdUKCF2jIs/nk0HyywnKRZJL09MsbWgR+5NY9etv/tWDC4HitubGox
M48g5F6t2ERQvON3tcVmX//32QlOpAaSj5XuVcUDz7FIyiV/wWNLnTSw6XgTT2ci
KiZ197xAqfopjs6dfiMrh1g1k8JQAnOmpHNhsqJwmaIFCun3fyA3qRGcOHJzVYai
eT9sKFu5XzQgQIiWeR1bipFotwH8q+7c5y2LI4BdFO7hdse+/xWvJrfR8rstVNEP
skDyYhgExOkaIDujqot7E9axmOqpYWWF1sgn/rX8FwJ+Eu6Q9C/9UJEPJEJ0DVdB
bq4PmIVtx1a5CcB3a59ovKzEPVnPVczbJuNlLeP1e6UVxDHd0NEyltF/4qTx3oM0
yTlXtdI8PQ8CcoZgKxfeYx+V1H5nXpVNW07Bs81+99rpE43oER4rMzwzVTUG1gVC
O0mAW7raSixQdlpZVmf6x+gsWZyFc5PbBrIUORHBMKSqNMTb3h30sWf8n3LFhcWp
qtccJFYMWspCGrrl4YWbaKg90blA2LHTRjT2pDrY8c7FL5hX5KpP0GjTxXiHtseF
0IpIRBHY5oVnXcw4qUEORy/mkghlrH2uDY4mEik1D89JYnbBe5SmwQuQbxRh2zXp
o72rvDqHEkFeHYyLNZkUIaOORmsdd9jJjIgvvnkBkSFJWm1zbeWdiBmG/1HQoIwr
XXai7A/ytZED8lP/eMTCsDuXzfjkArbk/MFAdcKMhLwscmkYma6p36lqRsVkXvAL
PQqvGZvpCQzWCGLMwFdExovAEMJglVzA5SdTkquHutnBDpwP+yjVBitLzg7cszrL
Q+Qa8jSukPRkSZC21GdinV/ypzhJ65a2WHafFYbkBdDiBOHaafOBaSraN8yDeF4x
2zwdiftwQu0+5ltC4/lZotF7k1Z4m83vRwNozxreDy40xqHaBQnnxgySTRLFNlMA
Vvt6Sw+aQl2L5arzsZhM6zopiLi0bvX7l51l6PiYfEFvjTSgxySzdTE1VAaxJMJk
tHM1bv61jGe0u/m3pAky+FWSdxpr4dX0LqKjNHx46ovRbcMgkSZSYj3NgQ1/12s7
wKufN43udWt3FWxZhGPi7rQJBzPaOXHJW5i/2hwkBIaklnesEUjDx+ZWH+a5ymFE
pSuGytIa/uaWoyOXgyFuQ7S3YaOA9J0gWi0fHOEjCyFelmaUJkpiuGb7II+6JpoK
B/rL2uI566rkWPoMoF6G+qr1lKSSbEavb7KwhRoo2FcEVp1ZuuqVHVKCs5YIpZRN
ohBugoYbat0F+zJF1bGqmEKsBbr2g3ZeVHSmdlVPiSSzQRrBeHZ+TscgsW2urm8k
Sd3YZMyTkRoDtIpNtG+37qsag1F7YSNdjeBUzjRzJMpDehQhH/6jGkNxMT+ohDX/
JgfzJXKekzKde8LG8UHNv4gPGDmvFlA5z+JqffmM6aiEvo2X9086tg8mutNflBX4
eSJg+jRLfu/W4PMP4+Xj//2kUak39B6s3QK8/p1VWPU5Yl19/XzjPjE3rdDUFyyE
nrIW0eX3d2k913HXyleNp2UkWqIRiyzIZdx93ISyeJNSi+bv4bHC5S5DCxQ320ka
iWgEchsWL4Fq+FGpmdrSn16V38v3X5AjOZX9sDYRCFthFlmi8ye7d/IIK/lj8t3E
Tih0F1cSypOYp7NWsH2cJVBj8Sn9dKIjvjF3TKl39FqnkxcRlKNLQC74GmSXvO5D
ILbQZ3hpVP6rz108gxzzRaBBwS8Brinc4UoGD0XrI9xQ3iL7ZmleczhkSPYfZHk8
jUX26JxpezzqkqvUu7GEFllOltkbMVCAjiVHnzuER1p/pIrcZ+9LRNhnqKYrv18p
Iqrtq8Q+Q6NpG5rc1QG55ZMj1PY/8/VChDBzvPsbLL9jKhyig7ImLae+nnkpDjjx
YyBqVd2GPwvrvWU8+KsE5IsgaYbEd7i08mqkfOE2E7Hok0X1/3q4555aUtUz3HPm
F7m3wOpWrCz94Raacm7KOTwW5uUXfQxN4c3rlaz+UVyzjGX+x6SFO/DIUe6u2XyE
OE7aVXLlHKFmoOxM6vJ7vbNMbDlHp/F1/gGDHwHvuGSDhiBZPzKOVWxEvHQ3HEdq
UuNaC8XjIesoqTusslRh6xDEt6xhjtwVZ5sqBaGkgzl/SUtadVBl+4Ru5Ef6GiVi
UvSGa4Vlvb/gGhoBuQRTEUfjhqsksayQ/yIW8JrXozDnJ19MNT+lF3vvDKmMmCXb
nekoyuo7ngtGl3eLCTUTQ8PUiyThmSNwCNEbDVzTOfA1ZvWai3Ab4UgGrYbC2FPQ
Z65b/fovN0FnmRTn60OgpaCM5tsuoV8rJdpHZRm4DUOv2C8zL63WpeIdUzFrxsdd
veoTTYL+pPoeoQcZFda79CZsEDO6wHWw1LjEMYwIY5hVmctMad7aU2mZea6m1AOe
SVgxkXkbXivo9/s1vChxdouuDPhwKuPPQOij09QTGp8ZVxIzlJ6ab/dS3LlagCO4
oa9IQZyrlc02anfPzz+GWX+TZKwMNbew2YHimvhc7JPGO/mO/63/0IB2EFyR2jyu
4RXWxnPd1rYYDESem2c0ftz9n3yJrqy67G91VHpk25Wht1j8znKRRBlxHIgR7fsK
4/IhDX72iIifdNRGN48/8uoVVIxZEfqQzOYxP7TlqWI5FcBugLtZdlBh7vOZjepk
LtS6B2YKOSCA0mb24Ij7lB0dAB4E0YpCV0Yl9S7suIb9ukQmpoDYpF6Hef1Wx2Q+
lRx2Xq2dMmKg/gkMLSX704SKjY6INkO7W8UYETZnGrAI+vyx28BJi9cTk+wBOHa7
5swx1Ze7+7rgjm9czTT1sRINiIUQ5TtEHAJkH44YFhO5JNPIKoubm9q3nRAWhqYg
6Y6xOpIPCymsAfH6Rhufg2hpmnLvZhiybbKVESMD+nXVUZWlMkcH1xaskysl0+lc
+3UCAsfyAKupySSaMujgtqhkXSJXmsnwSHsXuUNRRRIn2G9giiKb3TfkNhZ9f9Qr
oFdJdkUYrY6D13RtTtkT/6oFfwFn0AT1pzbHyXAIdS0gLk6mpRtqm9FnOHei2AkX
pTie5sDd4xSMDtF5RGvdd78SSOPXeWw1BhyypXmcAFkE7d1D5+oBP/Ow7OzdsxyU
IWp132AqsVht3CLd0EcCuPGuDDIe4w+9Qvl5NhNUNOLM6H7tCT204nxpte3v5a0S
QLEYpGvAbBb0+r9vO0+Vgh/uKSZHRgL+/CW9UcKi4QjRIEnYXQcKVWFQ7Fjdf8Ne
3Xz/vDRh2X0z536ibu1MvaF03viHc+RkWltJZg+kDcQaT6IhdEi4VT7rb8qwvpRu
irwm1FLLLaXqBpfPllPBL62zSqlyW4R7utvLCJ5k3yYmQ8L1Oc9//FK52t5zVhcf
uooYBDyXwe66BCnt3P14VcA0PWs/GbdZXueEeWhGFGm9nZKiJH0YjGAV7LWrxtIB
LtimAKlSY9J+a7P8tAYDb/BO4OUjTYSloa9qVZ9OPyBu8AH2Wq5EnBo2NUL/XWC3
DzQA03GPMqU1PmFF2F/zHeIr4AJ4Sxu3uWK9JvOGyqDUAS7RTO9opm+KrenamOQf
/KI/A/LLvjgoNi+Zd6qjU0J3/4dcCfdrgRHTPHhQiSLqYWPyqwRsiqDTcxE4sUB5
cvULj1B1Q40ymgviyKH3BezAKMnyrWNajLGDKDNWJW8wAJRgKLdqiGAVtPHCYOWb
TyxLfZzG9+wzJ1wyosnOOl4ReexFxsZIMW76aNXzT7uEcMdZI4TxVsqBSpPmfD1I
6ZeliYCRPIFnzu+SVRaA2cOEc+6vxaQQQFQ/guY4xXB7E6XvpOa4AzuhoFZB+O2+
6QOmTWvtORT+LXNqiL4kc0FHgq3RB41ZrnD8Pf0KGjHRpb2in5aljoyhwma560FU
n4Nb6QaVbPypVLon/qyQ0Q9WVa+njsKmNKWFnEKOoBkVsE2Yrme/xAM9sMwU6u4r
G/jHAlB0oLOvo2htLVXxnQ2MOcmoKenaUHj4YbOiC7Zt1c60bNstAV1BrFRQaEcQ
zHjdFP7A5r3Z1T40opKPjjBZhNMZYOWSy7RUKxlzmoPEmopWVd5te3OHBUArm2sd
VaJHQCv9uQ4vZMfzyAuZ4PQ8vUc4J6o35mGG/yYp9UsMzop7oMUB09uBFzvWRFG/
9D5ewxJCHwguZZMOCT10pqXNaHzNKecEMqqKbiNpfMq4PliSgoZpXMLUNMcnJiao
QL4cm9Q76R6JBswljXpmrzKvOJIwX6OdNIiRBzyDKFEW45mC6ARn0RJ0tc3XIQD4
Ddoochrtj60/7D/wRKDthlQTsDUk3gk86xJeDH/CYZmJVpz1KWTkkpfXOnuzXrBy
9iPrmZ0QQ4uCUxRp/ehVi+h8jWxbT8P1RbdJyRdqXSb+2hNvGLUvxfZcPttBFW99
4/p1/Zj8Lfxq5QGP1Ly5kZZ+NTRf0YHCRg1aYQQgq88H2EadAE3n2np3FiFuXFWH
kWU8ymaLsuHLAoKIWPMip2OOvqTtlkHG/gZJ/FkbadztGqZMcWbrsIdGPp9/bOXU
lJJJje4/eAC6tuuuuinrGR+zPFzAo0qlD8F/GsTghSDjARmFzNJs5H6zXn849QTl
etUzxPOeXCaNNENHRZNrOzefPCAHL077213Jj9AD36f2bSNRHllRAneZishkK2rF
AqJBwZ4vO3KqgMBM3oE4i0lmIQYT4DHkWF8lMiVGKfL8JP8ThyOG4oTijRoClJfk
NFRnjWXjR+V1peL/wSxDuYtO+ncbdQ46PO9pTle1Od/3ZddIa+/EiS8gngyBnvTF
yTQkMB2vNeqM8X05WxUA3EWM8ppbJvHzJehnmzgq6x1Kr2/8pUMsgNWmILuVtLy0
c9IHN+w9EmIioDjtyhsiBACaf4/f70ikN0D8jp1yPGKDdjHykQqUHn08bWh0NNue
NcJ7BnwNJoVUqsC2nowos6j1yUuhM0CXOA58R3ei3tcalfenIDpTz3zKFW+9cjL6
5McaFkWgyYi8JemNLOtFpNzs9aqxEJGww3MFwIJy2MBQpw7LPe2/yoUGFXcVBkPK
H/RrEF/cAFBjOV3SBMFM9GRGPOST6uLBChGzsw52e5jCe120aqcRMAOmOB2h37UZ
z1gpwSFnygEaA6tl/idUJGcZ1TMQftpfEaRPtxOJQ+di2deVUBtas4/I3vUIDgcV
6BZHsBZR4bPGfT8DMEVTIFOiBseUBrwkP44V2vUMSBsWjzk9BaOpYFFcFwdej0dP
zkvPx+pHFWCU2O98xdvEFsmBJCBLdcSxfrb4BexXNJim9gIt7tvVGK86zidvoWba
Yh8Yzgbwxaxd2fZ1DxWGm3qazPeKwOyL7qL8opWWJzvTqqZx+Wk5huEHF7qxV9x/
7DSrJDAy2tNhnhRmuU0f0PhQMzsRjIWo3+RYNvavG0HU2+roKCwjdUBRSSmbJ20Z
m86SvN0MwORAaCii36LosOxAhvxg3M+Bq/FQK4UXyaIb0AjBqFKft+olvhbgm+yi
Bz7Ys/7iMf1eqH20KrG9/STRm8tndLP4atZ60G2G/Ft/VR6mGuGMyGgPgC8gsejh
9JkgHJs5fjl7mO+BooIrzDArz7zCXfSp6k6MGoTfDvkP0sqgV/JYWl4DBMlE45e3
EVsY8wpRQBDtXopaCi7C6gJLCmVjCqMXtWEjDmTdxmPS9UNWBP/Sy48M3fABN/4O
5jpRjLtQClvNg4ogMYd3dHg+3dr8mud0UPOvosIr1K0QX4CyLpnJEtgTjzD4x0Xi
pNYUs6G1VRoNCqKav2snJJEZSH5+2MyqKEuI3glGqB24YOGjpXBxOUZ/Q09fvAXd
YBX/oYfFtPsbw5SGkKC7LbcrJabjwmqKrtuoWIuwhcuxoo4sVFVlPFWQhmOWhOVn
k6P0oOVuu89Tl34D4DYWi15BxzhDN9VqsGHp7dX3O16iWfBEMCPrm48edtkTE02k
fd/yPx2hV7p6L6ebJmbNKFkLBBmUGm/O4kiiOBLzYMDbDRw7MdKLmpZQ1ucQNR4I
ftPQycgTDZOCnVrbRerlQHco8cqi4SVVrHrViWQX5COCnFsKV1HkehnIG4lH+XFe
PsbuyoZpTPnKf4kvpyfLcJWabTJFYJDcOTHs2EIQWJHIxIvk6i3zbpPIjRZl23EZ
d17xuSCUnJZdBijeYzwRcnaXwieTbybt3E3g0W+ioXJlau3aR01hNpXgQ6ll3JUJ
aKuPJGiYO9Zr7x4RQvTaDKh9at0I5Yvq3reCZFSM6H5pueOMngNhegJRXdQuZBqc
3yG9NCCeyMLWqb+8iIhQeTd5UzD3eBeNtoB0d4azKky1+hlo9Aalo8sN3Dag2o7w
7/bD3B5Uf6oafdu5M3+d0eTjYGYopysdCMbt5dPMSiQwWk1XUDbrlolgUpdvM77r
BuiY3im4GT8ZSnpV0QMNg9hygUNTtrZiImuedxxdz64+5p6HZLSRz2MZ3w6ApLxI
+AEhLjqEZirWRrGrLhLEXwwFoeEFOIInmKwVs/CwvAJlzBZQRCVpZ0b2Sz9VqdpX
+8ARzP84DBmh/2bq1UXrXHWm6T66B3L1yzfAcbO+XsF1T6WfM0LxQvrT+gDa0rd0
Y8BZUoFshmUUkX2lj6tQ8RUQtCB4UKo5sxMRNr5OhDMwtkVqtjohzHnq+qdgIFVB
VrJDdFrpFtdhWoH/ybUB474K8QwWqI9sG/h7LhhcDuHAGKyzkrNKGllljlC6e8Xq
deefkTnK84tbKaATUQ7J7GFhS26E7e1Jf77/Cr3DnG511XWw6/18RS4FFYNeB6Po
G1HRiP/KuDZIxDIHz+7lEo31w5J/l3/Q3IOzjnE4JfWx8sU1K40rcUDxZk7F4e0L
n7niPjcx2V6z5yzxfh4Xhk/MMND7dMgYf+CTjAiv1K5FQAUnC8s9MSNa2SVGjGZ+
o0X9C5nQ9dvbkg8SwaNCMi1BKXjPmnm6O7ED4KeIOb0EgMPGjg/Oq1L95Oolc/MW
kPey1SNGU4SAKY8XGs+HKP/VO/inLZvrxORObwlDqL0g5TMcDvn600ynHEZgJzl1
ligRfy1SBu7+uRLz6w3JGSmJc04jNZNR5WP6UAsUkoTZn0nHL7IjVDy9DvbXtohl
05ErZSf9IQs682JFuBFWPHoLWF6XkhZ6Z9ixzskojOagL9BCUY4fidWMAlKSf7C5
LuNCqi0s6YXW2XIyCUdZVxD5xZsS2ijp2wrWMOvW+g02swyVwfRIhsSqpQvlcvbG
2VvBKaVshMgiWR2JdN4OHqUvZMVZHSabHonKJ3FZm58Tv/Gu1GC7OAPQQ5UArqVl
TIYacJ4gYqBDzJyVvKHr+bEfvw0M334sIBcHFyx4P8/U97fh3ok+RzblQfKdYMaT
FjIYxvJDoNL8bDL+ncj0Mvmj6/IBGfsLZM4aMMY8dGu9pZ9LIv4tvRnnM5As1M4h
kpLGsJ1vN96E3AoUeXtbGY1MzcXGmZ/ZqIsTuWBdYU48iY+ijcNVsN0/p78GrXeh
bZvaK7zApi0FtNtJiTlDesreo7gK/NVCEH6MMsPJTgzzx7T2206hmb7KpWFtTNzy
BMTMjh7ofCO73oQ4blbXBiOYCDiPorjTxnNWkLI6fskf9bJWI7h0CdYMay1ZW0HE
UzHicF4RHe6nJiytgFDAX24yx/gr8yIbrMlmGFZRtL+kjobDNwXvNTecOGjX9i5D
BC3s7EHGzaONFDtMGS7uUsz00RQZPKvsLExn+k6X4UJ5B3x8/4HTf/4ls3jHoOTz
6I3wTWDdb/EFOMe1rDwT1+ZZXT5yZPPLTkEQsr8YkMKAbpWzApHeCh2YsDGnx8dO
xXgq6/lxuMcXX2CjqYvhcYcnY/RjIVNW6i8knxVtpWWgqSRKgLskAxH9mbwmQASy
2/4uDAZuCtNkbKGg/ws75HNoyYCfTeROrJzEFtl2iFei0RRVNBh6coE8XXgt/Uty
cfLhm7pSJSZCofgoY6KuyKDeYsroewV5WPz/ojfTz/26u7Vcw7IEm0j4A6p53FLz
5ZxRPB6Ar1ac+CA0mbhjxNPGiqZ/Fdl7BSOoVLTXXbRhCUzBBu25C7jhq3+cuGDW
7rLOK5G7bd7AXT/16fWPok+XEM4VUcl0hpHPI2jtBzejFMHo6JDLjxHM+HLzOOcB
6WjBND+9FflEhQrrTkIbOjAg9dcsh+bQjQm1yP/UwI6J3XhpGMEarL76ZslodyL+
Hr4GqHWR6a1MB3yjYRjgycnii4E0UmO5dWCIho0y9K/37E3PHraTHw81c2T9cM/j
DdG1MVJ+6Scj58teWw9RCHwD2IS8nWyATViwCAwo+ba21Sun8kCibyA0hBfifHEB
lUOff0/OE681tahRwTK4+NnQbs31d4X8vGBOIkEmE9QG/uHJxKdDzlwVLbwhmbtF
deQA6mtgkOYqgCauMmMqpIvwI4S6hTVsPkzClRQJ6a4IYHkQgdI2qRhcQXHUf/fU
igj69YmQ2f40ouKVxNGAPIL+z+GRlH10QyinhHhULIL0pgJOtEDd/V+dPSFODOYo
qggd8Byclul7P1vF6J8LBfEAIBFHu7IxZLD/MsinuYGHIODZXjB+MKT4Na20q/36
Zw3jkAtVfIvJbVueSovPpmSbeGkjg3w/taykdAY/1fJOuHnpBl76BwqENrl14/QL
5V33HvU2VFV4fY6I5V0SKipofQ7LVsBlmPmmMW1M+vLM5Oppl0f5zzWUDweA4vxX
1D2n4YaMXMe92LxRtTdzGu8Nb3NiLCj/pxaIw4+8heLWl14pfzilo8YlqdtgBRzx
VF4I/P9ParDNSa57q3JW7eUpuXqmACV+uD7QVercZ8mK7w2h/b7nGZ4wsdbccEKU
2wHA2ifXezOiV81nXJ4cmOf9b7SneCSxWBkTt1oGKbW+eIR8BZp3rWMkAcraxnP2
mFC1np3T/eHcaTuQO7aSnxiY9ieDrereBqPy4Q2cdImEiZdiDvU9tgPKhOfcmDfV
PsriWztwWzXK1lMmsGe/IyDK4UCDc1sUoupMR01kWXsdSQhlAeO/xjw0fxtgcOgf
mmN5QeNLZ3BBkN+3EWE1AFsXgkyHH+AQEMNhQmVt07gOYDSqTsQ+sparMig3mUOP
S0FdRHCQRagf0GBcqOjTuRTyqrMPCPeAl4FhDhLxNGkYMaMtHNZmSeoPgOk4YRmU
9ThwAQMaAlhrZtW1YUPFLucqZeyZg703V3vVfk1nY9RFn4Eqxlks60HQb8BSkZCb
wfJT97CvjyJ2C7UJcx4ujg0jCg8hXBrGzuvhLUdcIBwkguHyHVbyygxxPtCBxGS2
J6np8KKduMey4Xjrpaiqms9B+bmDlz6/8Qi1Vh2Rd7I3iR0mn68GBet/hnf7G2yK
LD7VOnw7rRtIA8gWtmWR/972zf1/gLtKk7S9C3r/7KDuLDYhBKtVZwqgYDc5oI5z
PHNnKVuG8eH3zquVG3gyFWCblu3WhslsIEn3NNo0RXKfa5gwSo1fBv/SBtfWMcpn
MMe40HEwjOrwgxGrmGZBgCsQnwaTsKKK84bf4aq6cCEJIDZhqCnU4ww9CgC4RsQ2
IESNErbpTFdCF+GbjVpfdiis11a89I0Fit5dkaPwgbxFK7TTgQddqQCCpDs8RPeu
u8B3E2x/eh8hhORKyjFuej+IGXZfgLxPiXS2kI42Z8l4OtKGxhKv5pYPJD4LX41+
yP9sIx8GCVQWcNZ243pP2qTgycF4XUhZxHsNKk3u/V/kcuHxSMQCdv3K8IJRyvkS
zFxn772aUyqprBskO0fwKA3marQNWLLoyx0UW5lc6LeaCP/IkSaShVfLR+2exC0E
tlOc9P/j4K/OKAwKzNYGi/FbHJFzkARbi7RYCGwIy4Alge3kyyLWH5hVrRURjmxH
+JfQIE6wgWF0KVPJV4ooceJ/qtsJNk0tFEjvBY1lq0V3sfj+2ACxjON6TOIIlb/q
zpgcAqRA0QjSl4q2P4dc2xPETQg3jWN6A2DdKiLAvHP6sM/PjJbicOvflS1CKx4h
qVNTYxS9+Ycy/9atN5cbUDIfy2azddXRlG2WSn19XK/42XIcXEhpwJnKoESs74CF
pb/fEy6tqtuL1MUWMaNxOK7sk6zWXMWN2VlWsw8jhNtS5xpERlYwMloiqaJ66xvN
bKMuOrOwHwwGSvyy2Xq/xVFm0px3wuFpfmZsb8r5s+ftwUa8OhN19xBzxQJLj4xn
KYgME6YA9jNlkCBlBIq1Urb22Qr/mHSnw0yHfm1SuU3zlIroL2VuuBfqXcRotr7A
OXR87THeNcQBq00T3vJIQyB1838t0hnfe+q1QGXtXOc1m0Bmnua+idgOSz3B74p9
uBzCmM4Y5kdDbSMkRZ2mcNWLfdkiTHQznhc0un8l8PJxpWjlC+8c2IVnAC4uVkRX
15fDlzl66zIZGQ6YR0YH1uNGMh1Y/7X2rPP7ilm3YEKWRLCsnlFhkvHTu5S29kdk
Nlg2vfRGwFsrEs+/3GVGUM/GMdkG7vUihx/BVOwqGim/GiNIH9xqFx/9mXgEKVTY
6jBGw+Trby40PY1//zbsG6JgSeN/FT0+GI/xestBzSva6kFlKXNZL8+494HVBYF7
9rb5hL18GFB8QQ2L8YJy6XOyQ6XEc5sOyGEhfOEFiApBZGFbVI5dYDjFF4cQfhn9
LPQsBs4Smi+UGHVtUTnBL+tHHJptfwDGpTYR4dtQIA7DXzpdjye2GkQFhH2Qw30y
ORl+KrDxgugHG086QxeN+xgKJ1sse4xsTBkL04aAAlO2D3oh7ZKeycOTyPg3sQKB
g5iM83630T4uxFyG3mAJne43G09yDk7ERZaT3yh3vQU4TTYyQ74NQj7SSOs6wuwZ
Ehe2KbwCtXwobqhEQSs4h7e90z9LI7GQ2m8kZGMXD8KX8MknsYueYLF4kSkbfgvW
0ZGQEa5D6fZTl5qfMZFryMgOyQzvULslytUjFVKrI3oAnP5JPqTDmFitdB3l+ReW
YvO+++PoO0VJARB3bHrWlmH/k43A+wvCRZ4T0AcJ+mBfP7L4F9s5UdMdn39/v3/R
RUMSJsv6swTzJcY7gjvoJh7qccZ4T4/eAxKkEyFCk6Frn0tsC8Ry8ale0bNj9nvD
AGDy0re8SyUhfPa4o2wwJatsAFgu6wZ0dMw8M7yIAvPlWmnqWOaDl6tjAGjSIE/3
0kz4yIsyFlF8j7ASR65i9BOza5zA9yviCcXQB+ffNOIV8/VZ+E9YFW8CP3dIwWLl
bBIkavH7vg9FpttxqYxy72wkkTP9fmf5tSY4HloLWezMbOmzbQbnQwuAvRQxXz4o
G6LLU+6UvOay4tBRTblLWyKwQAnmIDKmDWbnEa+KWZ+mmQXORIebJdWDfNiUS18W
LOoBF0PrGg81VORZJDrTJOpnF2oxj94RU3pf7t6w21tUtcFUzzd61l5DvHgqwnw6
BuZ3tB0QteIP6Pq30gHKvJgS51qqfkqw+yCHSD8tAjYtBAfTtm9IZvGrDLAx0wDI
bdzm0Ewq6lpKbZwB32CyFJPc44YOK/BmYjKmlsTIYwaN8I/asYh8rB9XehdzINSx
sY+hbK+dHutOvgZIxMt0bZuoI2Zsxu224QvOWpXa4CuxRrt8n3uiHrCQsGRebLQm
PU16N8hWFHmsJJzCVPCZ15roDxELYyKsAyWzyac1iJEEoOIYSWf9/85ZHAPOaCMk
icaohWe7WcUvhQLS9KBjdB1tEPnYSyfR6spOVZK+PEPesi+X5Pf9Z9Z9ZghK2k2A
wV1rwNSWQ562uX3XxAj02MQz1rn/VGAbZb9/jBslkoFgrrN5k5MPqQC2yEHcDrdz
6GzSA3s8jd67M4wull+X33njKl+hjF2PL+Q4fcmfOiydOTkfhEfRaF5Z7e+rEn54
TfTOIab6NKLuRvCGJZwt4X/yZctf+Tl89b4eW68SYMoKeld9nC4XbNanlPg1WYoH
YERXpWfGS5pL2mtUpYD5RT+dviaHmNx7vh700xnQUFW7POLLeYM1dJbRkpmL56hG
S+ZE9SCIyEPzBr4Y5FHfR7XVT2gl0j/1wuSs7MN+SdWuru2a+V7vj2ACBdXgjLoD
bzFpIpcabHZGc+cQidNp8h3s0VVhS7yVpMVpk2IA4QnHWNtfia0HbCTPMDZt7Y9k
ZVIBiNDZoql4nDVdxrOQPXvRmsX4v8NxU56raENubk+tsodU6bI1Cx8JO7W2PeGH
czRthzA8EDiLkOxFonaNe41Rq3wPCKhIV9HgNqy93UzZC2MzmSaKcAN6Wh3+Q8A4
wR61EV2ctG8zMUtOoVUBUnDhvDtnLOPuE2Msz6jFkNGA9mxzITyGNAkCLauIEq0U
QBEOBiMIARKGcTIYaGou88F6FQlEOIn0a8TBB8L2FfY0a0QCI08tV+ETbHCaOGfk
0ojl9dudywjC2pafdN8D+87Mduuac1vyXp4WlRGXOFS2dZAKJYDyctcZm2gEbB1y
QWtMAwSxDDQJiBDxP6tOHtRAqmmDPbN0N/tZaEm3lA1cM4HQyrctdkGkx7ycMApv
7R2DGQoMFwJ4QoIB1mjKxGuLldfPF8J2XdRfo3ZW+FLFIgR0JqMkCNEMFO6BOn50
PcDxqM2LgtyhzSLvvXSerYwDFJ4vd2qtV9LqQv111CRkuQiOy8nUKFnrzfmm+gyJ
HFMsnraaG2EXvYkSfPfU9DaCiJcEO6Ly/0x6+uFYfnLt45BVgQXo6bg1qArJi74O
a71+9890TqoCutLIzNzpqbHvs3EPLZaxcMPaMqunxK1B+riARYB2b7qZqqA9xTxF
4EbfaC1q4iCd9PgApeLWf1rN+u0b6Ti2Ejwfx0JVZiCfTu1q10AwSXUPS67+tr07
nQf8+56Qf1TB8BYVxI6RKmcDAHULK0QOwvgZNFflLytWnoIDc7Ixxows6hjO5uSL
X0ImU74ZJC+T+1XvVY50cSglBGw6vxB1GZq32uOFYxEq9ofbxBQ8dSl1Y0+guM0W
aASvVA20pKT2fsGMc96DZ1/r5Oy8+5WTL3BAgIvvlLLL78tzQcaS2RX7OXqg2Rh9
64t7hDViko+YhnmS3nsfmxwHLAhKOvGBApQiQopJ4iN2IRE3XYyEEk+dnHPRvPac
EyRc2+M0jagBgazBbVOYB/7cPnDDonc/VsgN16jHkxaBbHELOgX5WakUFbUadrnB
F4wkRT1f07bVjDgQ7IYQ5o67Cw+EPS91e3gWOiFhGVCk3Yu0F/UQ040Uif4s57rz
eIZ+g8q3cmHCn68SLsm1pOnJMkisYA2OUTSvdXR0yZFjpJqVxacuUzcABVaWOQBA
jRz3sqpvnA2s0LaZrAdZM2q8G+wLFueNUdU8LwcMXdhlfX0gl2PZmiyQ3qHLvuQb
T84ZfcN9cw7s3dcTAzvlL9vOAbTavW3OhTczkOAoZgVg9lzYvLK3SxZYOA7Y8a53
68eZy21J964KnmTOu+1+4r+ssBQgLOwAw6G4G6RTze2mye76dHuazn+udR/kkPYF
asU0BXZeLTCQl1f4NT+jB0hKyqcp8xhQJWvHbYLM8zi4sm/U7zDr83mf3puz4yvk
M9Dlatfg+ifNF+RdN/54Az+Vnz0UvOuzl4FjzkCVOW6sOqLk0qJpv3C1WSSeGciD
6b3eg9GwB/BB74CBUCEDabdNarIOccA687J2/5MxK3WLq+NoG1RxkC/u4m0sWPUs
bAR+SfpEQNAjFOPdFbK65ggTrrp6Ktb65JD+uLBHdHcQ/hDGJvCMNPN/9yMoc+Sr
TE+vO5d3D7i1flSN6s++0+g5PKPJT0K0XgoRGRg7b7LytN4EZ2F8zBmjrz5kD+EI
0PM6JA7hQRvDhvhWH9VVr7PZPsNjOTt4o9PpqcsTVl1a30Y+I4DYUJlxToGrVnfc
q6tPKgRJmxI35eKFmMSR5LZuNoxjJ7CdKfHMG0qykt4KVNCqm/0mEMlyQWOJWN7T
ynqzjpgbWuDumBkx2RJG6oFw3BD7kmpb3q1+nF5hn9YkHH8Q7goXA63Rxb6+mNYf
01rcQw6utGgKLnuLD4zCod0Bd0VaEuTE+IWCncK6VQwp0fAVUBW10fAGlHLe3H4Y
/ooHiIOgJqfsvf+af/W33y32hDk3clzpXsnLmmvkjNE1Q9DOnmXosaEeDSkM57g0
pTpBANJyOvLQpkk3BoDWu2Vs9AaEGdrkZ7zLjG++IMObV1Qz5xnHXSe/2VRkziJP
9plk1fegQiqUzcaRF+XB8xcxYh9MEFavOFK+8VjjjaRzE/09/uoU6zDsWTPKhO4Q
LSnB4ChyWozHbnq0lomHBWdVOzVwHuw82t71VU93+lXiakQjL9ZL6Y8UCuWgZv3K
GXtmQSyFeHRXP7b6Ad5FKdCcPL8ke4HjRP5Fh+YvX6HYrhimETozKiFlx0om+Haz
zUwpFfLXqLDiP9v24upshOkRZyYhjgzZjNJpLdaTsAK+rd8soJcg47URpcO43rIK
42QvsNvpazXgNqvrH8bR7jFVlaQxSYi6jAEBYbXWGnwk218/gSwivkmu/CNOMYoP
rp3ocffilZIszwAGAplMfi5HaFJoFGPegDdD+1H2gRQHhULTheHUnkS0q3WJARcp
6I1M5JUwvCRFRzXFnmrOfDs2VoGON/IZHFaNFllxDE9gXFZjghg/qOogp+cD04YU
CWvwzY58lSGCdZkVvqYtdfoEFWcX7nOT1nZ9F+K6S97ZkIv0f8ltaWYabgD3w1LD
X3JCiaX1kwD7yk+DDDaYwKLtiwm2FyVL6rcilIqvDS71XF9uWmcnOEPlh4E8lFrs
BfmvuwhgF5IMnX4L7qKBqwRCWVpZgUVjj4keRLLBoraOX4hNMhtQLRrGkAJ0JBqM
4frsoACpTVep8yG23DrGIp5uPthpW7qw6uYJn0OYIFvKZulb4uraaCF/IGxWUPsC
gdvuJDSQaN28BLBcls1hb/89PgkHwkFardnF3KT+/Z8RUSKa6cEvZhOcsPW5S1lY
v4jjH/eJic3SB8Fw5nTEGz6Lo2dLB7kxvz/XyqgiF2TsboEDWpF7BEvYpnED/Eo3
3FLun2FOZt7bdo65uPSKqHUnvaQV5xLQj64dpwkawnrRfTKKNuEiP7vE9b/LhKVh
8rJeejeei4ggcnkuddcws1caHq/b6TG8OtYmOVfXtA+6d4QLmqQvjpR38bHyxS0X
8UOHDtlC1K8aVqCjPu0UbybkWvWPNp08q8cC6mAN+eQQ6z9JZLLIF/zkYC37lAYB
kC38PXtwLljzQI1+4I4jtTNL801riKdr0+5xo4UCU9OQvGlkhEYQoLnxNfAPtb6g
oihjo6waPK6g1NCjyXJblU3JW/+1ZpFdcm/M9IyQeM62PFrEIogYFCeu2LxPC15k
jh/i4vS1cI6RdB1fseBDzAAlDrFNMiAz9pcgrzwTYAXsVgP1335tQZ2u6PRTGZkd
oH3pYyLg1Af08CY51BW6KuMLw/UOepbvd+iGUL8HRqPaJCAVZuLdYg3N/f8XY2a9
ph3mkG5SasZ6YWMxuTSVT7zAehmEfSawWxagU7eGla1Zb8ngkCP71q+//gJMDDIr
0jHBoVxCrKOZS/WCG0QHGcZUba0Zwra1I0VKplkNbfYntD3OAv1cgP0uryyjycs6
/vqBlaTtwkQIhkRZUu3W93Fo/8kV9x33Uuc8df7C6sPWheOLaZ6nJoEAx4yHw3Hz
N3HsQeaAuGCaQEkbfFc4LYqLHIevMb87vQPHW7dj2QCf2DCWapwH087c31J79tQL
Lk9RUFZodfl/On6sIA5D5juk1yifCykc1Pf1ZgDS5DrH6qdpyKgg0bjd3Rknl1eV
afv8uH5CFkhD5Pj6AbnMq+JexRnz1C1A/87BnoiMqUXK9LyCYC0DcRpqgT9oy2vY
ggP/Yhp1f8mhshhncJxK9zP3O2ffcjuuOVlE1pAa62kH9iMnbkNUhA86flyFR1Ie
VYNf4UAxMjvwxq1tzPO9xOzAFnM8k/sdlEgfB68lMo/zROeTfbQ+JtaXtV+KhB7W
l/a0a20xVvfW6/xFsJDnPoa2wJVCs3O2GCv4Q/1BJbFOXYu8ze85WNLrDj1kvLqS
eP5ReQuVB5uyqavnXPBFxh0nfHeihUjD8ffBvnERAUeTOeWxzWI3cFSl7e753Gyx
w9osN7tjaPoqSv1uOmKOZXb5xfzZKt6Hy5xp/uYTukkY4CR1BpJSDmxhCBh8hrp6
iTp1xEg5276GTjx88FGFBvS+w7WPWJksKO8QmB8YKuP6D55IZ4i9Ly56mcD+Rt6b
cbZT1LWhYZsGkkeRBjz9vo5jaLns+n0LoddPlsiMDOvPQ9Il78eIYeezvfS5YmYS
4ZuBNrgSaaM/3KM0TQuDqJ1zGMVM0gUDgnkZj2up5F7+BfjXB+cKugB08pLe07qs
c6r6HEdciJVCJcc4uxeQQWcYPtVm7x/H9U2H0dsBzIqwcYIw86E6UjzwcBsaWaNW
SjC5hiEDVOuSNeHehjvyvYxzIybrlWlBnkVX3xHAVulHqwBAeGPskLFnrvvD7J/r
yX3f5IEIIeVZXnlNECcH8bsJnkXPhPaSIifPNfUxp4bXlcaK4yxwYy9+NBeGza3W
M0KeRceUcB95+yGcmuxpZBfh8VnJEbgsXs1RjLYCNvhQzXy9u65bfPZ30X8238zO
DfcBZZ6Iw1s/yKQ8pYfWMO2HG5YVUEyOnUsFH15oE3wCZqTH4CY7i77JBPVv28ms
wriNfNoE3WildyLj3r8Eg+L4SMYmF2Xm8Tcex+vtuRtIs8dz+4HTASX4jmX1Aj9Q
KQ007qu2Z5ENDTHOG4+a+YEv+NfiOArJfmnSLe8b4wtr+CTz/M4B/TG3jxkTKgsP
IKMpLgbMzDPL1VqZihCKMmkzDzJw+sT6ccrbju1E8AtpFJ5ORBA6UM3dYypiXDYd
cOZsqV4dOQkdeZxBsycVJKJ9gy4EsMSiS2d3IytQVCQ5W5GDWeRftY2SfVg4d4gw
p5LN/tZFeG28BkeUQKWGe2nzEk2GZ14TRf6Irkd8Bk6YnR37MERz7ROJ277Xw/gH
TmsHWEH6AnoznfFVI61PzSeioa6cZV4rVmAaBNBh9N1IWiQMbf3iIvcaZoggrAnp
Q5DOBP6f/fQc7IzcbkZONwTeT1nx0qcHAwCrT6R5Toi5KfHysptd/Tc4xLtI3Yza
RMN+08XyqSIqwLEmnKwkEi/qPBpuSZfxH01cQIuLg+00BbzlyWQgUSe4huv0sN72
Jk6fpal30ehA76YF9JjQ2vIbX65vKCnHnTG1l8Wk+EXQuq5cAUfs1QUrliB2XR2J
0K6dfChxWOzUOn1pjomGu6R5v34/b495kgV1cIfaJUxUUPjBMfBr3I3CilSrCnXE
wW1vNyLiQO7mQ0WXFG4a0QDDp4beywb1iT93ooWg8YfV73NSPrhRTTRbaPQPxl5U
PcT6jNTOhAcQBrnUHUWkJXxti/7H6XrQrT1/xCeF3AwWsC/sCeM+BtrfzrK8wbzt
oyx+ipk2vVYAb6r/+BCCorZ3sSDkrSFlUGCB0nMYN2t7KSa6OUr/7GEL/oUSTBKL
UdgMvWXwvSq2e3LQRF7RXmLrJqlLdtC6MLPK2AKie4lBpZVjxV8wJDz5aaLkaEQu
YaiSeT6vZTbSuj2LgboUHgBX9y8EaQNurRrJ7we3tlek1cIjqFPCEFOd01890xCn
VHeJXUbrFxRm1bXNvBaUbfvqrWboNcej6T1fG9euW1GECGYpE7QElKdSEVelY88i
tivJTcXfNHdqStZEnAwfoCiJQevq6ixS0jLkGvkroXV1ZgEw9RgvXDHI0Q/2ntAX
tO3N7nwP8civyhnJjNceXv1OHF33oxi8obCXyCQsXgyFJ9qN0safHtN/08qE9HBW
CKH9vsJNONQ2neDCp93IPSs1GLXsiFuRXUSkWbeUvqIrMefoTl/kM33k7A5IZbdQ
mpJ7yToPmReYpQ734Qv3rXpvTjkXSaX2oBPL1n9e2+W8Ee+7CwKw4rbJskKyZo9f
b8ICx/ZxP6RO26voKhxBz1wyUa7U//EWBBac5v53rwkUats1FeHPdTgtoob/kOcY
2G0b6SexIP16oXNAbV7stfZZ8Ok7IZ43iHRG+Q0sU83HevuLaJzTMH3HnNYk9HVm
czNA+7J/GDKZnrJjZmS//RvdsIwqUyL7P5eXA/eQVnDfoq7jsie5or72TNfIf/9F
k+DFG0b1ba1Mh1Zoc2l1i7G+JGtCDlxwryg5BPNfDtNPURhmP5QCsrrm0r49yJ3i
yyOCKInRsfQlHopFXx1KQK4oTWCeCievco4695jXRBdlPc8DrxxJ8jX577VSS7ax
UCRo8ovrs1+LVns5ffxvDhIz4GbtrH97YG/HJ0FLW9y07ga+2zyhhd/CS5tDHGd5
fhhoZwrphTjZ/rL/KtsRLJE8IRoHqRpKG4dqy12n+h/pjj4cPj3ip+MR7mThelci
cnrCFYEWrLlmA5G/96nvXIQrz5iViGkoS+uVadNN2mZ/Gt5D91b+20yKJvj3Adw/
e1vqC/r+df34woq+xUIwZWc43kL+1KrxFliWGGn9TYq8tk5q/SIbCuMceMxHpQti
lqvR44x8YpIgYU6+WPjJ+KzTIutEcUN1u9eUejTsr4f2K1NQ0yG5ZA4N1+wwme+f
e2cTo4WEDmcKbe9T+QY5U5W5/0OKkLW9UIeRjwC/Re3BUCV4umacJmr6J7OvpqtQ
jRwbMI3WoMOs3xf8OodiTI9AQ0Z6+Ct4kOq+t6B9CEwpkkvcydZBfyrGZpvEpTCK
EImv0QzEDTKJyg7k8J7xbJD3prxuNCLYqGmZqA/d3z+okQmayPuwLG/fw3PbwCwz
vmy5woHV4u8BaNaU6OF9ljSOj5ek5gklXUIQo1RYJVEYS8XNzrbS86ap3Az4091m
GQlzYISc+Px3O3QSAnt7N0xScImDHJPJx8WwUdYabrOMT1TPtXiR4yTu8TFn1B2h
EMNhMhlbjYSnfkZ0CKXuTJnKRsE1DJYZlK6yMLp0992qkAsM82omzbwghXV37HOO
Zyju2OpxTmcg2GrAjhr84mECiZaQnqj8QSYmOXoPwVP36Bcp1t4a9UC01qI3Af6Y
br9TUrChnIjKcUnKeWjiq/98HwJ3c4sHXMopQ1fgs0o5hnIbiPwB89pqlwUsPsbf
nCCGVAg8wGQSQUjSAfyQg/gqX/ckN6sX6NsHFfDvKkeOfXX+SdtixjeyBhmdg8vW
yf49nspixpOY3k5+fTOYlb7oo0NAx20AgBVK19dJybV/6cIRHDSGxt4wvP/pg88c
mVReVp2hdDUQtEPaHdSiV/Zs+X4J2/VPTpvT5lOWgJyC05dl4f7a0voh6sgp1XWX
dBOP7D5xYhNwwxFFcZWsODIpx1UVatdsdKhYKUY9P/tJmEqLHr/I2s7zDm1NFd4d
/QmVmf/vmaFIbsCF0qEK/jaVTmX5wprua5jYL7cD/CL1IkuaK3MEWvjSNz+QdQdp
iLa4pCo2dwEK3pXRnEF9PN7CIm2/vvhEVDlE6MI21f4ZPhtwf9OoKeb8J3MX6kuy
0Uhk/wonrAusCK15aczh6aujTqG+avnVednQJ7itOmMsAdbVOfkNYizP5ufmPa/7
2jlIb6Is6tt1yOwTQRD0w0mwd272Yrb+GTGwzsFG3UQjwPePn7SMFwyZeCylqimW
AXkky0bhQa0L2cVkj1dLv0r4TDxIG1W5E34yeio/RKruRuXDO5CDA0gHCLwwixYw
PgRPc2a0t3vdcG+EGlOicvWyi/aOSSaeEdWznY1VSJyolBMuKvJvHQ6N6Vrbehg6
mTpBoeDy5PmbtHIjmpaIWW1DMXIRdJCeBLtev8Scu5B8Rz1fXsYT7lFgcgGJLr7F
1wRIZqmTvodqrxaIIllU6dJnfRgRGxVmFwR+/YsC8eaHlkUv+0bm4GI+pSKGfqK8
OygaK+XuZzukp5DEgwCG7SGU0UsFYHc0oSafymkibgd53nR+IPI6aDvNlzHYPXf7
Psbet54KGA9JKBoKm92X6TkmwFvqqadU2YxXwCiDd2zXJovr+w51OhSxWs1pEvRB
qs7QPTeN68J6yk/e4dphenTvFcKJxPWzgut0gMnH7reojdY/pCgvPQo5vubs45yi
oUnSb+lo04FaxkB75nWz6DSn74mAZgAO7ngf4vVX4+LGWQg+wWQ0x5hf5blIO3YG
3BaKYqKSnOWZyYoimxelERT9MOwDNs/i3MvsY0K4AkhlJP37uh6VuD5I5yZOOhcq
LNjO4jyFuGWJF5RIZiS256QFB+MO5pbwd6mCCe1W1u7nqxVWP9HAH9Llo0c6XGOM
Nf9cwkz2IclwssIAL2oF0aDCZ8wiWqhdPQ9bRDN5auv9h6w8VtdPjZrMSeT9+T/H
5IYrsfo5wtizAQeaOxgixcc/Paz4dpT2y1kBXX5xOjEPc0tb5FtMthJLmZQmmPd7
rHajfAW+nhilBAlZT2uW/hY7162gZyFJMCIei+WNBhNK9752R7W4cTSbxonYOa8a
Xicdhm3y0HkcqYD9r1KAdSuKBbO0VURdC2N1nOptMeiDHQ34xEsuISZutXR6QJvS
p7335RcWhaB3WEfpfO1WnRy9J8GAAPDZf0kjqigPeNAv8CRNcjE0fAZk96Geu8yE
ZCHCk+FtaDN35TjZHUP3yNVHKvIt36PG2xQhiPmn+/sNXu36w14QuJXDQ07ESF8u
16z5Uu3rViJr0gLy9zvj+foZ1dzJ/EkvDXRgPTPerNLlu+m/2OsZcVkjz16Sjqmh
LdchiNkZSK0aAvp0dGAGYhnoSH1LC3IyTXBObB2Fu7HaZPbWKeDaz7SY7BnLWISq
Tx5oueFQ5BYBI573l0+hLOa3tmJLXHNv1c5yltvYjdzQf6006qy8kyo1AcfdU3Vi
6067gHXDdsyfRrZfyJibIDcdq0x7CPUEg+878rX4HC7eljhUH1uZNZy0Vg4MfDME
p9JI2f0l8P7ZNl+Iq5b+i3KJg21ajJvN0vB1IpJKxH6+eQIaahSU7hKBAnTUIlf0
jBEELqIEe874aqkMAl0atDRp9BBNXxdeWbTJMhtFVMhgzUqxD7rreWehlXF2/hD/
tmvz0lYZCb7y4xowYRvDXRIkscaroqN2GP5A1oGm3NBowxM5BR2NGm2pFUN6SEr7
vWs/JOcjwQ3NNNteRMxBr87tm5XsmYBhPX6ayDkTj5GGgP4VijmKk0XwzWTLWILd
3OuMx9dOKs3amgFOfk0Qx/mPZwbM/CRrZXUUNq0faJ4eU0CnuIirdXy+RMzWSuv3
aQBcwKvJJGlGyGkzPVG80Lwwx51C2mfd2xEHKZ/7x7SyGTjxTu51fdMyOc5QdHfz
I5+LyuqD0r7F6h39WUvgAu3s+j5UG1+Utp6KL+idKhFet5VHgSN6w+ZmcMoM2bkp
/kXLJHvNMjyKCgyabqpa/iKXENAEPF7CxBGykMBzoX8MnPVr/yzGANWa7XC7zC0v
qFsWwjssQCcyiCoSwnTHsNj5y2EBkbhTaMb43eFE7oStG46fnXcIIn5mEsrtidv9
Sj0TRI5rdDKJf4P+Q6RRPSkLqIJkSIdnu8RhXydtyENsP02cvgdPvyAI+nryVxWY
NVRFJDA2ai/lxSNmhTLLRqiuRNdY7JAt43U/8aWduGH4DHJf8Skh+1kkIi9kwKsL
9pFYxhW/BK8f9FZH5o4meUpiMMKfVWC0ZysYZF0i86EksHeuprQYxTumjHv6XVBE
wVbnbBMfeuoxPjHKoxcN7mnlhqdWVDZdedmhMeiMGTNb+hdgHmAZzOSKqNSbdJ88
SoqcB4fMaHA3MNbvXVtNlaxhqVvfQJkQm6UGY3/QQgsw6tpGEjsku5hVHjta1OJP
1Z3DL+kjju3q2NCkXJQt6BtyT3UjFzRLJIddjRPo8XNO/FGOtc2Ai+HmeKJvV28i
2DUBsK99P8r8yH5aMPLMfidlU5ctix6T/dd8eBE/uNpc+3vN+oyiwYlnKfPLj9Jq
PUyoOyycH6FXTrIeqUTl3oLacuViDO/tFcQpC8kKG9cfnwm3q1K2gG1qI89sOmtt
DU0tTERATiXoN+dQJsZEs3+J7vZWVMspXaCXWmoqJ87vp4B1tNOOJY8N3/4HR0X2
EPzQGXdq+inDq+foq/XD7JWP+DqVZ657Qr8GkAlv2DgkIgPnx3M79RKnMN5ahglW
XpT2H5CvL1plhJJ7go3cYL3RR8zRVxUa981xV5pYEd3uUbuSX2mh3ln6xvs6qZci
dm7s117pOkGZlb51WPPbHxIX+bZ1NvT1Ozx0YYQhsbLJfPLL4f/PDSnoxvR52Avy
XpYi5TYZdu8OrgRxHkd44+gwneQkLVv6bqXSM+fdA3rPYwIs08JbDaxgGq+DNnCC
zzKePJsiSd50bI7bKUAXuG+cmqMZvFEXxWUkUPb0faGo9m7Sk8PplNDq3oTvxUmB
Nqm4pRRBvGMpF6Rrz4TRXaf5Hy91gI3RlWu6pw8ZeKHpzY0ZqA4mJrDsRhQGRAZf
xaB03ohzKrsQBtyLAUk238IsBqYCbtRc38iJUsXeakdEIpKlBhFkyHPaev5g5E++
BKNLqDZOoVxzZ4AcTnASemyaody6jlgKibWHUOpl8/rSxx1e0TM8iZXy4SwmNl6l
xDUrlZB5g/dyUs4xSfYxKqaPmtMRArpGOCuvv31p7P1HVje+RC2eo7diB4vwGJyu
jpi0isZZZgdQgsJ0CSVuFA/rG6KmAIJ4v+ZaKp2KRD8HoFXfRNaukWbA00mUPbWE
5bhfPQE3oPSIQoQLYlL085pB7tjcM6vWYJieSSOw45HT95DcoIm3cIGrxvMXtvBA
iv9a/XVxFvfr6/VAZ2ZIuS1ofyf0/jwMHq9BgE99+rwpf5nOBmN5a9lvB3VHvg5s
1s2iueh3FqHr3T+Cr9ib86hVXvIH9NDh0t4pD+jddb5LWdsVx4fmr/2/eYyE0RBa
OsvP60Gb7BVShrGZRuI3ZWlUNSMv393fQSsil2yA1b2AO7pSO+aLt7OnaoABsJhD
dXa3SXpuwUmguVqnVUZLHSJivo4kDvG9Okw2lYb8cngrBKUUL4z42ILcFpzP44RF
t+X8SxIkOVu7nZJnSM3Fr9oLuT3QN17dTAhefZ32uhz55xC7DWbO3Hvt15zyKMfF
sgq9v4lGhYZgw7eGEcf96Z6AL4eGiQg5aYnmhwk2PEUsN7ubji/P01cr5NxdxAeE
cmpFBJtfBt25mv0JnlpyGJLCzY4pVg7nECgKopbmApqOZao+d2KFhmLBrO99gtV8
+snqcnr6bDETT3OiuLMOv6KkKuyIJXclNnppPX782TKWm2cEIgXqrKjpJ6Myzq/q
zJ4o7iMdvmcyNaavhxJni55k7dVB7I4BOHffPePRXF+PAv2cACbCUMvUEE4Ab7nQ
uKi5WTDFYh5wOVkLuix81650XalAvgr/qEoCBhVQ+QxOnODM5Jlr4UjSevf+0cro
ItH3K2ve4+9d+oBcLlb5Z9cyg5D+VwfTpwSKMgj2K+IHtarBgPCwFGXeuErDD5gV
Qh/046trbwa7qK2761oKSJe3gx9E0cz9DqhaVOil0gooD57RcoH0g3Cd1XgK9Tfa
ypPAGV0rcwNrjDQnfVxtTgHzTWsVqHdTBK43KR9ArXkzx7GDRI5hnRpSuU/bgzSJ
10aZXpvVWjzVh9gbFu4Mte1bu4bE+xc0/sXh5cl2tsInlOSZeGQ91JghHFgV8Yx3
9qTYH6AZywfJD36YYeXPenq/er4P7/jW91Bfv3NYuOFrFzKO5N8mO8nVasgjMdWZ
GPh/ixtPn6m1wUwyHJ9nuiGkLOxKWPD2xEfmvGQ2ki91tJ+tWfHZFcN1775fFhTi
OIgempIGPjYxzqYkvWmxcZoin2/cd8liSkapV5JHEYrWSl3PAYJ3I1+/pL1dOIOk
jpbmVf0Z14cGWfdnRyOpFRf/I3HAg9knfxNotLTFwMreTWh6gsa2Fy874gGh3GSw
yObD9KDsRgymme8sWm+AZsQSIgbeHs2K9aK52Uw6wpMcndtnlfnwS51koJcWWpm/
xBiDSbCFyEuAD7wkfgNUPJ81ySo316YJUO8G3y6D3ZDRWf7a26necS3aSvDKegep
yxbCU4Noz0yt2Nw2u+JoR1s8WIwT6FgOfR2mKljhr3bcsDgCeQ1dvi+r3b4RQOUG
a9AYyxrZ4CP9vZ/AEukkiayR6xdpPIC3P0fmyQr8gd+7WLjMxaZRW0dwB6ibJsH3
728msoTPH4rQm4/gNFD7I9YoR+v7nhSDQoPXW5/JEDxeK6Q1q/pfuhNSjvC5hzuF
BzBkvjKK4eg6wmQja3w9DaCUxhgaoCagljW9L0N0WFFn4WtluaLp6eHm+fBlQ0/Y
RPpz3ickz5aTSZHMHfUxWm+VFQS1g3Wy7k9XmvYv20H8mUSRXu9egVdnULxY2b92
DieRQn743OrB/W558YYg2uXdC6TxZFFJ8QPoc/4JTJXfV5/FgAnu7RRgQu6WmLMs
/77AL6OaG2R1oysly0j74Lj1cpOKAHhCC/GqnNWnltrmgoUP3YOorG7Wj8DZJS5e
JZpaOuJfCF4cehSY+6U946bNgbSmoRi7P+jGD6sTOEvZ9m9X8OIFU+MEtx21gctF
2/pkLmq9G+eS5/dRfTMVVovqGuLKueLOqwhUvRmopBwEfHdTGepqr3g7FDKprZRt
ae2XHSfhXwviOtlwKg1Bv4ywEan4Zdn0aChdf9Rruh/lwrxetTJrmZrf0WWLi92Q
mDDXq6xCvxxI0jCbQhbEK5wuIO7nah82X7UejgTYiScpQdMq2XeAbRr5jpK6v7G2
a9uF5KTel/o/eMetoO0jISZagCY8urZdCGl+m01zqACqtiWf8uWFonWGPvVRTHU0
LKXKYzKNas8XpcBBYC9YlesF7gpVIufSPh6fAgPWYHBdBIvI7usrVulle5q8tdaM
1+CPVH5i4Xe46u0xyqnx2hFHKYowzGyUM2dL3S7iGIV/S0xKlHCQFFIqBLXBXjwj
YYilH0aSM7rY/37nCCa5bwdbV3z+hgV/jJTcpDpcZhUhj96EiGJAjUh9kk7zpCw6
eAR1akeTO4iXUYdIf1i1Ui9d01rdQh1hZRO1WlWOPVj92CKmXBpsfQ5uc2jitGAX
WnC9ETKVKW0wUXgCf87g/GvxekZg5jADgWjk2oT0guo86x5Nhl1cm3dAFjcp3qCQ
1toSHoykGUBxgNjF8PXHuuKFc+7SW8dW3y/e2Stpe/lACyzCJxiwbiRkV86f5cfd
95RdpOk4rjqlm/UUQS7jD4InB6ocfsZvYelyK+56mQVsJAfJCK7cQfCJnclYdH9E
RrBoO+h8kQRNQS1pVfE476Y729O8i7qH9MtmX2UaYRor0+1ZQJD0Ra3G1svcdIDH
el3AvyCUoLCdwkW6Dm5eq8Cdy6BMzsLmKvFx9yvR/dZCF5kjjq16f4Zs5tARGZYf
K8JSW6a4+JPYDiHz3lDyOyMHJmAypUxV6ZHGHVPN3FkzJBy/bE0JLChVy/P5hBAY
gZ86TwdkWbcSadwvB3D87UwiQoan/BJ0blnT/NahJqKCW+944snBIHxBX5yfPQQ3
Sn50LsM869EozyK6DHiGsrrL5I5actU/uDPDhCBXSj7Mdzhb8C3vAYjph7yMF+zw
6h46w+x7FspReYIrJv4eJmHbLbmd8Jm3DfvulasRqh2ZZwnTQRFOkqVus9flr6pf
GeyCkH40MoAMakQTR9zyeSts8zkMersih6THgBSJHxHzVefrrBVtixwNg6jrniGh
qlo08AkRJs7Y7DDggZlC8mZ93rUmKYy9WorB2r7SZ+GjPbHOeRYOAMc9pyMJQVbf
C97kY3GC3dqjeBLqryJHtJOpU1PR0G1dFbs3DGGqqVqg09ZiC2JrB8SWyjh8BXhW
cCsfG7teybKCZ43HWK/mA+q/1M8OsjL0t7mtx4DZfdyVVukqJ6i0qOx2QfrDRXhh
WRdt7zfxooPFS6eY9aU2G3SxY8v9b2oP1amPVx++T85imspgvKkq4XCauyeZxo1v
YIbYCwsD5J+wmpcyO2RpZ+FLHYnxUkygkDCMjwL/u6jO5PIT/nnwVa1QLRNQDUve
m0U1dDAc8VfixCVSB8UDG+ZRH6BJcgD5/lUtx8ZvTVCr+7bc+VzBzOVFRctt55Dy
M73dTImNW3P+RkwZwBQ1zqjHpaufOTpElt+W7unPwABgSb1Elg1kzXnmKMqF6Sj3
4Vr1D6w6QFflMLzvXQxyjeizQzdsbcYixEChN9f0xjs8LxNFKfI0wF5bMaeLfCQs
uUd0IKcBJ3i7nqqIddKFTFNbvm+B9Ckrt95ZyVFAi7mXdzjzGfKjy7EaTE5Sd5b2
WtnMPBRV/H63vUifs7mcCyBTLttA8K9K7CEHAR1cChwjQbN4DBhqjAC4iFKj2REt
2gBJS2wVdMcGa5s3PbwS/gUlbYKwY+9XrGi5KYmqxjbi6HVDbUcbdH5vDgDgAIOZ
z4PoDcVZ1+ExTocPCkoj9ZH9ZJKSxqPehQZa/BYCyZ3CAU0/oIq6IScyEdWocIO4
uSmKQ2FZ4acSjsVMEPy7olh20d8+iyq7jtNCkASMyaMfOp16Jzl0kbGdMMaL8sud
NPRFLb2VX1OKSLrTr4+r5IR83Uef67MY2xt3Xiz7xy7TSYrx5FKI2UHJ2uImWQaj
+W/RRslCEuscey3H43G+tKXDMkFK3MuhyDAZ7msHL39E/yAIxAiLoOxf2BULl0r0
QSdBJ0nVPRP+4ldbAJvQeqiEY2LDSzSLnh49eRoOphUadl1zQQp1FbWaGnLRNIaO
Kbpw47/rC+TMem82UC4+zef3ceyIj+uKpmkBkagwlt+TuY6BY+ur8UiA7MU4CjwM
ADucAVRRdOud588ZR2icV2dynMldjg3jCw574JlG1Mkrlrnol2OwVsc2whYnzeez
I5SnqGc7iOhv9TU/t+mIOf9EVMWOvxnFaptUUWXNa79I5F+uOUYbdaY6L0HkF1NC
Ys+x5cASvRkKKU3sm2vvpoZVUEIdHzAoHph6Lmu1pxF5irs4t7gUf1Ah/i7g2/lh
e691iDUTfs1jaYLssMSsZzWyx8M5aat0JcOIw8TPyybkc/YL1kXqP9NdJk6xn9DY
/YmJyMbWUXZj7G4hG5He8UiFSFapFjvy0923jYTwUiw59dFUxgCe+stggmp5qv+8
kEbWj3CpC9goCSs3lhd/RtHVKqDUhT3B+Y2gLsb/FqCNGHAfRz516eRLwb972EpE
rmAAPn9Zqm971NDv7xXrGZmVySK3y6b51bpP5s4YkYz1OU4uo/I4WYvDjAjatxOK
2SxvOVmIbGTtE3jCg6B6aIFytIszZ7kS5dMsxroQFUXqkvBRuNG43hI1+WRh4VDo
arcK2PxtRYTPJ5Bsk5pmGDNdKhTv1haU6sqmBGLwPJy79jCu4UsSfl5XQvcQJSMB
GR7Kz5RxG8HEESZhDMPctGEwvQWMwIqL2Ej6izvzEQXZNF9NNdTGUj3og2PeVEZE
dlosk+mJauYCJf+UiT6EaxBErq0RNwFgXM4TqILbtPnNKGmw0uc6EWloMRCgSWyL
+pnTj3jXHguQfDlDU2SdpB5yRjuHEab5QhjvVsX7BOZmZXLb/W1ciCcokvHFl3MK
MjBnjHmYDVmHszshKDycWHHywEqsUcXJcCy5Th+8MNkIk+QUyQkAwPHta0MXgO1T
giVBeVZpKtlaHBu9KKoci0+Sj0gD7AcbWiq9NBpc+wCicTKTBop+rddGloGmbIvK
GyewY82xGeAwZE2A019CRTnnJ91AKtW//UmNJGNSFX6xiudm7bdnPmv3/wDlPt7F
FArhRp+gQnOwSzPMcL0yEjEjgNoYFiBTB04gXHAGF92KOPhWr3/84YN52mt4ep7R
r3RNaqyOYuw763Ruyp1gvQMaq/kHSNuAt/Xka5QPBkbVmji3kVeVYkdHiegXvdJa
6305MmFfhm/eh5EHkWXmK5Wcgno6tkJJAVnSOLZosUSbFtSB53rN3uIXVYavHVRI
FVfg3FI/Sm7pI/MdtPYy6yXMsA4lR6lKRqYETu6ANWYPowanAe/HBJGQ5OEH5TXc
DJFNC5lBqQq1nR2u74XeCHOM5rBMcTZ9q1uxX1327ymEoAHjyv7itFsPMlnJA7//
n+nbtAoL1LwmMqdBrHiN0HmF4LNKFGkpZFgTspnOAzfGXZGujF3X78M9cHD9/E/e
UonwmsK5Sz6Lu3fWoiSovVvoG/KCzPoOAoz/JOFTB9YprEZqvGp8skUENZ5TeK3y
doBXmWVyD0F47NB1Vq/6uXIWntvmCgRyvIf1Hh+MjLIR3+A5V6kTGBPMqTsK6Ps7
6HUO/lX2weHnWaYdbQAK+2GBTKC9VDuOV3+jlPo8BaRik0iHKXXK3YPO1KEIHRh5
zc1sm+Hh8L6WW1O4XTM+Lm5Pnp912mK3W4p58jc/U4AwJbrZBHIEy1xSGQ0Dfpc5
4NK+UruXwQO5woJOzb/qbb80qJDqDGct8xEk5jNbRpQ99sBQy9PsZm3wliyNPkjU
DDhrecTAc1U5k7tEKRPgwSdH1Rp6C7RjXBPYMEHb9TSiz2FhojVO0170xDY4Th5B
wMdnszVKNSR2d3XrOOPzLgrTpxXlhWgbIVd7prJ60tqJwo5LckbYDNe4RPVVlYDg
pwc4/a/OzM/F3I/3hvoXA+V5Szup38VwOf41JhHB77iXZfr8jS+3Y4ZgtjTgmKpe
GMhy3X57sFHWAMxZ7cg68jdjKiL9SnDgkGPZd9jcHNchbJ64yVlnjLu5IjmMMse7
GgLL5EY6jS2KZdSuiNqW5xUu/2151mpdy9IKw0zHgNoBI/NAmdIGZkKA5R9Fe5n5
f1Gn7FmEwF9333CRvEA2fo+29tqnnox+mpRaEvF+U05Y9sGVAykYmoJsYHCDa6Uq
/0udzQjLJWAwx0mpoHX9lqy6IwInDn5pkXzQMOX7kq9rQfBb1SfTA4Jf/XESbnVt
wD8wf5d28nm04706ny0+UWUXNZLkdUacuAaBnAPDg36OgqLD92PPDl6KcNPo+ZcK
Fg9Knr1a7Kyc6lUNRxQrLbU66pihPTSUHUn0UVgMrPk/UjJElm0eCAarY+GbxvrA
aquccJ7BCZgXhHqp/m7QwDSliyEY9seTrL+Z1sMmSnvSlzC9tW1n2Y0zfd9VPXK4
ZJw9gMLT6rfijme43zO0QDZ7Ibls0lOqsSHiWXpyx6Cp3HJBSQ6zDSEK1Pyx/SfW
vWK08RZ2I9n1jZDsCqCH+Z+xcT9L8VKQmTRu1ouu+Crkl7PP6bXDxyu3kiWmPRyh
G8Ntl2Bf7K4AJSF9nefXLsWbhS9qDN2MFUUZ220mL3rLSphKdXEapvVICxc6E1E8
XtasQ841c96lfUTXlU7+sI3KUpmCFwjbnDPIvv/3df7Khwi3PheI29ivQVCNHLng
Yj1Y0mHQ3t6tAQMLWRdixVVc13YBfAwT6bt710I5dyGmHuZ9qZHvt6Ti1WUoYmBW
6ev6gmmnleambUDbP+3ecw3m7vlGaM9yDiseWVHeGLXADy8uKWzcj02tDyPTOsnv
6WpIjiLrktZUxNE9gbvkUBGyALZqvdrLyiEEdeu/+KPEpoNt+MqYGLjbuSAqZmed
ybzCZ/rtt0Io2Hc/6zxr6StAoiJ7vg5eg4t4GiXnNL5eRX7/JFiJqXlYV/LUZCqr
HfKQxN7Xof0a05Yzc28CX7k2W/kNU/Eb/TqxXHB1qZthxaX0+7qtRLnCCvBz5Fu3
a6f0sOsjF1WEqsV1JHVA4hz62mjSSjtBroX1DtrNKifDC6Ls+qs1w3fGxi5Llr6l
eOaZhVemeZJ2xPvggIx7zjJAjb9wE+aYrpq7W+wtMRKSMYL4/+gfliFUH2pWo/pO
VF7iWot4ixiMUMcHBSyFIgMvtXZzNHEUWaAvMKNCT3jJUNmbNZLqQ0/Sn11IgI2G
L6Ob5GY/0VQO89VHvqpumpY4GjtZN03azfvnCqIDot9cvAZkliRNKEUHxE/4lhrg
IfYmo5e+rUvD9MlzzY73WzwqoVfcTmb/iybY7wRLe5nLU6D6wOvVo3q/c9LP2ZhT
65RaahZcntAut7WsYqky+fnqsLSs77uXxicxX/DqLBLMZ7J+sI6Sb58nDCABBeK8
tbGFZ4UWDNe3TaNjp+cbDZdPvSWPH0KHJR8WFcDl860uMewXiuN16DorOex0aAxN
KUD6c0gD0F6m5YfxPU3Tpzx042zlyigJyOVzFu16h/t+vAVhayZ7afPgrkMJsjq3
U3bGpLgKnrC+RWrvC9YZQfQgDRnqs7hniiWJDXSFu7p8I1WBR2bAUnqbOSh2WFOL
oXbXKKdtqGjNo21lWhnSf1NAAXnUQnEYOggVzkw0mHiFgr2fkjM1sgdGdsFh/lem
NRzi3CuctRCiiTiIgGoBZVGp3Blo3ypjKuymZZ/RgT2GREbZhYipeOAh8Ng+Of+b
cYpDTJWZCdCUYSaKTRSXzQd/6awBLYb58NgZDcqNgcwKa4DHdluk6S0Jw4zflx1V
t+HKRYgH1VgurL9JeZJ1IAIlZjB9Kj2IAwwslhiGX7Esi4DinLFC2T1p+64bfJXV
Pp6uUAeHqAarIq0IpkMKlzEgFEZtl9s0upLN0yBJaN7uRQWomiUnYRagjUxyNAjv
IALE0tjsscXxGnw9tHpxrQXaJ4p+a3UoW7/jxTP99N+XFQVCwwT7ZdRUlDEff3y6
iOZdgW6vwlK537fbfLTRjhAz6Wu4uTAQVXrx5SjPVVqIjFBuBneL8D7X27CyHnUV
KMspy/qVhxt1peogova2K3hHye8KGp4Js7tA5fbpriX1+XCb3ChmPvObDxIgWxb9
RvK/CRhk2LR2Z38h9yNEdtYoGm22YMmYCVYDo+UA2kBFKOjuh+Z82F067YdGMFpf
kGT53mGda+A5GNAbjKM6K1jIaAAJWerB8OMUbj27AB/Ub0kzxYqDP1oNL8wDIbS4
51EuKKjOgHfR9qhfx9UDbtxGo31ndGlFQ4/N2BHlNesBGT4kvWmh5aRTLKruyuHx
l5tN/3ONmlajBYs0i3wG3ieq2jaOR/idN3aD8B3JZuQcpfCZat3d5W8IxsRM6Djf
NZbee5QhIJ0sevgbKDGtZoAaa9i+LEjIgxg9Zgg0Y/zh5LlABv8TwvJwnfIVsv+9
i7bvJ6JnsYV8eJ9H/ufonPtQyYOdHBXMCFXTESwRAyBPQZ903R/IpUUNqlwdUx5/
+ea7XS3G3h0Wd7eD9D33KDHVIGaxEU6HtSDnNjZBbcUTtOZZI5vex/rZvsjU4kDU
7JiZC5TQqtf7CHKPJxc/69giHJOGxTewwkckYn+CVFB81vZA7iPPUDCSilNyewDq
xrp+Y+UAzLbud3aHgEF/zoM8RO0zfUr2mUvHsM47ladNStjLLNc2h3Z+3F2fzATg
XN5evkfvfCp6FPCFTjuwWDaKiI0ZXn6W9SIHbVdBl+TaEOQjuhnOLL15iOizo3GJ
yJmBwDpxNPcUtUFUzu4VcptXh4zA2J++Cb89SFUJuO7gqtevJOCmgcH697Jr2g4T
I4vCTXOZ2nLwKpMM3KJxPg8neJ9We33Qd9jXhKfYnnEq6knUCjN5iqW3+/cnT9XX
6FYxv4rSXz5xKPvqDMsKmzUtrQ9zvHsQHOifFIzqZXZpP+eiBYJzElMQ4NiKLHqj
0hLTYAm69y8kKmZyEbu15P25MoKqc1JFHNyntH45tjmzc+9+J8hOvS9PwzyU/gr6
8zLmlWCxy2mbwi9l51zMdmvlozak/Kf/AVzVrL4tJSa1eZfynPWRBWluOh6bw2P2
vhdPmp866F+fSlsxxXOGP7xhKIg8l3//ezhFlLas2fpwDLataTA0PbEMr5RMqHRZ
CA+4jkteDL6gMYeXmAOeJPKYheIXFCBnMTfsPzWeE6dg9n+e7XniCsfpcfWg7FsC
FzjdIOciuz1R5sMmJZVFLSRWCi34DH8NuLKUs4ohx37C+IpTb5h4Nvl+o2ZMZ/4R
rfHGh0DEt8a0QuiHoW+AaPk26sMRB6R/X49oRz4K6t0L+y+HFpm0fbiWFa1PGoMx
TK3CGFSeQciXSRLZAXu416MOrc2+3H5WspzRAroYtba8UYTmYJYsultKHsy6Yszv
uDFQPraco+7+/1lnltp1BSPML8m6yFhsGSP1Hvzaque7tiEm0XmkySYkEf6GzYng
xIxMUHUDxeGBnAQYs/xkqv/gtxUeVxnxa0lKPLBHYGvIIC4VTOOyB3/7BinUCwj8
xybIcxsY1GM2BJvfVUUtgaExXVDoVA4K9dCaPzllTULSfF3Vws3jXOesRCFdTtyh
oevbDVGtUqzQjTiIAcFoNBFlNzyrj+gL7aWLsU24xqMDfr3vzonEVBy/nQQomHoe
zJwRNtdpo3Fnj0daqmgjHYg71RBja28Yr8HpLIsA/J9jlyAabo1YDFRlndKc+JqN
uJSypdzxypRfTw3izG+EbG9wTR1ImU/35fSbVh9TrCTwfCLHLOSPNxYlOay1jTu5
yy0gzoV7V4gX0XarjvbyzWMAy+sasFqWW8w9R+7Ehh8XdX1d3zNJL5nqY2B65BCy
8QGCkDTy3XDh5StEASTavO8uJz/GDh4ovtrCT8bQstNCbMzouG0n06Wxb3l+kNWu
POwOMafgg+ukxE+IoIdCMLLh234BVfza2hn+Jg2quuUqI+DEd4wBL8/xNMAkgdVa
IjxGUwOuzG6vdZsqkMCelpB9QPeWBGKipPh55xnUxIxeULHD1rT4sNzUybw4rNDw
12b/SU7B1gjxKW6vpR0563C0LoeJzNGX0pKGzXm8r2uTMIS/zrGM/XCAvM9T7UG9
+vreYztT8cSA5hOcH4+QDiQgRYvY6ofA80sNjtyZs6yMQqo6fPRLGUBYNiSwbAjV
8F8w+Wx985AmQtk21jd3XM3Ftk6B/C9BbJAA2mM1lOcPqbAGaGV9elu6+/Xi5Ckw
+sNXSVT66rpukvhLts9jIaf6DRV57icAl8jwP4/DHhvoyajxktcBbrsNPp4k4yRL
B88hLL5ro84reoYwe1tr9I6ZgQ2b3WZ1LcDfT8cEI2pd5vSsTkBluUUNJb/KGavt
T/65MXSHqQae5v2iIX25NzYNv1Ox+Sc0KaP71KZWkRb8G6rjNEPNdGrj4Tf2lyb/
FJ9oRjyTvLmTXjl81bmwZq53Z5z7x2nH8o0/4hg4MHXsnwtsm2oa9Spqp7deThni
1BWWwidgr4Tj8Bl142AE6nRlp0HIO8GWB1atHJnYHVygI12ZufsniB9t1J4YXN5d
Ka8JQAUR+hFPSPGH8INgBmag9ppZj2hLT29r8szJ8A7daUMUOLVZIt+xxasFq7lZ
438lO1/GA4DKJtL0oe6mt0IcnH/ID2wsoehvT7JPFodniSemrNHXy+7S8IellJFv
bADbNB6VhUQPg9fwepnYKpGMuIfugKeIDkADfOfC72Tx/mp3LB4/9c4TMRbBFZ2u
KhiZ4esLnfXdWCVPtC0r5UG/aU+rrbJKHTl4jesfqnZV+w7k/Z1D1bNZcB9pWc7e
1E0KtyVXS5ZQLj+BFKU0Ke+dc1SsG4z7pQWYz56l+xfiVMFWSA65+UGox/UsXqKn
9fjuL1WZkR6VeCZLx0F5oJeXl1fBsMsX8XyLCklrzemmsFynKcx3vFWhgyIQn9zI
F0OcQuLRPiqG+z5UWONgkMC8yRxJ7oh8xc4opfkkXifI6rOwI5dV8URmTkr8EaSM
2BEvfpEGj1bazoNvAqMwdlNz0PgvTJ/DOFvOXLkWBknWx6QcY0QgtlILv/Malb9M
Ce4ELJmUfwqzbABiiFwo8UBSaWugz8EcfUp+wWjqjc0UCEZ7C67XYfVxMateUB96
ru1oWdnkzZWaz+ExZfeqFe3vr5XeOFdWE5gt6pMNwQWMeOsxxJK+RV7LP/jhckfa
cklzu4GVKLm+CJp8lC+rlQooqmL/vOFx6bDb1lcAi4VGiqz/HX8MWxkxxCAMQj/b
3ymX7jtY/GyGeS1njDa+81wqj9PQDlbGOSywi707nBUQDA1sv2p1vvq3AmLp9gNq
+2VGIXHmtD6nAEbqlHqIHDGIe49fsOCRQ3Lxj9smZbtOMJyGI1VqGrCxX9bjabPv
cBgF1aMaqDzl5ubaRSvGPX31XKYe/LxokuFJjMeDB57XwzO9Fginl/JLWyDFcCO0
zbISwZM1F53sVgGTtp6Jy1pDCjD5D241uUmXYa9vEiQ4kl6TNVQxNxyVDORRCpOb
v0V0h9SzSvo1ISkyklbGNmtv5WonwHOVC1q6gPiqXUT7IRBk3z3d3r0aufKrodDr
pzgJ9+cRmYOGNxGIGeCpD8xSL8zIRWQI9+P0o/2MQCALCXdAQrUjCKD/3SMzZqvT
xOACkgOZiCd/2XjYp5nUb23JLL4h6eUy+OZRMW3HxMbbH9q6HIfCTR9wC0dTlz4L
NQKGJbXsHHpcwSI8IeOn/wZHwqWGi+FKSkNGTI4XMheKL8JzLJUCsHX2cV0MLgJK
Iu4GDpHuzQUnAX/LXhH9U55b2esY6f13AP1taKxdL8NYs18LMybwVAyObyebFgnE
ZpB9IjQRBLoFzoEHkhR4K6WRPIllV1dTAgX0eHtoqTwKi/DkQyQKlMJI5qFngaGy
LADDILxpUZa5hUtLVbTNtp3JlpzZr2a97Hje/oiBwb5KoULxxr22yLlDMUeVPHkd
0x5OBg/9ccxM7JLATS+dt0pdu21siqYzHDHZlqiaXupSXUWjol0jKAqKNGByd4Y6
rDAHvl7Xxix34VsSvtcfT1hAiXKs1pkceYB+CNC6b6W/getm88zMyr96YiFktXQc
Da6weNP1hvWQ8t2XuGkSa3zBtDcRL/ZR9Ff7Up7ANok/UHoIKznM6Soqij258DHz
M4x1VBsoIKxHRVSK6M5ebqioy3ejDNooM4CThfoxVHNUWoRpbVVK36YHaxBByj24
U6jt2HXKuFputN2HTgRwrj2L2v8swG7+wf9FzJ3EC96Z3CiBb0lBK0MVjJ7krv1A
8oYujyUi9LsWCAdiTQbDK7pEEf4aoTj13QGZ8oRd6VA6c15fBdWMcCmCV+O4WoQ3
WeJ/BZfrVAPtDMKt4ImuHxNP7wTbp+YFgfNSkpKvhEuvYRRkTyldx6heRqDguteZ
B9TBhCvn7pN9WyCRLY7YtusdDRaoxlOj9mCewcw28DqfNk+E42oGadMz2h56lTbq
nVFPENinwf15ke/otBKTzElwYaRtoE5GzyiM3Le8vF2FMhaVEYgiCNrkJHBjJ+Bu
nAGjLwLnKSzYkhevfoTgY6GMc83ND2IgGWgzMBzp18qydjEvIz8orRBI3XBuxZlY
hNTjRRhLv5gJUZ0MhiEQ+ep+Li69oHo55fmK75hvOlay3plpVURPV2L+drYEWBvQ
hjJXiYHUDw8Nm8vE+IOORwAZYr4fcYXLJQAiUCSQFTzraH4kUFX9megRdM8jnj20
9lcklgF8S5p/3MrvnwR4uh5UOBCKRWbKwwblVHuQ+ZSkUDdMpIqQEtFZwxYvH/13
saZxja6QXxioKK6ZPRTGl/tEZkMHfmYXgJTpFk0fCEG8KLaWryoxEJ/9IJB3OeGS
hwYKF2z3T1IGEZJKKUMol++SHRL6hnpsrIgvhemDpsz/wEmsNIte8UF1A3ns5Nqr
5hnLySRoW4lfxmp6i4RV+7fVeutbQ0E4YZvTX8BIHaNWRD6ii0gQgDMI9DnVhild
b5FK+Wq4k2gpU8r/lA4AVbRaIIyz3zgINNoismuDAgMhBIojFAanHAmxvCwK0uFJ
oi6AVdB2oNw3Wbu+srHC9SotZNtPQfo7Gc11r0iDrsPVS0nUtP4aKvSUMydc//pe
A/XptMnCKlUha3P+M//e0dtTwSTLpjWv8zMXFCb/fQDjCElvAl/JEeT+06slkwRD
m52MUghFN4MvhD213rc4eAFCdA1Ug6L2w5WJlJPvWv0Rcs0+DkWibQcfeKOToZWp
FLFyiEBCninJFAVaXlbWDWAxmh7InKBuwNv034KqKDmHOFlXJzB/1MYFcHQsjI5Y
HqCMvs3byHkPZCq2NNlUceHKS9w85292JVp4vKYur4O4u5VxXlMiQYc3dlhuAWwu
IlGWtYMCF5p94yOiufoT75742FzmFMsO8LPHfKeWc3eXUzT+ConuiE3JPO7zV4zZ
QFknpi+lNtV90NDXiKExgvWzdRFXXYacpyvknMT1tZE0x+eISWYNFKV4dKvs2A06
t9us4egoeD4mOFPqHJ7jhUqMsFZ/soX9Becmq2alSibmMMAtMCREwEqTn90xj5tO
4ri7YCUhpHRMqGWRdbDY8IRGP0xI9EEX78il6CC1zE95Wrhg/O/2iRsA426a36Vg
Q0DrkEO3QIsoN05l4HiK1JfSf+SEiQ4FrlhwCzKQGAGhI1wsN8G+XBqU2xzY1rIk
7xtq6YkTyj2LqWe2X/OwHMn0iwP8XWnwT2MwZ+PEBlj43EUOM4rRNaOzIkBQjETm
EyIwwXsDGlO0puacAoZ92MQrPjEJq9fCZB0JgAjH/5KyWVHExc6j4i7gWvfVFC/C
mKuoiuB5tITSeKAtJMwLGvMtEgUS0Ql05kgxf3VCG6D0YSF7jfjrDbagM9MvwOya
rJZJZZnZ0i92H8z0nO5c4FOAN4Sb3nKVt7IXtBNYIG+6iRQ2TI/IRYMu9Q/BpGgf
8sZX44njTYhRYAPwVrauAhUc9HudKzrn1J8c+YPy66tF16wcXm84OJBp5J6uKevR
dMquexGrGlMlvcXDs2GJZLm+ucG/aF6PPr6og5Y2lJMNydiw36tN1r2Ml8M8iAuH
Tz8TN/mGfsOcD2hM52UZqAGFwes0PG0rFk7nIO/noyoP3VUme6WPx02atY47DmDa
WzrwC5Jfu7bS8umx+xzLcuWJiHxvm+/0DqYilPivyUjsvw/+H7PufV2BEkbSulPX
Op93Diaetas0W1ioIj+1m97RfcRrsrnr+v2FGeN9xIo3D06QsQLxiOUq/HfC9r6W
iMM9Mp6T4Em/DW1VMuMxqSMx6IB17o9wMnr/TSceHUeUBqt6zXQfBCspNIo8Dn/1
Htt5gURyZ9vfvoaI5r7hIiGaF9nS83kTgUK7fehDJes/kmLb4He3+TzNiDpnOl1n
PKD7npGmRsXWVYmMLW2/EYIIKP7WAcH1YGtO2yo/wNbRc7JbpIai0diKZx0FE3IS
jvHC88QqVrmBk5O3WqOfzW3vIKbBAm2SBKPlCTaKgd5FDxDHs7CEshrsSeWAV86F
r5t4X2eywX/EyTZJ8Vu2SaPWxxaULVVpMjrZi3rFsH964Eavz+MI7c1BMW2enmAr
RMJqHLeVKXTZu13AS6SJvRbosS/sBN+hSwffrt6YYiM5WQrbJXO0N1fIpiT11x92
83yEHZgmWax7EYpvDdjDkgHaD6rlg67/OfIlGvZz77v7iJUbnQP0vZlSNpEEG7mp
gRKhqTSmSSFz5QYgMlsFdaG5+6NIwHaQJ/OX8+Q2q4FRixbHFC8ZqpkvpbAb0ir3
RH9XggSht4IXw602lJE+0qr6MX5Yjtss3RdVeJyTiMR1j7Hujpidclmkaw+qYntt
EdktoGavTwHHCu+g/ju9Wu5sozjgsiJnFst/8uiPXVHKIIMdcPeyJe91shGoaZaS
homejD1AGspIbWrY2Gv2qGxdhgsKMZUxrRFFMwk7HV47m73JmAl1033z3y2gIyl/
vf35myByp4C2N1W5b/4oSXcQc7MtUgsxgarxxxt0yo+ttR8xNimIidnLWTicfWUJ
dEdPDFTqCgsHeD8jTvzOCbGQaahUXxIKllVWq8i/jHv26iIr8Z5g3lxGcK8QBjLW
/nwDQ43yeqkMz7ac6WWsQCdazMxPZowfAQOOFE2OuWann5kV4+zdOdbjaBTSgKml
2Zsg0Qlqoas5hzH4/4TGNqMFqqwkLlzeaR9pAvi4layYOPYTj0AvrSzbu0NAwqq/
NhFbfJyjKoRO2k3B7+fBaKVnJpp6pm9hRJNDbjdQvR6BijikAutrK5bQuD1ETfuF
GVJOx05q/EIGsRp7M7C2cgym/HEwq/b06+2qvDhAArsAMvxlJFvoVb94MLESMoQl
4LMFjFli6f92i8JfTnzXgTcaEpainPYPKpAUsvQEAnJNKPX4YPxUUqHkaPCdmTvn
t9KOrSzbGiGjLkYcwv0u1hOvNj9J4u1Wzu8blE+1rlNaQXp5oDgabFmcPdAebJ4d
t0DTmOByGPRMVExgXNMknCT8AXUc/5D4mpaxjplfOo+fZS/txI4q2ASNzg4v8UL4
xUXahIVjY9WoQxPIRpzdkSGU4NS3PdU4kdJpn5tOwbGvoVuyNsc46/lft8S35+0t
GpzO1UH7c8EZDMtqEpqhltH3liHQw/nvBmVRbQHzsvvbn8MborQxuIuPH2dFY3mk
cxKiT9ZYKaBN6CRjpISeRCiSSm0IHj3uWqtrKzu6Oot7qzH+SBaEvl4++urf6LLE
2xvxa9N2knnEUk/IJGNBdko/VXM+XAOqV3qr6XlYSra3P3/d88w0PChdw580rMgl
8WCaXERlpn3FQjbL1e0/20HQhpKtiPn2gdAQfrCCL0+Vsj5Qsmaw36MgPdQXF0ie
g0ASIUYMYMB4bSa3CWb8BpvlLQYIGmcxUXOwJRcIm9e+ggPoTkKmsuW1NpiIgONm
IF70xOVqPCxWZIxx7FV2c2ZlF7EVRTMN8iZhzzV/NaZuoo6LomC5a2s4wdZHlEM3
tuQHtZvSNey3eyfOdUuoD8dHviFrU4xRGqq7AZXaO8fXgGqyAr1N1lJuw5Uk4j8M
vjyFYk/uKS1kwECJKTSWhEVcvt6wc+eDBQrFOGuUzxBIcZNErBLoAEcLLCwBd5XV
/5dgABxv2accoZfAYYsBRtE1j34lTA9g1v6kMaKG+jJTWRRl3LfGEbQDTd6PuxXN
+Uqkb6qLFxV9bfUINrNHFz5JI1LtTRaR5BEOFy/45oPU+oJwdt+DVwnS2gG+U4p0
bIcyd9laoh6i9tYQepLxJ3VOSCt9I0w78aEtVUwE6k3aGjBezcYr+Ez7lVE+Pv9R
GamtfqKYR+tVwJ1itpv3RCgkXpagI7JeT/tuXCwPj9ycrXJquzDtxs/luTTADpMA
K/n+tnKFXLxk62VOyw41UUpEYzY0O7cWvxvL/JrvL5QypZSc9JxInur/rBMc3YSe
Cwp2c1TaAJn2bzq/oVr+fSp+mDKpXJ1l3SgKVjtCgONbAbnGNqT1N+K+bT/2xNtf
7eK3nuBKV+NFFfXeMXD0OKlBLMfZYlv5gO853vgYGiF44NCYofS2+v320Wm0zkAW
Mg0kNngEcOeaEyB/bTStWu836bAz5GV+GSCtKUzAGthH34NwPvCKzIQlF2YIp9AW
Bg+mSChAhhYxsPuVilo+70FrvXiWYXEezZgiaybMTHLZK87Toh6WgUnPCF8whubW
nuntcqjfyKTTAXBzJZAiobcLkaQmkSBEvbN+B51KmzsnFyPoYrvqG435+Zdelfyw
zexnLwLhzINS85tPdiIAA9TaZbbKCR0rWR2LiQ4tsFzhaDLRZLo36BxrSCgYcAzW
pEiIrusex52q0KY5CfHBR96qhKuy9TmAQJXxmUqgAa5XnjN+EB9vRga9R+0i8fmS
imaiyFvjIGuqFgcxvyIzEogWNdb1sBSbVTaCK/9k5sogtgqP5l5mHCheYYm8CDUc
PfcBhdvscm5Y0JFujeiYdctHbAe3RML/bJl8/6Dypxbv7iul6qvMfHkOmjpswUj0
VS72apzj0Fcrh7SUHJ80s8N5ggSLkxOjtATBzi+0klzIPP96DCvEQHatve0GIAwo
muPAIwJU+5m5RV2sABuJFvBSoefMwSYnEE30Kk7DSLltemRLLOlUs3QNgsjnjsOe
jDUgvtlTBvwbVVg05HgM7mVShy9Xa3zZFTNaSgDvI4Mvpg6ZL0QheJCHKbLPt2DW
Zw50/zzELpThfyPJbDlguq1u3kYTRYiuwvcb1QXPf42yxKaRBboHlmBxzL0sW7Vn
udpftUPCHXwxj9Gejmty1RaehynWbdBESS897cweFK0Y+5e0/pPeYVnVtcpe9uFj
a0dGi+ZZ4KbxPTW8GI9HeWi7FpFAyV9WHjsOQVwa0KHXZFCjHArGDMu3Fhd/p4/C
vRXKZplZSSq/yrWXUW3Wmzs53vkJHe20g3NebOtm8j/CZmrY80quZvrUHIITjZNw
KthI4UaIKFZdmIYCxPWn26ceX8Q5o1nm4SaVd4xBJMQgC3RqCjdLarLw0l7vzWx8
+2OAFSqBSNXkTyLhkHCGjJB9NGlwzrXtvxum6MvXKfkFsTpLYCB54mL6BQzNW14A
j0AHF4yoyTW5ADXCztflMRpIQpZws+YdIKPyusX/z7LENF3RUYhzNRtF2mrUHZe+
a64GfQ189Y4+uqjYYMidb0H4nFKehCCCBoEsbiHSPTPHCZPBEizmaPd5uyeSVIjy
xruv+9GfjyEam0GpHCDZWBMkeVCjuIQ8mPbDm5XRjoZee3IuM/R4gabScEYUHQLu
AV16uw+hEXDT5fuSffrEVhBPgWJTiJAn9kLUTMmiTDtzawVoVku9w25ptjsk/RdD
uVQBG2kcptQOepBz9vLsAGf1K5/JCYMdRPlBM712fdWczzhVSUFkNn6vb9T+v7Ay
RftEA4vlEMwS+ZPi1b55zN6OtJDVuvwRnxq/N8vUz6Kby1u/fLm0VhvgsmSQDwPy
pA2+WcNcgMDyOAf4Ogafi46s+/QtpjeP2LB3zw9j5PDA2ALxHQl+pG96S3Wk9YXx
NvbVTGNdF0A4I2cl7WO1rIY6hxWWdv43QK/JzvjhyjMwS5chK19EcJFJeeqft8oM
qYkXo1rtv3EO5W9LKEL5LOG4aXyH3QFcCsfbt3kijdKJDPSUafsgjPODPuFtm7dA
KUpR/VF/p4xDvxiZMJIqiGj82SknU3zvDU8wwMsZORPC59ycXj68mzacI8GFXdoD
Fka/zK+96XmbaOLMdQ5iIlGrzeYtiTMdNpg1h/VyR7vF8JaW98YvDeCBjq9UWNfW
JZgPUPfmdyLNiK0Que2XWaQVx9CdXM+Rxu0rGjd+db6DTOlwyL8BgW+WFwr8pA2e
7E6e3FQlS9WmxsF1l2TPexxjWMoC516Gve6rM+eBXLEUCkVU5U6NWjpiIOQll6MO
4UfrXOCZvb7BnvInSFbeqHJ3lox6MXK+m8w1Xi+aSL5JTdggP3A+k3xO2RGE4a2x
XW/A1BPSm9aIXh3vNd9e1QS1bthaRcBjimb0CeomoxC/FzggADGT+9G3PLx6AcjO
xabJ9VMh7ckC1vJ3k/K7JuJGvxi5giZc4ini0rCVUTGsWF9IQY0d3lyhCiwdzBnH
YoKgCKQgrxRWNBfv4JPsP97VJ++sVfL4BBVl38OCJCRomi+DflHa//8AmQIlAERu
X/8P16E2241vkGu9JAEhjQpiIEtmtukZXM1bhy64TrgIg75rbTKesaTHdnf1EcBK
7fLHKzH3garSrwJpVsx9ri04PJQ7meYNN3cAao6qeSrx1eXV1mN+AnDw55BaJaVp
Gfz/RT3qNdPRbRLy+wagssCUyrGnXy/Re/qGabtM3D66i65CHjin1AVw/QpxrBUY
3juEZw9tMw+6No1tO79ivluEK2I2fjw1D94FvIUugjWfa+fSq1h96t8b05g5nwwa
3+sJdyJywqTCceg7sJOZV9l+LC961rMd2yVkPptsRvsK7cIjQkpksLvIBEXG9g9k
tc+sxJcmAc0xVD3moKA1314dEcAK2UYU0pJ27Tma+hJXgk81fkdqhhm/Le2JAtJi
vtc6+4Of/N4VNiQV/eS24WEUCOAK317HcxbdSzYFsJh+vR3VZxvPo7tGKEXE0Rq8
PwjZ1tgVn2tewQeu8uKibkWntOoZEz4jkTlY4cs9D026VXxW5g89D8D15sQfJ71B
roEN/+H7mSIMcaWM0RQ3FQrzz/agmolSLIXXw5kpfhYdPeucwXo2nSNltx5amGNi
8VwKQmuevR9WGwMsJpipswkcsrCAFcsnL8zMAA5IScvQTxduO2RKP6b+jmTWL1Uv
dcOmtuCALMY32XSnL1Pcsbm1NfPgKUoZTTaD9qH7OEOTd7AGjDON/mK5EuEujdFJ
e0FSba9IyLOqfkQBzaiN94q1WyvqhMQE93tmu/vu6OHBI89TqWnzt0MFkftr+ipI
4eRBtxsAl05C32OR3eMwTSCU9YlHupPyWxyren6pem2xVptBvmPu1xs+0OjkEtRw
SalRV2/l2URKjVDTDgIqFSY2AXVXvOJDY2wrCMCTezfOU+XNauowPXhXOYrKiscq
zTmexMFnjcik6m1oOQ7ykwdSdV7QI2is1OqvQYYjUoS0YIyHHcCRXyqA2BYM/+Ol
c+moHZwSvKzN4UeoSm1rBMT7M/BBHGIuVcmBFzhtMI9kA8bdV7cgizf1I2cJ2oRx
z1D7LRvWBNXi8Hks9X3QeEkYtXOh2HlInRxubyzKPyGssfuyCTkta50p5APk9GDW
jEIkDbFpYdhTWKCULKHN/4loRg0GtDWSGnOiw/6t4yoQXQ8h+xYJ54ZHg9XwvhLp
upbzfXwnx+a7Jnxd11Y4rXKrqX3lZybfgeuUzaQa6j3sl/5SmAo1XMaMWCQiOOsJ
R3rtL2Ok3asAHJwjyRDnEWA5/zv5Z+6VXfraIIQKdOQnj6/gJriSL7R8cpdpAySz
tjBf9YMtfJh18yVOCLhi1LajvbSGoSnA3p1MVHNRzOrCoKtklL+1ab7aO33qtbVq
fMhu6CBgmaP4TPo1xiKaA1b3XCgLB99069F2M8B/HDL1Y1GyqqBuk094h/Li7g5N
wJ2MQ7MRIe00mhd+muyKndmTD4mymO0hM1vMbMyjYzkudo0hyD5kTua5jmFCjNSX
6MijEqqagRWmkhCWhAsjlOjK4eDZWZcQb5+QYStBOL9cvPYrlda4F6DRtiEBZ9kK
a3pFKaFmu40L9tPQlnNIN2aPleuuJNN21/mrA7ztmjkPLiDWENz6Uze1mtNFw1yD
vnvZDSk1S/3BGOk+Blhb8ZBgPVwMTa6wS3d7+MZol9C7C+ysUXZaPv2l0gFkTvja
Novk3GnekB1ZE6Y1uf9rY+COhtbFRGj89IAzwWr8yqbfz6ZIyyjPqC8vLNDTmOHo
3DvIsQa1GY5jk7lsQ6Ru5Ra3Bdw6MGgFAJaY3XZKmT/mcP5iHcNv3nFT8N80+hen
fXGeaVpTkphbfApS1gNv0O4SroknaSdWstkd8z00RGWqIxgQGHEI0MceWJ5hi5DC
22q2XbCOgUkRpWnoFW3TG0l1ur9Iuqm4TAwYre01Q/m5fnSURAA7SCiQsEQGXcEj
NvAsyrFunkDnCakm9bea26yGHohvsViya6jMeER7vf5E1//DOs9lAww8hReE9EmE
K0NKOnReSUC2pLzgrGffh7ltBvUOvdzD5FxqHIK/6YDo9qsr9PHwzauwFEqs4g4L
s7YQFvOo/8e9RoVMgkv1CbTvHNZq8bhJhQZ71t+JWGEKf9z5YPCnxw3pg2WpHOPN
lleRv+F2wQfaNTfvzzZ0fmd4TuVXNqNp3NAq4NMSPHokV7HH7D9t1BHA8kHTR92f
RvjFQKl9OFm9h+2jEQXgN+2QKS16Lw9yC3CGzlQ34TSMfIvdh5iFHkA4HC/IK4AW
LveFEZANbtPloOYta6WQymvcHpwibWjqviuvxlVgIdaDiIa986ZAt8sGQbrKD/lV
tplZLa+Lu96c2s6OVZfj36Ehs/uAaVhHTP30uvlOBtCC9hSVQ1uxyYxalS3h4XAY
1yiUbry0uHhBtVerjM5nv/PHL3DY9M/6uCTC6cN2hDZv9R1NZo3wpHgXI7blJhMY
Xun6t7mEmLTq2RDvmlMCHxlLe54NEIc8U8y5qI5E+Q2EisnN4bHsbFtLQgaPJNSa
ltMokaMFb2v8moL6UaPTnpr/kRpgPnnEVZreQVTmoIkZjoHbkOKWlARN9j/yr7+H
W3h7AsmLc5RxUyOFQOi7sWDIuDerBIUW47bR1zqnQowjSCp+IFVJsm9OTDOGRUJZ
f0EnFTiVUWWquCVdkNfq0FQYcuYt1+B6m1k6IsenR7nnChATbf/Az7JTTOBKtq9F
yDi+pXxIcpKflcaRden2t0Jm3+HPaZzmVW5fOcWFzzurNdVoPC6MPXH1BvLiC604
fW1D+5r1/OIrOnnYuQ8SKsUKDmoNlNHR4xPVsM+vUja1vIpYNbExTKbPG88k6OBr
lpTw5wwaCe1Ev9rXKkdXrGR8N/XFp2GeVmWe67vuivoYbz8gX9AkDlW4QBZb/keN
btP7lrA1+WcV82CkiBYbq+2v8lGx+oHVT4QJfHTOLgg8kxgOCxzxe2iUJa95hy+2
xk41OdtZh/vPKug43eSCDmKOokdnMTj/PplXXPmb99BUDIYdatVg0CahMRk1gR5h
UdVC1gNL76zERMShOTMyB7hSAdY4h8/64/cIHqaTxkQtrqkSZT8EsKzCAMlSrUHK
2SHg2egrBVmpzSZdLH9aazFTsD4d4wLoLHMBH7vGArQ9OIGN/NdnRgkDwcdMFKMk
9RSMWPJtbNqtT1LhUFNUKubDqcm7DsK9FTb3nl/+LvSIfX8ewqBQ1U/YMx5DuItx
P99L1v13pL6DiSQjTfP5pg1JW3vzcrHhG3lM+MUqtmSxghaoQ/tzQnHQ5BFWDNWa
WBIv6U7R7A+zdkXhTx6/QvcqX9z4DVTfFq+sqFkkyvfm9DunWZ3AGdGgaBTRLsJe
OzKs2udN0hjIHFitUYxrGAW/TBZizvtMG8h6CI1SSd4WkZys6xUt7DIFJKvaCGJK
umvDNIeqO1BSRdMKcYQ19tpWkmgFNY94ffrKSEWECuu0zciU4ARS+j5aRwcJ9xiQ
Hg6oVYudDDMo+5UpImyMckBX4qGeqgrmlPdgmSPLxzOt8LRNqCDDwMON6vl0BCTY
f7DUvBUmaAA2w2mI1pW3IA9VTk9IP0LgQmef/cwUVTf6eHwfO3jxCh1+1eNZiu5F
Oh9MhG7P7pRfhRn0KiZk3WdVNwIqcTJVjQSdzEqvdKPamnu4uFV2RzujfU+KbtI5
ae+3Xp2psWWo33nOhQZ2DLwpqDH53+ReNrxOwV7rYgcCW4J3Zw2PeUv+ZvrTMbwv
P7rV9k3IWFmsCdUerzk2cjoQ/S07PS9kE2FmENto2IAAaYen34FUaVacxurRrGbE
f/XCdCaOSkdKXISXj8ivq+dXdV6LwteAZOlCcKytgaIY4FuqkGm1+FWwnVUjLmsf
KP+S8TSe0RYJ0NR6AVbSv1DeZGDSmgNq+w4zFLd2P8vHWOSTYVDTcEUaf98VNS+z
yRmLBJ++Q0bIy4iAxe0m3m2MW7gUWB82ZTFhpT+Q8OrizY34Y4IvqKV6DjsG/OH/
EqbvbfuZM3VW+ALvgaG9Sjf3/g/fN8oQpu3NKqGj9gX66vfEw4snavCOFpf04Zsb
oxG2e49/AZ5Dm5rM73QJD47NPTN6QVzuj32U7ZRoqyKeqEjziMp7v8lZitvVGJjt
ihRzH47DUlJ4SLR7PfolrYLsH5Jsf1x8bUq5a6ulLtTYNdZOxF18ksh0lWkcdwOS
mem0MqVZDFKdFo+Eq+X8nHd5Rkc3jV+m641YMBp6nq17ni8Weo/PUaAL88rXgtAd
h1s3XALSDMSoJjnuecYrmp4bgbGUqfgBGeZemYvlas3Ito3Zy4whxYs1jZE76oNg
6k/zHDdwIgPb/5+gLQftkHda6yKNGcLHTRdNCeMTOzmhAhfhLr6zediY+w7Uzk8L
adydJkqV7PWlvnReFI+GbUxA6imZwYVW8vBukUU43XUV/5ljbM1XEWGOO+tECwuP
ghpR1FYyjfKUp49RtvVUt92WRq3LKDfM5KYl9fT6fePP7jzS2dw+AK4xOIpUzbjD
S8Q6nrQdFn6hFosd79MlUNtnpdJntyLC8FZnS24In+v2wp3yjyYh3IFpAvojeNYE
sNNjgltgVCgR6ygBsHKXCkfOPXzv2/AeP/v9cxbIpapV1gR3BfZHUfJj2V6hXK/g
9T8W0hYT9SrS/L8wDvF0Bm2RKId8HuQFJ5NX8V6TExDfXPh+nH7CpIe1IwsjRQ01
SdCqUUGMGG5HEK6Gvptu5IkA+LQ9TmQyd18LEMtg6C8qr0pOUya+Es4mHchpQEoY
KNX4/2zUbk2l14Ormndmv8Ki0s0JjLodHFf0wqXUcKTyzSwNReHEk0l6bNQuLshv
TUitFIHvdZNs4Bg7sVHYEnakxyYfzD0q19x/e6eZZDXRiblfbdtL/OOEHW6hpD49
Qd/pfJhrB1/+TpFxcXM+Wo21zbuB2batYOLpElScWoXYV4nnnU2U3JqMHXpU9fqT
INmwqP/UB4ju/3jXhzsMfkiNEPpBIkPjNSACWPJD6AUzjskZdEYoLw7/yINNJDtV
Z+JIBN453S6g6l3mRzSThgGKkQ3FvpY8NeJSyZceklUuKVO0+Lq20XCiHsRGGYA1
V+Uc+ZFaDidsBJ93LPaA7REKb5/We2/wryZHxwQ41JW3cukLsEvSUT6YvT5/RSGL
sIZElwdqdnB762hLMyRDiLQz65AKzlRJssZtJuRUHyXreQaT49DuSe4L3oMZTZOY
y1cXR3YDqNyDpMppb/zuIInTa2sv37rqegS/gS2QhUIbBHrbtn9kNTPwk8Mq8by6
MwhO1FY+DxCfZ87QhLCkzGttCG7AjudWC1lFfD1nyTqHZxoK2BqZqSdgbhIxEAkh
6Am6DHDqqfpwzrNVzwgfMp67yJt3lFOQeLPlw6DWkUA7FOvhENC0n9RoO/D5ixJT
IEdZcXMxtTZ/ng3eGoJkIT7FfVL32CDl08eK9zqahT5MguQLyupBnSuHOwJjjRyt
OeOMJlqK7PqYjYke1ao49TppZFKQ5i5VdnUz4d8x5jQfwgC2riEtZbWTJvU5G4q/
bzVCrOJwaB1AT9YjKvHxs4GoDtKNUOdq4BCOwAkkKiiN9j7Id+DJLm+PRMQ/D9Zn
Gsqof6HTSZ+wHjNQyKaHtDKbjKgVHPFsVea2y5AasL8c0EQc/sxwhvztulGCFudp
dK004sF10i87IIODt5DSabdmkT8LXkhJvvc0vnO1FpnpRlB4OAXFXnc+KDthBv5k
IocfTOpB/dY2asVgug3wy1+snHSpyuvBpaMjiQhRmOaMvRDCVvXGiTdB+l5qjC3l
y03YuvI7QtRVYaR7lyITe0W102dr+4KgIDqBnrLr1UCYg53WKN6wTx2q78DwAGhG
baP+u3LVb4OtFdqU/ElIjmEB0JLQ/lbcGDD7dFMSptmL0TK81RDzCUSk6cF6/f1L
RCkLUqLNXLaxF17LHIdjOBwgtVwjIAC67srEOT97iIezgufZUg2No+bOGt1lYGrY
zbOv6CjIRLb17ubbWwLZtnwoCxB6EEOPKh7aRaKWa6IgzNSUELjJm2WiuN+MhNhD
C51QA2D5IsYs9ZdycTw9I/HWbOEUfiwE5had9+/mixt7YSfDcDa3gxoj98g9EYfv
SQp80AQ073pWVhlwa6d7n+yrHYQIy888La0oE4ai8vtxuLngSys4N9AT9eHxZJv/
GbE/UUplag5sR5mvkHM7GadZDoBVhHEOoQdfalc2eIQmeqasS6r2+h09XnKffsEW
cRaGoMlREhjYjQri1G+hscmHR4Jx08wrF84WylzoxEXdsLSccH64e8Xy2igH9Xc5
G0T6/3Ys8Fi8m1LsjZZGngX8XgS40VwbKO8hyTBpidvrgsG2XeBiVZiWWHIWgThq
Lt2GnRFhUjvNp0Jsa2vji15os1BvlJyWQ1gcH+ozCvJkpnv7xtPlLZJrbndmRMTu
2zRO+RbhqlecbjsKuQqF7tssxOix0ZHqWfbfC4ge5RXjaV+E90Wlt8QLRRd4m775
ZKsmi9Iw6AN3Z87O9ZWbUZZYuJXo+1BcJJ3GFJQcKg6YyPIJWg+BnIxJeEuxa6UZ
06xBxAqmVnLWcl4KeaiRbDNXDe9MXp8wW5rEkMKifBsa8+ucc/UDLjxlXWnK5U2v
oSevpGJvjs59ruyRHChqmG2IyzfGu/PuG19zep2O2lvQHsDc4T0WmpBVSRNa4sHN
YIe0O9ew+pqlKJClVDCJ2LPTlGHOSzYGZFSyKRf3YvnuqFIJ1TqFg4p3OxJ4wcoO
YsFsda3kr8iNs43MbrjEJ3Utp8zVcusozk7nRchsmUPH0d5ZJqhzuLvuTpLFa2Am
D8nQtVzRCOClczJzyryELQgMeSBE9h3m+kFdjVF7YpUF8m7zSV6dIbkfN2XQmkjU
UVLoqj1UKMii0uPeEg+KE70dEt4+tvYSXcwHjOVOBw8LZdlMRvMgfNxvX0MFE/tO
M82jfbyqEGRSdymgi/0Ds/OjG7fSnraWiN+QhX//t4om2lRscNPKeX1o7KO5k9f3
tHzUE1vFir86XRlzCEch8qZddzynyHENPum2f6mUHY+LyKIbYkEYTWGmTjaTY45p
xR9OzpeXSnwH3XK6jd03V8DLQW5qdEbDmuwe4EvsCBzQgZ4ZUtzZOZZep8KtnsIV
cG48XbRZLkKuSnGJX0Yin1BC+0xMSbBpTchzN8l8/uUGbgFWg/KUw8bRYSDurkio
2GYET8OJG/pZUuMJiz5A6SS8hMx5xgbgCj0ZfsfmI8gBs1rpMi+xn1sCOe1jXZfX
QIYNWJ6hYNBmhgoMCS+Pda+SycrYpNSL9YpjhGEi5ZRUsqabojH4SnR8siCk21Z4
tXJQCBgdnp3tdtgGWZ0urEIvcLhxhLsTNQOE0JBiMj7n3Px8pjlaQstZCiPbXKJY
Sq5SGKRzzpORRElWxBDHVpVIdUXbLbcl2dgOmwMClnzT2clIcjd7h/XVf1NrlsG3
gAz/VXqid8K2OcM5l8MjtTYb8+C6Cf8MajpY5hCv8pxAuOEZyyA4wLvEshVzLwhm
FASHkNN4z6L1DhFqg76iXlffxtHMpCyo33jpiUeRdjUhAIlChMliAHO+6nnuvMnA
4Mx5CZjMKgyAGGVmnaHakUcw1PRZS3QvedLWXi7i+r4STyos+/h4FZ7L0zG5o5nQ
/pJ3BJGAEZUdgfvLo/DOv0eb5xnqqqzvWw6jroy4URALwEn03wc57mvltq868k9s
DCozWpevQ94GnIS0zRBzefSu8DJFu0kED+wu0kW+v3LSTlcOtKBse4vz1cjLZIp3
ColaVEtMbNEp1+xXokaediFEH+PzQPfnICdvLgSkuO3dYa00hds+/IBwHgZseFjD
XcDzSknUsi+ehY0OZx/OBiPzUUwwRGH/0dpegCe7F5cN7daNH9HfnSakunGq8dHT
pJGcvEJA6cN5i6m8C6eftdorH7OH1pZDJNsz2XnCX9f7ixvt6Tfzlgg3k+/zZ22W
Il0c3kx8Uw0AVn/aMvufl2ySfOcMkO/cOQIq7pytVjA4BoW70X/ujyXBKNc+iBFe
s9NgF6Sw/+qeyE2LL/KqVWmBG6gAGqJeI8aQtWqr2WXn0ylx5dXkFt1M5evr27C1
6OdIIcBOavqXz3OI6Tj4O/mEJz3FrXLt6qyWtT/TRYEz5B6jtoO1y+xOgYzOHwnp
7PXX5SiCY4TY5c0Z/NEgNrTyILM16a7ixsFIZ7oz+SgzbmcEKLksVaMWVo62nXFx
PjBAd1t/W/9fw0ak4oionxFyVsc+EooHYjOR3wBuAOGw2gdMmWvdgQhVa0Fgz5HR
BS9WvrzR9S9ZJmnwPcd96cnqR2Wuq5fYDfNvNCfJh0LLCx3JOw0tk428zQBuzn4u
unseSsXV4qCh3UbIeklE4ZZ+VqJQr2JK+E5CU6xCVTgmzirVpuDdk7OZMDNA4M9w
mInnmeUEWikbZ7KKIbQV7Z+rgnw8MyFzbpFMdniCpZ85Vw9aepq1JAbkkGJ099PR
8RbRHa9HhlqAUPynTxg9lS7w1xuEAThW7HJkd1lBJN6Vq2bkj8Iehpls5sd4G0GR
NTg9960GEuQL2nj9I2NdzZfJONWXYuVN22jkHhPow4kQyuW692ppBZrisUi3LT60
SKUoMLaDvTr0bQc5N7oxY4ZVfyKImVB+nsHnlbzCAcygymbWlKwY5nXu/tybGslH
c66VE5hG5+hhE8qm7ehj1+eJ9csJq/oy60JbMcGW3TLp5EucTCY4QXHv+aeJ9RIm
Lxf7Bdek3KvA8PyainRnsgODFe9yD79f/ycvMb/IzVvLORf+230KQ2QxxZJN+L0V
U+lghxDWoja+5odh0qrqRq3g6s3tzaEArmtAEbMLH5M+CV7Y28p40AMSFPg20x1O
4Cc2ul3Ch7Yz4lUQxNz/Mhki3LLfgfyVaN/WuTE+YoaZqN7qSwqlyfJCKO9+GMIJ
ftUYuDO1KPwj+C2PSKLmAk/vvBWXA2vJjPfqt4t/EQSplDPBd4SQ75x66QVrXS9Z
ear26ZsUZyRa9L/dRFgOexDQ8Q53RYJStIItCQ6MxewVnvWT81Z/DzbEeYwESVAf
cliQXDevI4USNHwCGxZ7xr6b3MXxH6CTbnXzfGWQ/Nabqk4GMYOV+Pz2AfqcSyUP
DWdghxxVJnVV6xEpr+pkI8atwOsbiCPGenW4WqYiyiQcAgi1hoEqjmWcb1VIaGZg
qd4yLq5fEgffZQMU/31VhJWbN9AZk0go8707y//QotlEqxPwn2Ps6DrrfRfEHo2k
f+8n2FchrXlSr79lvMb8lj3HI6NoT+IfJ7fK4RNdwz/xbWqirgEj2PDdDpJvtKaY
aZ1SLyYTIGxi1/swUy/XhorSGclLcVOzG7l0VxvqFIBylb3bGUNGYGw/3kpolR0R
9qJ0QoIfLF0Bb/41S5M1Qtu4/pSG9IiI3AK9BIcxz1y37C9sDqJguNg3xFaYxQxr
UhsFYfe69MvRkSgvOoOaS6SN8sVb9zaNX5m6kN81PkMRwQeBQ/gDxvTh1rNz0fI6
xftSG4+O5ygCUtu/9/aJJinGDT0qRNWpsyJbeHxfdZRrjlUVm3nBRtjiblcE+XOK
Cqe5S4TbSJZCJIIVo/QU0+jogy0EuLOpCy5jOS+QDV8lZx6Fg9zD+MPee/JTLgYS
ERU9IZd9MOPfGq36xY8Q6feK4MJv1eKSXsGG+c1nOsQAGf4KXWXIBjHyLsXitCTI
BCvHFk9wBqLyKxtcnWGjUFPGB0EyVYrNnaa01ArrMVz/PKZqbenyFLVv5dlz3AIa
d9/OsYA5jk++Y23Ncdw9fMkAQp6Dpw36nfkMq6dfwYfHQJOx4bKxq+hSRUHvxvV6
tL1Ko1BrQmZJc30XzRE9WnPmbZ5XXg4PVcvepnwDbIq434CEZEXyhcYj7KxAg0c/
MDluTuiYLkUygadCahJYzoi0Jw1k8al4JhggxsUzuQf8lLrYhvK45qUd3oN2530t
TOb9ogJyPfvKJDM5MXSVQ3h5bWPbGc64C4T7Uh+w+mjmc4Zwfv+hSju2BYxizFhi
nYSTPX55m/UlHMfPFiJQO0CgHMcYgGIFkqfpwyjksABfUXMNPtx8DiziCebxlA8f
bECi7SANz4+bGxXGOOPh+m8UhdRR7cFc9UdsrNU3QPUBVa1Toof/eXwpiRZ0eI/a
lb2qm/sCH0BNjQRUk8fyS4UvyYTxp0uPBvNUXI86zNM1KbbvoFaNlb55gVm8bgUN
JtJ1PhsxSt91LuIs4CSG4i5G1JY4TmgpaTqA2J6nedZ7A7ag9W4wjNoqZLFDFgky
Sx/RV8Khd0vk0J+aiBVo11VYZkofQefWZESSYLNYGkP+Yj6TJLjcuKjTvgQAFjic
pFcElx/Hc2uX18vp6BHYnpi9EsYn5vvp3QQCASPfzNL9O1mQ3r+R0Vm37gPzar7w
5a3ogccVtoN8p1pz35/0qDGcC3jA5StfqA7mf+otZS5K6l+LYqxIrCHvFZ+2TS4+
f9RPkCT+/ku0zxNuyTbEMSObIAp6uRhO1sA6NxDmjLGL3ZGcGBvzSuqcuzpcLiAV
CPMVPaE2qjY/M99w6zTd3jI4fQLg9xYu2V6ECiVHcLJ7jHKLwX/xyHbULWDqYYe5
nMI2UwLFVFE2b7C13/UxZjpY7xle6TRpn3c7w2JxHERvkY+GvLMzJotq2pGQh4ZQ
QlXg0nh9IL5xjvFI11GSDZ3A26FzKsrKb59AtkYg7r45oHdagdBILO5q1PcgJD/r
wuqCTq+eWIQL1LfzlqY9z01FIBYcdJ/2cOZtw/kLgwcxDnj8smTbpgPvVoZXKbc4
Z7lXSoKVLux6m4iZbS5gw4tzb7VbmFdYC25ngLRSLxj87w7V4lo9lk/+ptz2QhJY
1648dmDDuu0Q9dEjCTbQA8bewQ41iTjtyoz52xERiL2j7uNUfi7NnBB/bwY/AdKU
9U51AgcQiUWgBxtA+7Lw0YEhRCwKdXrkWsgd/9e7qLvKpI0uUBrAWq1DjmirwRDp
fJ5z9cw5JLcyjKI2Bncfk/LA4G01bABYyC4pOclNhYKGR5Ab6gV44U4Ik0kAsfjv
RPABjqEcnVp5JzNq5J3/MXOhsinnJQ/jMS/HjOmHvTi2kkr5BRE55rB72VmDpI42
/NsPi2QmVB0t8pB5WZUg2lXgS8R9r/wgvuo46hcqdRp/bnfpEhTj0jReU2wVv1p5
KyQ2w+7dGJVyKxWLRFGGW5VJU9i11p86xtBwTM3kXZQjaT7Qb/2ZlnYDhTXYlHtQ
iuqjDBjaQ6xFl0XW7KpNhjnON0ZmtPwg7hhUXz06fMuG/X3bLGYJB5Q/tAVQBsyb
QpowZNwDUCNTRdPmolLegWRTxMSDLRewrG2gJwTYY0Gp4r1z2Yzeb53H2VHCBwT/
hijGFPG5udX5r1p8L98kcWJgXzQ+fRaPCiIkUGxGyhwwAvYwnayx5BKxYNhtnsiU
djUOXl3Ar3LACVjE9C6O50iekj11auAdpFwZU4mp/wdBPel4AnyiPprvMZeFbrke
+Ntb4rrtPvt/QRb+mm9SoHPkw4ccQ2A7oGUtCZYZaXnIMZeh6MR59Yo890fgDyjS
gN3KMDykx+EByr/YDBnMwXBPv/5qkuy6UGrVz7A+bdeNvn5CdfZXFlvTk73HlcxN
pK29PZhiu8+t27vlMdmob7r2sFia5uYxC4OdbmclE7uN2aqOJHHRn8zGhHEv8f+E
HAHtW0g5k68vKO/pHeZMdJSO/o5LAgxkFhsosqbTSiIoloheQX0NAsKf9xG+5gs/
aw+THvENGeJQMisBHw9nyFa5HapJI9gZPHAgDCa4T+9w5eqNCVNdGlz2DtjX4pyn
bC6KKcC7WZ2BWFOmZFl/gvXM1q+THg29/gJu8ZXVZnYUgUfWNAR/5gBjKHZUmZ17
lZSLf1L62g42Qo4iqzlw9dXQSC0PYz4/B394SwSDiR08O+0Dxpddv/Y+pCHOYKPO
1/7fUJzZVkwjmPxlJ8tLijHV0gGpO6EhzJVHBoN2lCf+aw0Wxx8jRD/2Cmz/7HL+
AEZ0FCOHbihECwdhOhGPI23yC9uvTHwiUkpoEnw0ipgnRfUMh7m/K/+idWebtLwK
vvGDVw6AdesB9TJCp2pG+W1EpOnT33mev/CpFCOmysML5V51Ox0RSzPVUZyL1Y/l
YluDPPV6ftA/CuKqgtA/YqeVQZK6rzBnJj+Ow+2o+ZnL7ArRN+vZf+2fTcS2dFLs
lP1ztF3fow6ejScMqkusPoHV1zKrN2oiodJivwluWIJLnNcQfnV9QRWn7Vj6rEpC
c9JqGmJm0esM83Al5dGkpZFeImCz8ooHpFwxq5X+bHVhXdXphstuSdza6hYHARU4
VK3+B5qX3vbVmuIqvVzn+sWgkMuKu22tdXNTvCko7BpUiAHJDICUugufi+IK9lOt
m5jy7DXz0xgyFfd7h6dcza6mqanBA5rT7c/10PeH1zC/jXmU1+myKSRA4Y8HtMsq
rrCLgWdRvgvN4yRn9z6v+TyFjSPodsiYYkGGGekGEwA4s1/B+DH0zRh+Dz4rLtSy
2mLdJIvlAypWUmVh4vi7Ityl+ItA8SJTHtLdYuThFtooKyFUfFzHCRZfggC2bXt+
j7yZWfNbxwTQ/bQbNUUKzsLFbl+5tbKlXPUQJ90QiC0P7q6ZfS4cmVQRaFomVlwd
SHAn3dley/LyZPwWeQtIngQgKMgBLpUwmg1b9w85LjpNd31t1Y8feFCQjypg/9Eg
S3Y6fjvb7R7DVRtM0XQvjcjlK9OJypQ0XPbka2BXBpaAOzjR/izaRVaiaGdEs+Sz
/WLCh5+ade+VHQp99kluDcalfs+VCMhtibvZujG+PEBuEyFlTzBJCq4qkWtRIsTP
f+BS/0fEsVeuVbESRagxL8ESuChliwkUrSPJFMrSDmbE/+Luyyos3LlBUPqrn1aA
zRJ64wqM/ClzFiMx4ap2tzPz1p3zyIioF5fk8FV9ROj1UX9bkbab3Nn5GZ6sBOxJ
22uDNd7VZ7tzFhbfZriqsEgSY8TemkV5r5QquEKzDcqQofD05r5wtEMJxomjp0FF
BlsdXuDK/JiGey5LZVn/vFOzTM8RZOYUoKMlSpg8sEJaesRr2+R04ZDGHIXphlwE
5gwIcf+1WtVYvi/YrfUM5cPc2wR/WRtOKidsejNIBPcxSEdbFSv5Tn7cRbpX2ZqW
AEu+4SBlGSUGi9XfpdYxS0Xif2YtZXNUyO6RA97WEOw1j4vTbyMX+coaGEkTsgxI
ErR41bmYh7G+Z+Lx+58UpORfLytE9DdiFIg+d5/3/eC8wic3gyfx9YYnH1CwGQ6v
TCugF1SQ/KSg2Q4xgOmeJwNApRyIFxjrmthIKSpgcqZnpsZ31g6kMTV4Q1kLYBpQ
eGS4mgw5pPZAlQ2TAAYtbd1mYY/sJlgmTkZY1ubUHO/TYpx3ui7l+r0sOND444wS
lt/gR8qv/a3rHtRzqqz0AeFPVYdcvtxE2tOFT6SsodU+t6BJGv/m8gQXf56nPPHD
+jwbjVBIxzuZelgfxvb7UKxabsl0PeZTH/BA4R5ZTObtmQgQ5mWG51oaNtATUhbH
8h5bV4HQPUIoj1SQzHDAQHaGusAJ8t6053vW6l88aAAfNSlJ8/6WZqXgPMr5x0kA
MOxTU31Ubc5cJGO+3ZG9RMafKThZi87VSAQYvZvFNzDQJGi5vzLBmo4VJnBzdsjl
ZbBpcHigmg5Ff8XmrIDgII+hmNy0MiBCjoudxZSjh6fx6QJW9BLBdGHKj2WcIj5g
pmfymu7f98Qd7+uld5Bdc4y0/kcDYcbu3X0hIg6ddsHQV9cX1bTNRtHjedt0czIs
j0M2UmPAZk1KhLwHzICNhPeHQD3uoCXV1jo346p8RJSNnhRkDlBb5cgeXHDL8aK/
cXErx09Tn+FKrnrfuSdYo7uf+hL7L7Kl45aUkUJnNbW6lK7sGRx77gyryNUU+dqs
WG1jVjCKHJ8wjqS7JuwVrtArFOolPWryiO/lWGSGkpSNP42LEOKJ5a0/RldkOm2U
kYaGYodTv1UpG1/rt/cl3EwWoOds45Q/beqHyQyw+bVc4ipY2dxmQgXJkeNF6qiY
3vO2iV9Ex0zxsupbXDmgu+GkdRxRXQpekt7heSv6GNKSXPx35viUmH/jxYP8Vr0G
G1b+Qcn6sIyOM37ZVQvlhaz135fD08MhrI0GhiMW8FQb9wKeS3HZcLX5D/NTgDwY
HX8dM9olA7kRESntwEdlCWxNgix5CvdB5X44FS6X6x1rsAow5l0PlVdQ8ZAz0qbV
kHP5RbvHuEgJaPh0c4hpXpkafPJCAQOKca07afxXQYhILySE0XKyhDIXoHMTA6sB
DjIVeUMXApM2VzTua7jMis2Y7EqUxcuMa20mRdehnN1RBSKqqg0KawPTD57cR9WO
aL9nCI9ESgHL9CKjrLNIxklWfTSXY3v2BG4b7dqgj3pE/u5tV28gjLrNQlOKA3Qd
odcNrGLBMZcu4G5Q2NMcZkNx7z0RVB3KjhsHEJ1YGrXDe9dcUihKksZWbsGoRQSp
iLG63BZr714EfTksyRRRVk4NHZexXG9q7cD3sFEfaE+SqWwuWGc4DytB5rYJ2vwS
rU4vqPEwMRJIov9YTo0zC9wH+mwnMTx0MRWXEePdpHKJf6JiZ5CUX0g3E/wmlbKz
WOAhqZVwVMbTyjO229Re1985IcR4621eRnLLztJC2Ht3LATiPe4378vV2j38zibQ
dooJv8eltt45jytdppolLCU6l7xgXmIYsMx0kbuHAjo6V4yL9d4C9L0hO9+VbQBJ
ZHMHqY5WEAoCF9fh97wCKcyzFArWICpPK93TogjPLl7rMt5wzQGYd+4gmcZuy6my
9GTG6QL0BqIb0YJNcp1p1UlABK8pSiZp63wGmATXEi6r4gClvzlKhSti7/CK7zsg
CFUsoOSjv9YSGiLWHcZwDLG1LMeo2uUxpQacUtueNMpKmQ/HrMkahwBijWT2N/0l
hfa0F0iLn5f7fpx9EziQ5M8ZJQ77JZftp9L9vwlHzlnEl8CtSIYw7lzvX3PEyjSg
DSFVUZi5E3wuTQ9asjM7/Q6Z8c5cDWmGo6/l9FFSVltAY1kC/mh0XWvL+Hjm6A2z
AfM9/b/mcAIF2ByGlc8pg6S10KJNwz0jWR5rZFkVJwRbIGsLJywqC2B8rURSU0CJ
MVo6lFtRwh/mYj/T+Xhh21kMKj/qo33w/QSBKMB9uCCs3CuSKdJSLspwKGCjWQHU
J2xGuOMIuHDjB2t6vA4IAkSA/U0Z8m32MTHH2dNMv4Igo6dS9RNddcQzNQVBJc06
b7QtxUQAB9DLxj3SA0DrUu2UheyrLgbjGChpy6nkLqgzS0BvuIKxxmkmVqMbEkKs
BqW9eRQlygC3JA8x+IZ7hiy5GaQW4KXzYDZTlXPcy4eG88piYg79m9kQbxvMNInc
Tg7jaK7Rsfiwz/m42U0RJSEUpAKnWD5UXdA3vHvddy+cdjzC0ZgTV1WKLnkdkO/0
FgMreBAXHnTv5m7izqlnUJy5OGxwlJ7JnHKHFVN7yJLR+VMnMwbEX73yynhzmUg3
Lc0ACQlrTQQu9Q14PqLnw+9yFbsGcdBqEJ+2QFSVmSI3kncJhGfGa1Zk9eggjqVR
ARNDvXAbTbIP/5pdudrUR1mTfatr/S7VXz0EIMX2u0C1zhID3HchoODvU0fC/cfK
hTkPeks8aSphJooTItkEXdepKsonnNP4yunISR3TAMPmYuETqXAPy1qn1H+qPt2z
Pj1hS1l6pxksheyvsImPKABcoyYzfHpBLEyAeQXHyYMPPNsauwRF+6NJdw89z8G1
Lx5gFVjjwXRFO65J2bPuKaLgX1lFboQ8vG+Yh6qewZHYX7NMJDuHE0ZnbJNUdO64
ieABDehAuzvrBPyTFkuuvzyx5khrd4XpfOGL8rhO724K5tmAQM6fFq+K9U6LumsK
d5xCCcmFVMVSbmngvIeAna1mhTXlwe0/YcEZWuaehJjsh+hBcnGvhjPhsk4EpunW
F41aQ+41QuddsTRyoMtl6KDMluytbxBUr8m+BIOY8D3M+OgfeJoXRJBYx5g7LhP4
Y43Yb4wyLjpZTVF5bj8IwMnr1ERB6EC0wijQOn99/WYQCKfTsEGSDEIHlYCmZrWn
3Tq8cckEY+Cn8TrAAqS01Ws/VvXVzcZ86AvnFULCr1s5GV7yWU2dYkd8FzjHKRcx
AaRkQj7a5W29xwh/uIYjEqa8ks9Sh1XY4cSPSa2pwE+ZeIwDh7hxA3Ozqj0W7YnN
Gx50x/aUy0wIWe3mSV8fYCKY63BXa2MZyBwR1HWJf2X2fB+EDI9MnVPTaTgR1ewX
wtDu37JYLr7lA4j8RdixF05Gos9GLbCyueDyBz6lMu9V3BR7BW6kYCo/22mR+k5e
7kndWs2LqXp6njJeQ+ZcKe6ge/W4Dl+1+AQP52m6opAD0GpZVMZtO8ePkctGwNhb
w1wO9AIj/dVhnPe7AntSJhwFquxYNRhZeuh7V9NQgLEcaaZ52Ixqf9/TylEldDjs
ierZwmpKv0RpR6KNdYjHWQrxwLD3wnzwyQSYWmqB+vn9m+Ug9nkOQb1yJKMoBFdD
0Ii9IB0qo1BQvt3TO11JknhtjEod3+tbFZQuxhFNgclWODiSBZ83+ghzDMYBgXM2
4PKAgdak5zEwKV7cNwWo4YjEXQwRZ0uisJtUE6iep/cIgIdswpX03gOW9NEpkp85
nZZzdZBlxYya6lp5fePBp7QR/6MROA6+UjtIDiLefWBjzf8yCwJz9Pkdc4iEi0MU
ckGCBGuK2OnAmpROsBozeRv7uTZyL5fMTXNs5s7TAUoduA6wto18mAVXPO7Z9ZcH
9CP/3yjaFfMVwuAxggtI1iqRGTQPbQ91jha6FHCvRGlk7ee5fvSM5sYXmdm6loai
SvlaUu/EVDcEbGWuxQi4bRCzP7LB9nesH1gaY7D3bvhHKMEoIQjqyexmyTwbFXSh
2m2Hc36qOgVFsp3iRP25NRrF7C1i3SVvwDLDqJYmSZJJpwjyGkPL9rYdcCZJBCJN
CMn7cGhOSrCudOra5sCCAaLerS+Z/ahHGN9ARJ6xe+DMuBC0r7i6FtXNq4rT9tGx
n3hGu6+za8R/7oa/uh13QiAkYHSc39x1dMGXmC9ogg9LklCKPbT8PjzHVWKeY2G8
HtV5d4PLz7C2gt3NcCpTyorqCSfLCe1ucs3oejWG7LLwagLFkh075tSbjz1WOE5Q
p8lkhFK6PymJDTvmzXf0IkbTFnYzwKmFH+MpzWNTmSje5/rQpwFD8aIauKoxc5ef
fQ0L6S7PAQIM1UgeNeguNIliGwWx7wRcAy86R1uU03q0O81GYwJ15R+PIjYm1Y4V
0+WzGdOiULd0uArNQCF/eROjpMnjiF2G1b3jIYdZ5pUMTfULsdNtTvxFpFGPjceA
22WZsJfqS4+7VcvVBOHY3mpOMkz5eNmsy16aRROIAv+lnc4IvD/b253FLMOlCCz0
egfe5dWafHlhKYS+ITRvYidJHYchvR/WTsNaV+PImnk14bmqyQiLrqNopaWp9Anx
RXzUXLDvtgAArafNUKe7z/kwWggRtS2+QZMEw3xdkgLlap2CTw3UKIZhV84I92EZ
rH/4sk6779RLxgaztmjp6HalEURn0KoleeUPUIgBJPsgN1oC/4KygMuU8U4lbQaF
imvs/EgoT7486d315fzDiUYor8M1XC5P/Rln0fr0j9MDIV98TLP8VFi2pPEf3Cfo
mhBOBuGQCsbk5MPzKhMAi16RkeJqAsKAUY3xfN8OpJ6yqYl4va8VeMFagVxtlX1b
JLhC/jdFIhkLxilpOuOSKnyTy3j78sUSJPUbvpd8p4Z61gaX++tSE8ndL2xgHViG
kxMm9R8WvmLieVSPCboRz9NmiXgTi9Aw2sSAM3Jp1Fkk1HSthhp2rapROlPpXvT2
ksRmjb0Lr1HJQDTTWoSBpS69FeZFtL7tERyLj/sqbcNwfG3KdWLsMv/KjyL6v5EZ
7ONfk+HcNFs5NCc0IBlBe2z578y7n0Qv//+WVlyxD5FRC11tboAcLHTe8accU3Tn
vMIMIqrtGKSsh68BMzkeJpi/EBkJFfbLBcXIxA2qr2XxkAJsWGcDB5rf9LKeROAo
X01QCioBIWEQVLoa7MK5Z02m5BDcRzlyb8YAK3IyYwNhxwdIx36r6CmEWaAcYre4
eXmcO2Yu3BhuAhlWr65lcw+jv6tR6DO5FBn/bUR0lGfy2t+TD/MYNvP0Fj9fd5Ej
DsCzE/6gXifQahkTXkQB4j1209ZQk7Mjb9F0mfxZdkhV9QQJJhHnrab3NCEhBwPx
LAYEpReaA5Q6mNdFRKpu4JxIIlAvj5GfucF40CcbbJhLgBOcSet/RK1Bx8okD/Sh
q4vu9MZZ+hem+csFZRqPS3q+8tFDRAaMMd4NF3s+jkhI3+nRd2ROcCjkkCpqx0tf
nPm9BcVYNuID+rDXx6k9Jy2xCxzgEaQXExpw6dRif2ypXIybW1wFuIgPBq0C4Tvr
llLvbBf6ca9uIVb1Y4y21cF9U4paXusvnpgwPWFuNsj4POddtM+dfBXS8gBsQ3MP
RXxBSDft5MiOC27oRm9T7G9eXx5LcPIuylZAUvbofJryhuJ+6bRVhzKPC31AjHMl
uNsFU8YUDYj6PBqTmf8qEJBt8D9GAm1hbJWtOjuMf+Nd2U91Z2IfSBjt/8I5/fCG
OguzCDslhApyS0ct1JE1GsOJ2r+4Xu6+wUWl2458eDUqzOSVc3bnX0Mlna+LwYTe
yhcrijpv4G+cFhsa6fDeoSmfTFJ1kIWm0O3nIVEOFZpSnGuUZKUITAbtcovXlNpm
I11OjH8PnyR2wA2IaXzCsq3gENx7JouHtuDV6+B8Ed91vLLmA0YA7fZrxhP4NSyx
hXq6fLvUWU03i3NSOv1+B+//bjzIc32GEpsIC3ugd4YCbEJWKwXKNdjewEKNWPfJ
6s6dLuUvKWUQnMYozoruBcf1DRbc9ICmClumtqOnrkaAsHnHA9exBqCrGtAPwQ+D
nHXeQoHbrpn72StAVIDc/juouB5FafyDJS8kL9shO5BmVkG4Yqpow94n3ZJl06vE
O3dSBaESqEfr9JEKLC8MaI85ADL7F5aQpbwE4dKCM3pSz2NRaFipRtoo0oLJv2+S
ujx3s8dXQGfsM3Fmhj5Rk8Q6lcCgmiqohqzYrA20cUJzesbcs7v/J0XMiqrbqqX1
t6G6g9V6xBo9SckyffS/+02HsQwhGeJHWNWx442IewhACDsc+H/9nbHEVOZO+mjp
PgDjU3Qveog5KTvKbJUyW1ormop9p9tEx1PnFDIkfWvJ2IUkrmQi/v++L/ucJw49
3mbUQRkw9x3faOnBgWFSbONr8Cbyn/iy+YJtxS7wq13OaOhq4GPCBGd+xmj8dErK
1XWit8vOsqcuWxppJDNxRKqmO8Ed6kG8E9ZqaHh9ZM/CCPKp7IfDJpRXsiMeAyyw
vAwTyDeUdTQeN9FdwAiWnqpog08bwYoxdrN7fp6O8FIMIc3AbPGdCwSqL96CoRtL
EcNWx16bweZU0BFahY4lEe/RtP8FZ49Pdb4FI0wc/6w8xGI+vll23sfGbqqDDvIq
E9dL4FkgftNelLl5iI7GpItGotwEwjVRs1MvRep0F1pk+udAkX5Pr+qt+MfRD9sz
KYJPc+PpMKq0xEtQ7+aec8iKHEf2msj1iy0NW7PRkhJJ8e704n0K+afqQ35aJXbr
M6lSBCVgXcGSaYNBNLIkJKqC1tU35uwMCsbktSuNv8IIFlcnVqFXBJb/xgOS8ktH
X8oSR36Aw/O8Df5jSlsn55VPL1govCwmzmzZAx/f+6r55/BdAVN9HbyJD/E4bMyB
NlD8RYiAfDgzjx37Hn3dNX3wW8ByeVTJvnuiUd1sMRW215dTc3uNUPh5FicZXn23
uUHLekpsFUM6mTl4Lx/UtM0qS3W/1kKNK6oXvzGb/zCjUkliDojIT20+gOgO7yL6
04NrM3Ln/0LVs3jwflxU716TC6jiCEnniRMAmlHkTb0Zo6Cdl64vU06bGPtqr6vj
8cqkz+sJqOOew073hEsz2x9B/We3bMt4f5ZbVqLsTboV7ZbfRyxE6a22nR9T6wkR
vIjbI+DU/p44W9QA6n2F7cBSZ+LzbXX/cIYXTsn6vN5hw6ldKLui4waSvQsdQ2Xp
mIThvN8MtIvo/gXTfkwLIjdV7S/8vGZyuCrZabCjhhA/tdAqcYN/VLanrld8cRAz
ARENsnEGdHXFjMCaEwH3sVwwuK6KJ0OBw4b84EjNxcS7z+uW96g97zCUAZZuZ36g
inPa1+Afrl0c9cnmRnL0NARSvsRiRei1sHi+ILNNVG45GkX3v4LeDppkQd6FQfVu
c+xuIqWO7JcSj1/c/r8UyhQYYC5cIjfmyGoMRQrcPPWgBudXy3lu+IXwzuT6dQPs
OoxBONfHhuXJxPjvMc/lxYFemIe+Uc5UB822bEVLnmSEQV7JGTdFWDybUfZd2Tqx
LvgRTw476efsyVI5wVNYv2mnPr2cx83ksSGUONK0O0dFkl9NT5+IQVuezAzjCSro
v+oFT+KlZorr2oEAVSxfotm2gjaHag5A/tUoWdC9hFoBiZJM6SmC7qrt8xMGuDm7
fDEH51Y1KFLtyyfMoSxswvybDHhDY9FrQvJNN1MIIOyCsXM+EUsXR/EYNXoDqOin
IEgfJgJ+9HoZL+eVds1UtzmFSmbIZ80vk1/XDhRlfMPjB8Spszdkk3sTiIgkCdA9
o3uZNYBiB0bLppYRgvPv1DSO3jMyDXKLJp1ywrpVCAVl6x0bqqzZXJG91vATsz2n
ck+C2UCrRQnGiTf/XZeRRV/yPbKYE8HLfK8ZoBTpU8e0XaisuAJWlBdejKac2AUw
v5moGtW/t8xHYEXcuNV++DQrtMVeUJKgqBawJt4yUe6zJHNjx5kfx8QB0cDtlGyP
1xDesHPEKkSVlw1cyguus3kY3i9IWdfkOIbrqIFROxOYbPyAD6c5Dct9Q2b5lJu/
OhHHS9VRUD2hwQDboaV+pXfHyyc+E2ui5SYaDpXqHq0o+YoPliUICZ5T3h88BqWJ
oziA/2XnKUSooe3MyT1Qif14oCO9bELputNEUWL6g0VhanYFOxR7hl1MheVDxOLI
UmoEcWzkamdFaRqQsh9bxo062dFK1qBCq4/HJmMq28PECcL2ajFU0Ec/PuOd67kH
IaescoFVlpGU44jlbjtE3K/vda82HN53sML6K7kQI7KcTigXOF2YtjucY3nL36rP
FK9Yxrqbl8tOPRNiBmye3feQzhUQ34luYisU/fZfACu3H8WifrwT9zfsx5hSPdY9
XSGQVX2ywhoaGkV9hMabKYOOm6QGAlDSMfQ+x5L+4OhLEcgKHEhXX3GEl5z5Slia
lmWheFxgTAKS3oSDVyFxpHTxzHxyzmBedEcYt6n4pKVDZpz0VRYsqtavdwJH5Q9Q
dQ8rQi3cQNCSHtwxTEzRvw/TTqhMPL6h6R+QDoYhKzpLkX7kyeqjSBEcnCPRZCio
P5rG3nX5Gvaw+kbWXTVGTbrJgM/3VRUxstvj4w+pTMmzxl3lFQUaFLTOoJwWv/eq
sf36/00l+QoYiBoAwXk0xjn+w8r/fnfBt4a/7TCQEMYlmCZgLyKlrZ/4Hfd+AxL2
n92/2t7sPgubSJMbk0TwfGyguzXi6ZAyaXI4eeElKCpkZdwYtP5CrUgR0MNQKnRQ
FuQS/vlOUj6FYY/7p8gDCOmfO99xYq+/MC74gB7KWq1GOd6cBvhCL9hyxLa0Jp4o
bQj1SCTeqAnjRIgUZSQ+c1Kw1si1OQpqG6UNohRZ4FBdxbXjvx1Vd6/UguRfG2Zs
Abi8Mc1oDb6IvjVKUB2z66WdX14ZeX8GuNl5fj5kUbWPhWxty4fAYcxlHUpgRIxg
F1h3nzt6x2QshJE29cRPhwX1AXlrmy4BCwAQtxGS9baauJ4COHMRTNfsIXmGq69E
KupjdopgBiCrI1bIxwczkSxOQ2WeYLTvcRB5bsutvLJnlJtY7ManYe9GXvpHYeSD
ZNUiuvfxBOPz3hUh0nEA4nP7Tdu9m6UPAWz3tB+u8wLAdedOdx952dtsVoVKUxwS
r1utRwsTA+/g3MdyjKumQokCVN9mqRcMy1jiQBQnvOwI4aN0QQBWPRWgZLGXPc8n
1ilC2ISZoL6GOeAVO5rib+EMTZ0SLR8bDp5C6TA/1wQ5/b9sVd6rNyzyofv6hbiw
62LqmPSAn7bw3SCvSkuRDrYIi3n2iabkp/Y8WWaY4D+V7xte6UYExiyqxpU8rIbW
6czDxHL3JnMUv7Za4QGs5vkFE8IxNWgadSzBFFfxrhN8wxk5buFGDAfs1EuDdWhk
XhGYzYC4rFq3T5rwsNxM4QLSEMBHw+DB7PoNeN39EhCE4yCFWaBAu8H7wQa5bgZG
tv4lZItDS25TsABcsnda9VoHHt0m/glPrmxzsquD3rIgRb5Bhx5el5SkMfzVfpUG
aWZ2DD7Pfev06dXNPAwCAZoRlxcKix93zJZtQxhVgigRCMrSoN7pXQhbYRr3FHvB
p9xkK7XJVkCxsgMHhFwMTf9m4hLKRVNT0K6pnDz1LEem1uPmKr5lmxAD3i+X2GIB
g4eVqmmYlww3xFqNyaFfQHqF1sQwIr4VGC5vykmgUp+q1MzfkSLuaSV7ZOV19pCG
lcNLhJTIkADVEws/zvJKHAN5/BuVf8AwNF05VFQ4i2CHLoEbKElu8StVHA5eLdJS
qA/QwRQk7zQD3kuLXLNnkXBQ6+it3p0vVS8dUokcMS9nrJoExJMEiDxm7lwVJyS3
TXjtWOqRSjpZbbIH/vfCvSHB8C8/19AuBcCABbBPQbL9bbc/rBBTba9DZRpujhDD
gLiNHrgjvsrG8b2JL72cH+w2jUC4At5DwgJogqHHKg6n77pm/Y31/nmDVDo8x01+
Ec/i/ZUsiJnukjCKR17fVDUWEJb42elfClqE0wV9/SPI8WlFLnMVh/vVuDabMN2d
+C5hWI8QsRJh3VjxDQ/xbepdfPNYETtAmBaPwr6c6dUMAgq7hdZz4hHevpx+Mhjv
a2sMe4Y+Uc6Z2a2aAiaosTmDxyDMonmxw+b/IDNKHeSJOPqDPXuMB05fCLW0i0WV
HFQEKAbqBgmzLt7TZEL3s53lJKEunZEINKsmKxjnXh3b/brxKIft6suzpAEtda+b
L3+hLYJATBS1VTkdiM/+3a5o6iNns+pGVpoKg6pMxoFAg1rtpy7rpfITa+2icm+8
AtGxg5AmeOSDx5J4GBy24AyaLxHy+hjLRpYqB73YZakDsbrzLt4kjDIWIfNph4/e
CVnY7NYZP0FaAdFY/UFyPMUSE646QjnEVv0rB19bBquTG0SauC7PvqQQ7lpBnwLu
CEPu/LjTqwV/+kGr0xH5lIkrE8Gu5LCR6lZ8icLTk+S5EI16PGdE6xax57M48goc
GorixcL7LFt9iMH1ASBlae1yJAE50qpbhA+Qm9QS+dSgQeMTayn4DJ2V+HRMikoK
lpTRpyvxrGkp6vUvIc9Y8/xjkbpumsS5vqwQIRUcv4k+BZxhOj/UMioelX/aO1PG
yRHADXgdzDrKzVV+pI3p7HCAZDMKOMSwlW2+V5p2jcCLgwoV2yCvtfjHvluEM902
I7d5ba3Ve7FCr2HTbZBYdiUINp9jRzZ2xRpllWQ5G9hFZWXGlQ8pe81u4IpovpbW
lLwchvvOsZMW5kQY1SS/KYFT19+76WiPQmKoz8CeRDtbNwAXuQP9qVXolp5WmB4b
cX1HoWAVbbcolijV3RvScMqbHcHjjE+Wxjv/wqctRd2ROSKDfVBt2cqcmoj4fEmK
I4QTgTYr4KhUyOWm1Z7XrLA2xtyX/y1q7vtsRgYgQdagzSQgeUcAfIYx+/QLMsUo
sIAkkDZSuSTVwJGpOA+2V8hWcQMwawhqsB/Rd5mf2FG9dBXUkRyKOxH5e39zG1py
4eYQ5A8mxtY8O+g05LWJPdtfW9o8Ci8db+Rpd+enfmjQaocDK9wls9Zf83Zkj0yT
TTY0FtKPqCqNskjA73XNZb8+qHl0jcnKGt0675tXZdBIQcMx6GVuq6k2AaEilYzE
XFnsr99+HoW2br5eQXTsggCQ2BYtDF0Ffl4xtkeQxXqf4WAO9/9Etefiac3fX2EF
rwN9Mbdnpgt6NuQ9CEyi+fqNTVPrEl2Cu2pdPZ0Qlhx6S1qDS+DCx+NJ7LyLd0Gt
Wa5XHK6nHS1slXdYBB4VX9+ajxAnMcNtYpr0V+3ABypBg+y+YhM4CyzduKGPu7XF
0bFvKux7+ddJBRwTE7K53pNe2Aq6/UF77K4StlfulL7KNidNfk7avnl+n+quxKDN
H5kgGM1nNtCrAjO6tbeyj4NMQeA41qS/eYYurdARVFOGnvkCNTgQHzngyF/ukWyL
en+042rTGMDiwWto8opWpl+UVyPifBd2NJXitfe0km5kj7ViSWKHY2MtZn1vAyoV
2/rNG00zMUsMZ0Mu2+OBJ7SOGk1qrxkHUgNrKbWmJTVLAQ5f2nbGvsGtSClVY1cs
dM5zSBlcUkZWI/z3btPBEw+aDfg+gMcmk0MdfWIHPirugAUmJosLZDfpwJ82j37v
7BZbikl/Qr6IFMpvV9osy1hRoXGPDAOUVpl52GiyXzo9a7lvLPoNnBeD6KndbEJw
EBxaGpv0kI26C0SLc5qzhOP08KTeoW+XB0TyIfdFhEEY7f2ZzM27TFRmqSnT5yLU
fy9j9m2yzXRLtXWou7F9qKXo0xKMnwIgixiwIsfvEACQmhSHVzbRCKFWmOPuCHRB
06o2ND7v8kkA/5oh7ecMNqxTNTx+sqkXK6EJY6ADA31veL5k0agmHl4fDDUBSPVM
Ul+hwVsw934w754kyH5sdyxtGaY8Sud7w/GmHDOlkZKeNeoDGh3yPIuVnjevJxNn
ULigXF4gOIA9hLt7cm1IbgbUvQSEZx0u3blW24+9GJcrgoelTJ3pf4DW3VWdLIIm
WBbmxRR/8TPCdYdu0BmulDCjPjFleGZmmsQ2MgZriwujVVGvtxVoiQy2MwgdDp9p
0sCCyvKEtkG6QVyeNtzLkAE7PRVQphMPhC5wnJBfTBl4lDy9dTa4vj8VHT6cvGsE
8eRkHeOX/dXoEb+qNjnYBpiMqDshfL1CjtW113InWTi+Z+iyh101e5pBl1JgktNN
hXAVhMRRJP+2o6ngxra8jpbS5x8TTp1I+69bOS7jaLPqJO+eQf//0qFvzt9TsTxe
6g7CQWxw3Ty/+3HQna9OQF3oCD1GjsK4BdV3yYilewZcyyjAY6RuBiMveBespdTS
uJnFwXaJ8cBkmyNbXDE0VGJlz5sPu2q9e+f31ziFMZ3lwo4D2cNyplAF4iS0B3G5
cYrc/LIugoquePNf9iwx8z4Gw/vvAooA56xzP9qh4Rvvph6s1xGATlGMNXcsRTCG
6MLk0ICSKbuFdFsQDsqJgkNOsvV3MROwSd35q737BK//HGrZ9wThIiFtGcd61igE
s0VdAZ2Pi23A99GCmTeORHn28rLOC0uRYVznTzI2moxH16k652CP4KYH6x/aQcP2
ZvSIV40EbIKCdJFCNMbUDBomg8ZQ/xroGLtNo0ML8JeJcZTfYPkqynb9m3gFKqoB
+0REG/dePnQrR0XUf+IIaOfeFt5tNIVhwSudHqeAamPha/S6ntBlCjrdpQpd3AN7
nPPG85NkqGD75kna9MSLy7dHURRitjoB4fYyJpmXib8kFU/iP3p3b0zqVxZSHn1d
WwXPhxrrqDWQC4ADvAFE0PBqb4RlVAPz92wQcZom3R2Wb1qy3h+QchWsIp9SKi2l
DFOEgp+7PbdZ7Bi5An8Fee0nUf0Zk6/6oNj9DHJRbR0TQwNY8ltf+YNnzib2Ymfw
Jg4JqkoLV/eGjLliKkiEadJNVp57gqnQOkTtLau/Am+MG3v2C0mb0KP3fIjJruew
/76dFVSOdGkuE8Tfi9QAymOTT38EMNmqxxe+6Mc0oxKasbZemiAuiraJyS3pUk3U
iPoPa2MdTsjx3KrB4NkJfi1EzdvObVmhGZOiFhfd4BorKMyDgi5rQDVIDlkBAXlD
eSZ8vxF/Cp782d9Gey2MOgf7qENgV7aTojsG9OBpLVnsjVrso5tG+HZqZvrI2lLk
N0qzp1Jfw6iE6uGM370iY3zSHsI/84joJuyTxFxaNCY0khNQI/ndI/dfoZM3mzOV
0G9AAZAXnJt/h1PF1j7IzVq1PuGBClkgByZYKcZrGConC7LbaELNf78paAOrCXlx
csaCOGBWGkwuzQfHUARN281p+Rnx/VEXIQFCm1fS76KrBxApNDI4TfUgwTNgGOPO
Exfum1KPZFjssCskGUWUQA2m6y658V3Oc2xG/2QcUm/u11hHEbdeMUnnuaT8gahg
L6timdmYqzT7P+FEnWXm4Dl/+Zse+MTpmPRvnt+vNmf5HFcM0ETULq/wUC4XQ9GN
/YcOubLt00nl5wWTPGH10B1Z0OKBGqlONNBe9Gb19J6kJbjAT/VNPZRaX+nlwAxq
caXvv/71eRoi0WccHkYaqn07FQm4t2qPvt8XwlZTKWt94SYXNG4oALU4BK6rxNdk
4IHr72AmHURxcidylcYfd10hLDQKUGi35+yX/P+ZxsMYHduJLLlphnSUOInbnaGd
XH0hD4wAVe3vMWm5LtsyUyI2yVzNrjIzb99XO0m8dxeJKDO0lDZbXcwhZwK06r7B
YiVqvcfW2Ot6UYeftZmiS64fY1VZFkSk6/emrCoOszOD/QZajaz9SmUMgJr5vgE/
2S9LXR7O5Q/teApksd0SVvo0drM635lgj12pNgIa+kZMSbO914hOrfLOVLm/J2Oe
vWB8YUeX27mLzwDeG54h07eCYJDUGxmfk4BufAUU7L5CD6M9V0wWHx77/OujtfvD
oXtLi1COSWmUgmtpdzYM87qGaQl/H/4XDXDW89mz9Nnuf49/flLUBncj9jXsytEE
8/lVsdUqmK3V1c2DEfPgraNCH/Hnt3mOuPONoOwbMtbMWtU8ZQFPX+iNojjgyFSZ
miymM3cSgn0/gaV3iyrBYy7buuNyBkHsJiO0x/fNpgVnVp1Hnrm4X1O7XEZfxJDB
73YI7Kfs0gT+jqNA7r0E6gAXHgZbhm+Cl1+7cySdTggVRyXuNoJ1q9NFZtaLjoic
BXceurCT1lEi61EWE7bS80noC0wu9+BXULBsQaXgp0bLvnPpsyGYmFbKWnFGwyKU
dHi0QUqrtEndHeDlMtZvHHD+0iRBCZOl6DO3TDhiYDuV6o33g99fDGtx94Xj2Gvk
uPciSukrGd+wND80zeNnP9ytHUipz4qHzhW8MRUOsZ2tPIjFBBb1sWvVOAZpjacw
XVfVjxACVXVdTp75cKWWlAWPSQzbN1fTF4xPbLB9gNlxnYI9QopkNyQbw0LW/S70
Rf7CTy7Pa4DYxQl7/HIHwlKjHTyawVgOG3KFgt1ugAQAlBbIGKpL3OBZ6Ixd2Ezf
G2+wmAKYQ1lAfBrzlBQuN5IXzRiXRxwj4JPmN4XZnnfoVgLDKVpC78oH8uGoDcZS
WNFJ8T4cRVnjBqyDpJVINeTNxdtgfVuuw3PK6r/gwj9QP1Dg7O5onfQDfcOYtgJS
FstHPIdWgjznSGDCuHPWH/DTMsHgEnR+9xQBj9GWTix71snOeNSgv1slMSy4wkRk
V+jOprvln88HCSUkQZ8ApuExAkLa/ptA+jse/OqkRwT99tmfbI9HHVFlpJAWQIUB
eCBLgdNEIyuNil5r6r8/xtrNGiPZSojgzPny1m8TBco185HYODIRSnop+AEEPpmK
8SRbBexSLRPezLXNPlHBnrfcWWfkOrz2PPHM8/EWiaGCSbCfezvWnC2MpNU7NLRI
U37mST+5hNF1sSN/4pQxIqh51jmzQk+WcJP7YxRf8RvWc7vM69VNfzbc64NdiOO9
zv84digDqxH6JSLsig7kNAoyGQCpULeJJQqJNxUl1YqhUZn1fzMLwHOWAlN7NazJ
e/JPMxTbWSEpqdXAAuK7xoZnvk1qwaYJHGxwtQRxU7ph7bX8ogVaSFyz/BJeRQ4m
jLR1vkUHXyIAygu6LQazXmfkBYNjjYKuhxXeNmzRa32y6cHO7UAF1SKNOtAmaSgf
+YKxsnT3aqzAPPl+ZjS+3m8TPZ27fwGAEr/b3pfg2eZ6HfBRK9JeIb++/DvdDUYu
6WJ2NFWwlDnVacJ/Dk4NMpRTTyMeuvHJ0nKfQBDAouf4w3NVUnXd/s+t57a1Da1m
yb2tRSZ7t2L0WbY4Ffdvb644v71/wWqSkfbXJewjdqVHmE8qEuCChtl5WeFsScAv
6DiZizF/OhM04MlOm7y60MBkTr4kQQXHdmrN6jzzfNbw3OnTODZlxicU0sRtNLSC
r71sZ4lyu0oVANR1g+Tu8wIUEaTXhpCnz+updj3WCOFVbYOinyiXVdfudWUlpmL1
UqUcABO6FD0Y+2ZWMfhvMG9lnczefmUgSlS3lfQ4BvNc1f809G3FtsZYzDDE8bSz
NK04Uw7FujBRpvWV827kRFPnwGJR5FbC2kKdQaigd0w2K8+HtfKrVNjYzpZiKNeQ
y2IApvVSzw+sr6xClCdZziwRETxIZ6fScH+QRpHK3H/I9Y+MRx3Wf9kGqGXHNcZa
j8dM+g7pgXaWWYsPvb1DMkTbiFg4swxn7Mp0ZCkLdPtfY27/Aw4atlSZy2h7tin6
8XE69ESuSDBV9vyt1CZ6/bFuH76NE5AcVmKTsRTBAB1c+HFeb4PoNnds+DRCLBXs
uuK7C8tBvFM7Hraj7o4d6+yXWvwlgpsi8ljAHIJt2ju3OX5mEZCk/8xfhJ37ykWx
cyRTm9hDAlkbkSETrAX44bln4npFPMHXRIgxBbBkNVE9imRaeK+R0TEmNSd/4vpT
yAj5/zEuKPJg1uSDvr6dUX3noojNlwBFtU8hUmBh//mRJz6KTql3dTpueBa3Kwps
FJYpcqsmjvYM5GghFjoXJUCferXDoZgb5TlP+POtBqfppDTa6eg9w+5IF/Oj4iO3
ZrtMPmOOtT0cVIEr2FxFZoUMDVvQJ+3FuzpS7lLifHDuOKj3dSWAUwzUNDwYGpHW
QkRWrkfFceE7gtOLZkv9JSOMrzqbD+VScyc31ODJC90NlYyqtQykugjO6JT5PiJ8
DNoqroi5ppG7aNQGSTNRDMGY2wV1qgWjijOEKwODvMVLTSZDyTpPqKcj8Q6dJfKp
tPkZVW5ddOkitKZPkryz+OEmpFA9CYamKNUITMWfRrHKBbE1crE9sXbXABaZeTTp
HMW5CPAeSyhYfQkKhLr5nCM5Fu38PjPNDAP2rWyUh8DGIpWmQ8IcbQv4XrSpTs2c
VIeeZr+OhLNJID2j7EO2fqXaTGRhvaBlUrzEMGTWeV+u5YoWCehv2nT3NA5Dp7jd
ImaKRdOdESuXkuv+R1qzfLi8xDJOY/mFbaNYbWCfk5ahyRk7mktROrD5f8f9bT4z
zoMS+QI5aXZmkR/RL8N7UJ+tsCPjIlU3Rh8urXt9W57CvcFlKTtPkELNKNCEbJeb
ehZRJiYofcqiHVvG72UBJIm06ClfS7fRu9vUWu7vrzvPktgZ+20W+uF1Z5Q4lozs
6fwWQvmqzP41tRNB0F6BdmkoNypJSpheQe3HyIyA4IM5fgiQNTxK2BGKQdmH7m58
TbxOiTaa3lrvo17rS6ZR4lGFf4v/TFpHRKrlx/FdnOD1iN0pP40LEaiIf9aXb4CT
Vx5/SHMX7sx0RA4wMGh8x9LQiuu4NjqJfJoJbsGCZslE91M6+6tqBlMYWb6Acpkx
djq7jK5KSNnh62xJwBBEnaxB6MZRz+yw/dkS7VUUlwealLWnfwmnjZPGy2N2qDRB
OqfjUqF/SY0zbJzfTHAoWBsZV9s8zrhTXjN6RM6zN5yHu7sMieV/RKU19U0+4vTj
9GJXO/GjsC2MNBmdDcEEshCpDqFcuHsdfngOJkQgasN3r3TCmr9Vz8bYzzVhvJLP
Hr4qYUfO31OaCrePpMPOzAZ7Vje7/CtXf5A20n9SOztAMlk9y8Y/61rIXbTlHjgO
DYjbGVDSrYUS4l8dpd0TLIh2AxsF+p3bNN/nCRgzPy27del5zBtYI851AiZfyGkP
+zRdyzwcZNvaiLwRyYwcPsJyH8Vd7ujKIxdkUbU4fzw7wK8gKY7tK4JJ2vaFTNaw
blA5/BeI8wxflj/8oNUS1JsESReS2NzHdf/4vYrOLYoLqK7PI32Nqmf3x9Rg69Ak
dzPG8aQ+be0tCKuMHVEFBHkfN1BfDO/aN+24RSDamDuMEibHo2g3SDbI7VsbjByV
naoD3GVb1gYz4yok8cLfPb2AmlYhgiUxW5oegXTOT/cBMCC5vf86ue35RXArB5hr
ilbOFP73ps2o4kxtLa6qzrAPSbrdm86OBvmc4qqdKemXK71U1zj1xL6y0Jj6bE1i
17rwzbgnMQrc6+YTFrZ+df15XnBv93bIVjqCVnLJUpgco2Q6TyK28z2bFFizpob3
39cYZq+5i7f7abeCPUBFBKzKBMfVzuJ4oYkaY7efPebqXlHgZ7SzvanbjnE798gW
EIM4dkmhVyQ5mkZwqsB3h7n9k7vLMv9UyUedN5pbyXSLgpZIEEYHSLilFlBYIUm2
Haa6kjDBNEmv6MX4VRizPzwOSPMmctmnglFAHfVdBFG0yt2HgSd7NxtEm095OXBV
nfAQRf9+TlT6imaHsAfF5UvDvAcl3M5AejiNF+lMpPhkyVIe1nn5dgQpMvJCD3fx
DsK+AijmvMS0PgALl03CClBjN+Nz4voiCLonVON4CNE7AEwRVVFaAKIcDUBTqFHd
kWvnWvScVy4WTTMRSS0wWlNZiIdva+lMU/hl3tO+r3If1RpcVTC1d9cZbUUXSDt6
V0opw6uNdNEB198WAuRyttiwuZWEmnW9lhFE7FMXDlVd2dRDjW7b8GNsH2wb4H24
dBDQ7orfTAksD1ZF8qCPZystfH5IPHvbBX9XBOLqOYraVmCP7lbjPjgVbPc/+4Pn
eGHLKnEax0cJykbHaGOEX80jpgaY58tXnmsIRnpUkmoQ+Tj+so9FAxsbf3yC18qG
sc6NL7kCIbS7lovRBZSswMPJTVPQFuvlnSgjCbdyP6X6s33RqN2OLd/hp7rGP2Tc
zovPvxrXGRvR+f3iyq8oSPV4qWd2irAqfVYxjxR9AmZmJcxRnKedA1f5OfkZlf6k
mSqj6vr79hTa/U+HbMeoAj1PkpczkKDECx9VmiWn7FD8QZh4NyaOm4sirFPzzdvd
tc4og/h5cXYEIOy9czeSvX+OXZ26oNG2w2M/N/ya5gYy55twbG8Du/vfFXgrLoSv
8kWq3mmI7B77Ims5Bf+vCHbydYp9rN9jPOhY8Kt/uP1bixucM8xaJMMVGWdPpRwm
ARwbX55dNq5B72a9QVcoUtMKB9Q7lqCGalVoUWRIGAl/406ys+O37BNwQHKsfxrX
Rxr911X2fBZNuNcxPblr+1erIK3mDaJ5ClxB6WaFbbOdrg121l+DsDJ5GCTAaFIv
E7m247vnXtMrDvfKUQZI2forPYettBZ4CLlz7LFslBBbWijWur/7e+6jR6lPW5BP
DmtR6OYBcFmeXFJtCtS81wNCnKJWzZ4o7lIsWwHrfQQe5iulAulAD1FCRjmL54Jo
18DMTXaT3f/rco7CSk7OL/a4eG2EE/irrym/5xJESKGSPWa1UFrPINh1ve990Nys
UhkvNUtC1hEcwWe/zs0AKHY8wPnhXH9Tft3zwdMgBr+YdayxVBzNnQhCzVEIJwl3
aQB2ISrEh1gNX+7KDkPGxUMh81516juy5+l3fHVnLFyTiMMZZqWZskxyzwbdN9GG
0hJgSG8zCTNk9EEkrAut/GLvYrn7wuSlXMFNFdY0iuW3dyS4JAfMf6sB2h9xJFnR
ny1CLrfB9080XeTjn2VlG4ylbxD1LYggKwNjlLMxfN/iuJVeRfzbnLuvaBN88vCV
Km2sevL1Dh5sUDR5T3KAYnQMa6CKKjU0Xdxe8vBytZU170pxxsrvRz3MGGhcp7xh
H+bUInYvY/XSXGQZWHBSkJz6IDAbU55yMJxxEecoGssUskbeSFYi66lZH7FfoaNH
f7hl6geXVjL3p3ayyZHXIx3B18t2Ly+BdKsOgKa3HNr6wWucWEHY297dLnG203b9
o+7Dm3mDzwtoBkYyR9Ss/rF9Zw79L0fwfxaDCzYa0nlQ9HsZoWd8MZvl3BMe3gWs
SsyMRuuC4fHTJ1FJPY+9bMxJb68jZqN0AdHmZhfDXVNAIZkNI7PA5C/xmRSUMryJ
iHP5omMesSVyCkMK85eOk3hyC0NSWnBEPDTW5avz51GpzTEb64lZsOW++cP1bTV3
ClIoCsSljuMmacCLuALZ1mEQ/xzDmmIGg83dlrh/zS2yEOWrhTpFKIFzRO73xE6o
RykWI9FfSSIbNppQiplMaFzH9dgfq3PWn/l8s5ur8ooT86+qLGN3Hjru4i8y5RPP
nKMmSbjGdcRYlKwWy7E1mHxG+rnS48bIPU52OE7uLtNJGmuLQyaEV7ikinMfWloq
VMaQZjJnBPmb3CVTYyaC8FLtlcR9JGf8MrXhTk8lpOoGnej3fSbK5bJ/kNDiE/2K
1asc6ELNkAoFSalLhORVR3hHkI6TFpOrg4sbNzqaWHrAfI7b6vhONu1ZWlI8msp9
Ps5/3/HL6AarN5LG16k/iP298dG9uLiQrL2OsUu70YVg3XIooHgQEkvBYNvTQpGa
8CEoePVl85h47n+FDAmvv2e0ibhsQHCKKkGdINQ8qcT+UbHFRNfPFmYKmo0xjAHX
A3DCYbkG19gQRJSr0fXlWJegIpzpuKnpnsE+TvKJYe9z8x8IU2iS9aE13/ymAw74
DfThg8HbQ6xEvD2JUDKE9FyjP9E1qogYEMbNdljnPWWN3h4BGlxIQFI+n03mXXiP
wJ4B+HCtAdT6Yd6iGrDkUWTL4A5FzdKsRYGYutjFF6It/z2F1X931//L6gdRdwIb
tX/2wNQOJWKdNYv5qEIccXwAJOC2sZ3Ta2X7dQdtsIMcLmHS4Kg5JPYUtIpIINEk
jmsQdiViAFJ7CIPJ+6jVMJY2bYsYvy1RcG/eKvt3/AYGMTe/wzIv/axDhCx+jKtg
`pragma protect end_protected
