// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UtQOnI8g9hemEPDO8hqsyuWpULvqzHGfXfxobKT/FNDs0ieoj+e1dDJ6u2GaG9pskp52Kn35lYU9
961qSqcccEuSC5wfZKiUbiHNJOS2zq/wA6T/5mH596tAb53VVROU2fYkl1ELDCzi5+kKt7XVeXVC
nAn0EYK6WcuvOpG0znwT2hmriIxlFwxWUZyug5zeRs+mwWh+4f/mfy95J26hcLsjiUR10lc0Ep+v
mNgT5ojpIrIKvGHmuS2N6dfzKb3j6PiZkY10gIfaPZZwGhu3be8aWCNZSNaQuo9VwKDYJH190QTt
zoel9hYzJS3ZFFyta/zZ+VGP/c4AN3uu1/MglQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16672)
ho1/mAApjz4rQZY0394Nqak2+cKz8/piI2LdAda9advvrIRtHpYohaCPUsF+CIN/USHeeO9zmQpu
7qF6ONmxWYUjBqALyneNQJhF53aDZYNns8uHWChdlDELMavXwx8CIATau1AhBeZt+JIZ4Rxx52p5
Yv0x9W45/jAuAf0EqNFjlyYYdhQdTSOkbfLhjBPGeZp8hK5DJEZCsihYZHxu9LB4WQtAELGBFPfO
i88DY3UJuped5plBelb7vOggrRAAUou2eUECoghzValDW938xUzKLlpZIxo/voC/js1Hg1OYIyMy
9qo3deyZcQRjDnv5y5yheWXqbfoPDZxkCy8wd3WlNL04CSAwFMm4cH65OKjSSUrFYx6u2bAjEkI6
xKidmBL9LdA/xIFw/0K+o9PV6AVnMr84MvrsM15xaE+TF18/BJpGpI27KX8sQEzjlvMQWMU+mV4p
Bu6mOBn0vk8ll/XKjye0EoE1Dunam9/dN/DsWgNj8g86fbvv24gZ1czVZLs2UxpjRMvuqnSzGUMC
Z5C6QBPTFwlN/wfg056A1jT7ku0+uR8TgqCVz+o3sMVd5O7u6kAcAmyIpOgXp2QlemIKfPFXrMKP
2d4jjIRyrAH1c8Lrhmtgfy9hdEwPTWSZE9JpHHDWpN3HIPLAB54v8ztezb8SHLaMbG1Otbz1wOBR
kuGOYK7VsTMsqPP7BC8+XhTSDKDmkRBCJEFIjr/656YSQAY1hhDn00b8zxtm/plzZo78fyhPE29I
Z7oc/X3HgVmWXHjhgrw6Qc1uCgr3VL2YHueemz7V8CusZ7RY+VlTvG9qbyVjkDxjU6rhtf7YR1zY
r3pCh6E7zsS6zJ4L60mPu8dLAe8aKYgU9Q/xtfBoIADI23C25dZPF5NGmnHTXJHVrNpnfaqvriPO
Kf7PS253TWlytYiiXj6vNVDeW0gD8TKa0Zs2GABic8VxLkKHLlpPeRABcQLQDKnCihuyNkXfI85d
AIDNtLKPU0ncN8+aLBE9ofXHWJghaBTamYjsm6ErIDR+wlM/1Lvj4FvRIkbJg2rrrTvu/BT4iImo
cxjPSJ/DGrXxKdxChpjFcZqXWkuQd69DPtooeieebqL38kj7Dygs3NbW2RQHZEU6McxFIw2cE7MH
8D2DdQKk0am8XrqJmJyakljugbyKEEEfNzXKQwd8GyM1F5aej+SR69k7aZ76+z1+1FH3kzayY1Ah
cscv2EOkX57u3YdQ5bIXDCMkKL7fywoLdNuRlekTm+nk5Lu7YX3pl7a0U00VePRjjyAHSNCcdcw2
kj2XS0yS4kJ46t1VsihqipwS9tdHTrikoirJof/6TwR3BvJQhEsG1AwwTJ1iI5sk11ddCvp4UrVS
XizE2ZRz7O6ok8ucmNOMAgolze2PADXeFAcDub/YWEfbT5rfldEoiT2fehJtltLc3KsQQwH1m1vx
hIRWAEYgtMHknU9nf+GfAjPHBYSd6ctmVj7szfrOYKOaLqRwOpMLDdn4WnQ9upbEe25Mq3TUYgeK
U4AfIbxjNhnFvyHn/BJ2aAjKR3U0H7G3LNtKUqNhgZDGMO33VBZU64ctAqQYJd2aDxapR6Mg422t
gwEGDoHMVzMbUojkRpRaI0K6DTqwD3uf8HDHQ1fN5OHno5OWwi1eekbX1Xb1w1wfdaGJUFfm9y6f
F7qOA46nY1dhchcibN7iZDwHBnIA+0p0XFzt2yWRHJJHqq2Cz1iMu2xu89GKZqXeEaf2jBmz2feQ
TBDtP/TosqMgutuD4zunql0OH32aL6fSRggGgBR8XrZrlZSfxgPT2I0u6wfSnMJdSdQiyIhEvytt
KL6arN3LQTG3zTG4X3Hc9Zv8Dwr6LLw6IwSZOZMReHdac51tEARIp/p4sj9nA9FaElsyfQzcjoK+
sY5ehcraQglMpsa84qUyweDJ0hY2FH2ooRI7lsqhplRP0PgpKjc7QM+XlOESvXdwGyVZRYv8gJsL
qxxKcAL2O8NY2t26qj8wuGjVV7aT+3Vz0fE8j2L8VED2TrLyYPdwxxgSLdzEh9Xru0v7Fee3zAeH
vc+xpDciCiPv4WbAW1Xq0pvF8Co023IJfgoiC3vswS8QDOZEmScpnX6Ib4/InkSd4+m2EiD+7L4q
f2niGAc1VAi7Sax+sCqwtssdAGL3ayk+iJqZ24K9/4zQv3HxSFocOnSlW/fzhXjMnYt7dDosM1Zg
t/bKWAdm0ClCdcuhuPMYp8es3JxtVsY42nwaBnuSI0Tj5EHPSI7jK+x9iNhj0ZRoDmiY1hx+0Kh1
JgYMlYUiV+Ony/dNWfbT77jHc/RvVlM5ehnbIGwbBiABVDgIyDzPpBIVIwBufJSwQVDi63tG6yJB
9JbqzVA4sv/aBK3mUVUjCGhnY3T0g/IuHW2/n3QUhwUvsDVcPZUjipL1ORD0M8IHO91ElzmNapEh
lqo4mqtuaiFhZVGQDZYz7W4qarl8AiYPk5znGW+fobkeTR9frYCRxj0DogAvWoe0U305+6iC+49r
0CjnhBJAbDXv87jEEcXuOoSwoF0/KwUglnlXfiBU7SImRfrQU5sQvEGlcdpBv3G2CtSLeBKEvkRS
C2HQcttCvJn56xLEI3r8IzvV9F6LDdPTUOwsWXp/wDsu+oRnz3TdGHf5gEqARgy1BUHGIH1T6pNZ
Y4fRzdw4xJAblphcOwmMk0gfHRaIIypFpOB7E947mRbTAGl4vStNAP8u9O1UB6n+8RayP8mlHAIe
3h3le7FD4zXInIM5Ie8FHB8a2VAYoBXby9SAgOZ9+y5zbwvZyet69g2dDQ7cXyhIH5lCY1y4l3Wq
VM/E4gDjvPFFvrwweC/TE/xQIry/2CSgYP/snaioyGxqDX9aZVytFDz6CHk3RJLQsnDzV+zXbcsg
qs1W3yckBolzbfje9OJQmS2/GmjXulOShB6HEBPuDdhxZu8fkh4JXadSqjY+XJWaZnNMmAenY48S
kyS3Mp5oApwPVSHZWd4EP5BRukd1NujIJUeMZlx2akO13k7Eev39tLlN0J6h0iV+tz2feLdYqYt1
ID0FwGl8FFgOSMkOBBZlwL1i/hRjRsJPG7/ZXG6xjn8GpixzbJwzLm4limJxyXvyx/rM/4usgH5N
lD4xUmCmCijHGcEk5+V4b+5XdtpjIF0Qsln5lkVCIYC1le4PjG9lZw2HwJB1YxRo7xEulhVCmAqx
rHvasRA3Yc48Xw4gk1GqkJzh5dvkS54bk7aspOX1kn8PtWTRVkuO1DBGCSwaCcaAi+XunY40IrZq
lZHfotVqddHrIo8ZJwnx4IysW0MX/PancXaJUPAaITk5PyfbuPKvvJfR6hEsdomUdmdvrJ/g7WyF
mnsJdjU1yQEKBL42OJdBGNbnVr5w0HXFBJSY7iZbuNzBIIAjpbGLIeDmqKk4p8/LFSfq5oGVkLeo
/jrgQs6O4P1i5guXxDqQdd4a8kSzwwIAsReuRBdefjhlxY35dotlQjFkwIomt4vF89DmHD3l2mtX
XzSlVw9Xhkgyx5qR4IgJzyNxg7T8KGjUnK37Fz0l4VoWwHVhf3Q/KNP812xmZYVCqapVTqSTfmBD
xH59TaMIuwjFjiYLuhBSFZuYni289JwklQkcVzMMFAS0JgQG/4GyjMn811kU0RFiSRczCeQT0PJE
jlGY4BigaiFgS1I5/MKF57ViBgnE3fUhSbm39eF1a5OESqUNPJkEY29W2kw6iCkfLdVpBiaO/rD4
jK9WDAK5i/19bDCpQV8+7GAaS1Gla5xiCzQr2Y5eXcXYIOO4KLlRkGtmyx2t3nkjM8qntGcL7WE3
xOMlq+llvo09MkS8gyxNYfVt7kOsXneEc5h1BWGd4OcVt/fxpLkK/l+oQ+pc/eW6GHlZwj067xBJ
05M8RzBO4eNEny4HpG0DfsEfTBWdcXPPnLrkkOjOiraBjm5Q0WgIyOi62UpvsKKAxhPP6JxPnRh9
SkhpRSs5TKp+aacTBKG6DVXBPJxs0aziKA5A+cOJ3MLTprgYay82VQJkdWsr4YUF74M9/+kqJLZh
R31YfpzW/8o7S5Zc/iQL2us3hGIP32j9x4SRyFaDjlAu1P7l0iA16PgZT1FdCrJJHfaapywpnQUg
wWkj0TQIZeNDkq767Yns/DXF+4OeO+s9zAZP06X9WbataJlHQ5pgOhj30NnpunoALV8WKa1uYd/D
nVm3ySiGJmYT0u9PNINImGxBMX5EBImYSO6JeRWSUKtHxJ4jtc6Z6eipmm1I5Cl5xUJcKZybELPZ
DYdsirI7rh8ryKfuXMzk6NH7bgh+oNBPZleuGPrBSiZcjg+dOq6GQtQzkInt5nK8qIsp8Vvkq6JX
DNpTCa1jdzRduX0/YPOrNDtW2J8xL4Tj+YbdPGNL0Ekk9tdDlTI1O3NAmjlNkV6dhr+3GpJtXW8y
GtwBejHkXs1sjodkvwtZfcYfBDN6o7yqQWUT0lMebICwLXrWtoedbBDcc+n1MajDskXSandaphEq
KLqGcUVPKgN2cXEtdl9GWbAGduVn5BYntEadfphz6/xfuc8Ops3o9MKfT10T2I2UXtE9pbEcuXY7
pAqjRjW38V1zEBUg6ZIMovPdc2q8en2PZHFXBmgM6qsAyglCBF3GkDQAzRqcnWeKdJxsXZSG4Oc8
QfhA1VRxxeqsemOOcb+SmNUzs5CDtYD0Y8z4FU/Y0Ic6aVm8CSWF6rmISxDaauBIIjzKt3Ssxeez
U++ul6nh7efbu0SlkaaOutFZzvuXlHru7BAANENd8hb3pKAWP3sD3Hck5msj72KobMhG1h5dLejy
ORxxObByFTbkZ9aLcC1ACgl2LqH1XCUQUAtJYkKDa9b0iL+gMf1N/nsgFO9Zrb3Gc7P4Sh/4EcBe
zIY14oiY+SROen7ZsjZhpOsObA1KP4/H5T9mxQ+q1r1Pbn1GWpCdeXPv4BgEFJ6u+2VuU9ZgdUae
dnZpFN9VuByx6hiNqiXkEN2DsMxX5Ek7RXmtV4+oRdwTWJO8umpWk5zlNeuC5xq6Tgr/NA8e3X1f
XBy9Zw2x3emBJNa1YUTr9rVA+81U8ksvrw/dD5eAMaiPxe6kgf87mbc9gQmAOSdI05od/S1VXCkt
uun5RBQ9cihfO6r68lZM+nTFdxyLdIEClUHQndXuyS9tW0crYi7ijm3ktPGeq47bE1hr7IbWboyE
wj56d2Yyl7nYvEtslhoRVNRpsQB0nzpBPrOvCXK+0V+o4MSUHYPHXDZf19nALxMJ1vhROCGiSXJr
IBYAqJSGJ6/M1oyXjDRnIVhEjyPEKrs1w/KsD2/lhJyPHjOfm9706PpoMra9EVZjwW+TWb3K0ey4
4OaQ4LKiu36LKFVOfvsySErnXlQ8EGo0lACTwJTYk0e0RnXz30PXo/610oWejd4aEG5nMHSeR/Sl
3oYbMomlM6FU8qUZ1GQ7oP0mgG4TZPn8p8jEqX63wBIb2jiDySxFTJ5XjqKL8Q1XvhhddEgW5P9q
sSuM1Y1cVNGusy6bANq3Sw25ZwArm0uuV+YEgA9l6J8uFLfZQ83/eRKuIyZlivE+NUFghmi0vlIF
0NTdaGv7mKzLDYm6mUayTVnfLLcvyYuQyDM9uDX9jw2HXu21utVt/HZPfSmKKuZkymHUD7ZbzcB8
tadh4RHsJSYazVJEpjpIXI6N982iXHAcdzL0ro/309jnjGkO1xPriRm17FL26/pKW9xG+JkP3xus
+cvr9KEh3GB1NMAULLMUk2Uft9MKAt75sx0eXYlbolq551rgBwe1LTvkgmt0bJw6tMseQQ5eR03R
Rc/1PBXQ1oSpNSytLPINljfEiX2CrqZRsADr/0/6tfVOqLbR1FF/vM8PGaue07uDTNNak8qBks9R
py91Yp4Y++TyDelCqZmXg94CAv6qOfN1gBqpOQdd9r0fKw/zk6MG+NkglMQzSSZ0wIN80ThI6Q0V
mGs/fKOPC42yGR01gbE2rOFLmqg5dbrnAh1o94M1NV2WOBMimhhabCtnzznzmFuBJYGGIHM+L4n1
3UIseui4LZudN3rT65XCSgTUK5zal0MojKE0XoP09fk9X3HGrPco32cUoUnmAQna+cGcfGVpGVeK
IeN+DrFKRr5WoSiZAxo2/Uo+9b9DQN7+x2JO3PECzg4iGAgluy4HuvbMp1AVmb4EhkXBnfN3i9cN
puSmAQ2olQNSHxmhIdVyI7sD/PVjGHdzc3MkSW/F9pbaR/Bcwj8oV1H+AzoV+dFTquQGbxDYBgI1
gsWvnF1TM9/pjWw1WhLuJcEl9sBilCDdvBhFh3gVBoDS8Zq9XXdsXrm3kzmrjUGGT997jJf+UvTM
OpcOgu6HjeyVAVtIRGWkZqm/2FG4G0Y++PibGwBAnGuWbO243/sp8wrVRxZISzkoGSFyI0BTvHDp
ibVCJkqe6xOcSvDP+xZkH9K1JQIxjIyLRrdLzaGndR9vzZaVPj5nm0aBlpaBvxJ5qEFZtIqPugvN
lekKi2FZVmDNOSawIR4QX8U6ZVKsBaVBDOziAF7iTL7rAObygoJDSbi2Kt5Rqlip2e+uys5E5BPt
bTgIAdRkWLwOHeSl9Gj+25uUffaRLAe/PYLtO+05h2y0ypRPcUmSAgoasgpoks+o4oxBsbNORar9
NBdfYxKMjp0BHTquH9fRw2u2UEYpMkA3VLpOQrADLSQqMTiIMyJiVJqXnaPk/YkJ+yCsvv6nsbxo
Ut7dZkwZAFRAlRjw4SbrNQ/rAXs8Dd/n6VXpUt90TSMNgM6CzzuXTpvTKMAVnUGZunowMxgI0mq2
RMusruSbvlMVQ+UWzthEhEYfxxjVlc/HxgjxpYWSXYq1wmrBshUeTE7iW1Sg4/6F1q8WD/NQUn/w
ySBvO4dmQNQdZP/w7ieBXYR/fV3JgMlY/zO67h71J0g5ENEdKYVfKtUFz2l+RevuysdZME2uRuVu
AHmYQ7oUfO4XlBoFcRiQFGraGIzmUWxjIgPmEHw/58jFGNQNon2cpRfDsM/TQDxwmB3y8KUeGE4/
hhNVxt0fwmm135tPmGTZ5uhCv9PfSWI87JV1KF609h9SQ/aedwgi+rJj8qS8ZJNPZsG0Q6hPn8NL
WfdOJyqz9Dj6glmvsiZDqlKG+aVq3pL3p6CykKBc4lqsZdlJN1uyeFwUujvJ7aGnh/gCeXDCPlxw
pzhUFzfJqnJiPO84ta2iFQpT7suR8lpVkBw9GguZeQYnDiqG9MwAT1n9oOOU1TyBvVKh1cZ9P022
0RwjATl1lZvLJMj40lXmmNIHhhrbDZH/9zW2fs8ed+u/dmHAq+oGUCogE+R60oTTNgt8NUn5sUbm
060/vZAChYgfPLUs8+3NP2cUD71TFdlYhwhLQSLiPYvpTYVWopqY8DHrF86b0aFZk07J+1eDkuHJ
ispt2N8dXNVLMS9mtGKOuvJQ1KAEvA+8CzaEwZneJdZo8l4joeQqH0L7fSjSgE9wTgvUY8OnWgtO
wxx4ETgy3ve93iEywmn5WSMZQo1xY6ntYq4od54k/661780AeUaavlWl4wbCD9wlqPjJhRzYVIsI
gtOSPIOR6FObOx4Q5O60NK1p5vnszPTVHqVi8EfCHgOLJuVfPddPudtbw0WG+9gpgV4yxKWvo4jX
pFxr4kdslZk3muhmW0nNeh4SVUGushUngF+rHh55glZlkNPNRlhJo8g/bBNkvsvKnvqM8FbufRF/
b0Pu4r6ije6z0hububhptSRa/+TwyQsQMaevoDn7D7uIc+QaZ37GhKplxt7pn8CtixUL0LnverUn
Z/rYho3azKUQs/G6/3JED5R7UQwxUGzN5USeKwZN8hzhm0Shk7IPcGqED7Ybq6OvwDVo89iugtgU
TJpYU5kAB0SAsPs26Z6l3G1rt7cxp0KRDTE+Z2lImzhF9LSKAJFSfaOV2ml2h2U8iwijKoRAEjid
ZI1/FXnUm2xbcrfE3FDRCn5WdILZerTcKDQ6n1z1nRDgbVMwEbGZqJ70J2zRCbZeqJ5baVHx2EMV
RFtuuDwb9/prLlbfNhRdkYPG7iWzbUVgFUnX4z99/hOaqgYRuEWnXb5Jp+sz/xrlFuo5R/mHYLcw
DIX0szAfMg9GQ/IXk/ycvwRAeThd3GCHz8xZMOTG4S3khWvSlLcNMTLMvE0tvU9aTYOMICodULt/
6ETQL3JHk91ibfsn8mCNJU5/M8gZ+482ZrG7uArhvE12qEZKQAOFmVnfEfeLGs27U6vMi20FIW6S
bm8ZqK/XBTXJe5O3DvsNlFH++XBSHtq0tEzx2O+Aci4wIdu7etyJFp4gp2/4IwP8uyS4HwgocF0W
Vk2uQwNZeq53UtVPBu2vEAZoIXo0fezgvSBRaDpOuXyS3ltiWxiP/MwpsfwvKRXQ3u+BDeJHS5V9
mVQu3e7scrvAwE3QUndGVYJLCocEDvWU6vOO+GlEFXwIa8ZzeppWiRgeY8Qh56/Vx2frqYDffOWY
e0/vc+rxnIV4obk1m00BdA4pZaxx9O6761WNLOjmwwGgKloiWL42XjpgLd5IWeYWD/Ois++EIWyl
aME/it6HPVwUvV11zVl+TdQTVuSS1T1piLhX2AcfH3mvRYvTmq2sXCN96uhHEYFOr1xqf4a+MY59
fjKUh7l35Qn5dSvpn8FRaCUq2FOXwFdCGP6Q3W5OxAcDrFkAqFvmwrtLIrgglBubTB86rLgPg9mR
GaSmi9HCQ0jcciVthddCGJ5zd9I+OBARL5ITEtH5Z9et3kgTZ6TXwoS9UIwt16JwrbAKN/UQ05In
6b0WEixE+CZvi4yx3hyutwSbKxGpXFocHV34N7130hVpNp+Xd5CUVbdAD/oxSqeyyyj9HBNLW+So
BOIZAh+FFzCEqgtwkq0FIaVjEFq1o3FwuNxAIymdUQhdHwpSX38QKojsk42aOmL9tmTvJL4YOmWL
Q/XwNjTQwMw8xRiIFrAVpFP848Q2k/ygxtSU2XthZXVqTp2qchrUZYpfjBAyQFyhNk+051hO70Cd
h41HQSe3yFrV8QGwO55accsZxYsguyMFqFeccnfDQvBO4/v/cf91jV3hTauok+U0/Xc6PBeckROQ
AsKS2BOsHZ42sh1AizQapTqBIQTe/8taLVjzN62FGP3mdIL8cJ3dDunD4/DawGpyU1Dd+fILqz0+
1KUvm76I9je417Gi0+ELfRtwmpV0Ea2owQKTc93Yq2oNolI9lH4Bu74Fgv7tMjgEQgAU3H5J/ZS+
xYpZ4ttkYCDm76nKAuPHS3adUZnVWOFPVmxQ9vkGxeigwzEGrQvH/WuUO1bqOjifmzNMpoxhZ6CC
BvXTe+z6A3WIs/tRD+AkFbYqzNPTQ5Ve5D8zxUICrnr5zw4nB3qqKhE6ZplVtO8TKSpjuMlVOqhB
PrFiagA3GIvbLZ74Q640huX9pOX/AutHNekgmuDMQ2V3v/S303AnGbHKct5HgA7a/1MzKIx4nXrU
02NnwjrwMlPxbX32y+A1oq46saBh2laVs2OaXbSCvzNb+RdWWpeS/22XBCUQIWSqHS3ET7vEgF6v
6S8h+kppSB6Q8M+BE4y63wz64xu9sdglssz9ENOnEI9KOyEhRXeFXLX+UTB4ObLQxnxh6ZgxN1a8
sjTQvJ2MRdYECtqap2n1VTD2RcKjdt0SON/wksNZ3JMl3Lr1/VpkuBGCfBbd7/oINQkhkt0KtJ5a
t6w+xadRH6Nj4XuuLLtxMLbGlRl+KXdTm+U6G5/CzUR9eqY/uWylbL4pkQnhuv+nqVUvsv377p5b
Pcr3YhohFGnJlLR5okDlB+lHV6h0Cf7m6Nkz3ekXRsF+ccdFONXaSySEp/IzGmnSoUujp3fGzJh6
r4RlAmL9+Fpap2zxQUgj0vxtWyZWH1Hr/r7hjNlzShi8rKM+pirxiObslBw4uezyYBzipwwy/oyn
ppo6laOn1ceUYwPCaGfKkc7Q5AoqnLdk+p2DZwkQaVWWFi/+/hi4WhcFeFU+OKQ4tTMR/ZkW95Sz
psQ/WkHLyyy/28ArF/DrngR7CNKlI79kqS0ceKPvxNoW59yQso9jbvsNlgkSM49lTGE/MSiFgRSM
lP7hBKq0NBu3oHe4MOSfmnQfIxrJLrSuoKRm5uE1v/1nfgb21zucXLPTfwFV2Oob8EQzuroCexox
JUT0RZuHHCRzneyNPet/kr7UPsYzH8XF5Y/6uAWgFEdQ7iKvpmHbUXYYf54xGMVIIoEDF3pIDHEi
VjF7dKjS+Lh1njCQWYrTrCZqxV5OPMFQz/lLPy3wKksRW3vDtnRpTo61wfbbMQKzdJumkdS8GQ+f
OdseMF+y/ma/m+l1hp2+3/olVAl+ENxE4OdvIM9YiOusjFrRkRTFLzaKJLvOlc/UmmxkooYfP4GG
OFAGCVl4xnR7KFuY0yObRRgOstGz1oJeNkCf4ycCwrbxnbzOxX1U+srtx6JoVxYKcC93ksLIbBlR
q15FwAPzB1q7PxQjV14ObyGwEHdH73Kps3EpxdWsI3MtpN3cWYOIDNH7ImdTX6zgAXO1eiBFB1Xd
n0qNbPm6v57ll1RDkyUQBMdQjHRA9JuCavwp70cuhmSwSvvcHjRzZNwn4wJZQk/sdghajPJhJO3c
6Ia1y1v6Tx+lIndQF1/U9XJHYAKCHU4yH9mQYjNYhkDg4rBne25YIries8v37L5Qq4gAZUdSGXbB
H2OeTXE5ZXwO5XfUkYvoWpVGYrCgmc23uqExqC44PgTR73RXkLqMTrmkDJrO5fimBPkPEQbc3VDd
q6LVoOU6JpwwiAU1p8eVTOCEhShVegV8pE2GZE9qOQ7kfCodT+wUaV/wQ9xCRMgfXL0kt3xcaOAl
z9fjK55lRtrZcFvT4DfOBMqS9u0L0yXVUn/8to3qhoToS7YwhLZvgmyqdbnjteVH0/hgnND34XU/
UgursyxNqdfUmErDh9uN4y8Mi6cp8xp1h4fcQMD23j23uYGQcc5aXjZTAX9BFQkXCc/ax0+bMSwT
nJtfftVQWyiRuKUWfG1Ry6DoGpXX0lLKm2uzveZeQhip+kp9Buhpp37iMrkww3ybG8ubR5KT6QHD
lXsJWGtVB8zV4I3GTnJ2ZQgBWteC9SNOAdPKo13lIKPLdCjAkxtXria64O4csJ9DIQucNlbf6hME
v8BChOsVvI3FAR+rN07ujUHH6cw3kKfyAwcpiAQ/Un9suDxN02j7jxiaBH2XdduJNrjzWDrR0nw3
A3nQLTB46CB9BDqNAj0GLJO2gDEALuOwWRqxodHnq2eeldMLvf6XnBgV4E6tbC1NoVKWob3sFwkD
gVmulX7Q48g1xRWYNIvodxzKjs89SgOdrN6fcQ86IRHwRhYOhBlTEYfm356ijFXg74m3yad5QSQQ
VfvLIvni7OhYc8ViVRGYFmgndu8+3GAifTfjzQajlNSZGGL11fWaGuhuHwHe+QO2TZOPoO6rfyys
2QgQWH5u0prRp7X+vQaGuAZx+ygamVa3AMsB9TGtO+HGnO28TFmO7LC9o14mEA2bo5SizYwH5XqB
Hd9ayR8GNYPxRVG3bOpPz6PbOmDpWej8iJi5HTSfcQvCgdY06tW4bamJZYelTkg71GNFvJShVsPH
ikT39h6t4Xu1H7dbsggbPmLUCRlb4I/IStAjAbZvCwcJsKBnco5nvxWlb2y6HGNbUlpCBZCN8TZ2
2feBdqIt9E6Olpwa+1lRTLP9KZboI6Vzm1tSQV5VvbUcPpPvL0nta0fmQdJtmcYNUFsi4dffoR4W
sPqQ84IYoVR+qI6YN5YfTxAJT5AlmyHFKN9lTNuzDFKpt5HOOT5pIUs2hOIq/N8TzH8GU4qUVqTV
h8OdfJSqYhVt6iZTMjLFh07QP9Jv3WIzOrQRxQwqLEG1ZsFoXmABuFc679o/mVyJNWQJr5NbFKZO
Lcr/flT/Nu2ehVPRrn3NQRyhjRwd71RhAD1SSIDD53kd93iPGsJETgKBFwTZIs2XrN+BTgjds+Kc
j4QVsnVfh4If9mdkux73wLQWWU4aPkVDAPmWj1VEVfL/+7HR+kW2m9GS0tswZcDolvczBuJx+3C1
LydCdLdT2OFMI+UFIoCPhFSp+7T5KegKF4CYdpVLxy8Nh8Vpk1PcBMY5J07Rsf2vfDsWjcvZpGFl
jNz9DCZWuSBbk2xwN+b4dpGMQ2gvkTPH3NXWjZPaUI3bnAwJOh534djH8K3RAzSO0K0toMpA75zY
SzzK/1HXoIWO5bB1NkLnTWjsxS1ez9mVWSEbtiKbJ1+C+LveYqhWrPisHWdkU7IvLo+Cs59vWOse
5PudsFWj143Wf5YHSCD7EVrLNIhIw12XrOO/SZ6rjNe21UKIkFOgO1aQP2C0EEKQIsO1U24b5ogM
QkH11CRkFBnm/GsLr+TWe/JJZG2D42hxY17BMOJhE0xK5ccXaobLLJmAmMydXHXh204lJhIjIIIG
CvTMrHbcB2VL4aYSBEVceVBTwXiC48kXSbPaqtzG9kFut3qK5ClIT7JUXq0QkweHBCIrYh0fNU3R
spawESrD6PaSwNZ9Moat5NTjJMPQVUEOzOCwowU8UglczLNyHnmX20FvynWOirA5Q9gKEZNOiEkW
WsBcFZT7YWChklq00zoqTjrXY859Quamw93+SnkAh2LD6LqvhwXogjQuW7XoSHM2yGbnX6XdCAea
GgLhjKWs2JjhgRrgpkYeAmUI/427wycOj2moWcUsYuPmzg7JO2PxdzXl/f6cBNsnMCbZgy2z7L5a
p/QxtgJvrjGa59cjhG+Bi1/PiB4RiP7kSOCkOnaObc54wxh9r0QV2XWJz99xPEvl4ZPkufMq9fgO
6GaKtmv6UewC6a49EttZxdT749kYJA365g5oTXfWpQ4kjIq4KMf7C+varBKG0bzo7jYRb5x0XYtC
BQU/5+FfocVbTvYZ0BS+TW+0yoIxY/T7FqRaqLwnLHFA0LJzRfTAZISBq0KIFy3OPIryWjhtPVkN
HGj3Bo6MGvfBPVJMqxRqpmqqwNYHyPYZaNp1uJjFBIhl8wct9wXMRHElbY7dSDlNHE554FMJG14K
gXLsoYVbQ9jJ4duOz393BErMap/dt938ZfLmc/10MVow0Y7MCATFC9hKPixbnZjgp44NjTzL2QgM
45LjGOoy7JB9rugV1Mnm8YHZbu6+UChDmxkiwPnd5/2C9EbaiXcRj6trZnD4u5OwTLgUdtxSAB1I
blz3d5c61SUQi91S8Jr4Ohoy123nDOZ4zBZ5GWXjky6blKpQVgzoZ6Cyz4bNsDoAnpYV9+AlGbTO
XhN7sQfSaw+RkdbyPF4bLv/cmSG9sd95j2M/5y/GJkd4F2yz57adrpdPUAlwiW8IOdWtzsEoOfF0
CCpdDradP23LwjUaQNipWUFkYW3lzdxjMRZ86WkIYRzgQ624z1xJFA3AqlfI9cufvKR0FyEQP9vR
mY8fIITOv7/iyKg8ZYnd4fTtGmSa/I+h8T60vllGkPJELyJk1/H4Ekl3A+PTVxwn12mIz2/YoR6V
xoWF0hguljekRAzi+aak8S6mEHTlfOizgYMj7tnBNwYxbevY2a30+7gTcdP0fzfQVlDlhTmd5HCn
eELez6oomZkKuHWa0CCsD779VaWOi5F/EeKRWsOgJtckef/O2z3v9cQ9ZxsBUSK6F2fBq3Zltiu2
v6Rh1KCoXyh9aN+SlZY+3BMVWiVM/NvaFrdnFL0QLmJMvINJozikMSOtrqzxvbnlQPBE9vnt7RnQ
T91KPOjy73EbpTTK0k5Ss1An3S5KGvez+P7lj+TwcsgY29aZqHUqybVfOJXbR+Lne8IcVc9C7gFP
rDuLUzPW9Hq3+045oK9TByh8jb6EyDCRhVlsJRK2jfqmv3z8GjfRmMLeMSlrMM5qzTRy8cWN5RNw
uEj3G6H1GkBpBCJN7I2rFT8paWrCPmQMPhkgLYWV5YMu9FuG5HF4fAsYEkR0ejMeBfjYc/FbJTIl
zY8oe6uqM4trL6kWhy4YDsCvwqVzRLdcBMp9ETzoaClXK13Ch5bFcjOsOJY/G7fZS2FmPZoZg2Qm
mmhTJ0DvTx9EhqPFmBYZDNizr9ueZ7caFxxjNvxkIsja+b0Z2skp36JQCB2/G8vb4PM7I3mbkvmL
7q5XMltR6l2tuJ6KfUdbZnxb4pRXWQnIMUuQyMrYd71S278P2aUVLGpLQS0lhQZOYKb07qXACjCv
b6awQHU5ZjBsftXCTtH+2wdOMps45T+Ax/BgAN2qR4AepdX/+1ahgrS3tE0oakpLxq6D3B89mMYu
K+HjdWuy/5dpoQdlbu4kFw9msBbL4ZQFGPNSKUfJQl++EL6CcxYbGggfwqGplQ14FimL22drCBGq
Qo3mlYQa3+SVq5IpXwsIOCI/bnPoj+1TZhV8Cpk2uK78BE4fwz6SNzvvc9N+7eJgrCFxXvpo5WT5
sKtqFc74sYxjcNE4vkaU7/Hu+AYqV8Q2alA/Kd4vDkPWb5k8vJUS4IkJnguWW1fnTVVRDigVBhpp
cROUyLBZwYe/5Rw6zSW/UJvnx/Q+gTI9e+9Y53x4A71yZCcf1jp/rL0ybUI+/8iH41uHdVU/P13y
fxx1YiZtk54d3Nm2RqefiviWLe8rD7PIzuPcJZ4wXX1MLuTkLcurfBuFlmIM3ka7Oa0NQxM45HIR
Lkf6ZNFnZgVhqtpPer/XQU3HDu1/juiB9Z6hNN9V8ib00Ma/GJYFEosbQ6zih/vVmhJ3osB/2Pas
doFPPqc59z8B1dKxCzrKD22kUUf2EMtYXoN4d/l5Zx2e1BHMFKZvDZwh9Tk4lgkavZMVnlYLVXCI
I6hHxs16yy9/bY3I18Xdt1hD7nZN983vj/QZ6mgCn1jTJLRDALHCo3fHYRItcFH8p/WDkY6Nfjg8
A+oB+DityenKN1iNvIhGdk8dL8E7wYk1Ml8b0q6ZVM4m0IYsyXqvAFdqHaqM1YxY35XiZuHxJSi9
Oh5PzAIAJBZrJcdSAK6TKc/KpCXSwYlhxuIBTcgIOSCdLrlNRvh3Z4VqTFBCGYNnVz7dJ2eOzFJg
jBqEe3qVhP1boClk3+dCWTd45CJCN0J3Twy2f9O3RG3e/w/Y234YHYb7BJwcqIzbzNJD+EtbbtUf
MZNNEgEIVzexb0Ei9IvrBNUilgB8vBjj21J77VgIXooKCuFlAq6AYBVWACqlPxSZD2C8tEW+euCB
G0/80VDGuXEGzggnrPwOmUlXFGUCmqH6/kGfyKaBsKF8Gh5YxysVpjG44/fvP/ie9Mk23lVBSdmY
J6FfYE1oGMIT2h7K31cPbgHXfSlKBVrEfrDgABCb78H54NhlJW5O+tqS5dZKpeveeyrBmyYp5POt
DjaKTg45GqV+KdAhLog/EoTrCCJpU5mdGeSWSFqOuWXtnFBNzFOAf07mKZIlTOM+k5lHIKeFWNdQ
Z16USladH+qFypnQSGNVvjhReB0LVcF6iCChlgSqApvlpInrGtPYXRYP2m6imE7fzqiZ8DFtqET7
w6sNC1mVNXe0G+EK9WN2W0K5R2PYdYG5vcBzFDCHEb/8XWhmHzoIli+sCoNtusObxI/v8O2EEQDQ
fHqQQ+DDxVEtxoy/vcv/DDUqWFDBEdygksMgweG1k6U570VFrtWtssf/CYhMpZIB5ULxt+HK9jCO
IA2jt5W7y5FbchuGy8X0FDWnCYvx0g2nmfN8yr4s6apGMKpA0Mhnsq726SWh4qgEXESxfKrC/kFt
Rc860BaSdW4bpvge16N4tN15bUnQd8ccWuYfOAZhgHJWMake4npRrfMsUCR8bAc+A72r2OUZo+TR
jCu4aFPNv9QTu2T/TZBsFeI1uVrCxEK110Biv/Amh5QGXYPuE7/4AQQT6P/9fCMr21gZZSzIroLx
Zk3QvxU7bzVki5j3rpkbThmwt99yVLYynE1wWz+ycBhX0nuRXRkjffVuOzm4YF3nre3ZpEZDqZ0R
tlMI95Ov6YGAPMRm1W1zxeO+pgyRWc+dxx5JGeWfYbEPn+W3GTTR+TKhwLt0YgFMwFyC+kjL4EtT
WDiJhT9VyvkKjf6f6cWWL5Rgaf1EWciCBWG9dU4V5Y/eV644NA5ZnJbyrclOahEdUJryAjbeih8F
QCdd8l0qlP/8+1VE83sKCI+uW+N4x3YLz2nJGkwGXrenWTHpVeIlA/PTZ6Dqgm11GS5WrZmX6Vet
7x09QdSab/y5KzAVkLmwNXu58GxKtG8BNw18vE5Be+ypqU38O9GuZQ8WrGDYhAd4WsXmD3FoJB9Q
zubbgVEH95e+P3a0wYQIEUlAzo+i7+jzRgrSTHYN4Rh8fTRcyvr6lMOC9KjxzkYmFgyOjm6T3069
/jgcOu1pE3W26tESLp6D9dPaXI2C2PSov7WqjZCYyRWX742sOyhRs3Di55n4wi4a2vlK8elpZK2W
FWt6hRT7yWLBj8/exjzEUiYwVDhgPYNmWsIilnZfs3ysTc1leJUmCmJ4u0NqJ6l55nqN9iknIP6J
+9MpGuwfyP2hrGiHEpJxEOfPkG0r1IFU0gTv4nk1P0l7c9KvZyUEq2bAU5FrTrAblsI+QI5DJC2i
Wt4l6Lr4+ga1gvfwjhk4tlTkD7IHgrnDgnt/0IfB/XWJkNqyMIMX0GGJ9TDKLyNafdR2dc77dvWW
vn7gdiFFVAOPIufXMtuAx1Z3xm1viJsBfATrzi/KcXOWXGSAnxMQ04Q4I1q4gIel5uAFIbh/zhtW
iuNcl7WW4HUYc/PNjjWX2tewp6nyn7sHzNjht/dRuLd/n4ACm4/UhNgYSY2WDJCHpjVTB3dIiZo6
HphCs7guzU+KtS5usC/0qojSi9EuJ3HWnC5QxNkmQFoZcCfdcPwb4UR8MLQQtr1QvL40lZ6RhGNL
lq/3riU11fg2O0UirFnxqDR1KrF0B+kRuI80XoBPIQsERXEbHsDtZ6culQqkrPt3qqBM7qCHkqSR
Yguu7BN10DPMQYQuOFlTOUM3/pXW7Ahb9KoYWLSa7kaWycP+mxBoxBYCtdBWSXfU6g47ABhXF1Li
tNQAsmBjJkiD1+x2T+N9WGXKmlaH4PFt02MgYkhPcKZDjjmJhQefwQNbQGMQ3MBhD4kE4Olzmbkp
/pYg2Ir8D98up7GjFZ7JU34/jCSVUAGN01ierGOUGDpo2JOtFw0jpYZbrUQ/n8JH82aIDqybyMRF
Gm8CDWI/rT8uqcyzwTwsb+qjstekYmCEPjoI8V0haqc4HgRxipMi6Q26POACQODuLT1t4p7vlqG7
x34AaqvfseBWroJS+pinDBJN1Xgt9uwycwB6cXUJBqddkLL0mX1nf9GNxM2NFLypHoJxb++GSNnX
mrKevlf02srU4GCKaPDfy/kwxBdK/vyAh1hFu1rL0YMUAaRz5WAWI1PW1g0DE4zXMfBrIsJ50hiQ
FxetvwJ0/HLqgKb4Hd15oxJB60vUBbcaFWTFcx5Tuv18NL7Css8ybMorwjo8WYcfbzW0KLyFliiB
h9aty6YLR1NnJYV80RLe5PcLgudgH/Cdkjv3g1daHym19g/xx1f5Rd11p2bcTqNGdvhYdBC3MY0+
xpW0aXxpN9iWxOMzc3ZVy0IRzuQeldnOfNyrE65dpOggb3jvcb5KJX2XZL+7IWNIvpXLl07C2mVN
vvAt3Kr/JCKAoUF1Gvp5vO4xfQTdwDVALxXBjIRQB8zbhfwC1F4NLn6snXOJwiVoonkcUpX1yO8U
ykUmAHer1wMUXh/QR2JNSSAw5sQZgu+iMZfMPWWM6KKq1lpjUlPevFCD2HPJlYreKFZJWH/Wb3VB
NgNMBjpSARqpkSmzUDx8+mq2qf+aQWg9Rd/3mbB8JYnpSfJQRw4z/1VWmVU4+R34U9cX3YvIdrNH
g+bjiOTFTflGTMMjc++iVHtxAiDAKm8/KT1z5fqgf3vQuBG7y+zH039fDlwA6T7jIghrKlGdC3Rp
0F0c96TKvLJF2Rn5CgJkrrmZr/kKq9TAkaGErnzEOK60J4+31BpbsfeEefma3pyNHULbmUg6a/+s
fxzKDvsZhp20BwQ1Rovpqn14XqtWu6WOAoTW9K1YZxjNZo/ObI/gRqmztuaGBRxaTC7/MS/VhZnL
FYTqiMVQ8aP/3GUp95507DrBwkaHG+bJbMr/yZk6NvC/9EjKrNHQKbj1VnQGEx2xw2NwAUHhv2Es
aCkDBXPDFTb3wT0NSYUAJSjeNhRJZbEcDKXgyk03++0hot47Zo7nqG0xnkyOYg9A3h6CLwKT0L4K
EKNrDE3r7vm3BvCxBOXea+HYWd/wzBbnm7XgblaNzDmcvV6d5F/VPm5yPV35F7XApK9xisZCUhS4
UCj9ag/maPtf23Tzxoq8iV8EsVXRVvn0sLLDT2Ul5mX6qQ5ZZ0FeefP7vcfcHOsLhzaQ18K8jCDh
gQCTL2ETme7zQVAE18FXeML8OrGhOtxow2y1zcX+PBjLu1jI7i6lHecOVC4xTYcWlru+KZWrjXqK
sEPTdmBSb4J+fotsogb9V13hDOiw/byse03s1sgdGdkA6Mox+tHZEaDH0LWmfn33B41LtJ/pmgZ9
pVslVqlHiMxIiv3MYhUk1oZ+YevPAGo3UhFDtQzk8O44F48XjJNbTMu97LoQI+7svmh+t+ElUjQ0
6Wd0AmrgoSVrZCsJSPRiKW5OCjdvZLyp4XO5iJaqiYZEWQEcnP/DMdDb6lnKfOOMcPY0hNxe33O/
HBk6st8P5qQImsU+MNrvXf05aYCqWfWmJet7teYPqEm+bYUpO34kIDC1HWAyc2/9v6lZu0biKCUl
UFTiaJz1paS15qUTZIG4IPExVU1N6eKYmMf6W3e5LNbNJFD0pDvml0RSv7B0xXS2RCmSIiGWK9sr
xXKIuf0ysoVVY7nMPRwBT3BXB9MXOUFAJyWe4y2EFP3pUKsZuUapgYecdauMYmI6cDGH6zIPci8J
1Gz5z8sX52Cyd30CGNNVZnvCGqUhPUzI3rJea9zDpFqkqE8FBt3/368q4cVmZXqC52HxmbrkChjP
vdaR2h+jMLmcctQe64fTD5sLZVxFJz9Hh+RnALGbIG+HQrfmESXNbqCeDMNm9PNl2arFN81flN5H
j7iJYXvXOEq028bY1UYdrjWQFl+c2Q+9AZY5UUAzeSW80ncs9KFgh5zd71sv75Iac1HinB1h3/19
EO71x6aAWi/eOoy4GVA04sj/ZtMI9s3ejdYw44Es3MFUC1YcfK3Dyf7PlDG0VhqNJOLs4r5ciiQT
9s4vhk5jNLAtXQ/zPIL71l1h/vKgBkd4WNJM9e+Qm8b0qkfkxTPEe6/bpMYB7ySGPLxCdhiNP9k2
I359syRFBufKK1AWaw5acopk8i+RoJiuNS5HDXU3lFZg1bW0caHP9APvLTx0UqaPSMg234feCkfv
/46nuiCamv5Up9aWyikd4CpcZdcGJ/vtt6tHa6P/4zu88jUCnHF0oiGzUr1eFEHYDf6Ro2MJHqZa
7wTS/OE5hp+mmKpJIXQcQLOSan8tk+b1BRBN5vG7umRTUiqxcmfUKVXIm9GWzaCh0/M5As1BI4iK
l/Jz+LQk8ncjCAE12mxdGHVgrigJBO7mv5nDQvJlMUxr9tmc5HlkeLXLz0ny9WqFB5B/fUox11Py
HfyWQD8Gp17359JJOYaMe9vJeLI83lNoFiUxWI86Iy3q2v2JK73mJjR7PNcLLOg7j9qi5oRJH4cj
jr3V+aAc2XkyefQU73x1RHmXRc67sRYNw8kWKeJGvlexjJ1yYhrQEE859tKs/gH0uxjfdHg1ja/F
5I1Y+teGXqfSDw40jBwa3YhfrCQjPuOW1r2BYSsfZt/8uZq/VSV1VmeWtz8ulmGha5yAQyhN3RGU
UBx6ijmOyBk6ClGKsKbP7F5jLrxW+Q82SWd0Xc4FUwnR/ZDgSSUJTt3e9u8RHQt5UQWZhq78RWbY
d+D8C7NVcZKubcyCOaKNGNf6yj+LACvvjPcW6oWT8mCk61lFCR26ze1N6Rmk9wllLsTr1+GahP12
tUnz/Q+22Ye7QWq0mpxqaMGkfjnbmxXocLA75WzFoW5Qs+nM0MnXmWbguzNIwmDehnMKYUpp6duv
8HVLnsL5m9pnPaQAqk5t7b/I+7YbMgiufc4b6KL0YM/0r2dSGVntCbfUpnZzcHcOUlNZKCihU2tf
gnLfJaeQuXuQQFThvVtiRTyqO4V11oxfbrwdGxpR2H0fSTr70ykwQ5SZOm8iIAn/qvut10QSJOc/
njG2HsSZNkru5RuggT7FM/J36qtgdwAKX2k+Tv/Ir6J5Ljy//6sjjbZC/MM6OEq2HP0tpzcjrDGa
ufD01VOMgKbQhSrX/9ILq4F1S1aNmCnQ27YNM0m4+EnLe4kAGBzezTNx1KJKTLEHAALZuI+cQ4uA
sMcU4ds0X/OPREIr6AdIoJeS2eCCe+KVIyP792W1NxP8ydY17P6jQkTh2JCqRkkrqyy0jMBg0GOn
hzwlEHWOVLoxDLCc2CshWWRTncaGSsO7QozEQqiGaf+5Bw2yzypMapuUuaAkZyvAwfvvIJPscrMZ
CL/0CfjYvLR7CXwglNEfNFtBRpwP9TQh6hKQvH/t5psQbjZxt0sjNzedD1lNVLvx08dbrYDPVAZV
yIsWyUe8/OTmay7wMpfb6t9y6td4p9yLbGtiGuc5OPluaZf/8ZHw3UmhE82tgKjCNO+nUJzhO0b7
INj8R5L7Xcjes5/hby8DjGGA6jCf+uhCG9MRhSYHgFG0A95exJwZjqX7bACX9KcbMiQozAufx8WX
GO/zBdUu9ALYZF/ZsmoaiNArLLZojVDllw3l+wETfVqnVoug8Czz78SOaImd4xc3Br2D+CU8Ickx
q6vJEk0r9F0yvUOPjIkWO/Ju6mlzdZjEMXoU4pSC/x6rKP/5VhzbyD5PBJ356wCeG9H+tfbQ0pjm
WYqa/CrNTyXr8a5yEXIn8uo6M/GkBecbgP7XYXbzfLId51sjFcHm9yO0I9g3in9vstYGCJtFrZtI
d8qXTxh+5H0QthY5HHcdaUeUJ7wXBMgcf3hyi7sPH8HwzmswDqDrQUUVcvj8KVSKQjRqeSPFr/DK
FMNz+m52Ganif5UGl7OWWm0jMi5v4r7qYeAfWbjx0ovNM5B0A+KBToeVBxcDHschsNFzLfNSM0Pt
9zgTpH6b97A54juEHaKxfWBcDCURd3th4gAHQFDE6PhLRSyjCByL58rVQdi0O8upTtowfYPdTONy
H9CoT0K6qMjjU63FBp063ru4ImA0YX+NR6/Dw7RCI26IDpFblAm6Yk8/UCN3jXVckK29fZArjT4j
alscufVjRkWrahZSLvesS6lG5DqEcc0GUETddqpkX9QiGXhlay+ilrN5Cy6Kh/MeQ+9WIIxNKU3g
oHqLg2uEJL4KUuHfy5M557EHhhR2C3b9AVjnU8MwS9nirCq9lLKR8lXPCZuh778o1rny0x+bWHk9
1vLSdzFtwdCSM2tWhMO2WUvnd74pdxWvg7yH1jpYtZQ8AjlCd98477FbWLXq63l853WY99bQf1hc
ISsBh3PTpIhG9mwD9ciJzsi8AiY4orW3HOvaUDULZF3Y1AcH8uVgxxJf/f4TjYttFg1oGwpSn2qE
8r3Bc8DT6HNvFcIrHqm7qXi/bxEUGlKOIVoq48ut7yQVJXGscK2s29akYD05ofh1/ViEXXp7KYdy
IagUSCKYI+fwlfkH3TixP/+EYJ3l/WJ1atNqCouA+t49uX2lpiDKa9heKWqiu9A0KmwqWsIImVfi
SIiwqrTCsmWKvd+89ibMvzbIwQUGv58tqqpgpHTVm0So4YSkykr4DuiHvEVH7smAIfdQGEhPv63Z
1xK62HHHLhurATe59CpBiZkANT4ywWGWAdGfP1dykcfyf7UqhcPULoEwXjYvrNZxK/ZZdaUc9lae
AuF9JeZZMhr0K7Nda/sMkuUpCwITkX8RQH68N3iNTM/Y7oCnRXynJjPvVSMNCZ5ppbKP8TJbs4b+
RWlbTCCUDJCY+QoVjzMQ5VNlIhAU502/4fWH3cgUBJK0AvB1LznFMtLq+WL/uxKend/4JCVXrLR7
lHMhFWDY7967xCA30doTuRL6uxKQDL54MY0wKaK7T89yPLrxp6h6BNGiAdK00b/MF140Kp91355t
8kzzMy9C/QLTwRxYEnqvOnPcL5esDXIITZhe9HF/NcNEaj16eOQB3LpW2tsuonvYpEqD8eBMxzZt
Y2RI0YtW9RrIAL+PThKTGKTGS8ULbtoC4ds+EDt0vmM8zXszttNY4o6WLNFNUsfzmPH50qVXnvZO
9L5vuh0SgEtZEHnrGOo89gsN2oK688m9Ox47ag==
`pragma protect end_protected
