// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C2rAUL9xYIFmmb2iteT4gopFh6wXtIWchocIJbBC2qCPmwzqERQG4cwiCXDLEF9w
hHT0pjOuCDGQTRR33BFYVZ26oejGxgR7NNeQ188Tf01LCSlzajj65ILF5I3WYlU3
A7XU+ViyvjkqaZRg+YNNCqE0Yb3bw10Q9XEv6jTtOMY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14448)
+AePRL9PcS5PwquHEMz8HfLq3OwkfBW2kq62Kohk+MEFi2eXl7Dsm+Yj7N4ttbr1
+m9XMbfPgOe8WPocxZx1FsJ/3+ceZHnq3za0M5KrD6sqyCP41eRLnkf20gAdPKxk
rYQ7EuHtdqXZngMZBLcKwUzcpNSrlpm27mwtZi/MaDt8E77OeHD/51dzSUVfScV0
eboyhxECkjWSA1NzXwYlXpivEVUiHBO2cp0HPAeFU26ViW8swdavch2cA4ncFyEr
YLe4JpxsjjILZGUpfXwyZ2tXj7qL8/79OTpzlhpkhfPls/nddguRCRm4qGgO32qH
RUF68mxU37pgCuarYNrtlWlc6Vyd1QXLdTdtKQOmc2xUAyy6SG+J/3P6FhG5ZD22
D/kR99KGAOq5VurJxfRdHtmssafxdLr9zgH/nM9KzhBauq9TIYzus6TKayS+RQcz
h97CaYi7F6GLrFoaBc1ySGXfJWON9E24Jc0SK7gupnBYMb+5uz6HYt1kz1+TTe3O
m43xQZKp9pNaI2xjaL6zxspz/QWoKOwk5teku/XLJFefCPPCAT5oQcOJb+6fN04z
SgggIM4F2ZFRZsmTxgGjPSdCnN4AhUaWa+/hrvX/RkQNXbdTJjuPxeIkC3jgyDX8
bJFXwltagG28NEkCoY0+vF2cwMGzC7I52OKgm3PyUf2Ywf5WqelG+NuV/L2X0yJY
dGFq/THpW5UHzA56SNfuyR92pwqrq+lqJPgPXO3PDFJ+ehfRrI98Kqhx9vx6dsur
TwDkhF+SsOZ2hfwbPuhgWdnZ7dJ25EN+R8tINTgvNvbUxQevQKxAv31rNNppl2b7
/usvjEphZyjU1llYwt5LzEv6ozrJTITFwlZAupm0Yap2c0gDBzxRLxa4XtS5ijwn
1mXcJ8rBBWOjLiyQcj/CbUec5zLPJ36WJbDJtkEwxGcFAjIUw65VXAk1NRbA8thD
e08QlMebYicsgEi0Eu3NAJaDSqR5u2kXyMYbO8rCa80RCrBMb4qHiYy1YR79euK1
491UwIDThiQ3e/t/jnh0utvE/7vqz1J+PhiEDLl7bGVRUfiVdSKazaHHbvnGjycD
ZPR/tUJJtcfy+J0YrLIvCuf4TTlcflsD+p9QoglScLfWP1f9W24L2H6Z10+WhxVt
mHDLwy3uZC+xRMunTxMN4eQTHLNg8GiA0U+hzsHfoURJClgb9D5IecviQlAlG/A7
IuBcxtFczWvP+K3u6mFTARNq+3c+ScGU8MRb+FJJ8/ERXJJAtzas//115eq3nk84
mEjb8cyD/zVXpuNa8sq7f75ifGCnRLsSLsDJ6dJGsepWblrNMx0gBiW7EsAqsB+f
LAqcHoAKfWxw9j1b/wfgjssF+JpHzclQpOZMw01EMTaULXBXH1HrGI3LwzrJaFBz
RHBUgfhyQAiRbqm4Q5nbgZq1XFbnKjRv68MvPiK6TZ0hvoenFiNXyhn8vPRrHcpo
kWXkn1mO8wwBROBgHJFyKLZslQ0rb2HVQ+dcA6hIynPLDDVte5tVOA5ibRhq4ick
nITQfLLq869YoVR2uJTPV3PPI7x7wzfPCm8FGEuCWU7nzUKi+VXXv2LBGJEXaIvF
wD66/2m/I8x1RwAfRlWCtBr97KlV5P4OzxJjmQ+jn4hml0gqhxfbID4FTBrw+aPw
JIXpKUh68KqCu2tjRkDeYWQFKYb5HY8mI7EoJRwXEI1qox+15DMXxUqbYkHHhnSx
kuRgOXAcIdiE6Fxp1lAjV2EJBavfDHMMYr7UITp2D9JdtZzVpV/A4AqJRaFFwgMk
XlCbQ3T5r0RpyrzAF/VvPdqlevhYXe7EqWdr4fMZ8dW3fLfyubIMzsCwqXQa5KNz
hipmbAlHPqm9AWM+LOPEJ66dIkUocWTPUB+mdrttH6SFyJQzE08xAZgKNbWkSNwH
ZfpsuVcDti2LAzYsfAB1TdcD1fwoZa4tYd/XC941NMS8D/RCkPZmUXf03OjB2awB
+gWiNcEmfwtNM3ts+7TkMzlDDOBLQsHjpm+Id4eoTaB7xUmZJzKZGxWOPRDHDoyA
i82PzcSNzHTlUfjGjJuTYewkyGkoWhOxo49lXk1vA4AXM9eNqjKTxZZa7/oHLeyg
VKFdcK8cYECnOnNilOrsWvUkRolWqaZ1xjhnYq7F2hdHVxHAGS+nRzz3OVmUJqFl
FYt3wwwo/XffeaU11xVIIA9uMyQRfd1QmOt2OMjyv3tm182JKhKirNw2sTA/MED2
x1ue3ZdNjul1INj7jM3960pfqSZ7VasucQRHlR2BAZeP4gp6VKt1wEGyTaMvRmxw
A2KRYZrbtccz5cTJ33U0ZgFKockdvhUYUV9NHcyd2scO6S//XrvJcqb/Sgdf2abC
ggkehICpJsLcS8hvsLWrPlkmWluseaF5SuW3XExtJ+kx7y0IlCtP8zWn2b7rXbPV
L+YIHQiJabTvmIghQofHsRsBkauwFPo4D1jEiM9bNVzIjcVWSuF0B39vMmHIPtmn
e2lbom+kat7PLOD9ytePWZENZWZKd7Y/pmLGLE+NDcPsDdxgFazIG+5XoHwVjYRs
u/evhQQORtQqKy7vu5lDGt/UGJ0k9rPF1dTfOe8gldgk2REP9KRN3oNdwFx8TWry
Jl4G1Je8jFsJ+Inl5Tcxgf+Q8xfJi/yrdIKtWSRlt30IBeKC9ho8jO45FFrP/VCp
0jADYzbQ+jRaTrYnc5VP+HDYDPcxsdAWrH9MbmKEy2i/phk8XxO5CR02KCh1/ZY1
yoRGkgAi80V2ACo2v4fINTM31+vRyBnxi+uZZiJxPIf30Df6iLb1vNVeOR+0lwl6
nzBdBqYWDBmHhJJrgyvtljxldFoon/+GP9OFPsa3C1T+xEUGAT7bpQOqGZ6cpBRg
RE4rqxpRKBG3DYFAcFKwsmpeyGoYd5ycRTVmrZZAaTF3X+Vx8uOsm1bJ9lcXKC7K
FaFr/v3kPPR68nU1vYUVUM+3bpBXzd+3aZxP+1gErrd2COVTFl2btUpkifCJBd4S
InxuePgj/tk6WKoZx7cTPrURgFZbrdyIDBb96/KSSGdp5N9QqQ0F7ppKfgaT0aO3
/TSv7oZwiAPIA8+Oy/nfS6rLdZi9oMnZkmqXvX2+aA/shVcPaLss6jvsRQMLN8Tp
iDFQo+Mp8Td1YWcrKIlTYmFVsMq//IhnjZOo3FAlM7ovhQwz4PzoD7cJnMIDqKRi
MPGKMBeodg/oClKAPtp2EiZkj+2vipHVLezsXfVlGQIcQoN5UgLrayluHuMwvLRq
cRE9/UQjBKpx0BA2BHvWDnEw/tUjmUxNI7zxSizU49BgBnOlyVA1DMs8qzYqh7jO
7TE7sXJ8vLdSt8GxncxWZcSBMIomqDUlcppTcbD7AsknV/2gcoj9VMqIXVOiQoRj
qQfZmkfLFfeh8LJoCQoo2nfN2JGccen2XXp4vcrI7A4dl1gHqu+8YgO0hJ+XGyRG
CURmx5kQCPwOq9sZowWz4UaBhHvTIGEpuR4YyoYbRWW393uNrQCF5qjeuR1TlanR
t5m4aeSJP05pHNJKAA6ZtpgPYn1svE1OangDOCB2WyHedgfHjbj6Rst/PulEpa7G
/xDI1k8mjOJ+HoMfDXjDuoJdjvyzi/zm4eV+kq2UNbwGYm7a9W4tDEC+LE2xTs3L
7kTcC6OqLQVejZuhlEH/qDV7iG3d3OfGDEQAFITGf6JQ7TCYaNYEnLXTuGosdWqH
NAnP5s3YRvvAUglG/+iEY98l2InfyG4BqXOZu29TJ5P/azm1v6xdQLBlipogg/PY
Q1JOLrSxs70hG683X24FCW+B7hSWg/JSXnXa9lk6dKpH1rL0B5eTQvYRs5ddpQ+K
PfrSE3b2n9SIfF34Tj5bYhxp1QZ7lpy3LLhVNeZY7yFv6XIyPHFrEhuwTjMwsY2/
w6v6IJ9w4U3fdaWtt5IgFc4457WE71ITz+kymEBbllGTeth4XjeCbqlHKuwJyuim
3XxGLlWetUJs1/W+sSGHHtX6ILjGVbxhixLHrMutDh7AooQrvBb9Emt6iuG/uqaJ
clOhXwiOqLjklOfzNTiBSQt28zioWMSl6HhM7RJxJRgzsVtT5Nv3S24GYIPwtDQy
wyJ15TlQhnNVJUgMhYaIvf61bfa6rioIaiVwb3YX+IoBPQTY3ufDuPPwXBOD92MR
CnRQobwOf//y+dpC73GNgUkpCI/4TFJYXkfpn9LDYi02W5GgbCus7GMz938yMj8Y
VY86qNFONr4CMGmh9dwU5zjNM2jpsyWUqJByT1yXII/l81aMtdNJeJFQ+EUYlseW
kwge14E6Ttr8PRoecGycXT6mi840qE5Zj1vmjGalIgbSgcp46dQT3gi/ymgojgnO
uFG739PISYUrySdpxAYKFQ4d/ebhkqLRzTcO/UUsCNxtDsZn4GMhWy7Sgogyou03
FTMXfI2rXq50dDd56YzM57pU6r5cq79hEkW09k6cjf6160gieqXeiiRe6IwaHbcm
Fly9GnVJl6FApDdY7MY1nwMtj5n6/zErnfxWVvxk80TKlJb1K00cyV4dXIe6V/If
Lvvl5taraWEaicBmIUaFPC8GEYRbmo7gLXO5n7WPqIEXB+vAKdwIll96r5dRDBWc
J5OUp25kPUI5p+oKiPtvFFrFjDgHJxhDCNpmiHkPcK4KJ+9Hysg6oTHBi5+6Yup3
PjI5e1XgaqXeKHGoGASq6urRnji5rzSpxmDzNQ/L5q8zsSquSd1eevlc152sX1kP
iWzgNI18DHGTHBKn7yYcsxtN1y/Khaq7IihWssTU3HfY/AtLGfQYJIoYj8Ci/AXa
h1ZHgocXZZaGWaRvFpN3XtY7/29gZKJXd5tFy5xVDE5kULq3AacJBBpUJxwK25VO
11KMOkOJLMkDMb2N904WOxnj58tqQiASrDpVojDbb9UjNnfa93QlgNcYLFT0Lj9P
sqL4bIf1JnvpwC+Hu23juYhWfDe4JqXIPd/9mbTkrusuxdouEca9VkKcBuDq+43A
CU73M7nH2iDi6WECURzVDYGnK3+ehGAlL3xl2qihnRPDQAQe8zZTuHSuo2omW9p6
oKiVsfdDyocuDxTSqREki9Rxttsea2jwZ64mTdcFxCdK9SSR/GQb+r7A3NtuHIVR
8MsicXgRKqd0nU6n6RAZ4KzyUVupzu3hsk2Z2eTtmKKuK1c5vZKukaGMg667ho+g
6a3ishbnB1GajvyIw3G7mI/qE54jj3P7DTh0tYSGtqB0VyG6EJ8GAnCGGHBcj0E+
Sg5j73HYG9C+JrM0/S+hIo+sMXyH8Y45zNjeAlK1bXa3K5ihL1D8O0VVdV4qNMir
2FvU+4InuRigoAjmfg6rIx2nTnri+Wu0Qt43Z/hr0ocnSaP/gx9ORo9o4QkOyTsG
SL84mn9oD2DoYf7clR60tbg4hqNcBQD3l0jgeHONhZ54gRQ/ggICOU0uA/gKHajO
PLYydiP9J4t5SR42D8Tp0/2NeR28TMIAVlicU/LI8LOsVG55/wi2c/4P/UZUPyNu
166kISOMV7dPS6EqnG+EJIioCvgORvpEMF/1mBQ2u0qt5o/PPiqEjPXL2LJ5Y8zh
XhEPsakbaDhifeFfppAy1YUmC/RmBNMYxPIKAM7+asOSQropZUCnY6JKEGf/GBux
GoDoUQlIYUJ0XN1E5OIucYMhFoHXqaMdeU4fbH7pT41FIC0EB8RiI7ErpoHqlKhZ
SltEM+8GA2R9tOmJEstgK2XpZdysIrBsTfuLBoIVbRu74jfbTCnEJOpIyCzcqG0L
42KB2Fun11IWUxg5SggDz9EqZrL2072lGAt0feRYvhHSvSh9QBetdsWrUjMeOYCk
SdM7MX16QnsJEIUk/o6w8PWhuxxtNcbGqqq6puVaY+j4P65Fhg9Eru/hB7rANXib
drMiztQPrE/PsOGu63MnYw2OpQvREJNjHhLNlimh3qDnJJv4xtY722suhVEcdCuk
XXpdIfDJ5Ez8O81hDlqaFB8XqpIF/e9ysM4AW62DILYnjpxHz5dG7n/M05nOa5NV
weQnanUdJ/gSUa5gx8i2SXZaYRGDpwCGGKpvfePKGdfOneyYaFxWieHmqymAhFbq
hm4ltZ+nFEzcbiwqrOdeaU+RoVGSLn5n/XgeeyE8ytygx9VpOWo1Gojk2ygXS/h6
btIOuvrbk1GXIq0E61bMUMGCjuiKo7EFThgAAJIVmFYTOiKfGx0cahnsl2/TU+P8
zZZAtEe7VNiBzDusrLJpu24WftjnevSe7sPIK98b9E+bscHvINL3HnMK6YIf0SHU
+uzYD0qBf7DCbZWQ3edP5jEsnRPDiFc4nwa+IcxOHwAxF5QCxmzLyXfV6omGlo6g
V9W9LE8QE9UYWKnowjVpfRdRZuZzdyv8WVqjKWe8DVf9pm0vpOSb/J4VTWEhXMSW
yaNvsniS3lGE9Cwp9G63iHjHuc2xSoTXOgv7+qJmMpv9O4jPY8KycBLuRkVDOfT0
axxEm7b7FpUw1KRDFkTk8ffK2PG4BFGFe1DqpqZbIuUk04MXPe0lMmvwV2uMVuFr
nah0U/Pkmegk/tUBxy0JoNCt6Pm+JSH9Feve3Wwi1eQEI8XR5ZgLWXDNiW66wAxX
vPjIzcUlSou10ZsJRLD9Xg1oFZ8ccj6CJhP46RPiPtBeYD/LgcFNTNzjWDG45x42
Q5Ln25mJJi4I9qj55v9B9fIIENyOhtjSq+YRuQzLg+q2okxs3A5ng1NkzM94wycI
iYegD82AMbVpxlFcPGQRTTeGnmbHNWg6a98WBV8YofCMGDvpSEWxYtb3bsPeSxAa
wCuzLCqAwd8978/l0MWWTxeyslM940X3DguIQaCCjTz6e9EIv1Bda34lUaGO4VA/
7Gk1H0L8r5WvlCcM+tNyauaKq3yOWs+/XeTGf32MQIqAYp2VUhcOHJCXkLu/AiFq
C1xXGM64muse7qrQ7IDzfP/rFG2O8wESZ8oDuCKKKeb6q829QWDq/ak9xVJRg6Yw
kfmkGtkNyP0Yv+K6mcSY7r3wFBru8RA+bXxF0hE+JcQJV2BXuxDIVxL2v5xjwpFr
jrtQ7Ygf3y1nF4K52dr835HcYBrge/w0SpOmt33i/P5DtavYLnZ+VwLrZliQh7+8
9yDqNLiXq3GCvuwHpDagrdPTloeqzno+djJC7Hz6e5kvBC9RYU/UP+q/nTJKkBD2
YG46T6Y66lhrDdkN7Pi/uuzChusr1vkWyf3HVrn65JssPstJ/TQNjQeoFDNvzLDb
r1iIJeiTOmxbRfgqMHXLhc76b5NIThwBfVpj5fnrVWiYfBIlE9sfLdp84268dLUD
5xwBKJgWMrFyzZcMmHw/t8Dy2xKHY4B/iWUWluuVzkmZsJ/QTa/zhGlEMk/MJi1n
4ZUgZ0oB5KjD9KGeJ/fXQMpb3ztaHRJpx9oCtyjGWz/0DjGWRRTUwpLIvm9CAFGR
z1JEINQCtYHgc5/D2US/1OHNMC1BDS/HoyntylojckZp8HmLL9gOo/+RNuKNzl/H
oA2uXpPvboIss4kcvXowayecYN+kRUh+NzTcaWxHQEcne+j1VH7Wl03RUYPUr/YT
dKhkPaU5Ir0HRKC37Q4OVD6mkAavsQ5jTTgN4St4dnqp7V4LMnGwNQC/Vu/3AQFU
j/JFjaw2kUJQoXmNIrI9HUFb7nhGj9HZ/qnLQMfPLTpSDDwX1OfuHh9jsCNf57vC
cmoTJZnpsmQCZ2nxbhLdVgtdABPvufg1GRao330DAfnIFvHJ3l7mlgwOKocowMJC
83g021JASOmnoQLtnfeZ6IwOS1IadOccqSJC5fIcZr0VG8e77hr0tz+LKXcyymV0
wb6xoHxQhyyqymWkzLWb8vRQRPiaG7DOTRyC8iUOibG1ZfaVIlYc60Pu+kjQ2awX
FI2o+LAImdoSvneAtdWov8ZOxE9jSevWj0hrZoVuGMiv8BWENO7WcqiCX0ngUlqr
kGwahH85zsLahu5xuoI/iNfLn4ktZ7eyV0Eu+ucIYJkEU635DuAqZwfBwz6v5q8K
GKLaEfbzN/aXopQW7SJvm4qVtDOdLWPpMXv7EMtXTULiY/1JaF/7zzmlT++735mo
L/WJ++h1BLgY5zUeUftbUpM5BeyzbYdQh9GVJ0wtIKEPdz/S5qga2V4basos/d65
Td6mtTytbd3XwlrmfklLmHMuEl+d4Fp4qF9yPiG9+c/5U4Jm3gsK1U+BUipcPLLa
WtVpU09HSdBD352zA07zOsrR3knPxRgK9nd7/bKy6BypI+WIKOtovwuc1wlhb50r
iQfSEWUqZHaSylyEy9gsB7fYVwwzgym88+qdakI/pkUfRn9bcZC/1AD/16Uazv2P
Q+Z6oeOExp+/LQPOSS9+557sIi6+jDtFORwp0pfiQO85Uf0RfomExR729pJCNpNb
LiLirGo7GrXNnDC/u7Jp5HCESV7zo5OGy/CfT33EDOLJ2uX7sIGtpaqkTaAajgla
ss3AdqFZ72gHVZ6TeRokQjUBPhyQGifLblvor4K8a8fKBQELQQuc5H6qwRXsI4Ae
eJVkMyUJ3rcAKnjDhpIkKTAIB749MGo88wRTx8yydj+aZ0UW+K0I7QI9mVxygSV/
7FX1L4lCOy/sWHPGOxnEchh/kS6Fn8zrw5S4gFAjvYiZW8vHWE0Y/tSbGFKbjl0j
B/gTcsAxlFFgyZ8IVM+oJbvzDiMUs5v//nv9SR+8JKugJ7Cd+tjMnOqIJiiFjyS5
CznhwYR4pnqc+wSY/Y+WCgnnODnrP+7kRZh+s9aOMBM29Kx62KVg9s5F3hzasikH
953UUVVa4N/2O/AwrP1OqmePTTYl5xIIpkTFppdib76TxlVHAGrp4/4t3l0teBki
/uqpWxoEWtBBcXkq8ZFzU2lk3e818yYH0/9K3955PuWh54J2JQXTZpv2dVoqSi7F
2+itb3FtzLo5bF/cTeDDTPLGhwkyWFMEnK48BfwwzWrc9NPxMlb29+tuY3AOfGsM
aQU97cltVxbb7Hc7IrXP+i1O3xNbJxQcMYE+9LPBQVBoFgNEBMhFWQtpk2N7TNWI
OF99QF+fX0gVIZlilAOLgAQLo6uO4s/jFQr3ICdH+88lhMxKb2U8fEPQosy1coR5
qxEZNHjOlLwGT6774r0nY6LpKPziTlWB3sKtQ9bdTBRFJ9MNmvMoyiOWks36zB6M
s3LQZysTgJVXbpRk+6SlKq4p/t0dPTJ/0CvFwFq+BBOgq1Om9XiV3FxSeNu5UPxo
BpbOr0vVCkjUPsNHq29LdeGm1A2bl8+34mg0z7WLntH8cV+0AD1G7UUP0glLME5C
3+toJ6PqvncKOZFx4i+mx6KyTx5MSKEIuyN6lZvyb5mkhMnhc9duU/1SaaiOCAjj
pVzYlGoSqQSYHLM9QnDDFrp1EHwrO8WhIrFgUUoHPENFe2sc3ca/vu65Y80yhCk6
yn4yKe3Z0scf8yYhWKp2s3qU9z1yEoPYKnZRx0en7xNZjhyaLxQHZkoaMd/NLU98
l4hIgwP27AmOV/b6KNeonXshVEJWfwMI+5u/iDICbdVzDh7Zhz7GiFIrAx1ZAXDi
qr+gH+rv7ujx37u1Yl2ICFJYePRKXM7BYKyZ9qt1u/HG5ojeQDGMf3Frql9O5H3h
o2lRuq47LmuHth80leYePM/dWzPVqdWTakwuxg7yowRpkqjDyuFOgNU/px0tCtUY
ZnP6aNDf26MnxPGqD1hxeheEGWQOnxRgbX0IVuzySSFvPitEtUoa4Jp6RiDv97Uv
LDeC9SI7RXPmzbaErt4+0BDZ0K65I1fDtr1TVo2fQ9SKOyhcBVp/Phd0fuu2yTb+
CDvw1PrSQHcyaHS2MeH02cz1arhpJP/ZRK6MA5wf95pF3wwE6eCy7lDn6cp8KaJ/
0bG+bANq1EoIbFX37sHA4i3nd7cl0kQeVcPKNdyhKcT3SacIPp6sCSIKjLkqyBWk
S+l3QS+TNry2O5sXTFlANO/1TK38G/iMioM/daAQMvxa+GuKXoQ8eKd10uX7mDo5
ACq+udLMO3TNS/q47iNc41ma86Cg/c38D15QN1OmP6RBRLpct8yZ8JcDhpHi95sA
cm2APxLv7eDAefhqPctl0PABXo16SY0FQ8xKqb8FLmGAl79YrnJCbysbiEfKP6n+
NtxbnH3x1NNuvBEqnyQskLvjLXIonaLFAmnYKEFP9giOrovpkeGItyhtr1uF2Uyx
8lsQyfBInEKsArLuY3vNxn3e6o0eLqY+D0CzH6PEit+GMD+4HCAyZIE9aqF+mlIw
0xpmcigbN/RkKjgMcSoKBqAO3f4nPZSQhfqrNoP7ogLT/Fwoq86NCjJ1ZxyGd9S0
zIWubZjA00IHVEYHLYuXR4e1qcw/a1PxFwCM+PWrUFQRF4u720yIQkMn6nsLh7Lw
jWrh4NnijZ5it1kGb5qOTekOxS/uBESbic/flrRRASSw9KyNvHnvw6emqgFHdK8m
JpGgmuIGizALUsBUdZ2+usLKfR5LhOET20F2kv5aHY65DMDWGhGiUzQtglwGmZga
22aXf8uuV7uhvrLJtA7HtLArolKASrsH4ChS+YzeaMHUdR8VOzaLnCx5hnvMHQfI
iMuYqS1gLIck5b87SiC2Qx8yM9wxCgDH9+sCUE4sLSDEvHIn4ilhuea6nqXwj14k
ZXtPb5FEuNAQIux2Shf6mM+Yggd/ynGfL7Zr9Fr6NutOLxV1ZKZlLllp0IYV6DoG
IK0IJpNNXHy3rOjKPF+6xzN0JKY7eWDnfTSR9pT8fGtIQqsjgKZWQ8cWa9j6A3iG
YuH+rvcYEl9tjjBeKZxjvY6YM8w+/gGsTQgbyUsOydOuNglGv2KX5xHUwXENUDfb
k1rcb0lybYvH9yWJEV1KGi5MgEvIgFIzDkuRA410WWzYtde9JpgguE2PhLRG6vP+
FuAXfXgT8EXbQH0LnmEcRoVBCFPTJg3WRIc3CTMgEQvBlxXVecQb5hMI7jp9FtQd
6si9dHudrgZHMwTp7NvZGvijBsV7C8PJhXaScyXFjTHcHtdm0pVAK7BauGaG2ZMv
3dNM+J9Aae9AQ4InRjdx5Jl/+qZmSi/jxgdhpeSLv5fswabE0XWSPxxL8kzPxfe0
ZNHFKVQSDOYAIFO5N541Qlo13vKRuKlJGltiYjYCw0IMaArQoWigcdWs8jc+R1xQ
FxGDCR2O7UG5o7kEkHMcMr6G7Dzy8KeQenCGIDuoFtrK1xUeotGF1oBHKsGKj/aq
b3mMZEn6744ktfeA5F5OVcdx+NPpaQnAgdPHwGUmzL/ewZRr30K86OzCxlMgobg9
FEd6HXhw3l+WWaAa0cHJUvjk1gS1bd+5Mqst0wNjxClYO2w7F7OjkaAWHkD+eN4n
TWt0B9c4p8OooiWUHgmho25kYX5wXg609NQeoakfCkoR+jl4fmJYtN0skoVYEhCp
95mW1hFBCLp78p3DloZIz4wTnqj6LtdrhV8oj++8NxV5DrL3TrrbgHC33YIh0kUJ
BTwAQFFCUG5+D/4LwtkejWawze9amBnXO7/n9X8ev2D3CGnDtddvU3bBqjApXvdH
9JCAt9u5IeRO5tqRYVATeZtOgRoFFP43u2Dw6fHMVo8XmYKPscNbzM570BFYkYT5
/bSwhH86Hq/lcXKeRVKyU/sTWMa/17r5XuRA9nDIk2fZb1T2Sye3cotv057P1NZc
x9rASr2u+m1k6UCFgTFH45wRPe9xr9TWmUi6FWLbhLbP9fKwp/vuIQIpxDttYcM0
fh/5Jv8/a3+XsrZmZm90P4dkxDdInkpWGz6BaVBDUMKCiM1BxjuY5WnjOxeR0meE
sY6W95C2wbarNFikIU6bBczuxkDfPv4ZeU7WlrhsCWPoVjp1oK0jy9/ATSWeA845
t5O9h3C5LD0+qNlxzF0oB0hlfZXrUVdzk7JoqVNqMSWyyERut+jeBWNSN870kbTx
QzNNjws58kwC8N7u2iD1DTO2hlUas3jPF5BANn6j1RYhP1Zyow0uF+0xc1cGD522
BFkeBTh+SD9lGAAJpMI8CwffZGBu0L/0LmZM7nAKnse9mqqB+Z0gK0fsufQ6TXaS
ibL1SwQH9PNJKpwI7rM+TF9Vq5bdSv7ypNQQkQ9OGokNM/VFNwBki2Vh8QYqLg0L
MJIWLe75mxuftLgGmMNPySvJtGTHZFi5f0fXE88lx3URZAw26qEYqpXDfMEq/LVD
3CyvKbLlsMH4BLQKJywriDUtv+dDqRJE1aVrEw//DDcscX4aPkbtUy5bixqZTf1L
PRLAW95z9m39hpF6sa4j6F+VFn+JoDqn8t6kNiIjYwDh2YDh9JqWoOndUKbpZ5iT
rQd4tRUDRV91wd2mjmTHg3cVFrbit58b5blucphzhP9FXRT1JXqxw9RdzlObUuCB
g+oD8Fp6RaWplmh3imCHgwIKsye5Ikj9GjHS02EYkahRq8bQBB/DW/SnUA6w4YSe
c81DzLt2bzjMZT70NvRGeFH9lwkWNCoUtg+IERaIWYGSGhnPVB6UlzvW1Ok9dnj7
9kLIxbAt1jO+T86z8edA+4GeBrXAIgF82mVCC+zAuHoVypzDW9xXSjbGrA/IAaIy
oWw3IpcaHd7zEeP5yMIjqhtF0Dg+OsOvbtIuvt934E0K71DDG8/TSZerH3nIJneJ
bIBQXFG7GBvsIfqzfPjQGxXNHhuKIA35KNO+t/tPvG/dThvOkNArabzN785S7z0n
Me8ErIHPVsWZ6Qm+O5YZyMTOk+PhBAKfI8glePR4GWnqpQpVw5HJYIyqWfGOI84h
D7dGksqU1N0vC0wxCHcuQsgnJRXvIAyRgHUqqPx16YWJcBnPx5oaP8X86uphpwyH
T3aAjFv5teiztvJuFmd5E4YZnlettsyBvlGOUFN1aiDpz4oVY3pQGSIHx9QxUqep
WICd4lkOqp7+dggrMJFdfSu1ulggNGCeGsm++y1HNMStzqu6+ETAiLPOu3AeQZO7
Ij3KnGeGvUCZc3qxIf7ML4LoKHYTekvoBNjiIUMc2PJp1jd/LmT/7xRltWuNrMXz
0jwoVdZLX+UcX4WPYjGm40TdFvVJ3IGJJv3XqaZIb+rJlCS0e4K/AIrgPwt7Glup
3lgW0d+AkcFM3PNODsYJq5QAmHzqCV6nTBltjNxGQIepQU1uy2Ns5JQufrJAH295
YyO3PAcdjWFs+nVpUWHHkAFBKAR1YXDVw8GISAW+R81x63dHZ/3U6oSDOjbMfyJx
orn+SN3iNNfBkzdn+K5tuX20+rCBN/C26FM7IAmgNMD9rhobTqwL7Qp0wkpOQJht
lF0IiEB4OC2Zx/a4Q5U1Grcd1jLFfmHbFuW45OEtfETZQ3SveXehJ5QZh5MAJGtD
iQNJJIJO5DcdINkeGtjN3JF5kCynIt2P1NFMfKy/3NXkvCssWjrLzZ9jOt2c22q4
uWOWX2z3shq382puSQOe2qmB1BnBRy2Bajn3NYd+jAi6CyehUn3/iQD1BsZJ72QS
HaGzxr0gu0KHzD9O4k3sViWpq02lp9gOfjzR+39FSQhWt1KUtgE3bBSE4hJncqcz
0I/4TrMhyhD5TXTT0G/WFwXCPjfS9oqHlxE5Ybyjl1K7O+R4JiBJfV17CUDr0TOJ
qcuBDbR5dBmGmkSpgUFcINCUDBMfiA2RGjGbORip1kImEKW7wqHVo0etCwK4AD11
7sdHVFWo4nAIMc9PV+AedPtgDfEXlf8uCWjzMwJo01wYHRKrZ4949xI5sJnfvcuN
4G9AA8luVw+l63se2I6r2Gx6+6cU7mqhyWlNOzubfy/Ot72uEPXQepSFOqJOmVMc
HKswgMG+FL6aML043UyX1ZoRH/pFUk/2mBTkhh8vIj6VryDlQ/4MonVTx9rQEtMQ
mglpcLqzT7jkRRJJoptPBgkboL2OM9lex73F92FvptTlVzV3RWdKAd+R/X0iYcgO
nvyzR97SJrkhL11fQ/P/vyk7v2ZLEHvN/y5c0xxL9dQkwS6wvqp357G1SBU1dFBQ
FbNg7jfBCYlcZ34XfsvCnIco4Cke1InMiwlfrYiFrEQpbvU50XOQAGjBcwKmlmHx
UbZ4cIdXRrqJFNxK7uHe3Coulou5ACRvP8+5Og5PYE7I2DL7TV/Dugd5psgDkv+h
1+CuyA5f9Vw7f5Z9y6px0GOClrrsMf1jKu1KASXNLyUeqsv44NbpiV8jsEemQukv
8muVb+3VuPnjF8fn3ycOHCDGtRokLAr/6k4RdmQT5MgjauKMxfRV0zd/83IQ4Xpx
ZFQEg+CqtM9p4SkGNgowCBZaNlbiIpGwIPo20+11dZG/juS2ri7YfqrYRQ5qCDpX
siaBxLZTJgSj7nk8WkR9rD0r4Uwkmp2+oDelJpzrhzyTjYzmLIn4TDYimA8Q1R2j
fxCRy2ncXLBU66Okgi4QbUIURHWK0pMP01m5ZCo9jZ4JPfWe48RyggFP6OPxnkgd
JTlCCsY1rGCCIUbE2OGNyfr3VHC2oxSRMGvlIL/eOhmTSuInZGW1ckhSHZL1dnMn
0Evf+2BqWDqMtb0JpFUqAnhPSdwXYza/dFjpBw9/s+WkRgwKmoQBliFkch99Digg
5INYxBCERA0axNo61AXg9h5b8/TNY6XxjjF4xXvK4/87fLTyYJ2FtWmHjbIqsnJ0
PvD3Rs4sm4AYuc8BjybdGo1mOqIt42OYxUcxB2MkHdB/UyzIx5REvXL2Um0CbolC
u1J2UzxxEjXknojyHlsg/lt007LAIbaHN633brBS5j4pDfeeCikNeOLUdtL/7DiA
0f2YHV52Xus63YWFFfP0MkZrt2hkJ2sGkobAOD+kfNNNsO50m+YxA0oEM6wfq1UQ
3gQzjMDHv6Qc6e/MGMNfogFg9ZQvq77TFtGBjU0b3SxuT2H7fYcvbb7xhtdJc6o5
xA6puzp4m/JrxTzSwU8O8UfpW0ktwZD0CCeg27hFXIN53mx0rwu8yze+kxvXqFAv
1Aab9pa0y02v4RibnNZ2zKFPZ91zmhXB1z2bLCc/G7bNbvgx+eJ4EGOoit8ldbG5
WtCm1+NDsPcmhECaMWyqZDCE1IwrBXHpXazgwY+zV/z8A+kuLD4+mh77//igZ2y9
yHPj2nFnlI8ku0v9BS/1F+rrSQGdpqTRpLFsA07RlOG1hlPQn0PAXE0M0rgfHixp
wXyb473M2d560c8QWxqyPkQACaL3qJYnOsGydNY5fz02Q2+Zlo1U1c7Vk7VjF+tp
nanH6CL/KX9m/4LagH7ERa7PxfDqILgEoq5RvIW8+/3tbogT+21tfsiRtzV8G5Km
fesJpKNprUAZixFXbvHTG7ZJ2v9i6gVnwwdEwebVpChpWGticiVAQ3HYv07rXTZG
U/gi3HLjewqk+XTsyZh9X3bPxw1FdqzKgfHaYOzXu9sRYfehjMSqKe7fFzUgrdGG
jURKfb0lwjHDz+COX4QCJan/Fu3Tqb2YpRGE5rN4fsUuohQcTsn3XjHVWtvnCHy2
tYeBB8Nt47RpJbJcgaQISIl4zDuz+RVJypfbG8jAiEFbKZP9CFbSrQB2HnIrfnOB
wNhe/48kIbPRVYlQqC+tmFwBoCmFRJI01ZnHOPnOaQV/qvCk1WsZc2impSqdE9U2
8BMv0DPuQC4tbhN15MOGLfsoY+ZIaS+K92wSdACUU/rsXQZXifEwrlYQ2GhBDJJv
WE5hombfyxu+bkJJeO+RP+0iL2y5TQq7EUVP1xjKfbgN4m7WZiJplSwi7EMfepQB
5QuhCYdGiAO06/S/uzxGG4hF6GhJb37v0rt6BUhZRYgF+RpOZUVmqMmNISVg14rM
WuYX+a8RWybqRHe3DetvLv+o09IihbvULyXcN7IEAoiJwHV7LHqHPSQaqIS1LEt5
Z69oDRpO5XbBW9cg9gfHDxI4xrx8JMSLGMG99Em+qnb5vrMt0ph8az14kmIwEZnW
CrsoyPaoTuOCfMUS+I+1Ofi304DHn7P+j2Gn1qtV+Qdm5wbZLO0E3Op0Se8p2aPg
3oF3wR+H4kyiBKawO4jPaXOTOuF/95pZod/ZLZdxB8YavefMDxySPgCMLVCcJWep
VebYsVHfrjOaQLM1RbNyq660/VL0hzt+6dW+xrIVyhkxWPbirKvmVom+zHnFhKhm
8U4A3RWy+ekjhO4GNTb7H+mNsDnmQF+UOjXd0+BwHKy1y/+9LDLPDLt7iiGUA+yS
noWpKppe1GvBoMpK8eYHjktw5BZ5V3osuLZLAfpBhgEIoq2krhPSVJcWbLabbX5x
4jiSSD2/gBChKCDW3TO3/HAxOqtyq8ljYMVGJS0KwqCZI/dxxN3ZeFC5iDY8wDpe
b1UvMoFIiu2Fyqdc0Y5GHzkfTMPjWo17gqrzNsCqmek2Xn4EGRzbjDsmZ/lmcvgI
OnS+kIsM1zJpxZvzSjVEUZnPNRiKD7jDH9lIUPPP1fIuDCQw0lA/H//ukXg3ijhy
PlExm5oBuFzuP3uOcqH/NBUefqczhCbA5qH7RH8moNtIsN/LqLUUlpe8IVBYF3yd
ZJVpadMQrwvg7t83Z5Pp5LpVYAA88RZc+gH8SDvDKkzDWdUeujo9Ca2Ylh4FH1E3
0e8l5u3ePshIyylG9fnDZG8gsZBLTkiJ8zQ0p18a17mDetgn7u/bk8m4RAERcnoG
ItX6/3+x7uOihQXD1JJYo0ubJEXcy9mfAIx6Xj3V/NHhQ+9xkAqgaR5iYAZzUe/2
9tj364IrBYbXi2IhBHiECy+tTOMuo4vMQ0mvjt/+PCSVvA9gT3/0rh5x7zUH6kef
gGP1mkoB1VcG9XEKtXFqisyLZfuAfxYC+YtAR66dPLf8KBW5blstRjcietWPNVGS
OGYc6KujRO/c+85tpWjHu4LefYvr3hchC4R5eZ1Es3l1B6JAsC9noaVLxSl9wiQN
rK2Fapexv2JSU6H34q/MPbsS8OFQRPHwmzejeiYOxP58pEJ/Gczcl+muhijiazPQ
g4wbnNMeyBMF1WUPkrrLkaAPQD0KVExgZLiSuMwFYV6gmQ7TxeAlDhFAKWPP0Wwa
BhoQS8G2YwrSY0fg/fGc7c1K4oGpAxCNCH+OwDTRrGJ9QZNJAqFDxLbyG2UTJdUs
id1pSrezpiIYSL8JhMs338HiZNLtCHk3rzpgncWXw2fdhLRUEvbevypHvjSZ+pZi
NGQkRHGrlrjRIjoTG1CzPmLChe3IFBK/QCrQgO9uk4AuxOzlyXJfXIKFkjN8ocG1
pTJpFHhuD8LNptLooZrsA6iOLh5dsRVGnuFIBS9BCi62bCxJJTCBEVHqae1SuOJ8
ojpewbG9StbSZr6qCAwiSG2+Abz58+oepC3kgXioQhTJdG8K1h69Om4ZZEkLCUQr
2gwWvuFh5KGVwpPE9w9ijiwQjrJXZSvmu9KFVi0lJ+y/mK0gE5t9IqHr5tlmqqeN
USbkRQ6hwVCfe1PqSMwATLR7HrFftoEPjktVpTl0ahq5Ruuu0uPTxpmyoXd7wSZ+
EwlwgMLQ/Ad6jcic0Bw6di6tCLX1F+gCOfdw8LdsOL7dPwYWyzVWo65rukQZL3Ro
baX51d4seux7K3kLWuBl1E1xZ/hoCJI4mvYTnydIIvCu0Z+Krh+wFmdOm23YnoxP
XcZfPtNF8FMNGiDu/QWYddaZWcKLRe2MYR6WkVGpSciOpQrWMTUk27tOBBK4icHg
9ZZP0mIrVdL15gn2JIATbKOIBksJ0d0pinb83j9HdnB5Gz8eF07fDkkVpitqR9Vb
rUoyJGU9Z51dPIBiO3S/okWpdc8twfR1iOm2P1Z0QSEbxh2yyyRNWU/kdStj1Lmk
5b6hVMKMM2BWcq6mYqNlrsnEko+GYAhvUjnkvVyfJF9nFkeDgfAC2sySGFK/bNyf
R2ozrIIxja/85zuFnU1EbRfcwNrxvZqFyHL46CImAhm0RSFJ9m1UK9gU9yWa+2oO
actXNKIqfd+EqYm8I63hB01MLM/+J1R/klFmnh9oDLYDqF2Gt4yDkUeg/74w5c7W
V/mcQHQZmFMF3wffK0iyuv2DALSn/iVWsAaUmfFuwQQcCsffPLGeoaoTYrKxjKC8
E5UAtyNhaMwugYy2SbiXLh3a4VuqJOv+OUW/17BcmnIHb/CWSobDoFFq7XN5FE9F
jDFDP38dTkp+t8SXA+DPELiSKqYWPbcyj/eEd2Tx639VKFh0zPjpuhXxMARIX0XH
LWQNsCxPsT2nzDPfmS5yPfd/Zp6EvarWQ6G8i9plhKQ9pl+4UTCYwdyggbTcp0E6
LsbiULEnY53Df+K0JI5TNSc1Z24a+0PkA9AE+exe+qjRBsR8g/MN0eK1X1ckaRK+
d27M973ZY5SCFT6htzY77+iCQjpqHFjogGn2Li5y3XPocWrCvcyA8XVb9V9ryPA0
RCj8yuqNH2yctnnTqjDjj/LF4/1SCnL8iQ36a1I3w92flQ5hDCEL7xuuQf/km/IE
LOUGj6OdjPVWkSd4yDgUxpAtKdKe+2O+bVj1DDH70UkEloJeF2R+vw9ekG/R51Lo
6wiD//pcDzD+63NSXkQjFadPmjP95yCvBAGzBIrM+RbQ8oM3PydcL7WGCqUNw5yv
4mmsQ/7aTjfhmHXe4vAoQpJTYxzZapUHkcsJ9urAu84iQUoXpmxxKeLptlRqeir3
8aEvROIpaKLHMl/NcFa6koUpcXrZJJGm4Bav0WYCavLQLHWY9cN70M2t+pbvaPiB
ZovzRPISraC9VKzbsLPHrgDuSqDEi94dgQgUD4EtplWAw1xo2uKIQKWtVz59Mp1O
HWq+wzS/EvY246uPm/RRzqpNLw3Sq8rmeMWbhWImAGXdptIEYbH+1DrC5QMgsvg8
B3MShWBatJKDUaOjYn7G3qsTDDpVeLGZP9C222Q+m6uU6orF+MpMjnJhEIHTjh3v
rTPzX7Zc6toTszSBJQVXEwiPR5ZezxlKjxV5PDT/kUStYfwGU2klDJHUxhBxjYC2
xxXYZd8erIBAR44/2SNs7cFPxHHlGZSpS+jNkAyKF0Qq500JhGSJ6sqdLY1KQOVe
JCKgaGRkkIs8QNHgof7JFWZhDrRxCf+sj/NBFuPtUcG0lhUH4bcLiRxs1fkDhSTo
24A/vbMYJ/fu1h8U5ZL/ZhqXB+0sTxtYN1Q1V+kWoHKXeQF8sf0Iri/4YV/AdjAM
rE46J1QCmUt9/6NpFRMEqaKBg97uzvCfQBpuI50sqGU/611chg/Sp28WC7DthABf
mIV12u/d8e0OT9kw5B9qOJIngMEJrxJZeqHvCdmwhVAFnALKCcJTm3bXl2f9VRD+
T1MoI3kvgTqjrK/DrBJtyLXqcRq577Z2cLYry0g5RLP11Z9Hcn8lwnYj7xzTa46U
`pragma protect end_protected
