��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�@�w�4s%�mH䖹��F���xd��;�]��yw��`��� 7�]��>�9CV)��H#ڡ�0�����B��T���~���P|��`4�U����ׂ��5h���{�>���� �3�{3)*��B�\�����Y�(�0����9�����Ӝfl�*����n�s��2�T=�`Y��)�>���꿋Z�O6c1K�yAf� H�LT���6���o��R��]��8X���8��|:�).�Iv��w)��z�G�2/@��C��j���\Ko@A=ͣNcWa�Z9k4� \�F��0�a��nV���Kn��F;��|�8�*���n�Wr�;��Tf����"b�df�s3��f���9�ɣ_�wD��z���ӁhӨ���sO�e�Ƒ-\�3���p�r`W���\<��0y�B���놝�A�Tܢ��7
�]�
D��mkjb�M`�F�TG�UІ��-<?�"����kiX��:�╙f�(�������W׍�s��]�@�
��m�����U���Z8	��3k��Dt]Qp>]���8�qy���(6��{"d��l�tp�8O�E�����evMLK�^�]��~_U��}��_R�8 ��W`J�?�0ڣ[
D�A�&��m`����H�q��ɷ�@R#�K�,�:�;3����MRed�b�L]�1�I�NM�@`��$S���'-Q�7�m`�f;�4��aQz�F�1�E�A���G�,�u��L�Ϙ��nU�<����2ya5
ZV��}���<����oa�n�����ˆ<M9N��-SL]�rbO��lj6�P��h9���u��	�p�P(�e�>��)Nm�qb�g��}|G��1L,((|��"�}���,nJx����O�TO]+�g�����'���GG �X�T�1�����w��7*!���M�������K��x�i�3&SO���]���7�H �����y1�&���hZ=��؀A;� �Sg��GbC�	��M��m�a�֌E�-���0сU���h����pʴ�B)y�IE_����;4��{|�'�x%1|���X���~jۥ˷1�@�����`�R�j۶�Y �"wOh���b낆,8��l�B�h��nh�z��i��J�'��pQtY�s�Dy�≕`��9YbM[���)���%ZcBTS�KрQ4�H�zG�]�{}/O�]���3RqA�Dfc�.-���ѐT������Q���k�)aD�z~:����X�V�4����z|�%�N����i��8H�����kE��ִ��g�L��E`iຑm4�`�#$ر�8�u/�_��	�[�G�9Z*���6�*�<�;��p8`\�N������`��8W`V1��h}��ɦ�Rv�,<;QP�,��<���2!�nvG��̲5�� �~���&�LD�
v�Z�R���^��ǔOo)��dGi�t[>ߡ�_�0'�p���Pn �c�U�����h�`�S4ݼ�xH�~�dC�|��� �2A]9��,����@ۧ]_Qq�E�<?u7ޱ�@�}����qS'2������8�0w�,)���.N���۹�t��b'��ڍp��iX�em��"�ω,�}����}���ى�}��5F`��=�p�ĩ�r����:d!}������b��kE+�g֥B�־씣ńK��r�jw�����j�fB���lsj��zc.�Ҿ��1�V$�DTW�~K\B},�ŞM��6Z�#���m������D9�</��J�>�����'(!�MDɬ����GU:ͱ�+a�������y����&s��D��7���i����Ƃ�r}"��W���\p���	�,�u)���~��5K *	o��0��6�d 9��<��`����q=�٭�^�|�}�t��Y8�96!���c��Qn��ؖ�
d���6���^A��j<�v���GꞄ�-A�u!��u�����y#�KZ�a��m��[���>���mb$������H�+��Ö�y��"<���q��=P,�B�����j�N�7�Ep]������1�Nq��7m�T�+�^H�$�'\�y��TX�lR�ύFpY�1�����+җ��Bv�_���C]��w=�U¾����l<6D!���%1�ZOA��5�kp��~��h�BF�`�0m�],���C���Y㝄(�\�F��ϟ���e��j�rb��s�R���R��`L��.��NE�8X��zs,%��`�+�S)|%�u�9j�X��T�>���p^�O��p��%��VΔ��d<���m>�
��uZ/F��@2 ��N�V8�5u�0|�l�I��f�&�P������,M�P5���$=� >���}Dn�w��u�g%?��-=�]r��v�I$�?k�s�s��&1*oܯ 9)�{1��5�}���$�U�!ȩ3Âd��v~p���RE?5���'�w�KY髲��D����T�K�I�0�"��b۪_2r`�<�y��|��e{�	6�o�=.忕2�-ͣǀ>t� ��2����O�>��we�J��z�2���CI?�,�:@ڝ�b��tï�]'Ȩ��eL޼A$,w2Ft_����ԑ�6�
k偼� ��~��ֲ��4&�#�cIH3
<ښ��_�{A�񾳇����DCc� �}�����2ՊeP\�<}��#3+�v��hʲ�L��Q���b��E$46-p�R�m�8�d��a_u����&s7��;{�o�Uc��&��� �*n5o��T<[5���r�}I�Y̸`�Y+�Ap�Z3�ш��[�E�ZY�>�z/E��'7�\�j�ү���[�F���� �+�>�f�������ir��-S�ڪ�uM�X�����'a�u���e�za{OX��PB�`�Ut*�1����w�;pmTp�nGڐ��:��ǆ����-vKs�b����giݳH:/%����S��5�"�p�$��0,���53��8B�@�ͧ�A�y��g�G��N5t�h�N'9�
E\="��Ѷ�e��- ��8*�+�x����)F�>�3O�x��e�BUYu���D�0p6����E��{J<�h[	N�1u/s[ِ�QK��C�cRC�%o����x��h�3AF+��	��]�f	�>�qrN+f����x���1K�7�ٰJ�nt^Ì���l�)�K`�p�:?R_S����0�S<;W��:?��
R'VLy�.u�.����bd�4)Z��"�G�S}.眱 �T���M_�i;\������i�s��u��v)�n�YP��]��T'WD�k?��@_}����x��!i��M�\\���"U#�ݐ|�nhܸ��Yq�|T@��ga��l�z�g�|ȉ5:Lo,��=�"CC��,��6@�|�D�봷(V2�Hd��΍O���x����O|� �gtD�y�R���ly�o�e
I��[�j��\���=Z��C�f¥9��bE3ۿ����[6\�	�A\_�I�m��{�����W(O{̰WI��uڻ�=�.G��!	��Ew�S̽ � h���)�0�Bc��"���j�V�q���;��s���`U����l���C�����Ⱥ-]+�#^�ZW���%���X:�o��M���㖨��5揽Z�����ّ?�]q���/BȺ��ԛ��Q r�1���Y��y��M�+3Aio�F�f�cPڭf��i�.�(�iC(�x���'���\gǺ�t�-��0���|A���:aF? ZHəvܟ��9�i�3��&x��00�$�S9�����A$~g��%f��#N�J�����3����I�j@8[c��EJ���J8�ms������{�ݪ.JJ�U��`���s��H��z��;����L����4��_*z�R��Y��B�)� 6$�\JB�=���k��>wQ�%2E-ٰ�%�M͊�D�4�yPc}Y���1$a��%�S��E�v�T����h��4 ��"��2)�fGd����Z�M��g�b�Qw���T�c�ǐ)+*9(2�x�?��m�w�\P���e /���	cd�
'c�\�S�Hƞ�,�\A9n�
8�A�n�����m����Qe�Zk\v���x-ާ��L�6�=~RtY��&���r��|�����.�e�*�/��)p^?b�p�zm�b�jc/���٩��[��)xu��5���m�x�"��WK _+�L
��׷a��+Fd�e3��h���#;����LT��,�p˸���h��=���l��?���"�����I�*Z�\��F���g�i&ô�L^���oB����XL�A�t����m��`� +�$ݶt�5m��L��z_�,*���V0i �_����'�P>ci�m{ ��,�jO�gu�]f�}*Ŵ*�_��REm�ײ	��T��.�C�(��fg���)-��F�2���"Z\ꕱ��ޣ���r�n�Zn#�iw�&am�.ĉ������eB���p�"[$y2q�Q�5�bN���q���Dd����$�^r��@;M�s߹�l �G닍i�K�;�m0�Y��}U����}���{���K����̪A8�i��r��%	�5�G�q6�����Y��&iV|�,x�H�iqBTF�Z���:.[�fo\1����/-���D9h��[���p�Q�a�`΀%���Z��(୼P����Y[��\��u�\p~%�1;��
���+��
V&cU/�<Bͼ���i��Z��^�5�����M����'�b�YXW��>�DT��l��I�Z�hi �<�`�l�%��p�$�S�:G��2}�4�	����R淎U�>`�NAm��{ſS3���P�O/������3i�T�~}�gX�	��|Q�ЋV���+��(�"W�/�#��l��ݗ��JeI�G���W��n��e�n[��R�>�@}�%�n�#?_�!*;���Mɍ��i����0��Md6��wu6�D���7�C�Q���S��.wt,2�����! �eUUU.�ۙ�m!?m�D��� ���ІA@��n��)��*%	N 6�� a��f,c���<������|�l"lfT���q��CZP��X�v�6�Z��	�8�)���^��Dj�iK���7$?f(c�o�P� �Pa3�$n�����{�I�(�,;C` �@Y,��<��w�px�a�*�Gq��)Vn����.�Y�M|��$|�k�r�=���Z��R�o�6*����`hGS��O�߅�n��堨pab���B�#�bs
@���� �����gHx�+�R��̧8͢�yR���ώ��{\��C[��~�;�0HJIk!�ANv���]��Wk������>�������)�� ƭ�֕0��8,��8����`���tČ>"5u{�j ]:�?��͖-��)]��٧$VY�RQg���~�gY0֭�n�?��ܓb[!2)������JhLu�n��]V��⹊Fem������Z*	ok���yk)ҩ�W��-%=�R`볰����Xq�/Y�|���-��ޑQ���/|����A��s��`	qWD�C��)�Y��s��2hXNL���B�6!pP�v�J��ZC��=6�����P�����켋��H�w ��.V�l\Fj�y�~)؆T�s�������{&�0H.<یN�ڀ����k{�UbZKiF����eL�P,�����bWka�*ל����!3ڨ@����ɂ�����%;�LӀl�p���3h��wR�[��m�kP���-�R[%RUԾ4qMx��U���]�]`N��P^쟣�O�b?���TO����M,oh�u�����4�)B��3��	~��R�+͵�b���[���3�۰�uʈbS���F0�Hh"��p�c�#G\����t�QR�G�ӝF1\Yف#��ř.����z6̀�D�����ǧ����߀y���d�Q�ֵ������r���ыC���'e�,ǀ��d�뵖P�d=���FV8�Ǌ�g"|=j��N�T�y����qA�+�G��c�=��xD��\n��y.����bə;AY��;Q�В���B��xµ������f{��s�8��kB˾�TaYX���)�c���ݒV9��T/�%Dlt.+�m�����z��eL�J<�CƐ�g��8=�Q�&�����w��:��<��vx��q����}��AhL��fq}y2�-1z�eK�b�B��W�p~��?���{��>\�V������4��OA@i4RX�S�IT�kAcW�}�*w0�*` �P��C_��܈W�N@q̄.���I�yu���T�ڱ���l/���D�n�����E�,R���Nn�Ƅ�Y��T����-��|�m��v�E�t�űb����&��C[&�Č��@4�K2* 2��cE���n��D-�<���֪��gv�{��`���1�x�{�̧d5v}ڦ`9�~�Hr��R6g �ڂ��Ƚ#�����1�\��D�_��yk��il�xD8��k�yi�p0`�d�!��%A~|"�ix�y���c#x^�� 	�"�ovyTGc'����'py��O�Rn��'L�<�C= -��Px"���5fܘ�V��ƾR�I�|�e!b�s�����&I�		��+��܊n1;�����t��������W�;��{b��e�h���?Q6�ٲ#d�����K��m/�4f��ڳ�?�8���{@�]<�b����LPv��I�v^�۞-au��Vd���ı�|9�!����ɥ��&e���� �/�-̵�C�����΀� �dPY�mH@�R�;_X�=��)�V �	��s�+o19���� Z����.�k4��(Y.�A��5���,�\(@I��k�������a��&�w��;��b"���\�x=����v(@�O=��h����1~`v53��1�b�`���@U�|�h��`E�����8ا/NtK�Zy�T���&=e��7~F��9���uI[|L�Qe���v^*?��R޲�射}ؽ�3bus&k,p_{QD,0��j7��e����x�7�a���Z$)!XB�/�ȳu�5&ba������x.�r'���y��*��!�0 ���>�O�܁�w�=����u��AT��-EF�k�Z8Q$�8���i6�9��ݲ$��X ���%�hA��7_��G�pQ��U��/Z����0��9�5�U=�   ��Fe剑@����}��һ������}G�1ԝsus�%�����O�e"�18�KҐ���1� SNm�Z}ws����$�C�^��x[ �qE�@.j��~�#4>K�l�ۆx� j:F\�S �''�%ʐ�q���K����ͮ���z��� ]�Ͽl+s"(Z1������J���'-ȥ ��	�Rm�Q�~�;Mt�.2�\��7?;�bPa��M�΍�y.p�L q3M�'�{7����y�_�jȰ'��+X���V��{����N�L��.�/)Wؔ��2����B���������}�}��޳[1�n��~v*A`C/Ċ����b?E�O4Z9*��⶚?��o��m(�6�w���� p{��N�2'a������:��e�-ߣq(|mmG�Dhh붴�*oy�K���͚J�S����P�?SC{Fhy[HI@"qS3��'��%�S���[��A�o5e\�n,{�aQ�_eL��7�i^���i\�k��HKK�0?���{�����ǭ�e1:�k�A2q��$W��&�[A���Ů���N�s�0�����`�2C�gQ�'9#+L��C^��W#g���-J�~s=D}#8O!����	�M�U��0�VR��a�f}��o��u~�����h[3��m��:횾T���)G�<@�P��Α�(��Dٟ3�\�9{��n��iw3�:�R�z%u�ܗV>��n7-����Q��72|�KKO[�9�!N�� �!�7�$/s}r��[/�A�|z[O��d�3���6�L�r�:G���Elj���H<�,�W?��m�.�� c¾������m�w�Q�(%+�K��-\��N����?۪��Շa_�&�>��o�wA�6��Tx�\��n�O�а������ѧT� �顆���E+����0#�g���,q]�p�H����R���?����`:؟^���k�҆Ū�EK|��X����=�=��x��Ϊ�i�Վ��P?O��L!ew����r�zlT�`�S���47���m�ɧ$����F��hok�B���T�=1<yQh��&�%��9�	�y�LP�j�M�_aM����6�$�[h�A=_�Оc�]N0�O��U���	hp)���ư	5�����K�����y�C�f�^m?��4�Ē�������LSQ��8�(�D�ފ��t�M�DAk e�s�-<m�t��i�p	b���4�r��C#	(�o׌�<8KÆ�ک�	B=�*��f��ͣ|n�|�R��F���;�T`���r�go�N��ح��(4��(��`~��@���c�����K.e�~�rD�8΅ڿ�)��<�(���k�}<
� (r���1Df�Wy�f�A�. ���\�ڷa��
�^L�ѬF�IS����,��yg��?�~���K��EĲU�q�d�Zm*%^�E6!�b�q'[n?I�q	'b�&�1��p�����"��p*�u���E���?!F=i8��eW�#
۫eb��9b��?1Llֺ��i||�=f���}{���]?���fU�5�Gw��LԠJ��:�2��/BP��;�k6�7P������.����4�� w?�5p�o�z�?���C��an�6�f0��˨�ұw��V����+mdʏ/C�K\��9)��}�r_��qkE:أv!$���ɸmNF��04`�R<'���4�/m��=B�-�0z�?k @��pX�"ص�6�-c[Gw�lLc- ��$�f}9���e�ێ<ILF�Uy5�P�CJC�����HP��.�G9KI@���t�S@<��Q�Л�����8��)2ʶ"!���ŅwWb�a�`}0)h�^�Ph7jZ[�˚Vk���B��J��������d �����Xf�P'ѮPZ	�W���.�>�Vb���@��`���f
k���z��N�Ĳ܋�F�O'`E��.?�K�C	Fױ�;�X��O�@7�\�ӔP�I�#�������z�ֳY�|����@Z�;��/׀�b�r5c�Ƶ��t�j))b������@���q$Ks8b�`ҿO�뮟��%J�
���僇ȉrdh$���ZG�K�������h'Ֆ�3�9v������$�"��f՞�ci�H^sD�!e��1�� ���3��k_�J�f��W������W��1Nr�â���z�Hm�t�ǵp̲[\�5D^߉�2�/4�ʋ�����Nf�&�G��Ӟ�H["��:=�]0��ޘTu�O�f+\r׻ʢ3?W}�M#���eX��0�ׅ�E'~ M
􋝬<*����9�)��sN�kӁW��ݚ+��e��\I�E��0���7(��p���<®�	��OY*��C�^��_*�I&K�o��wy'�In�W8?cq��[�Xcj[��ӛ\0`�6�,R^� zb	�W�����ZX���u�g��//@�����|:/�zBJ�$���o՟י$�xǤ�s>���pȖ!�h���%�o��f�j��RMg�7�岏i�4B�Qf�(��&���@�h�qޜ�D��-�����ChƘ�E�[��0��yKQ�MN�IfIn�VǙ*�4S���	�llHgy/�	�]cHuy{4;�]�p�k_C�p:�]�4'h�<�Lx�"t�:Q,�w[U]� j����4�QRF̪7�������4?�;H<�:,﵁F�7f\ip���ո/d=�>A��^(�ԽGGڲ@I�s�`�Vv�bU$�S*-~,Pm�	��ݠ���&�V]U�[6�Tv��$�iL��5��M��_�y��hr�T[�A>~��Վ�sxߣ���bL�}�M�����|ܺ%������$�s	��c�Jl�<�;�=yp��T$&Qu�&�,��ل��p/�mJ�
;4�������u�z*����g� ��m�Y2=�~_�m�d�n������׊������(�1���q��MmpPi��?�j+i�t���$�į���6崽N��>9r�u�	t�Ǿ��Ϣ6-󍣇"����'�v�C���9X)�����-*)n=x�*)�Yc;�����>��9x��/�J_YMCoK�ػ!�hl$�ѽ����u���-=�	�ĳ�@:�̻(V�[�R�sr��98_^��pg:[�QHY~�=n�(u{��m	�(�^щ�.�M�J{.�׃�����$�<�v���{y�(���Ѡ.������b�[�t�i�����;H �A�E�e��ˍ]U9e �I�|�A���Cw���}(��ʭ�!��.�H�r!�4���,�H���@�9RNm��Qz�C�p��gʫ8;��ᐉ��V^^�Τ>W/���J�.qzϩ�m�N>�t�����jܠ�@7�HR��*���/�Y��?�P���-З6�5�~�=#R#�q���s�1�׍8e90.UhgP���.�.��W�Y�»-͹�� �-�D��z�Q,JY]�@)d�N$�&�E&�鬇5oS�7[�=�95��ٖwF�eWͿ�/>�Z�I)��[��!4U�A���"�H2����!���ӯ��G��0%K���Q�h�<�_�I�������If�m�������]�WL6% 7s�A���I*�Q�Z\����;,�8j0�Ó��u�)�gG$��Jz�a��.�p��>�P�T��H =�$��)B�	QQ�FF�n|�5J.@�������S�M]��qqp�pҵ�1��)r'��1��W�qb��M^�W��1@�9�N�Zom$����/��������]i.�Wz� kǲr��%ؚ��q7�%uL�<ݡ�6�5�V$������)8rs��c(�I�s�.��[��o���;M�h�}��(3�W���<?�0��ܶ�A|&�R�h��d�KE��Y^��D��v��T��n�KߠWXj���DF,]��+��R_*��o'HQ��J����Z�5��Q	�=>����ǹ�Һ���qH��sJ��HIp�c��c�@��<÷z��-��ە]uҽ[����t�\����������g�C��6Jl��G�D�ۏ/�/���6#��;\����9-�Y��\�R*'��l<�uNf�IBو9��̃S�PP��?�.:�=o��cTL���Y���S��FnS!u�C%|����e#�c�D�ت�~ik! �l��������x��ZZŶ_�{q�gK��n\t�&K
%�\Ӹ�Cԕ�I���]N��#����x'ʖb��=Lx���t�4�XD.>w�����
����]�Z�fO�j�js������rm4��%v���~}4Sxx�o�~��B���s�z��{a0�%FB-�S��Z�|`Sp��?��s���:��Q�m�˃K�y�ph������:sGIk@�2�X-@VH.���8��7�Y�b�Ҧ�#NTM�ʲ��^Hǈ7ـrO���"� n��xk�wx��o�ԥ����5w�n�67P�Y��a� F4��h���q|6��#�"Z����Խ
�{2W�i݄��8$zhd'wt�]�E�ޱ��5G�N*a@1H���"�@��Ϋ���5;Xs'�.��H%(��_CN�pk��Ai/R����������5T�]UlU�P;�ܫ�U�ᐐ����S$Y�;��}��Vh�����g�9ޠ'7$��O'�Kju�������A�3��AC҈�A��DGz*w6�XzY��+�k_kW����m�5���ò0��0��T�&�$:K�:�?O���&��\a�����r.9(:3�+��2�N��Z�<m r�C������,z����PRz�-��섊R�)Kg�:À"3ZQ�^��L�"vv~i��8�T㭫���o~?���������|<�Z���U����" b�9i�p6`?��YN��iT�9!�r���|;�*�����M�k	M�r��)���<T����n��f)�l���#�jrS��F[-��-A~/�ɶ4�uJ�3uF��F;��1.֌�i��n�T�K��
�o$�d5JD�]�+.q�o�9@��/�x��`�͓���1A��^�Q�(�e�j�6d���_��Wf����`0·���{!���������iWkի E��cA�΋�'��1��Ot *��?�1��S�Q�Qc�XA�^95�̂��k:	�-?�8�q�j�>C<>H��E!r�
���}��>\Iڰ\^$ �݂��[��t�T�!M�׃Q�t|�+&���S��1��.9L�J6w�����.�%ai
��.�*�9�Z���Q�;]@��e�q<����xr��2Mo���hG����D����܌9�e�J�A/�[C��'ʍTB?�RTxvn�r�ef��T��qc�~?W̻��%���?�]I�m��:^\7�U_T�-Q�O�[ypҸ��TE�+
S��R߯�["��+�On���S4�}�������6>Z��
G�fU�e�,/��6)�$�?R�Ff��x:�q��͊�;�UE���j~����̋o���au8��l��Ҽ�~��2�J���>�Jj�a�S�h��G��u�(BTL�]hS�:𮛂��\�� @��d(��80�ŷ���chs)�&�W�x�뵽�ż���D�n�I���Yea��5�U��yjS=����b1cU/g��R��ҳ�nIn�O�3d���i�s;�M����iZ0�7�&�04�;���Q��:_��=,|��𗧟�k�Hn�oZw �jL˼����:Q+�MI��$-ײ*M^�څ�C���C��Xs#�3� Rڊj�5i{�p<<�E��jZ��f��-��1S�Xf�M�*v"u���BTb=WϤ��Tp� ���N�&�)�VIE4�$��n��[?�������d�UYu����˼k2���Kt����]���&��+���=p���\�.:6�Pv���Lְ�����2Ľt͐�')�*6�i��@�I��������g4��=��e�K��,�b�(,��-�X?�<^4����D�p��^v+]�H�;�]���ĥGϊ,R���1�`o/8y�+L��S���	e�*����[�e�E>T�&+������7U,8t�Jw�xndˈ=�\�o�pU���6;��O�3V�dh@֘��$Z=��r��ؽ��C������G�k^U(П��]��3���o�Zk�K�q;Q�,%^�Q���&�L)OT�vپ��;�T�����=+_b�EC��վCu w�������D�S�ƻ\�,���jvLנDю�8pӖ�O���/���ٵ�5���8��!N�Sn&��~�>�3���P�}"���O��e�����	`+��$R/Ϗ��k&{o���dp��o=K�7���LR��D�[<t��:@��$(�]�r�'+�P.��	a�Oʗ3Ȟ\n����"���M��{�áCJZ���*P������!H��5��3.`Q�n������Qp12|����G��C+AP91��O�p�(ϭ	62���˘�B��H}E��"	C��*+n`�X������5m�	��z������E]�T*k���6�����b���o�W�J�ޘ&L@	
�{��<楎u�w¾e꛼	y�6�D�M �]�,�2�ʵ0IS�L�Oo��K!�[*��\��6���'\P�:����p^h��|qD�!b|3���R�\  �y�r�S�B���l�'����G� ����j;���~�a��-�i�2���Z���#�{�AA����e/��y��a�z������=��EIS-������z�o�s��Y�j��N�R0���e�D˴z����k�{+~	��>�A�7\�0�L� �^O��T�@����_� o7����"��N��n��o�,�d���uV�i|�1-�w/u�En����_#��%v}<q�HH\�����s��nh�V�����8��H�[�g?v�	�2����.���3��]�D䱪U*�2�
U�����C����g�g�qu��el���M��`�����̯��2�
[�1����Sp,��,���<Bn�� ,꠺�W��܆�c{���j�?a���=� ����$"^*�4i���>R	�S�iϊ��j��2�Pc��"~�;�0�El��r��4S�����t�c*����8w�63�
��c�G=jq�z�|����f�+uj���}�B?���M@�9���;)iǆ̲��y�����Q:,-���WF oo�۳�UИ�k�1�Æ�_P��g���,,�=�$~�a���D�ҙٲ�pݢ����~���_d��e��"m�;^���U���&��T� ÅSj���
��!oYZ7M�ñ���"�0dq����	8T��'���o�8��z��_n���<S�+�<��� I���E$HY���䐎�)�S�E�����ަ��ο���A�Tɷ��C�b,<ߊn��3<b:��̻<�^)&!���=������\� zm����i��lN��zF�mW&h���3y@;΍�K�觲�� R!XV`u���	`�����c��@�s҃�}
�������7 ���n|hv�[�'5��m�F>�LR�I��E_g��/�Z�@�����9��=YG���g��kX�uJ�̭^�dM� �85�5��֗1�^,⇩|g�#`�o����&�t����x�WA���$>jnl���FaxӈA���K��L:;g)}��^�82�;�0�J��4\���g���j��O�4�o��k'���^�!N!	��t ���Fp��$[݉Hso�^�����u1#��Q��ni�Y>Z���	��l���"�*ޞ ��Zx����?��.�Ci��������f
���&ŖV[�<��'�K��D��&Đ�Az�V�6�����T�M����#��|?|�������[���S��c�,�̈́��r��@�����(��j1[H!5��U�V!��{�-�Zfw�����4R�E�Jol �4.;��;6��%h��������8r�huI`xx��0x�,�|�xy�<��PL��:�/U2��Uݧ2&"�y-�G���쪎��m7�o���X ���������R��8<�Zb�(��A���}��������.
E���Z6��uM2�n�\%�ʬ�����9ƱP�8�B�&�>Sw�y�	l����f5z��u�>X� ��(nw5�[�����x�`4rG|ƃ���/E�a��]^�W�,�s�g��$k@bPٻ#�e���'���X���u��"i��H=��Af)T������f'��y`
M��5C]B�����51-�ʈH���">9���k�V�f�ZVW	�_X�����JU�t��q�j�5[g���Ý[���w{��zjf=�2����e����������0O�֑ќ�N��yc~+o�ݭ�qN�SyHl�J�1���K���*��7Zr®_=�L��b�J�T#��ܛ���*j��OP�v�́`uI��G�k���aUe=#Z�àp��Z��mT�~"�SQ2������I�|�4骬]G����i��L���B��L�c�s��6�6<��̫eܖ��++����6�ŚЛ��(s�bu��)(�e:JBSd���}3Rm�0b�/����4nZԍD���̴�<���0\lE�:�,�J������I�<�u��M�~��d���d?T�7�W�8���*=һ��ح,��`�S@4S�F�' 	��)��ԼK*�L�%k��dI�0�S����I��c,�x[^]_�����>P��N\�F��(@%՞�6�xD��Krkj[�e�$��-I[�;��`�&�9`4��K�"е$��'��N������(���?v�$uvX����bbJ����BY���vi��J*��4T\��x���9�@�Z.�Ю������9�-���oM��*�g}���h��3M�ƗN��!K��P���4�	���LƝl-��!g�X��Փ�"j#I�8��_�"\\m%� ޿P��S6G{k��A�n�[lk+�1|���笐o�][��1��i{�:�� ���o�)|��S�ol�׆=�~�G���j�ã����8�+W2&��e����0>g � ߻LX;��|���
 ��9�gvA�Н��uȓ���>��r�7�WS�FTה�	}�����zfR�4"n_{ꖓި�Ұ��d*�?(��L+��P0-�
A[>$锓G����Y���09n�?f�W��g�m����BѸ\�Ŏ�v�p���GQw�94���Y����}�PAC�=)���Ҵ}��T����w�v��km�'h�*��z��m����ۄ�&@@�$�xk�a�O�"�!��rM�H:����t{dxL>��˕g�$
0��.x�ݔ���b�@R���f�D��HD:�����?A ���������V���CD�Hs��߀��	V�b����%�������¢pP�^�>�t�

�:�/^5�1_u���	!��t�N�>���Њr�j�?�_�Z�%U�:Z0
E�H��;
 (�V�x���b.�X޵̕�����v��{$��o�i� "Q����`5��'���ʒ&kyB����Z���T����'Z���o9j�/y\,I)��Ӱl�~�|��mU��2�B0�_�()fP�(L)�4�>��>��&�Ť��=��j�7�b�9#(t�:j壌 M0_h>sH�r�7�P'�gCy{��Q��L�>(6���<�e�=VR�l�(��U�x��0C��1p�#F��r�����]]G��[ w�,�00��S�Ty��9ha���1L�3!��^Y��p����~�/���73�>c��7�Op��oB��f}fr��E4���oʊ�//$<�i�_آ�j��/ڦ蓲s<.`Iu�k�D��_��B���Y. �|S+u}�:�C,�i����?45�m|���#Lz8���o1>_Z��"����o'�_�XIo��Wr�8Xs�%.$C��z����Rm���^�4s3Y�;j>C2 (�)��짅�@���>���iZ�O�t�����8ޕt����D�-�0���o$�E�bg��M9]YӼ��-�E�>uwE^�����3/��T���v�gbw尝{�t���(m�dR7T�॔{��<��=֥�.7�l/C�� -�_�cN�3��{��ϩTٯ d���5�0��0f���z��yyr_�[��������#���\����xߋ��Z�;���˧EX�����_�<�.,�X>��A�Ns�,*�d;~�t���"�g��La�-a��"����#��T`AZޭg�� ��u��縲��푷G�Ӭh�i�� �Z"���F�x��{��rh,�8~� 9u�1�t��@%|�D�
��w)�\�O�!8�N���Ԉ�X+������E�e?P� �w}�򫐝!����S�6=)���Q�N���{ݚ|%�_���Z����'�d9��
��	��@&/�Onyb��0���Q���rp������],� ��֥����[� .Gy�k��]��:�`�ؾ�����Ըר�lO�j����P���%濊���#�����ML!B�1Cr��M�+����4�Vf?J��L���`!��kzV_���>]���d���6O�.��С%�hF��D۫�V$Ke%��F��N�VJ���d�0�]�eVa7T��§��=�bZ{}!OG�_*��M-,��D��(�&�?���yNI�������a��o�}@��h��#�װ6�p�ә��G"��m�GÍlF�� ��c̶৭FZ���X�_2��=��Y�p�>�p�ʵT��s騘s�Ts�^sOWh5r,��*��Ƀ�韓�$� �#�DȔ��F4����b���\?�-tR�W�Y�ԓ^�;�'�K��c��]|.�bςϛ��{��r�a-� 74����SIk&2�EmY�vXUc�_�=B����Seu+�%h�gE
�&ݜ���^�P���\���
��S.�x��-�O��?�H����Wv�S�p1l X�1��>$��=�aQ���I=����ϋ5��Q�����V�|;-Y����5�Z��}GŴ�q�{Va��U�*�����Q�A���D�IX���|�Q(͸�r��26k�uaaFo���󳀍�?N������ꤺ�m��l�N��c��$|�W!��c���;O�8a�%���p�GKd�E�`��Ӳ�:�#��~�^i8�CVoi��E���D&��7x�j�Ρg�� ���\I[>��Ǒ=	Vð�/����a~7��pƔ��49�^�u��>̰#8��&޷��>"���	vz�1�.yOSb��zb�\=�֭a�x�w���璋�(����ɠ�L�_��21�k]w�jT��'_��s�)��2��ٽxکե���	)�l�j��;������#I�V��
�	R-���W�@"�����{(~C�,?5����E�a����X��a>h2�EG����)�)S�#��M�Z�Ak1<�}���!�N �A��j��)�b&!��j����=�r����Lw�\s�,d�X4x���bFQ8G�xW��6VH�$�tJ#]3��	��)t:��ϭٗ-�qyǣ�.�idN͌�v��Hl\i� 
r#���i�<m��J��SJ�b���\/�n��D��-+uW�v=�Ԭ��mƉ���+%�Fa֤��V���g\.���v2���9@�P�!�Y��#�"�O[���ޛK%	�}l��|v�[{��p�H���Q�m��O�Q8��f������_�J-�G���*1a��\"�2�쬁3�'��^O���@:�y@�#����w�:Jp>��Z-����`���6�߫e8`Z@�pن��f	Jx.���O��0D�J`�D��̧� ��x.
9�����l�m�z{��,��)/���%X�K���ߢ&=Ʈ��M�zH�3��L �jrE?��,�S�t�&B� �|E�L*و���R���8J�d�K}�V��g`U���l���s�_�:9hڵQ��V�'�m�_Ӄi*�����l�v�(��8�;�Bm�ӗ����LFB�?������ʭw�5]�2�ཹq����������2��D0���i��㬎���1k�8t���Q	?�b�>�Ln�:��"�#�|U�����J�8��7d5V������8tuR/*&�&)m>��}�]����CN���4�٤���sİ=�b���e�l��Y��\O`��wc�Zr1�7��{����樂�"�$�8���s8�\~���@��׽�+8�J����全Wk��ur@]i�b�"���U��>$�~E&E�Է�����Jт� ���M������q'��F���Kw���o�$��o83��8��:f/��_�Q�wvP-,���9��j�Xi4�7p��#gj$�nb\oD�����o�ɪ6E�aҁ�Lc���`�-�0�p�qx���(n���X��~�L���blG՝�����6֡�!� ٘�(3��Za#���6��h�7��~j��	$A�*U�ӤG��b�
]�Om5]Y=E�D�m�������G��Q�߹��p߅s���3Y�7�xR��pT���-ޘk)�q�$G���^��X�u�Wd��)��*..4�Ay-ü2�>i�����3H��s0�.��u��(p���@�~c�:C�*9uF�?��Ħ���>��B$v��5\5�?Mб�3wWkJ�����
�8�OB�&��W0��m�>,9�X.�B�]�[�K�������!���Wi� ��l�80Pn��nt&WDk�|I?)�.fS��y��ώH���Ë:�ŞC��v�؊;;D����;�0C��3nzt�e�b������&OQ�O��⣗4�o:�P���� �
����R.3=\�>{����Ԏ������=2a9�����@]ֵL	
<�_���I����[���{f� 
X�� =�el�6��hX&�(�' �ѭ޻:4L��Y��yY�'F�k9�d [��lO�f!ђ�)��	�BG��γ���Z[Ը�Kp�L0�3��bԚ��0��(�|VX�3�m���{�ļ-�or�a2-���C}�\<��A��+�a�ӪϝN��)�Y��IӠ�W�����6x�q�2y�� wq�̈�H"<����<ε'ѥ*������.�@m�&" �|o�M܃:�^|Pˊ3A�q�q�3�h-Y<Xb:�~%�9�.�JyM��?N��2��j:���I�7{�m�4G{<z5I�D	ɰ~T�O��Qٓ��ˤ3��.qi�S0��m����,�ͥ3A|ָ����;�����Y4W�i�3�r���M����9�۲`C�?viK��RXU���A	�8��6�����^��&^��.�H^H�l&���)�m i�w= ��窉�b���Y�n3���mlU!�`na��t�y��8D���7� ��'�^LM��"�4��HU��WL(,]��Ĥ�3b�堔|��E䎬Y�����t5M`}�0��i9�앢�g�o"/��#�^���Ɋ���0<�W��=(|0��_Ħ�������v�k+���˯��p���xg�c.�v�G���4�MnN�'�������=v���>��w���ݼM����0��|3��Zb�e���W<��j�K+�Xh��i�Ffu:`Tjl���c@�F�PB �p�[CN2�fa���[�E���BY�q8��O����uq��e�������[}i�r%�!����60��@��-  ^���*9U?S�P3S�����V�ω��N&�r�K(T��Wt>����w��9��q��n6���ȡ[IV���|�W�n"^�`슛@u5�MơpQXs��B��KM�x��[���[m8�g��?]�)[cxYE�[fw좩Yu5��E(��3�
� |8A��dR���Ѯ 8�b՗n�~����!!K�PIā�̬�Ȍ`��Yg1RQ���0�c����p������أ�a5xcb�����Y�҃�}&�Ĺ�t�l!)$U�D�2"�8��I���}���L�<��O�;����5B�v��jHk8�R�C�����))"D��+W��z%$�W��kq�H��>'r��1�4�A[nTY���=GYV���H~������	캒�5���c�r�MJ�<,�)���K�jY\'򸴃T�FH)���v����:.B3/��`�;���5o{ǅu@k��}_K�$��:�İ�����,��ɟ�W����~@��>�7zK捍J�C�!���kP�~�p`I�lvAc�C/�cb�^���yU���U���\p��?
�ĨU>م����fƋ�!�ï���~�d�?�@)�ޱ��֞�¶�.�șr�r�g��v�ix�Sޜ{�L�
S�O/�����i�o�V4����8��N� ꈛtp���D&9I��.�uG@;�n ;��.x匧3î0���(�#�8�����n��f���9��<�$��r�$C��_�A�چ ��t7�N�P�.���3R� �a)�.�䕀T�%�.�,�|�}.D�=�M��Fە���lr�I�uT(��a4�s5G���1�t�U�k�44��%[F� J7���!��4Ʌ��2v�s�$A	�Y����a㉻[=�y���S��1������Y�~wq\��{x�a�~�.��m��ȋ��cc�ۋN˕l�I��ޏ��x��L�P��T�_�1���������ޣ�c���`=�˨vc0a�Zci�`�	�6�N\�RTV�✣��)������	�aj�<0/�
a�%�o�qh,��9>O�G�P �ߌ?���QO#c�!Q���C9B'�AL�����gSmVCB��2VW��s��Ԛ�)��3"^!C�h?�?Y���U���V�o����z��فtG	N#�6���:	N zJ�ķ�MNJҝb���\O����h:�+�6l�rn��KcT{�1A*�@�����;�7ٯ,c�磒�vzN3s 
2�4?�9 �GL�@�t�ѵ�#M�aI�9���ʈr�f8����O�"4��Q~���s!�T>��T���lvnr.�Vl7,
M[��@�k�V�Mxg" �	�����ᔠ;��M-��mq�
��>�B�7�!�Ɏ�O�M�6kl_���N�b V�ă ��=O�䢴/2!�����u)9�K��8g6mH��O#��]}�����*F�m�b��t�8��O�����Hu�17=CZ����5���2��'�t��_�S@�Gk�X��-�ȷ{�ơF"����Iw���;�bO���ve��YDp�+6Q��.��>����C������VN�:�1edV�㑺�'Aq�r^ۉ� �.���{��"�@lÐ��YI�@ڬ�}��c��õYR'�ӥ��Hk���5�K���sR(���W͝.Ń�sޕ̈́�+=��]�@^���l��ϒ'�2+�M����{����W�HJ�ץ�!^_�34�-jL�hFuš@Jp���ʝF4x7�g[�H��<��/0��>4�Y x�|�N�ׂ�!F9�v3���r����gI͍�b��P����9��I���5�2��r�O�i}T�� 2E�7����N�im��#��c��1�X�P�WX���_�	��:��l�z���h��/I��G���{#�́�����b�4��Y@��#�8BE�b��U�4��y����l��w�{Y���G�� {���M�+z*�-ClCm-a�DB�e�5,t��ixwj�dȞ��i�SI<�7�����-[��FhTi��K1�jn��/�!�&j��ݼ��5q��1r��B�*CM ^T)"��6>�կ����L�$rގ14�=f�|Ʊ}��1>[�l�������\z��b�̆��ixx��-�%��E]�s����+9m��//���xA:�K�� �0h'��3���$��/�z�@_O"N��������_�a�h���D8P��}�)#��q�[�1%3�a�!�vU�v��=6��d'�ZH6 j��?�/^F���:X7���<�c�3j�I�Z�^{+V-�
FU��+М����R���6C���F��bwE�?��hJ�zk�bU�%5�U��o��.�¦"�/��A����63��\��C�BT?�gy���"E��#�Z�#y� ���{=�U��)�<ͨ����X���Z�^�Gp%�����J��	kW�iL<뼿��UIن�zayv�7ˁjTTͮ����&;)�a{1�=�Ǹ� 9�o�x;.�\����<�,ϒ��#&-��/!�5ƌZT�m�k	�-)U�gTm��n�Q��Y ��y��?%$�@0#؈�m2՞���"�7ȫ�j�c�Ax�(�~;���+D�k�Lmw�"E?�O���8�l���Ūh��b�ҤKh��$]��R�C�҂���ێ��n��霮X��r�U��mw5���OE��nG��2M�9j	�:��vn�)_2Ǳ��I?�a�M�'B;�,�;���Gy�E�+S�h��psT{�P�,����>BL�Һ�.�he?�������d���eM�G��2HVF�J]8#�)
WdAQ_]��b4�'t�� �0�ژ�q���dF��G�L�g�[i�iZ�W��E�0�j{ ��
[��sֳK�����)�����w�EQ�2��Wݲ>�%\\/)�N���d?�#`�+[�Q]{�z��j5U�olYl��o�FWXo�Th�[vŀ��IA�8i �4�b����X�&��CA��Yq:�?���U�9}�N/�g[���@�g� y_��R��^��Q�8�
��XDL��b�?P��ܢD�r�ǿ`Ld�E������T��gF%�^�f�sc���d���	W�V�7WD��g|��z�}4KH&x*c=��+Q��/���z��їHj�~0z7m �#X����C������Ä�Yɲ+�j4C?������)�|4Me<�=T������x�L��6 pb�f\�C:DU��~�e�!>;�Rt�w�|&���PwN�������%XŦ��\�h�����)[mm;�p�F
e	a��gm�H��?�0���`<�R@���X$�Z�,@��H�APek$e�!�v�AN�J:1T�5�����?o'�7ݝ���ˎi���4�����}2�33=mR�e���J�\*oȏL8	��=�1í��t���-q P�_݈$�m��d^�)A�>u�,� ��D���s�q"";�5�EQ�e'����ʒp��y�m3��J�~��$��^�������Vl�;�R������X�x�'<7�H���ځ�*�)��nTY�ald�8�Z���i��/��^�/�uZ<�1<�d?�)c�dΡS^T�u����N5���i�8�Jt��� ����6+O�|F�+���]U];��u��=-'�͔�&�#�u�f�U�5��'[��wY=b�8�{c�y�5p�A�]A�1�ɴm7$x����M#�w�M�m��V�@���29`��Pb~N�y�3vҞvK9� 벓l|�o�-q�9FN��0t�q�JA�QWK�(�l�GA�>8�yk�e��y-�X��_@��O���������Q@(֎��b��V�F�:��_�n�"ϗ�I�C��@B����6�b�<��\�]P����M��[[���㵠�dq��N��'�[���#����%}����}ϳ)0��:�G9[v���*� 5�	�=�,yI�X���_j3���O=�Z�����l����K�������d��e�[q�X��ou��B*�P�Ϟ?��x���`BH=�Yv�L:���8mwp%Ũ퉒F�f�m���
���Jx

�&R>�n��kk�W�7:�u@)�WG�m�4h�����$uf[?�9�&5�]���Scc���@p�=Ts�H��Iecr4`I��W�ː���������}vp�vg�M��g�Ԩ�[:{4J���-Xz�2pi�:��;e��
�^�Pk�p)�_�K�sc�F�ڤ�t={�Vl�^_�Ђ�ѣ-|��]��*3?�� L��h߹t}C�ҙO����֑(:��:<��P���_0TWG��Q��_R�i-D�/ �,�A{	�ud	,N�b���ޕK�lxH޳V�巙��s�{xT��>�r@x�r���;Q�0�ʏ�pY�R��HʭĴGLo����O{���_�:����ܙ>�s\Y�����d���*=����z����cG��Vk:P��LBh$�7�D���c�ࣚ�뀁��6��PQ�F�L�:��;��F�OD�m]������G��w��a���_�y�*
�E���bO@����k�( �\��DS3�d�]z豺�?ӿ�8��s��.d�KY��g�h�'� ���گ�u�%$�Y��9ux�22WMZW�OvL�ĕ[�?4 MWk���uhn��A��Q�� �	i.]�	�礰��o+SǯG�P߲�S����
*�]���B���(-�)1SSb�,�_Ѯ��[�k�ȶQi����<��R~��(��}�f��|����������[H������˂(A��=���|g�7���̨}��?�&-�6� ����_*�a� �\�[x6��ޕ9M���
�4��2�'�H\�#�K���W��f���-���.���zϵ��{�����1=z�:
� �J�1�r��B���C�X�z-̼q����O�g3�]�H}�Qs�V�ɓ�����1&�T���e`��?G���L|Ӣ��$�Er4�r��+���9�|�1�@A~:�����"O���aoOA�-)��m�Ao�=w�zR����/O	�\ Nu�[V�[��G(L넘���7���d����^���&j�����2�������x����&1���S��O�pFw,�%K��5�Dsn8�#��)[�ҝ�eH�;dH�Y�l�<�I��&GxT����}�ι�-�qA1e��Q�Na^�k�H��1��9_hM����`���n�̓�]G�����k�n1lƜ�+����M@���/WTh�3G���#G_.Ш����q-�M�8�����C�0����fA�T��/���ϲ���O��ik�B�w8!�����oI8��c�3[jP����K����b����R���g%���%��YO��P�����j�jQ�~�U�*�j�ƿ��}7��.��_�?��u�a�a}N�F��lLѝ.P���|�'�ȜΠQ��S�PșA"�a���0&�B~�gW��X��8b�u�f�xS�TCy&��6���+mZ�0f˯��p���i���������^��<�M<{�0�V,�M���&���b9���C+���D��,���[}綵¸+��]�3�ډ�B���zɽ���[��t6*�k��e�ЙV⼌�[%���rF}��
�i�
^!}
��ETp��X-�-�������W:�,�6m��������k�����Ǻ�sI)���O@tW�{I��Rl`c�yq��m���
�U@�IʈH2��J�A���1���@���Tz��"��j���;BQ���7Pu�� ʽ�L���԰ ��1��o�ECI:���9�mL�9ȵ�\��%9|�΅��W���l�4%;�I�C��AP4ã�/���W���6�A��YYTqm0Tƃ�];��w����)V���e+��>��sb]^Z��Op=� ;�:qRp�S���t��C�t�#���[n��4�8�{���N��ɤ�����Q=�+���&���Q�������(`��ȏ)�B�Y��4��O����P?���)
ّ�5rx�.���AvB[���P�����$Gtt���N_/n�@H?�৷��g��C��BQ�ax6h�T#�K���>p�Q�z[u"��&�!���?At�)�vذ����B\���əJդɳb�}��ʅ��2#QC�04m����R �ڴ�c�w�U~r1���*�����Yaɛ�C��'.X�6ҍ����.;�J..#u'��Ϳ,,Xn������x}�,��s�=s\��{B �rvB?,����lJ�� ����.��
x83��l�Q�c,3B���-�ʨS���';@%�Ֆ���3���λ�o��Y�jA��=T���:���تjʍ��Ӡ�$W��<�+�)Y�,#�}8U�	����*�M:�E���t���MQ�$ؘdΜ&�ե[�A�/���a��)08B߿:eSmR�i!x�.^��*��/�Z�؊�f�ɘ�j�^�<@.�IZ4�� �
`"a�Gg�g3���'�+�l�HtEꞡ�̷*Bפ3���dM�W�1�74y���S/Bo�*[�.Ғ�f8���f9~4?�4_d�_=M^�5B���uJ�h�?w���fw��Ѧ���>�P�S��I����ݑ46Z�9�u^��Q�0�!���r� GL�x�8�l~���o��^ �aǏb>�B���O�jx��Ô�ȶåX��>�ϗ-���S.�+Q���Ci���ަ/�t��(��>��'jٞ<{݆݈����)���7$'��ş��K�5>��CL�3����XC}���I>��W�$�b#{ $pD�aE:;y,�O��d=8����Я�`�-��z�e���zu��h(A�(�s �f�5�LW�$6q��}�/[����P�
���x������A��<�J��yS@���$�|��=���o�NK�m��6NT�8@��n��u�Er-A.^���z�Z�@-������J�h߷#r�m�����(��2���X|I� 6�*1!�^��ʹw1z!��q�w�$��4L�sq��b�F��?W��+b)��a�C���I�n�R^ʝ��/R@'�%@�&��CG�X���v=�~铢��� ��S��
�Ӻax�ϧß�u=Յ������l�ˋ�~���MP���*��K�(*�z}����ƕ�Y�;j_@��Wr\�֬��9`hʜⶄ���V��rnXB���t�Md�d�QI�:U��\s������P��"����e���I��y{o�wD��E�#�2�����gN���.�i�t.yi�� ��d�/T�Vn�@�PS��qЬ_)޽Z� �����Ԧ�F��1䅎U*���5:ɞT�Hv$��!	(,���Fx���WD��=���ui�$qM�\�c�sN"��h~E׹| M�v��jmg<ot֖�2+�1')Jl�*��I���T]�h���1dZ}*�ٟ��$1���(�!��z���1>��>�� H4m?[ݩ�vi��I������96i��}s#�ǏWD��)x�Ȍ����Q���h�a,[Us�]*2�c�.� �5�KCC�=Nw��MB����[�vߘ�X���������)�N�;J�E�:92}+N��?=ZN-I6��JrN�v��ƨ߱֍�P�0��c��G�p�G@q������^*V�A��O����_�D�s��a[�^�����_�E��[�x�:���fe�k�&ڮ�a�p~J'���j��(�t�
��T���g���a�I��{)�N������o�j�ҷ������'Ǽ�7���`�����y���` 'H�z�Ċ���Ǿ��r�A�Y�����f&��\4��Pּϳ$I��b�M��
ݡ�	�PʑIP�Q�-gM���=Z:�&���X/��f�FL��J�P>=������q1��;�U'
3�9�;E�Y��2��˯�F��Eǈ
;��)YZ��$ge�q���c����{���;��jn4��%�t�%&A' ���������1&r7��R�a.W�GV2ȊA�+R�� K���qr��v@�o	݄���W>r�c��9�V:�gfd�o5��˰"�})��ǭ`�ۮ�b�A�(z>�}��([2�^?�\-xhINY��~�O���GN��Nῲ�y*.����4r4>��tA)�8��Q1�~:�iix#+cn�&������ν��:���ؘ�{�3����M�y�Ӏ 7�j~�C���Q]`���B�%�%�T�P�ݙwքW���ծ�?j����:K��9Z�mFA
���+�,^x�~���#͂�cz/7U#r_y�{�Ձ������:0����pf���aҫAMJ����t�6yC=L���W ����9���5��E�;^��Ş4�|���mS�c}��I��%8�J�A�Ğ`���3GڤN�&�)��?��{������Mʗ~0�vM}�b���E؂u�B��� ��9�5���+O���A��3�J�.a�3��G��1�H"�)�<M2B��!�i0���dM��=y�$l��!2N37o��ᑘ�6+:'�-L�A_�\�5�T�14)��.�Ơ�'�H�F�QزO�&���&'��AP�����y7�B{�W9�����96��/�D��R��#�6?����-�z!�q���#�+H�y�Qf���쥊pj��M��~d��A<�w��+�0�.,����eUL�L�z[B�����$�{���!@��ܣ��@9�g9	�xI�d���0�L�0ZY�k