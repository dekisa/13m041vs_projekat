// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ywV5KnYdk9VEwTQYNOZ0nATHQn7pmgYuQJvwbpcK2AGxtyEFSkc5TYBdU7f4ZBqZ+dr1dXPzCh4t
eXWSybX5AnUYIMuJu+PkUJSmgpqsh/StwWZVSPlnBD+EeDQJEYORnujyYkihKsY+cwsB2M4Qr75D
tzdH1JgX+Jgk0DQVPiL4A4Qp9MPCPrMwK8pIU+gZ8w3aEU11aP3j5BioO61OXQ7BzoUcZ6vRThWE
q5G7TfDqtCRI6ISS7oVu+XRJdl8F6RRORmtoVLO9llWkbpc5v2B+ZDY6vRmoFXn3ofJM9Rt81+r0
ykdcUJTPK443ebusCHhNpnJyja6xgf29y/J8qA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 42448)
fMWlm80Vnn9Mq59V2vsaGcqttmk5dp0w/diS9B5gR65ZO2gOyohnlc9Q9bwq8MLPfj+9gbtI88cb
62RueMTnLEYfxNSLHsZ7J0DhOmqWRMHMs+af9pRcgFG5r3MWkoqpeLkoaEQdQ6VbXA2vYNGeYcPk
jXPWtEjtgKbluseXDtgACSLbAwZzyD84tPr8B1HiC0tf/rkGzL/SosI5c1MqnuwFXYyQ1yRoetmj
rjWkI1LqbCf08E+WyuruiUkoc2jffbBh8oxZpcFTtg1KQ7XYMdBc2W2cPXTzW8qwEE5H7WARisDE
aupL+v1Jx6cQESlTyYnAShJgKpV1df+NtWnphNFSGnK+JStzWg8+dnR0kK/CYmLZLkFb/BtMb91P
2gbIDH6jLQzbigRLMZqUc1AMSatYcgSz54+NfL550HLNbaQGFIaW0dhRCx7htmHwuIZjjhIt/Q8v
rMTcLRDf0Hhf1w1NjrjkOSEr7Kgii9gRa6OEW3caBOzrNb8SGSu4qhmGpPdjhJuhuobTGDhO2EaO
2buf+5YZ9HQ2K23vJAgxEb2XTlt4mlLhQsRiRn7UCgqDYGwKY4B9rXFTr1tA7LUaLhqpqQAzfjaR
21J9XjS+bYlzz8oNo2ZuxTy7gg2yfYivy4jep6wipMkHEgd8nNR55ddSRbyIzsLeHQJveKJr8Zv5
fp2t3DFiSjLfdyDrUHDmg78hkmHIsIC182qNn6Rjt4TzRdiEEkIJUSdbEL8ujGMWROY5g2e93ioj
7RKP/c99asv+vp57SnsjIQMASZHWuxeTcvAfFYCXBoWVkLI6IAwfsSN2AuQelJyOzWX1PplFzZ8R
yeE3pKadaaf8+FpgcTpKYSp+BqnPqtZyTUkr6+NK3CMT0A1attGTCtULYQurJxf6pTp7a9V8EPbJ
mBXPZSqQd9FZ2gbEk1kX3ND+qGr/L+3/qFzeG6KqEO5gvXiRZgHAtZwGPXxwlFVDZsB088WSE3w1
lQGsJmKZPI9hzLUVfsWp+6MDsmqi5/PBijdAlc0rMYT/NkAUtY95UBMi9jy5WQnFYIbqTprG8Pbt
vBE2egO/S09zC535Gy256sZQ0RubiRUDtZa0EUzOnBHk4yn9IPitjZ66JgttLUtoH4/NusHXb69r
QJBYJmWnF6YSg/6LtyAsMauSjrUIve7N3NBxu985vZUbdLPFUgth6u3YMonExuzvqolkKZ/YJw0y
V9h8H7GCrLPXdJ8r5upw/9sJvJEFJNsy9eLJXujLqur051Z+XdtYcqEeaPQCQojZJhw0Oaqx/NW7
0V6dfz5n3GOTytbqqa8LTdkypyb8qpUwNlUZ7mdnwH2f/L4b1/g8enYrMDc50qaUxVrnGMkwfN0Q
MN+y0GXNZoO54cx83Me3Bctryx77oDjlJFVXE5RAx/Vq6o6J1PfCqzI1p4KZ2+Ook6GPmfJLEY1v
pNZUigbqy5ovOWWhTLpbOb+97O7OtScN6pr8nvA1G/ph21iN6Tp534opJU5KXHSs6861sjebRDmE
ZtYIqQGAkfZONlRMVquUWU5gzX8P6u4E7h6Cd5PKyI7Hypvbm2A39BWeeT84duxyvzYOUMJkh7UB
1RDwtyWRCNZxmD8vkkqXYNzit3fq/K6NLNpGvlGLbh2IjZus7jomKv2wwKzX/cqeGq0SFsTtgaQ2
rLbcmLqw3P8XhoOXJzRAAaJuAgYA9XcqyafbfxnyVJXeTz2hzyPZPj2jY6/rQI7PoI7LojLGbXnx
cIqMHmNeHe/txhRAse3+//SyTMpWqo3LKupNkfgaj8Uvr5QC+P7lBSMu27hfj6EEnuscpfQRjz8r
cctWZLbJbVNXfJ5BiTeffOuVpj6DYFcEF61LBsXu7Ml83JB7Zjalz5YTGaEefMzQHWxrUNnxMIdS
2jOPj4wEqv/qa3gsI2UFS/Ov2gGMgTBUmgrkQHi/puiBperI5yYfcra6YgF3KBCCrjwZb5CWa68S
kOged1ZOPM5JIUc1KZS15q27I4y6E/OEQulB2XjRY2T+sxWosS9XF7v67STVsglxjgNC6nsX9QJu
YBTAp6h58oUKOmJPbafNEnlzIt0kog8w1LXXqdRN2+CwE8cOnIokAhy0iW/3meOYA27JW/bJyS3D
n1fVclF6qcJC2Vm91N92XhcOKGyNQEpO2J8hM0FJjEOFmPMJn/6RYw3FmaTx0CVtNmt+GoAH4eEa
f1z1AwIB6JuGyTNMfepl9kaCV/rjD5MWQtadxgVF8+vWBqden+i8nB4QUcMI5ujo2N9wXBD/+yoj
H+uqnGwzAsFA48iJFsfYmtOB6f5Tgva5+v2RyE8AEodohSc/VkosY1a93Xj8gl6KpB4z1RKdnVaJ
bdSACDyPDYKpwyNdduW17p4H7YYlB28SoVFO7C7AaeGm9vABY7dskNDkrowpw686IQpmlT1zudPU
xIf2ETzwbqX7ruj94lDPPZ3JOyWJoDrSvR6Wqvn+HERkrnlTpBMath/fvVUQ3ko818n3YckrO+b6
8iekkwucGT26yhVcmQJmFw9cTlHhYyH5/6Qp0QjKfAhs4Yt498g8B2s8haGrdZ5hVSqJg5FJ3tEX
Xk7KFNtzx0+ROKLfLtCxWYxIkJUbro7U3Ej2RsCLauOYj7Lz9fIEq5XBONsUlRYKyFbMcXvNcDlz
CkXfuUePhfghddL+0wzVhDdNYSOWdhwsNZXQqO2Kbw7pHywbCHtuwdyPStuYRWXL9XDwCvyU7jNI
caIsazXLNIt6hRwOJ0DOdv1E1rFAFq9fwJzQUzeZY7F94e13LtZnCP8OMdBCk4lTG/xbbXpCbBCf
+vQDohsKFpfzfX08bOlwG1bbWqDq+xH/8Iy69/gn7Il9UPy6mxl21XrNb6JlT6k2kiqma7kTIgaK
4Xs5XJkzxtPwhjB3XvZU04UgBg51ngVBxefYewlZ09aZVz9KdLNdRLT3SRZ54f4O9iFEA7RoBtDx
NHJFhws08aAYHKAXfM90GPkDondyCGzYbR1oKdi02CLE43DPDMaJBGzmsd5F8Zi3jjSJNQ4pA98G
EKf0lxYFkP7rUopuBxNj8zPwrjeW+0Y4Tsq3F9ezeVQsa1qSiJIe55beBcyimpIF7O8T//vF9sZp
65pQ4ZwbcM+VPscpm2SNAJJSyA5sivocOpkVcd1K8wp7jMaYBCEGeaVVVoWbPBTrz5BxHT6UH3ca
dieS1Z6H73nWVi/GpnXXPLA4Ew5bDCcQVuDO9h0sSpyYWRULuhanNvRIuZ4RWRu6YN/qjxL62fL6
zuNAmaw7hqLtcdhpn78gHKVKQ3DxDUSBVsyYGmRYt91Y3iF4FlV4Gqo7gceOrfbTIx9TN9kLB16M
41Dki/mATjkTNmXW5GAjgEzF4cYRm7bYNZm53goNsZeIlZommssxGwWTSRg/8Hh+V3FSlniJrFLj
dP9poxUh73zVDZCQNwRlXons8pxQ961SdRlzEXPyygYKN7xBO3Cc3nXTLK4SOcnnBH2PT1Tm2gE+
NDC1H9tYcX33LCfEbEeYONc7f+78frZUsUAc/ahkVjFABUCGOTGMEPgPawvDy8yo1haWXN4gCP7F
b+oLBx2PygN66pufZuN4W+/arwy/q/jlAZ3oAel4UGPf+qF6Qm6RWGlWx9G3X1A565+JWxL6lqFg
+Y3OASApCQ+OE4JfrCKGRspym3mpL9TEgTuFWMB2ND/KSyh15y3ZoeI+Py/h+1j0if1IJtPQL+Md
reXV9H3r/9SBH6y2w9UDgPDxnnlqSXTm0t3Ti/a4MHyrE9nu0e7nw0BokicKwGEVvZHi2aU1rn7z
3wULMqorSVxFtaZAGqzjmrfCEo8a9/nw6IXKLH3RaHgcvfE2E9LUSa7PRGaQWCbc/yihwcCXXlsI
CPutS5PZYy3QfVX9wwy6gVVuprcMYim4XwOAwjWAd/+7re0uRX0fc/jKaigz1Iv4n9AcpRq0Ml5j
124p3Iz3kmGAE3AYFr1JeiKFQXhoSkKvwayP2yb3inv/yQ7bv1JVBFPlKM3WCsH9j/TURCi9yEIl
siwuCiBo7g31pYVpxSfifoPkhtBEiKOvMumuA1HorW0Dffd8WtR4lhTOCUuvUq7uSYXW5TvQkwu7
r5P2HspD2gZ+LedgKyVRQCFBzY+yq+H8pQtNQf+ikIu5nXGlA6RgB2DNdLflYQ0996D6mXrUH2R0
S+08Nj/fyCe4r0Q1VHQzEvd4EbKg96LcxchyGIFhTq1p874UR2scHptjq3gIKUjEysJtjX9fwn4+
IT74xEVF62W7WR/aL4i750BhN6Q9rb4x3D/Wvs3PGFkrpFKIuF1i+L3+D647xog7bi0ig8OKi7dP
jCMmSUeXRYF5317TISFh/i33xik90rRdI0OYe+7g/sUm266Oyw4u5/bueZ3AWgHspEVQQ8kDED2+
ETEDwtXoea5CMJnuRxk8ss+GxaQugj6SPpu2w6eVY18cTbnxnOJB4ckacSmec0OauUJdYoHVSV4z
yUszqMdFyhQnkOUR1Svm4co26tNO94yAVFoPoTkfKb/vsONnGNV6WVSlqOxrv9G5aL1JQGF4Y0JX
nzJcuqdKzBkkrV2dINvpGd0OBuYH5nmAivz4uW9IKz3Yaopq01WLjISZ+3g/ViYojlh7wkUW+g9S
aXWbo9k8OeKHOMqtZIg4JxSm9LVVmxf/7tFD/bY2FICvrJAEJ1ucRHiGeutAWgPW4pVzy6b/ye5z
QvgLAq/UsQWV8qiQI+Tg93itIUsv3YfxkQf6jzOnNnNOoNgpM5xshlz57SnCI9CrOjlWjFluk3/i
7rT8yoOcZ+cMYxhYopPo79Ygc7KHNaKC14sqQJQANhs9CLcH6zZo5Eln+6ruJ/6Q6KxR439iPywA
g/18rgaYoNULZASftL3p1MAkD+AOBg+jAHvdC/+6qCVyf/YcZZNECeNGfYnlVtmf2Dii6VWg5oyl
dVa+GpcW9Z1Z3GvdcUNtu1ggEmzQx45OnXype4Gs7Tk1boNpErB4wCozexiDM6pj+P5kERBupV9K
9VTmkCOvx5v9I3ZlXU6fkek3Ahy0CwTu5UzZoCLHQInz/p7tyTmJzbF/6cru2WnMcA7MbrQGLERI
55+SDxF67cdObJnyzAxlmN32919WQE5jXS6Yg/6HldGUZQ3k6qU/C/uoA8BhGVjFjZGxqPLSlNUc
34Tgm4Sx/NP+vIEh7IxIYrwaoxC9t6USsPWm0OhgKjt9x0ASK0k9VWYBzUl2WfEG0hYgxw2CabOn
ik4ixsucGZ4mE5WSgtPOHn6ihFI1KSi9TSn/JC/QjLID6i59DvTS3Z7YMlX9XLZDF3gRIgSjyBAY
lW7v/HkGqa73tP7vfIUdKEUX989IK3SwluQwkr3h3CkKJGJJr4tnMlXSclOG53+m0xPIyeRj/Xi3
TSrW8ixq3WgAFG0hpps8vUVH1UYKCHOGAXBnA9GKhu8crMUHvfUNPIah1XG+7vQRTkuwlrwvcgIF
gsR1kWBILemDZ8hH3iQUol+lgDKHki2aDHB3m7OjFvx7W5akdHCT8qKYo/o2tLFCIFMmHtmAuCcc
+P15ZdUAwj9DkZFHWIEfE+Ubaq98H7dDFiXvFxoagKSdXp4hF9gJwNw3DX8jlmw2BkRjbKVXWMtB
8BR0fO93N4P6wvX6Sbb3VBCQJjV+ERHITNpY5SSOCS6tQtUOyDNow62RF1a+RLKOdczJ0uqb6/Pg
gn5T5n9uo+48YPdioO+zAKOrSk/YP8OLb+XRYel03cxjr6eSdUPeikGP/6KMoGIim7WMqF2+lr7q
gSAS8dpfR1NvbPsBqA/U0h1esresyiHibg4O8hH25vA44MoXEn59SaCXQn05bvIHL+dWoXkxn3ZD
6R6Z2VHIaxFxi8qQml4mWf4tlOVJ1ka63aWIWYF2zCzZVBl0Q2ee9ziXwLk81PUAxr//nX+4sAJ8
6tDx8KezCAjypVsKXUW2sZc1VPfN8+U3GxPt/iDGrCwHe5EQD4rUVlmxE4eEIGhqCAarWVYnBGlx
3kkqiwCSwslGbSiCxTPY9ecT7/pi6VZFZFeO+EAPaaPHaYs0x0R74SjQx7A6gNB9gMx3N42IjjEL
ibRmVsuR+MLD98+ugEMrQLvBwZr7mJn0m2LKlPQbjimCMF4O/FJFEr+5T002IWWuD5lCDa5Iacrl
fjMH+LFOw+6ox0Nr7WXfB637L4R10w7Fc/mx91cLRfow1iH6RV+p+1r6UNInhAJgfvgDlaPOns7c
3lXkcJKlm1RWRR0xk+0BqA/bv3husu65exbKDZ1grgwRo+dXzAailx9v1d1IgknRlDIMTmYytX+Q
yfd8V7aB6M0c8wLGcBgUjgO4upzKtb8bNFz6vdUxnx/U4zgOGsMqg4oV05GN1GrQi5FptoSnD2Hn
+m3fBC4BNlL+Apk1FHt8+DjnUS/9W22a2JXe1ssYafTaReZpn6Hx7vr5sWgJQ2awM3Au+MFJUzfB
PP6bXl+4ht//0QVFtqjP9r10koe6tIN+CA7OqstjB3ZF3C/SR+YAiMroV2D8Z7DIlOBjioQwhqNo
74LW5gtu0VCMrnWvjVR+geihY/Las6h60iC6Xh329BVTBTtNOsLJ5VoBq6p8U6sbqkYSGqXrF8ZX
Vxr6hinJD/p/taLKomETBRqweLWELG1dFZpazaw/sA2ajVDBYAgM47FjdFYh6N7tE6bFIivI1Zkb
LmatDrO9tHTKZ6i1ibUz0h0g13ZolTsrRuRsj3OV3H8whEqWgmhjLewhuhjHH29sFLRKkL6oHQp+
VuNuZzp8SnLebKlwWDehiOPK9VDJ/lajB2u+DMzinw9zNJrErKUCszkundDxg3apwQXLC3ElzKEC
kxrjVLDaKDPABYsD0b+l7KLnH6lDf+tosCNR94gDkwerRtNtALpsAOu9ocJqXaSoAKLYSTWk4RP6
LCRBpHBSflpmiLBE/xFgq9Z1pixRil34WHW6HP+myJnuU3A4QEGoAR5YpHyFJ8H2UFwkiReHWHR8
V7a0Mpk1LH7236mSe1rV9IjrYIcbGTJHIcYaeNPU6ZD0zZadvsdEvunpQdUfBSOhn4x6arRn1K66
d3SNWk66hPDhaJym4m3OZ2ZD6Osh4zLiD3qs8Tpv2RhgRKvcYF06axGDCx4fzsTVhJlNSoybu8yG
mhbd66R/V1Tmh/s9mmZ6TL7JTFPHPKoTJInLBGtSpoBslJNwYNOsYebAl8g1BNyn9VrdiwTucJQY
KXHsBIacZOojxzEqEVvl+I9HHV5FmALG4NhVC5stwXLryevIZri3wAPmaQIP5AN5rRIzACbMArrp
8SErKXZopsaKrF3u9eQWTBu27N9IFA97ez+0Xj7paWsFa4iByeHKkNO1YJHA9sqr+M2E9KcC2x4c
MPn+Tng7TR8nTcOt5UmSKqB55BZtBKPsQQbLE0SQ5DNsVaQtoxcgU3KsPLg908xuQAeKpqD4NL4G
SnOQDbncxPkmK86irZ10Ea9S/N1SyuO15j3vaQLU3EdRMpER7QFOqc/fI4sMLOV9ZePfuvEg+WEq
hgQC+nRu/iPdc4rHRmfMJ/NVq+JyHu9/CRtXTOQLhKCEucknHbRbsTRa+s0EQCgAT5AoAv0NHcEf
tV9d3WYyraouw/HmzcmRmUNOldJBkpNx2imJ7RBhhZpNFSc+wMsvIvZM0Wcr1Y3mMbkqx2Dp4Oo4
dkDiCvQMIjK9Isb2ZFiLSFW8YPhYxStHu89kNPocpCevemajAQARVwH/6Z/hpb58ehucbKl//Sbm
jkf+V81LTAxJJ3iwZ/rVEmUfxJVBZFiYJ83XgLvFRrtfsoD4hNZBGxrrrJtlp08LB1hPgWmkw2X7
tBlmSVapTOOVSGG0tFO1m3ydIW9cepcy7QDfmTnoTkiWqf3BMnOjPb9rxyi/yqUrOS+W7YUFC8pq
DGPt3KuK5Ylh4a+DkQs8IC+sRIuUKawiso3EUQEysFn6mypB3E3dxUJukrJGMwB1DaSCrp4nEF3A
354dXbqg0ZY3w1CO0V9/q2ctsLbbW4a1yWuwSb4a18mwhSxtL4DhH/QeZQsAJswpS3zWa8pUmqTd
ffaf+mqG5rExEC1dUqqqdbRkqYuWveg1bCk9OfJofag9qFdYQ/F5z4tuSWANmw9Ulf6ig9MoLuYu
QMvqS55/XH3UWuxXGaiAKl9cZnXehvsD/CanJdFJy6ObV6Y2RGMq6TbJB+eEp2MzbPaiQO4xwlGR
y8Mrobk99AE0AkSKvyU3NGzyd4igpsXSbPa0Dr2+6LwGYPfVp6Iu/cRfGJ1jzn4enkWR4I+ek0X1
FwVLV40D6zlpeqU+08aUVe4lHRS4f74n2uytinfxSA3+mrN6p60z7e/plpKBV8XwqqgXglPqzOV0
1ntq3r6/fg0ZRrba6NQ1jI3ZGnICkYEAQVDNUxDe++anwXiWPi1tpJiih18PDAkJn+gC1+bkHNMn
iYgSQymDsTY8b8yk3xI5f1l9lK0rHv6g7C+JrTC6pdN7wkc/GwF0H9K6IqeD3PXjf1N8b7yA5d4j
xN/99lakYpafj1T8CFRgdfvJ4JX0jI3JYjWK0MSkx6P0n/mTZBE1lvARhJLiV2Gac6Kaa9gx6EOl
Z69YPPYJBiMyhSQOEvfxVm7CE+LRvT4HUbsya9lNIfZJNXdPJzzzZZaNRFG+UbYaaM6ktfonQmH8
TBQDFVc4MgZmN3m2Si5ZnZUf7GBVMRZD+dW8TJYcyu6zbU+VkMvzGs47A1q7ZgVllBicIUv9kgi1
bio7m+7xtXEEbWPuHxxCcahpkdwetpqAjSgd8GNQEfVD4bJIXnu9AhrW8tuQNM3b5PWDN1qCL1BX
hIDK2I6KgocCNTBcpfJv8JxpXjPsLgVXIv8+MKQSiP/OKJykQg3dQuzNEuP2tbQUWKV+rF2J8XcY
dMcHEKQBXwtWTyFiG5EYUwaqBhjD0DnpgdKUdX529iyNYVaavwhFK+RITkGyDtrZx7sCrw1Vgch9
g0CEwgqYXSVMuYZI9lIQF/gukPIpA4QHR1DYUumndk4PXF0MDGePoAXygz0vtQ4j6zYH0QYaRDxQ
nWLWfV4PwwAVbgkGUd3RLbBpLk4Q9SJsx5icZjS59a9s238mrOuzGkUH5OJnkqKmJCHFoMnNGGvJ
G3y9ScVzxh3x8v1/GycIvrXVpzqV4kHeE4/xCrYM4myF2SQX9Z5eEOn3YWcA2hAUAO2Cs3i1Ao3h
qQRBSzL6bQHJl4/1dhQqxD94Wpgfr4Xiwto3YJqXcV68TpD3gdRo8wWRYez94bBSgj5/mMf70sxw
tzEjLHT3iY3Hb5/gdBD30GVnw2UAGxCRAKIABf5DzzXzPdaMcvZ1o3IL8MjKWd58iEpublevtfbP
Azx+NcIt2px2+mufOslE+g3lKAx9687u4ekHu1IfI6QY2Xw/xPQMhDh9qzQ/zLbLwT8jRVdfzPYg
iM6hcPAByBZo0Zeczfum5X620FP+Ytn6WmgwsZ/ipRfRiBS2VDFctquGnoIkRfOwbIVrS8Ts3kRE
fZxhKdJClYTIESXYLpZpoqUcn7wiRuR/h5eKWSbjzcFue8fAfhq8Dj+cRLJqgfkVunRsWJNp81Tt
k4vF6DRAUrhUyvB2fVktmYtSaMcSTVhVaujav6IqJYSU3VIbJSxYcqkEJeXdMHe6uEmELpA1tx/f
i4I3gkK3QeaQAY2WYuhGM800B9K4wB5/iHk2Ayu/iiNGamIMcAtj0LyLd5cyc1w3scOOWzDpmVHQ
Dihzi8gRv17LxinLv06We2Bq0xoVtTTspzDk4LIiPRP5/w1WWo8jVZp5IhrIHhNloHpKiBBKw1JE
htNNOTPWLB2vehoZ3O0g3SjGywcPY5ZVrNfZBTukr8B7Ag6mkSvL4YQ74TuHkpx/SNQo0yXBOFWJ
H6mu91L03+kA9z77KcRjRFQXNRx6Zj5hJZc5hl+98lt7ZbbliDkrt0OtvMiDjeuH5782bTL02GkT
Hs0PuWQCep4Hn7Z+ZOz9P5iUT+5sJwjmGQ0DmmHcX+pkeHu90eTSg5YO9hijHKGotyxoXj2wKJoZ
rfrRSqamf8e7GPpVDnglwMsThPZV8c77KV9Uv3eR47FMZoT9dfjIovCcRbfTwAxONkdtO19XkAJU
KIzJWDhlkeWx1cNsJCsJ+Vw3vD+GPqTuWVn3l173n5NzMH7d4Y8Plr5J8Wei3TnLiEIAcIEgqu5/
eKVIu1Hi5GZ9PaNZ1BD29XLWxLTJIHoRDORaJXk0R7Jf6FW0ynBRbuL3Zaaxy3h78WMCSp2k64CF
V18rZZqAWag/cr6qG7EQ8QjzSB5mlhDBOzjT8Cp59o3NTRfdSZcXYwIwsRiD1xS4Zdd0gZdf2J/x
wK1v5M5+jsbFSC8LSUpxosU+6iSsr9JhP5DtZKEwydXuFwJAoR78cfpEL2rFMjfSMw9D0Jv6q1Gq
esxmxLx81yjH/mwzcVs09ipsYKPeklHHhVKZAq+MVVNdJiREkmi50TSthfgjmGFrWxd5Ikc/I0pv
r27v154qXuv+2fugKpHe+TDDNtRJNMbzucEb86bx3k2E4FF9oPuyJXcnycjfA5WcsOsj1AFoqveY
mLWGiApA1wqOHxGGNyC56sUecUX59Hb6MEirJrO9qgjvR4iIOngPkWMCQz/u+6JjLQF1198gbvW4
i9+FdNTtZNvTNJEsHfX+AuMr1ylatT96hwGrKimA5Qcm5g2FLR4+RuMfoo65D8Q1+wh+z2bkY5EC
+tvlQMMgOzjHCb2z3dXrCnDomv3KifppA+hI5vxCB/Wiytp1iHdDhInkT6xrga0JuwNKG0cXq6gc
0gZxLYsevNZEVpyJR9z/96R0dykh4Tcky7RZEh0b6HqT8PeT9Rdd36WnZPOh47T3bIxlzkEQItk4
ipc+aQ4gC5YIOT6QTfQ9Rn1MOuqLCoqLTM+XnQ5GZjoFAvxliK1ac0quFIR+nP4NnF9pEbY/vMkH
fgitKiJicCbLa10iIvzH/DiIYyFBO1NKKswL8yJaPlT6rZ+mUZCtpjhKyBtgp8v2uhB8LWO2gNVf
+kKBqhSIjNbiDqdxcQUpYcKYeotXXzGRTQ/DHBkuHizJeRX/k3RDH191XYXlWbhHvgHccgx/Fooi
KVPgKcRiH/Nk5hjQANghmMXreUwT+Jet+0a0xEuyMY7NH2igkuukj76Sb7WrxI+Xqp5lBaYwUF1a
+OWXA821upvZ9OVeu+NJutP3NwmupEaT90bBTFf6x29OF4NX0VXwj2im2Icfyu4mNEmCqtUiB9co
OipKn5W5gsERDBui12HRffSQoJuzyoj98uld+JoBaGqyRX21JT4hPbFpOeut2niK06/7ycq37Saa
mJmdO4jBU7AZowQI/RzlQxhSg87ZUeparH+B/eFPb0/WzacWSl1MAYT/vZoUIdq6UJiHnJoerq7J
r5pnSWa4agAKuM4b8OUIRXWNNfgnUf2bHTVCT6xlRsg68AOP1DzbYa8zoD8/yG5Sw1JvPjRXWuyV
u/IbHMPr72I0eNNfC9zgRwXrpg3L9JwzVO2u3KS+imi9dArtizIaqjPF+xCOkUv2LRN1031g+UBh
wJXwfZcjG2Jxajh3AewObpMGTLlk6Aovp40aS4Wc8R3YXgcVY+V+fWNETUmfDDVr423+YJQP2Yqs
GG5id0lmaKupsgeDawxGfs+lHg/Wd2MZjFVVi3eFEGvAinSkeX9DaRkmubm/vqDu3FcyXPLko4As
SdJtgJsaWd7enJoJZNITvmo1nrqQLHBB1jdEPYSpmvVd85sVI/heSkRQBK1UCRfZ62O1YtzE9f5Z
6s9KPcCMnEpO72E38+7UrBFXYZ7qLiHc26rzbH/Px21R4Nruc2wG92MtLoFql5F7L9Pd9evxkkAo
u74J/5lckQaxN3i774cXIrprUoAAhVlbUlZzGgjsjFNfl2eWt6967ysegdrLPvX1IsaweggPNEL+
wm3vE2+NZsVmTt3eMq3N28Y0kpESN0UQEdRWNnov8CqrSpymYLIAB4H8v4uVb3J6gEDNzHL49QBY
t7CriuFjqctmZOq1BiP9DtOzrl6s80a/jqkqpGmhcOseTV12FWq36TNt5TOHy/w14XkZagHALSe+
44gz/ARAdiWKoNnXsp0VRqXXjhnTEEslx6oeiPstEKHvKZzo1qDKRWwoLYZPSTgp8K1D/5J0a+9Z
gLYwqWgD4lf6aeaTVj19y4Eo+XtHZA7DRRm9IZgGT+/pssFAYHqEWHzXu3lbEglw+oNa+ZK0jAVi
ZVoxTxXX1AExYb5H85xNN9GTggi9v2pIBRlUecXHL1bZxsR185x0tyGSXtAvPMDTYJ3D/bljBUfh
weO/B0+Ai/4UY9lFPX2Mufes2AXuMm71rDd8CRXCKz3sClKKWlca0sjS4GupUuE1yH2Nq3gJWlXs
iQ/L0GqvvwPDlCHg+/abv6STCTe86sH1iPUO9oY97Rd3I3mMF9Qs60SkaH1Rl+eZo6WtVoiT+1Ha
q/6YDb6xy9+mkR47r5V7m57ng6esCBf8mlX7sOdzjFULgn9ymMU1lCilP5/sC6ouwbydAiYslUBN
DG8HZdSqAMhH9FR0A8JAJD64hb2RK+PESO2PfajJpuzrLG1wlj9fabv1q3CotzugsnnAzijR0/Hq
hd6b/+up49LM83F31R8Q0o3qDB8EGp/TE1Jimbku+dv+Vsu8iOH3XBLUeMZe9s3Sh1mCQ3gacpH3
xEBnkfaVT+WWpkmJ/JUVAynzkNrHIMRba1NT/M2nJURasZPsvz/DEVXzRuJb06+X8Dm0L3No5oL/
TDVDsl5BuAZhhCuqupGTTT70L05AxMstMd2pFaVrJQF/CA14k+c1yCbRJ4q+iscrUQVHFKXUiukx
5BocL1TID7E+zxe8ge06sn1qhiuCdmqEfpQ5P/+QJhZ5fc3MN7ZcGB02gcEy88596XVCxPwlowHT
niphUM2wEci/UKf9OUTkBAyexXSq4QO4PRbkLif3dUdXPBOXvAosShGlH9DKoIHxbam7qF3Dn6VO
/RTdDqd+hfQiZma83NXD2PF1KAzQRFWRNGBWxM4duGv4mjMZOFpukFV2fBgNNLdVOHxAWX3uKzF8
8vscfi2aPsk4FtbAG5fh2lwpkzXE3UT1Llj3WhcZjIfiamFAFqCTgvYQtjpIHh7+jAMDd5yxwwwo
w8ZWe+pnHDOFSmRWkVoEUkiHQAmSGn/lZU5FWlrgXbjOK7tMfZK4TyrOI00s20uQmwVq8rOwveMM
kkNem4t8lKvOCar4wuMBZ8LOaBpYR69ty3ReWuBiEbgAChJP/rYZn22w6XHC9SLukzj55zpVsY0J
NwXKEo7KPjZ/hDSSM8+ahONxmCyi8NyAyIOSsrZM68ma4bHAJSlGq3idwo3JiIlsMhDjCCrLSEcZ
PTF9vH8NIpgoOh/honaeF1G6AUrDq889YdN7WdjY2Evo3fHWMuuHmLPJX3AW0YGNQ7aWGCU6h9wH
NUbZndfw089UhgGUqTOxf7Q+k7haESaz6XEDMyOemH6nxK8Kw2pcm+r80lbUAX4deRxte5K/Vo01
k+v5mzq4y18s7YEAXXZpVsjKZp3JwibWskuvjcrbl4zQvrKGgcQ6090VEFfQfn2lPxfzsJZGlcwY
PrG07xHEj6u/faGJCXihWmtP0PlgcDpSpghakpsCEfzM2YTXSqMwYPnHSMvExN0CuIl6/1idj2Cc
fUOdETgfUcMEcYTHUIa5dWzxFkGs0ZWtN+WCvCP9Zu9ryHHAS64R1bEBPOUu5DCyDfiQFUFSCyMm
+nAA6AdyM0EOPN/GwnSuUBJd2UIPzWHXhD7cHCq7CB89OJbWl2XMYsWIAUyzit3RQv/X2bMk64Q0
BxIX3HoC7gOgRU3QwD5doG9thLlpOFPeRMICPdmRg+2JHDoEQUwG9u+VlgW9WFhiTUQaESMU2Xrb
mY41BRYhBhRroc8mx+G+I9m7mZs5cKvYxFdysYQxGkKQ+yc9KmZgIq5KIm7Joha1EEFhd4XQ706p
aYi156gHryI67VbqDz6Mxzz1HSHE71FkOjiUFMTI91EKUEnzsC3ItJaf25ZVaIfZzXQppOw6LPkj
lRytIFjOSaUmqoSxcWHmEJq/5GA1sBvk8nzITyezUad59H4/DAzgle3BTC0N0AI9xAuJQKet/c20
jFw56aMr792igqhDy3JIV9SENEaoeOGWJMFMx4kkrnjU7xmAANKjO7FpEw11I1uUxh1d49wHNY34
mNzR3Dj04zo7ndxjDhzfbkhPDI3O44XnRDHUWs/P7mvg9qXLcjcVgGCpELo2lP8g3YirGxhonf5X
6SWhGO0ib6Ih6rOHqcgJwmKc0XEmqWULzYWBTqvSVvoCLcl3/5OGYq14JHOZtviRaxc5vfQvluZB
bRSd0BT+Cd1W0+hCDNyv9rZM/Ys4+o5+JzuU705IP2UsxvAa6tbWpYGmBHVR6PnZqDx7d/jihcUL
l7aCve43g98kom5GK2Fgw4zJZJf0LzbW3Q0Gi3wkCl+dZq6Uoqe1M6XaB/hs5MKAMBMXwuqVRZv9
jE3KN9+ezUEa8UJOiaRelOsDgR8+0yq7pgORKphNdZFziMGkxCGsYhnMUp/Uu4272/OFvj4FFYNZ
V67M88Z9IXQa9G3WwfgM5AOzzgeywQw6S0ZsM+7ftG3QcQQBzPkobh2A9ygVXffkxtwoFR6jNPYI
fHORlb4F96s/MxxS5u5ZnoxvcfybKgHPxJ5NQ4tLxjxLJEHd7lb5wgQEyn7nIBPUoWQz+uRORdtt
cqDHCejHpJ/5pU2GbEOwnwrfqTeOM5bwsfhcOPXVXRNz7Oe8kZCXxCZoqxbbITbu28CF6jaMGumj
EsoTz4VYX+AWdMf9d8GK9v6pT5J1l8oEsJvg5dF+ET4WaitV+YoIy82ODmu2RCyqnDAXOg7RnJfq
T9jqooTeyKHhOmTdO+akup5AQ+geBkH+bo583c60Gosp4Oi+fUE142YHYTq2OYLIUFMmpETxwSdJ
xMiVqrUrh+rXXhkb6BsErmBULhZAuwufP8mhF6Fhz5ZHwvPCIgvEsC9CUR3qFKNgsWvNTTfzWheq
pXJGiLcIuvRjzbwPmiY15ZPF5zLPFTtQYdOW+Vrfh6UUZJjoP4M23du8rIyyAV90n5mILiMpBwO8
DAwuSWwwgQUa3Rpunj1McVKdKsGRUq6Q9WvelTk1iXprSEyrcM7UNnITDYrCFXuVniSM+3lz5c6v
uDag5SV8k1In1bz8UtTa76AbjeZFgyJRSGf3lFrYCe4/iX8yDsCrizhrBB3EfP3apX90FQcm/gyx
tMz5COblgVdE6q458HYc7c6i+Q4w3I2HOBljhY3QhN8vHvDMtBP/vdWqEI87tlpcaRWBUGDS/A4H
YWDQnm/EJ7GNq5MmlgYjeBVanC5O8n4H/pGydGcC1d+w43PKoRdSjSDtBCLhy52+Okij6+Zuefg4
8oJ2hXEi9WkujI2yXjuhhPNw8NDHaKyfG29LuSRR7ow4vodxvjWUoUtGTlvR6uONHf7OVjnIB7ge
rICCop/tR/m/U/hvm0SeFrCgJa9tXHO5Lm5ijN8gc8dayk9v9e7WoYvVhVTfU/mZYOtZCdveMUg6
Q8Abhx2dUYekYimciiMWwLYN9x0YpcKXzlfXzmPhkncUe8VTPYSbePPeELjEYde/b92QxjUIEbbs
2HN1vJT9eVthT5cI/NNqi+1SPDLa1oCrUXFtlCcMVgBLVtDP11jE5NuBvbHLNzaTSmPExRRAKLYB
q6UaFyKRrcZoIJMlObDutZVpcenXDdAUrB8NrWygF56exBeC4yBLxWK69fgRwo0zV88Zjwd3vce+
P1r1N3p37yv6JPqog2Ffius61zSuI6O40Vn4oE23wu1VCaDECc3SQeErlKWk65qw+0ckJ6/fChyu
FdSDgckAmSO619pJgnelYadASH4ANgJFaG954UeKD4diITRTto//OkJB6+olo7zePlp2DOw7odv8
CX1LKlQFSZlLtHDHIKyFAyy1Sn3tgr0TMnzUKDDj8Jstd91zNzI2fnRLSZojjBapP1qH9nHqXgmK
VsAVzKMIH6Zr68PveybjiVwy8WxtnkI/vOkaGaNF8Yo6Menfm+naKw8GyFKrg/o9QvXsFMwcGDDf
oDMFVF6VJkER1SgKApNKgjUnLPE4HnxDlOsistiI0ACdjdjR62OxPzzOqLk+3dkjb02E5X82Xx8T
OPle+qFfeKm03WG1NqSgoB5qIQPxJZWIaQRAu5WbjMbQYQNiL2YsIdoed/ByJEFyB1BcGhT7KMZH
5fsGjf35PQkyt4fDpPC4paC1QbWThO/cCpLD5AxS4WdXuzR/qkCcg8sAFagpZLPFp/hGE1xdfSMO
rYktzx1hJsXi5pMupOQDOA6oj8BrW2BwPuwpYWV0nz4H5NgoIeP5Tm2jdSoIhGc/UQwvQOPJXgFy
qsJC9tu14g0q6TrnHQVs4WRTeWPWgSnpXgBBqCLRSUPj1ivbUtM44+eIRaFYYoRu3VnTU/c7wmD9
3oQMhnmVW6EOPhTBoBrNcY0aWOcQqqSFICIBXNTL4Nj7X2UCLaHg3iZOuyKgyfg0xErVZsM4/Goh
5TQPmmxNFVYN6TlDR5Fa5Hcsh5+E+mfoZrkdFf4wzKBno70dnBSkKJzHFxRkrjszfn6Jw0kMDJIp
rr1oM1B1LJCRuzeDkv1gAyXbXHjciKkwlYexTodjT8EB7nJuUqYC43MtZm1t9aUWnMbKybk9Gdue
mpHVPYOwdpSGxqeI0g6suM1yHDGJEf0eQck4JsyKtiKKXAA95x6PiJ0C8VM7h3js6Yj2L5B0nnAi
QgA6eLuKQclwBmFd32x0hVfYm49GsvMQ0eldz9O3w7tvtvVw03L2V8oovlXIH8yeFY/CKYnhAJtx
h/PoV3Yx7s+SV3PWccMBIWJAOnfHzB+BSKre0nhwEXLoXVXxykGCNxm9hmFsOr8YNm53qEXCabLS
0K9rImb11eTEo/N803PYWS9Q6RRD06JXYKTgUYw6Qcx6JqHaMACbZvcbs/Eq8qRnA2SQTZs9Mx83
GTOH41GrU844XoJQ+MjjHjJPzPKGkSP3IUxtD1aVujZM6K1BHpzLUQ99mAT9fEEs5VakEm7iNCj7
TfOx73NANXTaT005KI7nrcOelAZBY04wu+mtHP02abld0ic2WQ/c5+VOX9bhGEWpZaVLSFKJ4ErJ
jPxcX0mZfKduJxvy/m8fHBNCr343Chmy2sc4l1wW8FPmqXW/Ng9HVzdI/cNKcsrv1KUfgGTzXTbt
oe0B6WTdhdv0dyi5vUuBiiycGVx68yALTEttDsYvjcBuiwMv+XfWu5bmfFRuEh+PRGZIcUn7WmXn
hCdRQnjd0cNYe1P8p1ZC01lvKAaVZWbVnIwSoEweed4icXgtqGrAYWBmYnIeb+azpy3tl2C5V2J0
gpdcvNWB/9hSEWnaKlHqDhn1AQ9DJ5Qmq7+Sq9nBVIUvz2grUbf4YU3rvHLv481qmDHhVGm1L1Ql
sNPSjndzCUXb4RTYdK+xjZn3vzIajyBXDSC/g9Z9Q90yFAMJOqpNVjgtnLdZJs7N2ZmZV6LuuD1/
oNV9TLVcHzc8If/2WQeAncGeROCueIeKIJtRSgCKhM9KLRlrAxxaLb8M2b42HyRTRUhkEn+rUZBS
h/KD53J9kUGlDAEzljhPNBAHX7LtYDplU7ZaDSyazHoM2gSWPRjqCFnGUesQcPGdd93KL1/VLMre
3UAreIj0oUqBHVZRnKkA3wwv+6NKT1S2jmf+F9BSQXZYgUtt+fCkvD6KfVT+p2ixqwu/j0Soxodd
AmhAqbi+MGSGq+218V70z4TwLedBgqcQ2ZUqBuLM4BtEKn4LXZ85BgAfMth5noEgYEAvrbsBy1pO
Bm8s2uKgLNVTkGvEe6cFIWCZGrIjFu9YvxQG8w1W3D/FSueWXi/pNqjWUG15J13fb6qihQEpOiNi
RGhZwhetULE0reT2dg/Toj/WAR9FdkasCjcMXypSvDdC/LGgBdzKXqXubVdF9TxzFuyit6FJWgaB
R93klzRZ334UwJV+IYfb1QLkz6cZgqirQ/ERoqcS7jPD6Osw73NURmgzqVcDtOocKt+JUHmJM4BK
EsRmGEnBgkiGSNxpU6GbWSHT5HcJkKKeHMAXECAhGdmrlgM44lcx0wpv+TgO7JhFQs1SnF7WcZTo
1pamKGGatpUho+FjVGZgcc+TC8YXKCZgA46d+sMQQe+aXZOFLYQI6tsZZK7GbWUTvXOkqQWF5oMo
iJQa+dacEtjF9KOsTUE3xT2ntvFNZ4GjeKSq4SlcIi0/BCnlbmM1Ui844U3rk9lgulsTmG6jZl4o
5DyikmCCXaTMlbBgPsVTluRTHPVAM9ElUHUz5BApdAx4GV288C2NmSqhK8YvykuT4eNyTLVlkHJV
qHejLeJT2yYUQAX8YV6MKIUiA6gP+/GiTlbMvIhQPnH9fPptVo093DwRLfb4YSjy/3RFXgzrkb0L
tnpx/3U9ALZYILuqf8b9y7rFPtMewqfeiAA5vVKI2ktaOB88znYr0sl1qgirCoT1yHYaEdZOxH7s
QPLTaIxUzADwFG0f0wQ5iwKnUIIx6SjwHXkISYBD6n/kPWdPCNiDzbYC6qKJVAd1lRj9Kmb1H+CE
of8g6FKDpRk73ORCSP3+Huy0uPGdGNMGSSOyp+US6pKz8GDGQjZKsCidoTmLP8a7yaLptiMvtzFX
Am1+zNQeBcnYQ22mcXklCSXvxIyjWsqgXowUDSuhzuOXicm4mJuyrGj+bpr+6XRSN4oPSU4bMyWe
Ho8143XL5iedXE/Nofq3lad4vOIULtXvAAgOobIq6FR28dpoGKucRWMbaNJplfEGloDewLig7fFd
QAJwW4FQh+kHaj3Wq+DGUg+pMe72wKf/FVpDffdgft4INOns4LmCnmULqD0XvoJPc8xpCphZYAbH
q/M4mDU+4nj0ZYt6EZMO7/UJ6Aj/743WotKzQoGIjyLjqNOw0E4B78lnU5j7ZGfLolVGFNBtevMG
NSC3d2d9QHubGt44eqdSEBqOXYte/Wb2Wp/8m58YLimc38B5P84eKRvlN/DNPwoMlS/iHYpRN/bi
75snzKblD3hu/o+Jw1X8qzP6a9wSgn4PIgZM8LIPHwXLyG1/odedGGb2IJoz80aKj44ut9gzzvnG
G8gjp8dSYXuEpR97936fDD+yV0ilTx0o92HxTViZmcV7yuDFah7/7XFjhXSn8lePJumTPq1z4BdB
BsYwVIhahzK9graIWQJ6onBneH8RMEOOFw+/fRSCw0NH4UslK+93LuwkDDYNnNk4ept2G9roSMTH
x63I8ZP1oRzn/uv2X9P4JkfQ47iItmZgj1CBzHoY3OVQclmaniodHhR0y6M0d8AFfg7px+haycna
RxB5Gz3BlSY0lI+lSNR/8IHL/mH92xu6vbAd3wUvGhv18fkL8IChLkXhWGM6njVI/+nQusy8p5Na
jLdJEZ7azMWvFNmsGiMZzSwkmG4K/pFivDVHoi5ohg0zIvbQa/D8IRkCF4dIErw4/sLYr4L91qXo
KXL827bLvcmlwH26uKPw4JG976zTIc1r4N1fgu00cqWgYhtrY9LJf0gR7gxYOCg81Px7DRjdmyoo
ZbFI7nse/Le4jqFkZCJLr2UZwhnD3s88oBCdWugl8WJDoh+wkTChjxMBCtlBqFvMqGohpaN7IpLi
GoxZkwuYfhzIWmYv0MRWEZ1Zv2nADr9/igsyKOr7SiZFmOES/1B+zaQAgAyFLMToOy9oCW8a877m
vYpFerimSTm3AAoCkq4U67AZBpdJRTvz3IA7xxhOGw5v2U5obdlL4GQkdJSNh/RodWOl7oh7orlu
9OvV1Q4lpJztN9dI886hNF3ruSaDzHsVoHLrnPHhHCPSnobcGZCwq/jMpcGLyooNzS5VlCqLCCnA
8XgzEcN2Q85oHleuf95YoMZmjnO4eqPwJEt3t9aZAnKc+mC3RgXseKzSsCAdnAaSV+nbO8aPii35
s0NBYJ0fNK5F7oWU8Yunn6TT7NIIApc64MmgcnmFnPYXC+TPmLOvz4d91JTt+TZ4S8aRldEKfnid
BMuokISWARIH8Qu4Qgi7e5hJefkZpbssaLLyxH5vrKGN49P16e9JZfaPjwWlpeM8/j2ImTbdrvN4
bGfXOcbAQYSY8wtenubfMliYZlBCd1Pm+3BdCGYBLh7oiPlA4CtfFT8et8OULtTowU6m0tFEaJ+3
t2XwNGAv9DfxHY1dj5ZAq4YPztsNFryJKisZg3oXGLW0Ta8Gh29rmVCwhceOOYfZw/GALM035thI
mOqTPOlYcYmAtKS2Sd262vy+xO3DlwKNI8Kax5aEmfLlMqx5mKrwkWj47RCqc4AUXmeGFNqvA47q
8TNGZNG6VhHirsTllHu3D+fr6PfX2xtTTEZ/jmEsj0hyuJY21cNx7vnk7agEnYx9lFZbDFYtoduI
Ef/W5NsjFPfKm2iBvDyJBW/lKPm3xsinj3hCkPEPFbdDHbwTApMMvGa5/CCYjskIyIWiu2sKXBJW
lM/kDGRAO0DgnlH2qp3xGwZfJynzjDTSGi38I9KRypOnTu51x0X7T7RJhAKe8pdY8x5F+KgPrw41
dg2HtBhHC5pVH1dvAzmxZPdLmLTdh2OWdNR/XV/SqIKSxhxHpmfZMqBExAkG68dHTjCOIY0mvvbN
/vFCMhKZMoOAXPPI8cTcWxJ3bFSveBnThj9dQO+tAt1Go7vxqRqjGM9FuwKP/JoZdu2MIoAxqFUg
g5G3nk43JSRHFo/cygh6usNpCAJu0MMsEPvFK6pkhCTXq9bxBilbuROKFhi6GoGMeLnsCxmy9NYc
9RNVOAUqAeU3PV/0v+sUB/yCYinZBoV1R1bC76lY3wzHy0Zlvj09EJyTDQDSWhdXyCU30bnzLaet
+5v824CELeFN8oxTqXWpFXgSDj1WGMwYSwyI9Ovu6yaa8ClgdJuLVHXQ4Je5+rChsUkrciIkCzCN
7YYU89C3uY98TkdFVdL5xsLX88no7CLQH8pkoY6WaWvKsqhHIrDRI9XyKfrCMiL80ky29qPBsj05
HRuKjGe59mKi7yHb7wz9VksxPewQ0q0Fj+TWXVd9/A4LY3yI4+8oxb3duMhl9Soz8tIiUtaIuf5y
1ZXo0+97uBeGxlJKw6539LjWZ/ih1mVwu93l1CT/hRPeo3lMDwvv3q8bf3YVPrdjkG1rCkbYEEcg
dcbpTqwPFqItGph4h9rEr34bEy2qIMJRnyl19g1X3YoKH2M4U2fWXYyIEBi2r7S5UWATCZRSLUBs
zUd9mNQVVyH1mJkvjE2OQPQQtn5HOvC3ZvAiqJ4RFloHlv5XAN7ilvBh1isYe9gV57oeAnpW76Wh
FUrjPS0b9SdZBzHsTM2l2CiWp05fKYCU3oYifyEmsw6EFBR9V6wvuy1pULpKxtvRzaeGZ1KlYfJg
h3DE07w2Rg2uZMcU6nseQzDLEa4dTBsQZ/EVqvwhZVQYV8/QFXkE85XXUaL1zQ6Pwoe5I0Sjx9iX
6fmMbUL0PdTv7z7S4jdG2qYxFfTMUp23ADXx0zfqIk9IojgHC/u5hoNjAubkUJcfUXWEUx0dQ2uR
ExP9TQc62efyI0sKvbbuyBgyJUs0iAVU3dqEAz67qvYSWwmcNjP8wM3wnqFRAiID9wSwMGBbuMSG
52UL/JoCRYK8B4yTYhaft45NJr6wIOoJrRHJydECiF16jpSzTariGpSz/nLVPmbbrN4+FXFOnc1b
HE1ageyoLwfyTeWupGx5ACnI6xjRqJcQuJgS9NyzzSNTLdIu/lpmUAOOAtdbueKjB/mEJx/MUhAp
cHU3dO4XhNjjdZ0WeICFeUQtMl/nhlBWSPeuYuq7s8TNmjQo+DzyyFUEjCjNxJcoq3dqNgRlrD8z
wRPXpyZQbpWyA8IK7xD+pMauxRl6jUzs9YhxQqfFeEvyuMdhuGGHb/rtw27ldqDQcnyjCmYGHUXS
yZArhR28pYFo5gPXzIqxYXdwm/xLN6ohaBcIxtcxi/CKkwZBTHyIEnQVznGmEUj5xe4rSSlUD2IA
fbQCtsAKTCEx9PUU38bAxwKdKA9+IGGbAFu7XPaHjGmkUvTtzbvwOBqxBwQVzSUrR/7Uw47LL4qI
1FvQFLc0jqmin2yZ5OkOuvwZYj72DvbSoXt0n+CdqwB0BE5iA5IM87njj633SQXJasOOHXIB/Tv3
eoKykApFkix2jecA1cwRd6WW2MfIeMM43H33SyPPCdp0yJkzGfBASqaPpAZcOgrQyBgYEEV5mDbH
L5GpXWnoThpa2OyKDuEsObgLiCCfoAlOsN4fkM432yQiBE1MwJxLTDd0t5u4i2NTyS/WGv+stSZj
6t7e7qHExn28HqfEcW/ywDbaT/JOjxJZluOpjINIBYogx7VHth2qOi7g1LP3BJ+samtgvOEFCeuL
H4XNE6K9OAcRpJvbdy/ih/s/J3fDB92SOPFv4KURBRjvjqM9TBem+AYUclt5RkYL7nBHzbY3RmDP
7U9d9IOTnbfatdA//oNFiRJQsVeDtrC5KNApKUEWyaikuI/fvc9MRlmKdjB1DJ2t+obTPAFx28jz
KtrQqg9tYgjwfQwLOdL0FxzgEm2/rz7pfInxx2YaT38peX6F551H75w5T5cZy8yNhnDQPguhQzW+
A6D6l+/Uh8L2rNXGWBE3fCz8tBCupaq65I/0RbPlFF6wFZztRESCol6/C44VxkSMzpOSoEOGssyW
gXMEbs5QiyjLNzovLYhM4OgPors0qHmaKBqN2Zbq7dsWb6VUT1i70QwoFW+wIo5iC+xGmxHBSl0t
rz0xKpH/imCD8lnu+hfFgLCc6g2WN1ECqrZ0OB7nKwe+EnIXsc6k/wZIPTrsJlSQJFyGOuo+jaFy
Uoe2T750mWCeTV/7FtLuwozhs/TYJLMsDyx+CKWbuXfKrKSqaZND3VcfIQu26cvg8Lz7vCMM1SDy
rv4JYfFusZ/fZwbfBOOqw9YMk88ANoS95EYVBV/E4W0sv3qOHllP+yWLMMlyZg31Yw5nAIa89+jB
wlHqJq0J7nCdzq81E4k5QFt7nU1118R5KekEbCPfdBF4x+KVBrMEYnNkRlhy15W3PhOobhUYZiKN
UJJk9VPZ30iqGy6S+oL9Z3FBRZ4LwycQYdnY6p+rLnXbqweYWI73R8imcopira1ItY4n04ODGfnm
KcC3HG8BcnbLs+12omMdXwVPyknJe7CoctjBjNp2guymapJeXsXLY2fV4PFuIwrpHiKnSpRau4z6
XXUpvelTvzo9w4YF46z/huzT4GBPacGfNWHyFyHJJxzXoVogkjFWOcKJqJV/Nxv7aUt2JlRVByJu
KhQmafrnqcmVe46P5TL8yKE0h7L4IEJ4DjY+p3K6EV3q4aL4OUhm1hgobdDnqfei6+M70wPoHlkA
gK+D9AbLqEtsAvY1XzZjzyvPhSntdIYxrsXaHS9rpcZZ1Av6D7gTtdlD/6Mbjmgj4mzIerkUHkWI
ylUQaONmkPEgFzn8PkaGuIA2/iIxnrgg7DOSF6H7pgIZAmYB21KFM08405ct2nLDkY2mwnFyWECw
D2de41eEYxJZFLItIc3HWk3tDKyQninZY913jyqrl3KlrsHxh2WSn/MP7kLeYkKdaOSlAEsAvKQb
E/awoAkktUu+YLqvJne2++V151bfhbRvns2g3nRqfmcY0TmD+XgW7Lbh5JRyrDJFDtdZx+QfqkH1
+UT4gde2wsUKQaixCVgXFgswyD1/xTnSTCud7FkWa2va9/XloIQu7qucC2GQtvjcrdrEwJpvAx8I
bPbH4fHMGR73Ux3YQsBeFiD2z0PUqdUNymCUuzCkkORpZW/4c4tSpcvC7Fy/4ZBSHGgSxseW69qE
LqvxNv0qrCvPU1bdTywe0tupuZbW0H1F9CSXrfhojm+DY5zR96J5b7T4YJZ4rTFRV1rki2pfJxah
TizM4pfbTNc2cEht4t+h2ct3UxJGA5eOjQRsuke7a2FYhVOtccZ4R0uRZ/qK/inDWYnP+Ufm6ZRG
qRXTNKmE668vY6x5OK8g9OvZ+eQKjVn4CsjKHNxudgnASOn/hV3QIDRkz2BaKORCK1oQa0TQ9Quq
+rULODvhqALt0Ym9BTOTDemdYjaTGaiZRqvC3EFrKWCSp4apSNaXhn31o3I83eNAelkxrT0dAxfF
VXUDF+u+yD1/O2U1smChDaWaFJqurw7zMyC8g+X5isrrx3wsnADQWXQiRgy3Z+mDDH+8/SG3Whhj
vMh5SxLKbZP136VRD/wd+1MEuscQDRSPxXwN/KcElFrpSeP0n5rxXdCLRNhueGMY32eXDELFPCzF
5P5eB+1UZPJdoPK/0wZW0JKLkr55ej8kvy5R/fdJUmkYv96wZA4tFJsVvGpU7P/pp+2WxhPZQPZk
cFHxh7BjouGOXseHqIfcBJk8XmlVUnT7beHOOMvrsUmei5wD12kx4d+OGJER+3qMGKHZwYjJb2e1
wYC9Xwe9+I4H8+IsgajbbchL4QC5OsllFM2PypEsN4a3i+8wEfiCRYRKiXBmlCgCuaNOneG+uj/p
FuDX4Gs+s8ry6tCsDNDRib8xgGWz9Yhf+5LP+gm9DaHU+6c2WpvSaFjfuqVzgMLNRgZlgdvBsP+B
jvZXmVdLJ8/v26C4Zq4RHwwQKtGdW9PUJYmrOF2Kd+KIlvrSe54zBRW3UaR05P07qKs3vr1Sx0AX
QCklkgxzk1gsOPueAId//Qd+jFnuhZLfo28yUQVmEnEfW+2L6/4okksPe1D0qUQ57nfV2JvU7O6y
sIUvbotXyIK92MU6K9kmjpzKntJAxMg6rafQssTl5b8MIDzGzeSoHYJOq0+uiK6JxOD83rNBuC0i
btXY+2SeJctaa0OJiqTGQzvmULfub77/y35UKL8sWR+fex8PMhAfCSfuQTlY6ZZBDAEBken+ugdg
DmgirO4m6bTORSGFQaz0MFLqLYrS4ChHT6FuhRUlmvCBCbDd3bDHJ1H2uLvJycLwRDE6kjE5qCRe
ftfakO1dbM2XPoVqgAqXdR//B/bJw3ZI99mh+GjtbAvDeK5/URJuuFrygoKyENSQ2DPj7WYMfZjN
tl0MJg5w2ddstgClGOGH5sozY7AFVfy5C0VI2LaKClg0kBbgWfpNU7ctqNIWSTamxJKP9p/Dhipm
Dss64z9C9nSFQ2CaaibR5l1n4L1RBeK2Ta0IyGAJB3CBRiHDA8e81CusU6c1FixU4cQU7QWW90Tn
5E4qU71w6ZeKzo+mYAIZMcQlmX8IQFbLrJv86ypuwRBUoYTY4TqoWWGqHU99OythbgWbEu3bd8f2
xTCoA2bEttIBdMSFNnj3k3/OFHKF5bGZ+M4Y6f57Lkx8pX6WqMFQ8xUBlqeESqeVmcDr80UYaOyB
iAvGMV4pQ17z3jyBCVQBwjhf4XGaa3tLWLxyW0sA8EhwBCLLStnIq0LRZrS7OgNX6stvldHQxHrs
gBGL14+t/nPP+NiLz9iIFS+W+yIEO2tZso+1Sqg9jg3MmiYPKfcyCdt6dMG/tu7Qa0VDZX29M8qn
yNuhq3DeKPVCmms0DgYfwlCBK7wRxA681TbEZ1YIZ3Yn4T53TMZAAr0kam3xkCaGS2xDFhfsF/EN
ucpLzew+drHNmlvgE34bmgFH2XIaB5hLqeYuZDsuM7axu7fABx/551elZa4JvjP438K7h/AQE2kA
XS94xRtGNIQA5NI0urauuyNVToj1e1QB8KHcAa5ImXdz6bAhXaO8V0r7WXxrd1IyOU3N8tDtlejt
SkoYRvnmJuPt+IFBxvgW7mLTc4B7ULCOv4cRo6spzzvTshrDDX3flwxx81EFb3TG+bzi+xSdXzVp
3jVBN/VJaVAgo2akuRZozBBnmNhPSr4ESidj2JFJNfSq0elE7NQj4LUgtCy5270mu3RtEFPz8nmg
1zKBBNEtskhpAtQbSIQxz3IRZFKLlDx6PS9YLDv5MyKCBHmFZwT4xMFX+N1DUaBTa0SmSyYgu50c
gPKIiKDd90XuTx5+lozVZ+JYSZkNUO7qQGHGmFdQUxeBCcsOxvxpeNrW0yHo0uzfq4NeEos7Wivd
M09jEv3GniUp9b7A3f1maQ/xtYndtMQXaKEZ/Qi86pT0rD2bcnNIQm6W5+ifdsbAxN+ikywVP3rp
eFw2wMh59czZCI3tlD8y6Rik75ybySKXLtwJWkgkX1Q6Y7M+oujtPOFNU1NJDzbVs02wqyVxQB9T
bL2ppQSMPv680usFDLvzt51cqWOFweolt5nb6f0Q0bEq+ldHxkN0wcPvVWD0Duwt0PIx1vx0jPb7
s7mp53l92n9Sk2gxDKdIbfTU6WFbjKLnNMcMFVcJRCyvrI8UjKJ+mswPzBnTfmbFzzbcNTvzVdh7
HDbAoVB8h14iUSUTqZWS+/Kgef5AvsCf/M5xX78sRlY/RBWZe406DmhssmMqCTJC0WCgWYlI+Gca
dcvYrCZp9z5t0kFLVFxlv2x2Rs19x0F4gQfUnZfRTqjxoAwquIT+uvd1Q4nFU+FEFR9PVe0MTb88
AYbleiQq7NRAlDZRj5M1YsQQw3vI9qGiqoywSTK4zOMizz5XRvDWFyp5AGZaUFbvQxDE/c6OH3cP
4OrYeCiTxfZhfrsE5vnDZ5xMziF70eVZHzPcdPv6o5GLZ5vFktFNxM6qVIZlfxQ5GeI1AjutHhiX
tdIEBrQ+uuT4LaUuk04Ln4px9di4S/vuhqSfo9U8h4Oh8boYaRM/lwe3J4nKWh92Kcqx/FpE38RI
t56pOKyJrkNvhuIDgNHW6kULmxesjdsxa1s6/joeNxrqozdVGuMJTUdEYjdC0Tr2vjBBdHBD043Y
u8TsOSxg47alDC8JWNZYMT0bh7laF41XvjK8a0TpfJxZ8QCcsyKWGUt9Y0/dkrYJHogek2AzQZWZ
PS8SLTg4zx00Owym7slxOTzgUQgFVEAgGg+zuKhT4XNfAa5Fd+2wng7RIxZDJ2BwPA2c26vNrfkB
iNB0+XTpwXX2tqpDoEgwnufWqVst6sunAeltDvugWsnjMNIdglGZ4J5oqoyYNZJnB7c1JaNIqS2E
yGMMIqgq9QJLQq5eSS6CnsdOwlQMy4+Dv1Fk/JUdBGs4XMwO1sLwZTDVbislGx7tD1x0AV29pryA
UaSm5LiprLXIrXi7+lVWX1djJwMIT9zVCaYZFqaCAgtCH7SMmK+fP5O+d7KXC0H+NlNoIZg86UOA
eVzyLzKgzq1C9p0YQPF41Or4AGd7EedW7LpEjrvdA+C3Kozpf70zDEmXUQXcCBGDrnLYObo+Bk54
+HvDikiBFG453xcdXMN1/CrybTWchjtPEtM0Kljjde95ODKdIBDAsW20DQOLZwfqtV+LmKTXg8Bm
/RORuEILM+N/anjnTaWD7BXbsxnsvzJwAZ/NRejEPUqNNavshx8nPoWtOoOuSvuifS8lMOW184i3
MtM/VOLGN41QCr0UVTEO5tCOztQuWLFYu1KnjjuRosAXLqwS1zcgxpXzkdspgCIPtsI3oQBkh38r
kDoqWTiEUJ2H/tyGUs+wMf3TeAXibpiD9kK8U6E42F93HPqrJM7e6zat0Jk6tvDVVz9QbaFoXffi
eZl9NCYvblO+4ivKl8brikjSl3a+gFqPKp4ipJVOYj0Pf0GD0HKRN/NqFva1HfqKQ4VXwgn2LPSs
vVjR4qTBxkJXGIDVxbNN3+4MrK7YehH1MpsTprZl6FVY2NaO/6YMWQfK+uZyI3gJsZnD2iTmwphC
37Wz8FxZk/cKWzDteq49nPQH3sDxtlgO52JpZHIe0zSLW7AFhDlc7CEXsrLsZWrB4ZdCyidP9S8z
uufLd6vZmitBRkA300lez7XQi9LFZGBxyenyqtKUpFWYrLBlatocBIAZqWHJ5YO17fqhowibwWba
j03wqyhzDHW8kcp+tlr6/IQGK9uH9XVDG7GLI/cGqXothbWfcOJfDuMR7s3stFX4NeHTzbXT75tq
ihL1btjX1hEp1m7zJcddjaZnFP93vlp3LZTBsTf2yguiU8G8X6PJZydC6ttIxTw311xdv+p2/ud0
X1H3uLhp9bR+WU8ft2n7RBbT2N/QBSTfOgh4lqF63Mj0NmLx1HpjjXeycOvUKHR4y5baDacNypbT
p6uzf3ODd2LQ5foQ7dUYMajhJvF1Cmb+fOHzgu1w0KnVdEE1RdzBHAc2YT65aLQVW2oHr5Bjh7Y/
QBLssgT/in04RAx3xYeW6NU19vqTv7/6XgJB7CDicuRNsU72qqc2a0H8ihtAU4MCXE+iP1Segu5F
bK/uG65Q/rO/Vq09V0KF9G7yLwjjd6zB7DacjRBbErjPNLQrrXdp8t9tSFz4uGsSLFvH9dJUt/jy
ciJ9BgDYrj6TRC7gTX87kAHypJjm/4iwTK5i9pEvi/2XcsGE/RM3zlnk8LDN9Ism5pg2XoRNFttY
VlZDUgKxh/KkvdR9e5GcSVrJATi+yqWfKlQKlMEwr6Kev8OFhpC+KBM9mwVBg9vCjj4ZWtPqn1oR
0mLXMYCPUQml65TTYJ+ap3M+xDS9/iAUwkN4P2DjdNEuI7nypM1RFNJkCT0E++xP+2Byo9WOMvPA
K3usfQfC/i++fVjQrUxCjpU8La8KxPFwWvczI40y6i2499YXD7S/3JXJSn7kI3NUVc31vsZ+c032
6duUl5bgRq3WWg+GWBWbqri+2KH1KqueEqo4LSbXikTeB8yG1tQJJqqmp8k39DkwX+/nLxc+nZEP
QXjyM7VsoGqeY0HtVlvwkpbaxp6oWPBpQh7AcKDE4eU3T4eL66eDBatOMMOx7ocqMW2kqcNkyM0q
7GaCiEseUwV9zXFNgHlao/Ixhwn/lqONK6aeEq/Skw0dpJJIXqZeZ+lgS7C48PfXSY5L1chFBM3q
aOV/hfswWk/JFXYKdg/5/KvVObgK2hVhvgVlkEc+0TJdv8EOrW/ysnkIgiZsZQXUzXNFSZqttCLL
VrL+pFoYYcKHzZcbpP5GoSNWo2iM/3tW27Dnqd88KSKY9Acexi+CBaGTMpG/nP9zGzVJu2k3DzAb
JtYsitClvN3GfKxZ5dLDq208I7Y/DcscodnIFwH2vxCOhdr2Pct/N/ESLBXg0/fQuq6fdS8guXhE
vSw5Jt1p61DhusYmN5gRlz2tyreGq0txd/ZylJrYlNhq82hwe3RdxkNvf+HIkpbgpfYIFQdl+yJ/
Nr96Pk/VJ2b92hDy1f8wNRKNlQJMUcIjyB8oip99Cr2bH9Ilj62Ox7hFgMtBAkQJY5xfLO5v1IsK
MZDNFmTRlxe7vLHSORy+S059Jd5ONb7QhzN1RcZCO15BLAEqjnxeWldD12TvDSFMJmCu+qEtdsJo
K9KRhtSUVKtKaXkc2Zcm8OvwlNnbJ0KqDBLcXQ72+gn6USIYxgRyBo9luZLM+/0olJorFKAMvvY/
AHUjSjhDfwdZOAFg7Oyx3/YC60wjxaQ3d6qxSkFr2qFl+S8ctf6PxH9rMph321OTNYrZZaS/bidH
glDuOosXmcO7+CBtMh8qcgkatPjA8RWPfafaaI8ld5s+KlOFf27PdSANtyQ1Dh+XCuRWciUcjdIk
HFTr1bMtSy0OBepaREKhnszjKn6g2dBQ02goveJ6xEz4CHmLtC0WnX2ncCIxQXWkmaeHDTu2s5ky
pum5HjcTDMIoNpG4eIpz22HSbmCwer/bIM5W5GUYGMcEP/gS3QRuO3erN6Fr0XpXB+izJpOzaawN
VQS9DQveh9tVyz1PQLvnPVyAdXeiWFamH598XykF/josYC4GgrtMBfh8OFLaGD+ATj9YG56CYVsC
zAJGDDlw7gOUmaaJbFEC6aTk+zijvRkcDMrZBaI14fuNE2umNzPOv1vLkZ9b1eU+GIZ8Mv0GbEv+
MH/eaGN8ZYzOs3gFJrhDrQ7xg0w4idFfjHCjvAAZOgHO0lJD6tl8OKB1XLvjVaCmHEyHyHge4oZB
RT9K4VSOe4Vj+1t0XnWq4tkAL4p6Stw/LwU1sVzciFtNbHsgiMo4RfiLy1LMpMuZgGRUxOME2bsx
8A9w5i40lPT07iXQtSxKvqXbQkdRF9Eyndb+4YfQF3RKrWLMNfWHuq57LtvhFuvZxtTpsinMjtpy
7nCdG9s9qwz0v2YJUcmuCUCLkPpTUujWHvHDeTbQxmZgltYlGHpOKpzj29U91sfZmDJzImTcDItu
LXFRwyj6cqhtYTrLBADxzti9u+FyWeY+L2k1eABiWpAASkblMe6258u8X3fJQqNQkpUdkpRp4JT0
eW9/dOhohqWbT4kRlgHCeDE83nBo/kJioUaeV9Tint7GhM3Puz/VcXV1259CkthbtVXpWBYY1iLY
lr5uJFyxMAyoTwH6jSivRp82u5ZfCMxV+pkI4zztirtxajCMQVR0AiVwn7N7vRl0FKi8PTDb9B98
VSOOj44upUgjF0rPHrqss1T2XmJvxjRoZweYxyBF8hKw0E9pl4Sy0zPVn0xttUXzJjcKMR3aaxIO
uUpEp7s8ajwGapMiJxm+a9ixcNgxYwvvz8ZCW3/YLPzoJSVrPRAxhkXCSBqM/O8E8fsX0eQFiHDY
5TYy/fUjpUK1bWruc7uzoVbwJPO+YkzfaRJZctJ9vFYLwD2avMk9iDitVzb2cyR5dPvzZkfy4hqU
Ch2jePwmB5HDrhq1MzzHh9dLMuffW1KfEnQK2JmltCQgYevOVPPcyptllKHPabNO8AmOCDqdDDD3
p8/tb8jkWu+DvtFdRRscuHcSkiMBjmepbbIr4nATdsCtGjAuenirW/mKUIZiJzgsOxjDg1FEbYjQ
dRtZD7QMJJuQTAj0EAwt7+ZOKuNs4AbKx8HChCDPEd/8CveLIpqAAOqdEPRYsR9WD0oBOlUd6i6y
WPqib/U+hxxfHGrC6Qt4BcQBTwF88aFd4VoJhrtoc0UyMjmVcz2lurEX9mgg303Jv2Zi+btfXbqc
TQS0/noGmhYpk1XNfP4dXd4B5sVdPdual01NtMhEU0g3UvKrP0dbNSHT1L0EchLGV0kcSpGMxL5J
hRUY45KU2STfKYdMrZB3KNuXbb7u6Nj0pwJTfxbp5rUXPHvixY0eSZD5SeYtmEMSybwQU1Y1b++H
CLq9KJ4mPU0gr9eC+eJT1PePzIhfaJXffzG+LbUPis6BOjTSi2Pz0NDmJ0pOcpPtQQ07d2Jv6y6G
jXBipnwA1f9szkwJ80s+BgDGrTFPmHasN5u3w9muux1SYoBvY+YYGWAAeWAOGjT4gM8zNvVlfwlQ
c7UkdXlabWlH5dXVVCOXIXyIQDvVAJnO4oRD07V/nzGjceJdPy8XvgiXV5tCISJ+cF++vXR5LFHN
KO9TP5VHe9AU5wzsFhpQIswMOoYFLWuWrVbiF1PDFcblzP1pHKOJG4sgRx3IPuTKo5TtCuNFvDsf
WBrFfPOW/ajMzrtdcZEz39Q54BHlNJOooW/orlGAYMK6W0vqvnQ6rAxz+rrDW0rO/cc9DCRLk1mN
vwM7pajtWxN7AVjM5qX3qq3icLT2hghlmsFvHC6TV/toZpRIX6ayaa3cD8Xy9+WfqXeZXHvgY5P9
6C2m3w7ka5l2DJJ/auTAfUHuaEv3M7GVHhgZWUa1oA4gv0WYmsNFiWCcPy6BL7nWOjFQskBqk7Ae
v9bwtGz8GHYZAVd8jJx+zLb8UWDpCm5mPF57niD3WWjN2iGAvNj6KISzjGEM7j+TI8n6LKIvCC/o
7pRqwdKESVPhY9qOxRDZHkYmAK4a4bhlv94Gk6DeUIqNMEeEv8/I5BpnyZR7Wmybs5+7js6YycBh
YEb5TMcfnrbGg7/aZUfKAekw2jBQrstawPXzRzedSyxf8K7kHPPhYSxO2SDtcbTi/xlxpEZoTW3S
SISXi5bW1W2iMczq56UkHKBM4N0tDR2tYV7I+6LFrSdwbXDyAkjYr6OvOd2BmV9WVEaP087tsKs3
wsKJcWjWCK5cqow7kJidajVTfPZqgqH22LBSpkmMlZMMqG2XlUHBf+rCFnwUOxvGbA/k6tLNqpRV
8kB8trnnVzcvjTQRSnkSEXOyaLjnwZ64j8tN9SJwmt4Ydom6PiRJW0c2Zmo7eabpD+O5sg2T76O/
RG9rjXI5bhsKDaBVFnzuAMA9zowOxn7tBk+gXiptiYBkzvyBWmX+C56B0ud8SwPHe5wQTyGbKveO
rWnVbW5dONABM03C8ccd2gYL80/MWuZXNrBIqGLu6ysgB+3xk7TEXq3SL86sBf3n76l5mpgA9TQ0
l/z3QmHW0H2aPkMn0J4BXHzTjnk3gP09Z7xFGUC1mxcbVJK0nIvXC/atElLES2ySSm+qiOaASHJ2
GB9vfGHf6EieFv1K8C4ykgN0NDkmR9OM1WPfmQQnda2KHO6n/Np9VsPUczauxCHPi9CsaNWzEjtY
gxGrDxyZW7NPf8RHbgH/D9y0Awc94BGJjY5gihv2o07IFvzKeeU/RZWsnbKfDsm9xltUJcyhcwRr
CyfOlRv3By0XooW7OQbxx8hSms5Ur33wtq9CQ/Y7PLQfIGB1DEzEIdOFeeMo62bRvnt3m9sq+euu
TBdOU/Jp/3+SjeplTm4B4+691nOfJPAhyyqq1ZV3UIt8ZaEyLLvRpTULdODqMiSl7zmr9dfohCEv
bt5KEePOpr82Xvl8SASXVbjPrJWvo4pJA7mcvytsxpIId0yhnfE1BCat4NoyghSirmngNThFoe+q
U87uE0xhN44n3toSVDqd6As4/7ygpHnBLfKy+cHhjBdqLSU7vFrOeleheUDOnt0Ihv1vhe3OyU7/
MHn2HU6nYnYw3TmUrdFcDoslOhaD4SW0nKFXIk+MYBYmXhIKWfhOuPN3rhHTYDOsgF8lS22Y3rJt
NNKvEAqgu2ZZNL8VCsCneXl/vcXJ6TU6VO1N/FZfJ2AtbaqtM8S/xSWwQjILI408ju1MupX21Jwd
t0MPDqzjAgIcDu4WGQTCkrc0r/YzXKMwkoYz/zf7LQAuBo/t8zGpgio4OgiSDT4faA/09WaZOsih
j0C+sutOtCIUXd0VWPq3z/9TmOImqDxjgX1QomoIJdPrqfdDoJDKmia6TT1iKA8PjnKNBC2wIxmL
WAOZq9+USgZfYTbVnhOGIwb/9/LuZfUNyNp2OtnTye9qyrFVLcBBIMYbeNB+rdFP1pp97EfSQ7ig
Ht7nes8q3Wks/1oiGrmxZIpQosr/Y0N3alLMRaxglrXMLjq1dlLHpE/s8Gb1QtqSfw2v7JB0bxmi
rxKyPmRtBQZdoalzylTB7YPbWw39UsVMPcBFtY+ARNXABdywAEwZUdEbHZYWCv5+mg5v8Em1cKRf
AS0EcIezTk0mdrRBLf139InM3nxk+Niy7itU3QiFmxheMF66IAFyaHCcfWVVapl3A9CwOj1t8c2w
kdZmrwuHRd4y/CRIJUol4DxWn+j/VcRX2MNQLZE0SlhWATLhBYK+h9dZggxYtt6Sytvh1c7DpC68
QGEX+mnSFCgmpx3C0p9wsEMwtpDY+ANUAvkUoqeuk0mhipR3UglX1VVOHwB/oF5Q8oS51fL84lxm
RwxlBchOTlOfDnOo5kH1ePBAgghHTXa3g8TFtzm9J+moPw/de6ByL0FkU9b/IF431mxvzytglGXy
adxgclxITFJaLoI6jIrN03Qa4nsBsfsJ7XOjzTaDK2yvb60nYKXcspQnnbZXquAz0ThgQofnusD8
LpsHhTOXjA1K7yFwjV2vGMl/qO6CWJlxj36XqQjlnrtDTpi8JxgkxnF0X6EsdKxLG1oiLU4L224o
QQKxesPPg/aWfnLKrPWVY88JlkmoP/qxeEtjbvLlKgry/qVievaMlNOrY/tXX7JAnBis8Ji/wsyZ
y73on+vOW2Izn/0zOhvev+xLaTNkJss+UStG9mers16euzIW82/rtPBl21MgyFbaB4PLwYK1aqDp
6ViyA9GQVkVXSoVrjsc5Ol30z2jJF1/vO8uf1H7L2j5zWVjekYoM9UPS5iDLAdI/SgNwZ2N510Yg
pSGuIGNfFg/NR4W/yuhEeBHgUBdi+7vXPKA43VVDVMgIOWSOSgjD9Crm0ib/Xi4y99ya/ADLpIZE
dBcz8La+jt66YSyJ7/Yqf3yZvpChspo+NGo7RjIPbli9nZ0+FRkRwNXR48n5Kf5TSRRuf/WSeQ4Q
pWdYYFWHtfFWiX0gfD/YNOZEO4s0qWECHHYd3Y1lsN1EsIRVYOtB9gd7gj5BiWpXf3Mkl+GeThLN
pujVy9j64XT5bWNR71nAh4OpfV9P00NHGnJsM8lGszg5iIHCWvUzP1m+0e5POA2QpvmxVCmUf4ZS
M6ilrA2HpDI7SSXr0frsBR2M/dxjosCEI+Hd42T6lKi9LGTQm6Jd2gIugtwfDd/ShkU79bFUNeZ9
WEVgl2MdX/jN4cQACheARCS7XkCyHS6Iqi4ogNN2HSATBUfYvc+Oxt3V/ku2FIDU65D/dxEpUXMr
+8PiiLaZL2AxD1HQAWHASWXmVueVMc9KsQDUWIeiEde8gU+7O/Z4V3bH3Yo5m1HfljtDsq85uFgo
xkacvmK/In8kE5u5tVgw8m5+SEZccM9GKJTpiOSrlTiNAGrCjPWRz0vuZaR/MQp6HioGDJTKyMRC
4v2xIdZdV0yziffJBOBo2/O6fauhsR1pWS1qQLIyDxvt+oYn6w+9UpmmZf07ASh+0CkrQj6j6y/r
vD86Fm0AETLBNOU36ns8SHIfPlQ4eBpaXluoK08YVsqoBcp6BM9m1Ec4xEcBiYTnCT1+mSzuvc+1
YiT56zUd46e/EE28qScvB+0cMHBJWtqWrEhLCUXCryMFR9s6z+K9MoLx0b/hLr/50N4HkMEdlAgo
6ZJxU4wGLAI6kbPQaXTcCTSAaJ21miuCEqxIwi9mR03VUNGicGYGfoLxikJAfoQ/KOra0wDmSIyw
E/QL5GtZ/VFEMl38nvrpSH0pfbxwHlRjhQaznazUkfhcLhoX8OTczzgPtD6fm8F9Mk+ZrMhBonKg
mZAzX7iDm6amfDiyBHt/txMl0elWNbN5XqDfDpXRI7NY8W+/pKH6oQ4KLsiUd0dI/4zKyJcIbhHk
UDu2rKWwsQZe8cr7d54KQKGOYPC6OgQqD/5NsMl5h0yrjPzDkYAD2/e1PhqlXCrLURISiQvpIVr8
eHVit8CQgHATHLIKrZxCX0zoo3036IW9o2zq51HJu9kMkPx1eq0O4jNMPOkXUUBLjY5TXjwlGud3
pB20dhIehYIU5QsvsLxyeNeo9SuvUs5elBCQsO/eAWaXxU0KvVJrKglXb6FWHMbPKEF2oHPUGN6a
KLFuZKcMJIcptlgp7UKp9rmXpqp8PosqLFfXLJTrtCavZOp8TqS9VvcT9srX2W5E6WVN4XXAQxRm
9LA0qb8yWrTzsC1M/m+sMfuGH/jZjWJ4UwvRlPd9ApNGk9DWhm4qbuyQhl6ut/VhIpGRlwgxlNo1
CUIM6nrMaDZ0GAzPEk90EffLQ9ecpi6vaUgF2JqM+w+LWSvFum5w8Cl4SnYZQpFu+LQHI97SkrdB
qgl/5GB43uYjSweUvOJ9hL0t0CDPjA01oH8eXL1Ac2+cH2xb2+nXBIYRz5I97vh8zWybs3Khi8G/
hL86lbPGKoAort5NPXx958a7iejjj3n6XGafOyU8KVixycZ4Z8Qem65QgdtvcIsGMEVxT9CG+2tf
LnCOwlJNFH4180UR7Cp8OFpgJO0Ecis7JkTSSX3LJaCLK3rDeLrWrTFjIrRp9eDVBKzWkpqtgQtf
ycRm64vlhiue+/PU+ceU1UGJO8BcFrRvYX7i1eJgNwMyCFhMaqfGgiZ9iehlI2tZ9/kuJvX1gDnl
N4CuL5od9MD5kBumUy+HKvyxB/G6vgPBEXDde5MvL4MtUhy2NffMPsuGCer/WTowVqTMmHXWxFWS
gRFSuiyXYFRm97hbcQU66ApTq5nQKZTMjwfN+XI4adKro1EQEHWlt7Sabs4GEvB/eaZgN73ceN+h
pIB8UU2ZXQh7zf0ZGnf6/0A+CrZqC8oCH5XoBIqDshynuR3Wa4kFYRPnobx5yA4e5MlR7r1ZUq8e
0Pq6jnuoqUVp5vyReYdTuaIvUD2ztToOVftdJnr9GantP885yCuOMqk30m2al8D4OruIfCdVhzuG
0kwU+fKHI3RIlTvNI7KxDmOTutcQ2uh8Eb3K03tr2SRfULxirJ/bSgOJqWKOxOKjfh5szR7Ee+zK
gxRVQwmA1uEPfcQWkEnh24troROSoeZS3iI+kp/UkwDahK4KGD2Gg0uu2MjjW9CvosWJBbcdrnWU
rLm8OY5gKzSwryWq+SqL+F0HfBk3QSY5VDVWLkrh1uYbpfiqls/eKrSRl70kQVdw6cTYX8VHM+fU
Q7XxGzJYJ9F/V+skBTupC15zryimcLcfXixZovadjW5ve+YtiFaPb7AvO98yc4ljdVR9iZZNqfg3
jE5V7TdBJ6ShK2ayVcaLOIWIAK4GZ/OacykOR8WifWGN3YgMmiPJV2SKYwJINdXsUe1KGQMVYpXl
0SPBCYsXx2wu3i/ZhzeZ9XOK3Rz3TWF+p1DRyFdpUn/dCK/qkejO/ieOiRLm2NPVfJAwpXEzVB/A
/X1Tcjpor+U9ki8MV/ezQERsJkJCLKrdCbb7NCaIic2W20OnXxTIvHyGTMgEb713UpQXv4aoetwx
AImeHtp591Deff/uqz+y+wHCaZ/YZKSxPuaipFupbr3IuNCZNt71wsd6k2/uhAukO/cQPwbnFAf+
uEgfSUDL8cDKqbmEaVAdlPMz18z89j7azND40Cr0zEUzchtUCSVNB0nBagzxsUJ5MsnrnrM2/Nev
QqIQsJuKeUjqcuKjb+sVb+TXCAMHQ04V/d+rexCwUSrqf8SKlxDGlCzRqUV4El3URWMoS55wPCyP
yuKiRK2X+IQuponHTWORuMtuoX2uhhekhpRb717DUjrLcWBO5JbyGASKdiacPYF1rhu8/8Kyj5xw
7648yPSvLW9DbiesVkW+h0tD3uTN/Htb1KWyaIbHcGABAYa75jBli7pLYJHMBiz+zT8Kc8Pswtkm
nujoNIV4NX9y3CAU+CeJItjb3czOZd6rFYzPDXx8G2agN1WXVKs6d2VOJ9q4QpjnymAlmuc+tGE1
jFiQsXNpQxF1cwkoTljpMgez3Yr7fk2Ss8lauWxQkk5FcDtmSso9jbugP7mnMfiTMH1M0uZThxN9
KipYIuvsvxzUsiooZ5YZ7ocxKaBOR+f2Ir75Urxy2+p+UIipXWKBVtmiBWCFxCTBJb859CRYCCLp
xqRp4RPoWvW7WRC+gpawGlK0LR4huP3PvVTo++UAXmUCaIBT96Sh0N+U5MMqdNumiBTIp34OR5/m
aE3rg7Aup4MSO/IFZ32WRYpquwsWHlwc04av0qL2kkPTUawIS4hpw3JSc/MOB6syrSEhpSZ9ioqg
ybCzKzxz1HVsj4J0NrzvLbO7NBWOWzIRaSa/X2HtB0pYmtU1kSlcOVrZkzaetxmI7AFzMOLElkIE
uvopl7y+dwP9x6HK+UputW36/UFTQu+aG5TqM81Hm1nF1+txJlugLqLxWJ6I61XJPO4D8kkcDud6
/QSiNT9Mbm8fUcW3i7dXWYxCB983HrV4cKurv6vR6/i97xMN1GTgc1ltLK7GfBxEwnHGBNR3ed+m
zsa6FaexSV6ii+mFjj/1aKE9smGvXA5sGn8KHCDWjKhpwZUMDnkseFeKr6jQM9Ij9lKSClLir5KD
sthhcPOIt3LgVw2khD4OA4VVPaAxOey01sZ6kca7OwvkhSepDPB6GP3OizjwfxxtOCrBN7//zJqb
mN8x8figtKytX+Uj7FoabCMIRXb3s5d2kJJRcZZZfSdH8rn3Iz49jyo+iDnIlHmBMWoceCiqbXJp
MTDLZrgOo+e7DjQ27nRaXi/yLr3touxMe/PzHjVKyg3x+544/Y/gCaPQI98UPL3t37B63Sbd9k3I
U6MOtKVyRsACfEBWZLI6pCFoZ9WISrgSZVIw06qGP1Rn3V8gRBkTXK372cFi2rXAWoXQ/h1nIWcw
ufLCPTiSg/dd+NWgkuOzl779Yowg+qyCctwxeoWSZWp87pCuQSQsYU5+GOkWZ4r5/n6EzaX1UIcz
23EkYgalOubJOBR9XGK9NZiLTf5tFeBcW0fS7yxa6A69k6oMDglviIDT1lEOqHcY3NIs26FvwoB7
+z7repMlKK2euggNgu09oerIzK+QypRKXmd0Xq9Hs/CBP547w/Ybr9Uh/iU2OwHpZinAuW+pXb9m
ou0H8idqKTurbvmd8fPQUib9LLQFsXVwCrCy31tSRF5Mn26mTWu3sbmA5qCXOf4QArWe07JimKMG
VtIvgRYptQupykKFdFsPzEbcQvdntiX1vK5i+2FXh5vvq2xp/uPv7AaRzUhUW1Sh6OhL11eI7CDN
dOO4dzTGMLHmDWewgN74SiFdWxUwHvErvdOFRtgniqmobQsyvXiiXHsiQr+G0uMl+vvUAOnsDQDU
DHhJf9lt4DXUlibADkakZBSNB0Rwm+Qdx9s4pg+eTVWc0aHBHKerQfxTPZ9h/wXPNKsRcBK22pfP
l+XRxa0DNoxPtaEEzAI+DOXV4OArHU+eT6ZPhAkQ9cemDh6XX+tRjlp3QcxMZ9H9gz3ZLMnF0wsk
JgJfCUMxWjgK1NWLoSaOiFZDrZYB01liqvthEEVw3oX9aLmQuUwj2Uq6mcLWeK1PKUjb1ukewxuf
yKUdy9ANrhLouNOdaqQF9OjvVqzN2WvkguUdPAASz4gx3RQNf3qoHjP23U1tqBPhqTvA58YVJbeD
WfKw5cqgrZoDw/zQGxgDtFNyTR/vR2MxrRjK4QffbwkE64+NChZb7OQ6Z8V+1QgKHTXhZOPrmsad
HovzVplc4eBoQ2BcDrLEwH+nbjvD7DztU10f/PPrkoW0V4ApDS93ft+iAY3bXPH7idlHV9rdHMS/
vJEvdhm7Cl3rNBXn1DdUO86G8wzrk2hndyPGPN7vsLtKrywkQ8nu4nJyn+wV8dzk1xFJefZ32wJM
nPBXokPB+0hbNMiYR9L4HdHlTXwK3zGpxghaj7Qr9hIvESkf57IYUq7yULudkqXj847YBxKHRmDX
afNwB24ndDlHdtSxTMbVWJXXTttw46PAgbVYfDVGEuemZT//cYhPkR1/jG3jKC6VxQP5DsOCCzz+
MH+aKHFs3vnijph9joYg+z0Tonquk/giyCs7AmQf1G84fYlyxUG3qo19DriuE7IaASsvrGG7d455
GLSuhq2vswaqVBU2uFxS7qayu+VedLVK8xR+jLca7hglMTd2XXlikfs8yJSiBRihvT8EOm0gqax7
KVKik/DKuuJVD5hSRZMAWqz2aLGpsWFIFdR19f/QJIrV6DpFiG2cDwvSOh65B0lZRe/ai6Y9K56J
LBDfkco5HI6emksaYNQYSl7lxqtCREaBRtqCt21x6NzIzCrXf/gydC+D0sjFDjsLC4rmbf/LNgSP
C3/83SZGeh4oNUEHV4cTdRQzKLc+QVjwYdNfkHqLyK9XCT6enz1e6mybLliSjiWSYxJnJ6mKl7pQ
a54V6DX0UcysqmKLEZB7VJsyut8XwHk57DC0vIkR2TUkAGfgyeOrFxyKEtqNpovRqd0arN3OUSoo
yT8PbISRbdm4VEvLcgwvt4NAwh8f+8NuGdxDTiDJrKz6vAsh+A0pxf5RxHcyntJYFqMjQd2dwrnv
IhWhEsXxgkaEFwWHVaBQp93SXGeuOmjlo6WX50wK4zj70M6zk35GuDFM/zMkO1LjF6NjGoCJaowo
nGFn83DCEqA4SL9fqyQp/VgIfy7wEfgApjCNIlflJ09KG+NWqD8gv4WZER7JxdJOJ0f29RAPGlmy
MeFfwl9+yRWcgN5hzh7qs5xn87RuLxZYKrAum4sCyKRrocrdVMhXshQEP4E63JEbXRxvQ54BQAzH
9FdfZuIlNpJi5wKo0z0B4Fgi6Fq2L4V996nWA3LrzuvQGWZqAP5XDRgh3s4fASA+A70TPuC3VpE8
Nh1gGVKMCWpTt2NWKlctRSIDem3f5LXk6FfwNJmS6F90F/IHPDhTw/Cm8U6VHdcAxtZhgJJsy02f
eOKb1YzmCmTKosF1cntHKj9dZh2yy0zuT0S7/x6eAOYHSEeKG/AeLMekLfRHefdDsQ9eHWdS6m/Y
TRNNg/q7uJjBoJ7MGscQaDdIbv7xr9k7tuc74cj94xMDSUyY8N3EO4u4+khBn7kAK0dPmUalwisz
+CJjEpsM0bUj1HCffEyqdiHBnu9/iqvaF5i9rDyMf8fEPnADExPiVww74ytWYjVD4QobrXkzpOSM
tNsDJ6hz4MkMq9tb0kEoJYly7lPbQ/j7PcfFydnP2G4tO+f5hfUQlobCeakpaQsdbKc1gY6SwGGq
RKWReDARj+9uNzvUGvJfRroIm7GZChVNw42ZU0I0niW7qzlAlVUngqmtLOBNT6wgl2/BDKDRYf96
7rzbZJtEq9StMWSdZKZ8j5ZK5z2q+y+HtP2PejgBC+Rnl9iL+Ug2DbWtiT0MGO1D9dJGyDTQKH+f
N2bJMnAoHkxKA6meN0KE42b0sAVFTOp3/Df5Daef7WZi3cx3fGl79UWBP6G+7Q5L/VkrnHetDnE+
4OzlE03iweDufuhhRIwp9F4p5Ua4/6htCTS+55+HpLxFxyv6att3fK5+XJmSxIpqw1fW9kZun9Ry
44ShLXfIjzb24aFBncpP6vHyIVXdhhTCC1trmlpsZ8MMC0UUAWreWAYStvIXHNDuNgbp8C+HvGDt
0Kh1EX0MWOQkHbzOzsOPzjGybOdYlqoqAEFIufTVC364d4DJC54auoSebi8eiHB05Q4j0HvBLG/B
qYXiEtD/GqFhfIsZGkBuuXRP35CVOKoDa7lzQvhz6EZ1kdjG+izHVf5UolKDY9gahdGyoFKMJJ/D
MedCEQoj67nGZwobQ9H/pOog6n1UlXmo4HbRZNp6ZxnEmift0+/GaK++veaqRK+dmO+AyDm9wayW
51F1vIyrezxWe49gItXmt/DLVwUb6rnnBKtdHc1m08vBuyvBwqnDK7WU33w/rFN43Frs0nNsd8uQ
gahGcCAWGRp0UkBvbA//0n75I7Mqni31Rn3E3a1T+WBsz3gv+sEa2GFGmbsvlIKTkhD8X9U7aYOj
U2GoRJ/eZRFFKhgjdPps3jg4u6YwyLXtMhU0k69gPCY9CW81WJfyx5rwPZ5NZkZ4cMW+omn5OtSA
7/tUBnJO296p1aYXORDTVjheCHpJEibCZVPajXrQUJyagQEEWI1aPLi/DdpBSmVKPs26VwS+arVv
2ziPi1ZIDgXEK0XAdkvNe5NA+RKJK3YQHGMBsCLPFt1l1CpxBlGhmJVK4W/rSMAmNvIDS2qISE0K
kErhIOxrKwNU1smRJYtnzjl/tQfr5FSZLWo/CEK0/1Ik+JN6tNu9O8Omnn6eu0bIzO/Qe1naFgXS
kr9zcZU0p/RUYf3kZqM74wjL+KJaZ3qfs8T9mdd+vA9+5WITMUmte5BY2OYM4SG7tbJ8p1V74j3q
oRWVTqSLnQjkidqcv+O1cpUKow3K3FOq/l5nzvahIsKxgnIvyDRwXtHR9XahnvnRlaN4YEz0T+SW
TG8EP7bJt9vAoGtZ3CZ0jc++6blDxtTEsA2ab8GGry6jNbcJmAssseDL3n6cbJZFziq1OVymxYe8
JuA7xaHHMV/TMrsOHOHpS3ZEforVUJx2kenVeOQddpCTnQjedYEVBRI1I5K9h7ctq8FECPlLtHVt
zp7dsNdqxthJCplTNq1LbB+DR6xV6PibnecwVtpByF75EIDtYr0zN6gzyQCAqLV/CQuj3cjVLK1g
TFM1/UmiwKv23O1VKiKQ+iU1A2vx9OJH8XkBDke84PDFA62qdvE8TNuUG5UHbqogbuHhrOuiU3oG
yrfy964xeDK29D9/dfbgfzxX3COcbFBDOwSEI/1Dz/4SmuYsAaLEmDUy8hv5Z3AfGNfO4KXjiSv5
ARiGeJOpiURrVn3xjVhh4/3tSVEqn7xMVq9+HyJrERxK3MwgJU/7cCziftk/selXRlQrvvL/anTW
ns0q0WRDJUihPvFXHF8uBj+m2cJv/5hhcHugDUfy5wy6Ahasoen2YZiixO5A5+txlJldnZzToBv3
GS6PxtJ6uS7wEPU4XKnYYkys/yPOwNCzbqITvnPePkWgAnV1BXyq/LkxXNSU57zgolRkLOZKGPrg
A5wyn/2VQ4YP8+P6icgAgI/vX/hgwqeo6w5xuGCImch6qbHflRwW9H5otri5HIzxwUMBemAHu5bQ
NaCt8Xf2XBo1ifyDIVrRWqcDIjIwx5linnFwMhnvXOabzUXMmSOrK2Bfi3IaY/YD9LrVeUdbHBBP
dmF8lwdzHHzGtYRCChfvwnokdNprW5iXnBFu5dNxgwpt2XoLM3cWRsTGNWi2cgYMNUh079qOPEES
LDi8vplmU7UZGaqTZ57hE6mOch1eKENDBUA/G8G1H70TP3OREi9eVgiT12YCPpLMu0ytophhSIRx
lAR4JzQ/8UkOCOYVubUrEHYSvC0Xrk4nEFV4x0Lw9TbLExbCvuMaW6XAVm7WDSTEFS/NUgQ1cYHo
2fKwyu7frz2L7USgn92TTUW1oj/8nq+1QVFuHo8hZLKayHwBn2xPzvzM/uOpOPj80dF9CwH6xnnJ
ojDRs0d1PlF/LvkQbmEaC2mJO/MhssBRuthKvYePOlazPDCfqJCM4CvJXLJ4dMyjOv1rhV1iSdkR
svl0PLxe+gkcBqCdrPhGka+bSBGI4aHfOo5PfzGys9cZdqsxZvNzA4gmqwMMgD2OB1ySTPN2FTwh
Rv3cd6fLw3c6ErGbkE1WtH8wJs1zpyZVeVTBnxUC43KkV38RMA85bcknLJZsU2p6vYmna0q/UVtD
ST5BaojK20MKBd07utju/IUJgbKk/KDojvsUb79uASHzzli6qTgM67oim0wHoardBS4oA+YNyVYZ
sdC6MdeSSs/xTaxoTz9E980i7zO4PXc5XR5a90mkJgTMNvG4M6NY5Fmw6U9zW3ibmq+p7dBTZqK4
sHI20F05OOy6HsIZiu9Uq4MvZcLRppxRxEwYc1/yPjt6sxyEgkUrgZ4FJdOekLT8S66PWi5gl6qu
/uL/e5T4Oa0KJtwQHkL5jngjLIvQGSkHJj6PjyuIcoh0dicP+hP4Z+Y9uhXX1GbGb5OpmeycxKqf
ENh2Wr/ah1XCDfH9buSKU8IjQCZrV5QKdxaA0qGNXLsojJ1weE1Ee/U8PGbFrG83jXryz9s6KsEz
k3b/X9hM6BxXic44XTgz+OUheK4QxUGaz2GwHScFM4T91PL4ljqbzmbMOcM/eEG074rfWxMt3y/L
Gn3/7JZ9DEg6JasnKqU86Eieas89pUXFUrtqX0AN2K6YBWGf69PJsbNsPHud4hAfoQeyAtCRsGrM
gfs8rG7wuv6aVed1wmGhiXnNyzUDy5D2jmfWCQKEegdPOMnxyvyE1tc4Cxt8LSD4svxhhbyiO8Mu
mAixwA6mvQn8NlSS/XA5NWhKST5TCWtvySsZXHnQuj/z8UEOA1w601VN9ezvN/dlkj6L7prNBv8h
GhH5GEJL/tqnWMupaOQaSUo6CrifDIuLFj/eMQqsSn/GhJrBdbZFziJOTZDiuV+/VxGlsHt3C5ti
vCNUiry6FZrKV0WKeBl92YpURDruheNU3iIRTICh5FXEuHtc3ci56K/rqunLCUVBNm5qQpYGwp09
xirL2mpgVsZSJjKwZGT5N7oCLlEsHiZl+F5qBmEDiZxM12i1WSCiJ/5Bg6V3Ut7BcnhQjwdidwzM
7Bt2on6u+SRfjrC0vqjr6qXWzql0D3ElX5Kn5IqgwbhZ8SwfmZsvMshf030JOukGKE2tnxc2hY5w
mmjhNdmLKzg5VUtZP1hnZGcr3/TnuvwckHJaBUIiv0t0xDtv+ftP+mD/YURWeWkF1L2LUtn93vwT
kU9jJcWzhKno3QW4auYK+EbwZEhb+9aheaM6wJOdnKg+9jXO72h0XEexbrG0xOcIggyOVCU+eT5l
GMluMJhDcR8/3aYYsN+xrATxYjYjWdi3Zkil1Jdl7otec9SLTB4amLrmybMIuUoF7sH9uIcLxVFT
4yOjSZUIDJ6omS+vd7vyv6uS6rsW/IpBpU9STDKsh5PDzE82nyxzyZaNzQY5vig4+WHUQ5KJtgeD
KFanOLd3MlekCO1RYXJt9M56yf0HiE6VWGS8FutiHSZO3inPSqqcBuAMeNnczZY1cqbZo+6EolUj
A4mvmDedR6GZrrC8g5WKZDbWWw6zGekHCMIY0YZgP0T+kfRgkqGfnFQm8LSsq1ccwquNdeP5/HCx
0ybpFUyHbhZSb30LUpUu/8sgvZJ3bvl7rugsQEkJvlKXFjz8E+skXH/8LkFCipG4RW5SXglAw7gl
0JldTlHJlkp27mWKNUNYuKmeMbOfOWdQe6dx6+ZfHwagSua0pt2B9xLPqSG9/2ZG8fwFPXypM8g3
RieqAxV2CaDP+hfrBvUpblYEV/53Q9EPvB4lrythcUeiDjpO9Z8DAOkKJCVgBn9ftooCHfadHM8c
Oc3VACh1xizO973EfKZyFJz8crTX06xq8fRxG2zLl7WzHoMMRiWTjy1pVA4gv/QtTqWNM0bPJSYs
uFuY8BGT/KWXUFkvUVaTPVunByLhIEvGUS6EYNCvxXP6R9UaIi7rkTnfx9FuTeK1npgCOz5hWXOq
9M/dlfa2Q6T6ui+gTJCM8XgNjpujVBEPbeajAYZEj93t7ixpuIqoIP2MlIsiSegk7eB2RBddy14V
8fva50EOFktanzAMJrWhcT9CqF3bI/2xDCeCr7z+TlVTtXTSnuGjTWhK3hn4wBFHou+ZCk9elLPl
L5wgxsRr9Zj1n2//p/3up/0vztQYDyf9iv3LpBwKaC8p31yF6UsVh/ZHgEBJDI9Hl6MM4hAhNG0l
qmx3zKomAb21Nn02xq43fMSbnjrpTAzngh6k4oj2qEwaAfXwmLKAxiEb3RmS1ueBgPwVeGmFbe+W
NdxXxCxru73PmXRSkmKM3tnPM9hA+gI72fdNUUdqK4dJXbmiHl9uWxCkBwGOJMykpo/uyvLl576G
X1ujG2Uo/AFOBasAuf1ZeN8qHva85tbChzBj7R7olyE2m3jTwnJxDKKgdc1hx4wQeP/7nSFpQavG
uLpUNkA0QBLdTd1h/X5KHUm9AFA00/VruOJaIMTwql9AoHv3aDHfV84spNKJyZyfaIXTfs6NpL39
7AHleWRuph69o5Q3gF5uLp+XiwxKjuHnouI8k7ILYbE0MS4a7VecZMAJOXnFvxyAJGIG5MQJTdoR
RdGqHw0tz4JmYnosKn3d/I0iMlUCNZQOE7qu5q9iruh9QtvzJpbT8g6rAVfJmbheQ3OVRGyjb2wx
xFc7yCxsBZjwGPTSigLyUNQVwTKaijAinTs3eFfOhkWgvjhbHP3z30K2SJUqEvnIuDQssNYd4kQF
SGOGu8bNXAeBUKJ/MvHJumTu/7LpnvjNFGrKNOZLzHw3W/5anR+8qGwiBgv0Jl9nR3lV4cnCylBk
z5ASYeid8T8jJ45vU61NRlcmBH7Px6wWk/6TeiwJwAuX/fUFODsftnjcsCXN4dNS680p/QXAGrA/
w6odFvikDb0Dk38WAj7Ia7gFyC03jY1bpWZVpGtDF/xaqrcAaimPJ6ppmEDiLFbKOkxIdtCo1ibG
gCmtIUU7YAs1ANzNDZ3wnMMdBQtdUj0MFCvpWs4wzjCbtbtw/4SlbLaxVL5bkUGVXFXF7eq94GOn
N/sxe5UGlNdN8JuBLQOQFbuVt1qSPobFmR/Ni1O7zIpqZCnYAc/oC3vpKVwXQPmnOTtAkwrgBaML
YjREMpC1iU/tYNuRqmdb9uDRIqR78mmU2GVYj6ykCiqtAbXmROqaTs7XJmUu6YA+zwfpNrMrYm0X
3HOWm5TdNENLbiyiDt582Cg0VUuKOiicMIuPEJI8qU+BACqxE6At0UuJWj6k1ruxXnAENuoCBgi3
FzOjkGcQ/zKW+6Ljfazk18chqaACNohgb2K/LgKK7aFIsU9xsxLrwckCFbae6fKrZ34Cth+w7bM6
IUOY2jPngU/R141uJyf0Ez71smoRNiutC5j6awxw58lfHxQzAWYUyRbmybecI8pY93d/ChDyYiwL
7RqL2N7IdEd2i8cnH2NxS+9NqdQ1v/FUsP+7cfrQiYmcgAsq3tfQC3/gChDy29qRrdJ8wt/BgzPg
PWpurB0KBVw/GaflYPVW0AG1FMsAjVGiyX4hijWsqX3k+Mrj97Bgdp+tfjPHdetMJowUOpbO03Qr
iB5xauldAzHShr91GkG16tzDidN/n35bDtSBMeS9eznT25ahLwgCKl+FRVgH/jxgtfizH+CkYUyg
DJqq5Gc2gTpWIP+5oL197/PdgXCnEivkDc01o8MzdH5s5oW3AW2zbOy7/meHciUi22mXQGKRoli6
I/+mWsdflhnY2eKivI7uW6GaFyTtoXxaJ8e3H39Nq8kXG+Z2iDdttibRzT3SjaIKp79jwFQAGolt
qby6AgdYX8PEdY4JIrOhfr201ohJD8jojBx/waEVWTKNUIImaQYIOcjjQbf6WJf77SCsQpXZxNlh
Pn9LYUHT9/C+NzcQQ7Da6lrVMhtM3b+OkOfSrSSWjgLL/bmL3XoSgvRdG4Dn6QmO0/jVf3vs8c//
Y4K02TbfzKFxXgoiHLkWOzoQhk+BBDj3ULF3A8HkEb6FeIBASMJ/uEO7MvacuqI6SFil0VrDYywB
uRQs6E4ju3KrCEcOj3scW5P10qlAajcNSsrPQQ3WBiHFocaUhvAYc6nQjpO3Zv3lxWsIvkAIdIAl
z6NPwbSCPHhOiJHr9VzLq+LhHDUdJw8KWiqe+PVfBRNZdvSM3EkuZxaRR/q5gzwnKNtTEISy1koY
OSwD1mlin5KrynDwehKWKrWBvHyjxWNctZweX7eygDBF4Tvu4nvxYOhy0vCVxmlTWb8wPy6ZGWrN
2Q4JkclDCrjYjRv+CRVnwduF5WULGAw9bfDwsgimcFcObyeytGamFoa/0dls+syPPBmM5DPbxcI0
hSUvhNkyxcKIf/9tyX9GwtJkP3rghB97SUCiEJxVJ+/ochNgNXifn43JUbtUaZQmANGB1R1F7E58
ejArfECrIPiCPThGcxawqafYYz9t8K6vTynfEQBdK4HCgE35wKyYG30hUEUg6oXzMZW1Occ0KX10
ii8foUzTxEzvSZZpDHzczJJMIGAXZhba53wiYaBb4Dl9yQHnhx99N8csVajtYUcIBG8fK4f13WqX
phc17UM+2Pjq/eGOHXmBSkTkyryRiyPiJYl6bCJs3cBlWqc38IFHvi/MuUfF0l9cZzdK9y812H5h
OmxNKNwJA18DSFGkCZT3RP30v3EuW87wKCbQUE8Iy58bqHzrpvfhVUANw5P9G2EeMhRguPvjc0D4
hd8/cIojrLfIwWKuZfm6MeGDqUcZ9QgxWSAnOZIM7d5pvForykFPjpLYcfiTNN0GdBe4cWFVpRfA
w+6LTX+6cXaxmXP/2WxHFalx8nLwYRwUt7drMxfnAUoZlzwiLHe9ZhG94wcPRg8OUR7PVEDQMNz3
3R0CYagi518/PXPsgsD8WHIEDQjB1BXHesXXqLH6UV9vvUhO5tukTWOWtHox4T4ZeA2ldm0m0i1Z
Ow7JWnY5mi5/K+S55/Lh9shYkbj5uALAYFEbIE+OiIWEHufOnkUwP0i3QQ09KZRDT1uZY5bMSxJk
G2N031s2Q5rSfpGI970zw1xzNN7RhYRMmrtMm3P+aKZauWMsrnebrqpzTf/x/6ouw9EM73hJfJjE
oYdonP244G4xVRarT6d5sh2geXiRrCFjpqF5BeBNTADwRYPPOFzF02IGt2z/LwHJP8EIHI7PoApN
2rlMh6e5IGib0eAyTS+HLPRaMV26Kgk19AcSqoVaQEZvZw2Fc3N7CcB98wWPUJ6ZqjwvD2Phwmny
p3OAAVmxQSvFS4b8m3sKG4bzjwOZx/8mxhoONwFAA3o5lr8ij/rRzfC7AHSsBDuAq5EnM+fUU5p6
XY47NskBwlAbJcmWnxH4nTxn6vqwVqkoJRo/tag4Z0DGZngwND0JVEzMLyUX+T0t+IUV0MDxgM9S
vJKi9RJatnHX/ZYWYCfHJQZ4G7rV330wspAfz3/MOtdmeEtF84tEF1ePXThXp422kJXowVDex6uq
oGPp9lU/6JkYvStXsy7PIPcBXAu7UXdy89lmFcUbPdEUnvythqBDiNU3m7zxKHi3jmCM1KTG1ZkI
kQQgYe7B/XJ3Y2Oc7nJjsjY0r0XeIyxeP+77L/XUJNL+Gv31mKYpAi06hTuk9plXgeObft4jwKMB
ydqUuNnfggImOSgNrd2OR/uROFWqpkQ6H/GX0MghxeeFPBHWZ7waTRgLAfDLzucmGXGErDtn5XVb
nwAWHfRFO4Z4iYhxHWwdZ1DabLYh4n5GiYmpccbO6NrIz9Pb7LiwBqcnWzwIeENvZuxsA70PntBP
0CNQ5jePN8KKd0d2tv5MT5VDDUFC7ggfEM211b5U1HNW3Bn9Vz0X2An3LgMPc9QzoFZlbdpU26OE
1ocugCH8IgQeNVxp4Z8nAvqZtvePioQKRJWHkBREvKY3Cqm55gipFNCOd/VTteL92VQoUDI+/hKf
3eaSwHok/aTxw9OzFmecHhrh+LaKuPzazTYvw/f/m1HWqziR48ogYbpEt9MRL2G8MhuiorkaiW7a
nu7rgDfDA416+eME/WLG3/mK1XyX0q70umJpSdJrylJwSMOePT9qFEZKuNx6zDpygy26zE/HHUjT
NutlvloHJdtDYBYoJ9JCMhDPHgJmunRcKz7n6PCeDidqZvvRbmC4LjjIkM8nQIM+X3R5YfWIwQV5
Ew1TatXjYc/597a3zDHcfi6MAOPwq5RR0zo+b3r1a7M1GbasyJgFLfNujfTDyI+yoAbFGc6jNeI7
m5nnMdeKrE66Icxl8psgEIjoHahQKZ3hBkMWUvixXdSqu7EOYryG0AP9OwT3ByvnFLlGIrJlhTBd
AtVJ1ELU2QneXqVnmHgRRtdIccH/p7WXvmnNyPC8NLb5n2UosTjKeZBzWGPxJTcAlk17SooUEm/y
1p95SwFiq4smbh1vVlpXrFM+760dAZz0rrUsjoVGPyEbL/E8dB7l7C5Up4ZNIuBjawisjiKbWvop
Sj//oBnLJO20Rt85Ngm8I5D4uSG8SjVOunIkIxsIPs+9rOmBz7p1Bgsa/M+zhOQoFV0roGJstQVS
CMPo2x6wFDINarzwZklr1hGU0AKp44/2/tE7ENmQA6GcI3rJgUCUUL/jUI/nS6/uURmotlakFoMA
z5YMOiJmCbkZvsKiIub0E3e6Z/HKCE+5t3tq6g+xwqCwgkphcsYgnZI6KJcR8Fo6qQt59xsCu574
uWQtKPFguLATgg1D6/AEVNUsv/JuMnmYMidUcscaXfki6FNzIh8xP66vVRueKgnWNNRSI/kQPjM2
BGOSG01b66QJb04HvSSBjLh75W44ncza8+QCol7GWQOzZh8HDkGT+kRTuVmY4iRG7PGliMXzBMeh
qHPP0EfIZLuCVDNw/mvIV7J8uS0frmHYHeY9j+85IZdMjkuBzmEE/WM+73qMUK1ppLePui3B0GLN
MTHr0sCWXbZcyzryQ/4Jt88l5dLEEKJhwI+HWCcSaP2o2OWqoDZX3XT7HI10Te77CE+bpmva17wb
j4sB3hnSoArwN8JmzE8sniJlrU5RLJHA/A4sEthT+LcTgDxXuTdvCWPqQgwZ/XTy19UMAecnjqJp
s//HpQuYd0jlgYIT3i4kt8RSH/URhGvyCa/eHMP6/1Y0ECqVedCSE9pJInOa4vN8QKMmatLtpvdv
Qpn2HxZi8BLY++VsiOZWwIr7mv81Dgq7sYhgFALXaem5So2JZXaYVGXiXFOY3nq7fVGCJ7+qw33q
+r06Q3I3WKJrhkNwr/5DLF+H9ykiiGr8xLkjrD7WtxFTCiaL2f+q9HxxJDn1gLvop73URR9o1x75
ycQgEFWVwc4GvDYgANF66OCGbIz7yGsC8I9uPab7rC7UIhW8Faf2DFghbn/kP7kGwZOM5GKHPcGU
ZScQUckaaFkpuAoteWMaDG5oVdHN2aMWvOJWJTr13/ds19NaMkRo6bNcASJT9Hc6BjX/tpOYFtLP
Ls7nW9QKmL67j39N93r+HKTA7czNIo5d0M0YjXrr66cIb5w0SSnrHYIolIabdODtAAUjtgvhfLnT
YtG3M+yAMGmOZXWLNoeGp6Qlf0uSEFxRS86fP5LGVrlmYGUZ0NvlyjXKpsayieIeY430bqZaW8R8
+Bl/fY1hQo2sGdlPysH9s2RCoc6SFML3WAkaXvORM/riCJGKl7Dfy+nfrZolwb9+wglYf26D5rra
ylZs/Kmw1RuJpxvuQofLDPGQAVyXPGQu9dSioGwU44qnjZUyyTKHMESyMmwErBsOoDlupqs23Xos
dXSi3j/KD5az3KcxDDZIxI1usxhSQOux4V8l0KV6my4JiAZhkqsXXRGmJwaQmY5nHmYjYKMdy45h
F009etNsDzDlsQGnJhZP8B4xrCNRaLkH+o3Feb51TsJzI7rZL6vsWLi61bAFnkUSJ9ynm3EIteBo
8QvTqUzgZxEQP3T6oEhcxCqagDpJCWRSVhrjgXAv5NvRZ0OcIVP1ie9W62rziJ26370uzcVas+gh
nFur49AL6AAIr4nU50XxdBr+o+KTZQccqmjQA2/a/QBzYtt3doJqEM0+UTTRQoFOJie+LJJ7QJjV
fbj1eUZ9nvevqB1MBvYoW/eqO47CxRYgug7pq3r4qBjatLVpzp5LTaA0LOXRUy/PbuDhDsbgmDco
/edt/WqUP4VsSwOlwbhXS/FL8e2BNHv9C1d050CUNOaKm8vEW2ra0oYYuRuhvaoRL87Ldp7ht++Q
3WM5VJyUiePa+YMpmAxlZUvx4tMyJ9cQyG3hTzYBJtr/aI9CVMMBkEOzCX+Fgq1mPPUrVZjdoMOj
dDZfjIRp6w3HWQ30pq/zYtz0FWt38yWAmZNDhr7+j98l3qmFju1ujTepEkL4UeF9LMKdoQLqBy/0
O9ZnMhEAeQXEC52e45xVAl6GOTTgLnnmPpJZZy6Kgs/kIco1VwXzw3Foi14+zSCzbkxK4GNQtwGp
AKR9ee/2mOkeirhZ5cOupGf4dkoXuyn/dZc/QRRUntYr+25n4k8FA7/AxjoX6XPqcpS+7wt1wBy8
EE73JblP92Fa2GHPCFW0+iOGSHMe2UFuBt81CikV0MruANQj+7O7lq3C2M4D4To3h0EFgFkWnlec
6GqRogE40kL08WskN8rQofp99mbZhZnwBlV3lt4KwdEgZcRuYkcWW1V9bfeUIfbJdemohT7hun7n
IAv8RELicuP+A2R9lR/QEJQHxWUC7GMs45GIONztTBgNpBmkSMmVvx/PqkAxbz0vLMpoKIktbShd
tmi9gaVLkhSDgvAcVJgYX9IxIHgU6N1J85+II8fDyPS3Pkbsa7/PHhok1ej/RWgWn2iuzcFE6+IA
TP6uaV6HhiW2P2UPUFUZR2DViwd50/g/Al1B305yrPJrEs3o3xjmuaMCU1Lh8OQmYilbUrruEiDC
Usc49OqvV2KYqexjqTB7Sv2idQSVzAaORCntK286sugQzxdSuXm6PQLRq5kUmJ+47X5/Z6r4KvIC
m6kW1wdn1En2s4b2IjTkrJahWz1vxM0dd1BzZmM9n51QqXzrpv/F6OBFM1F8KKWU33MmovkKUiQJ
DwnshZLMtE9pNefdDGB9A7c1U8VNxKAvj4137zJhAtMOAVqUbk//sK0KeaSCx5WzviluoYhRCYUT
GYs/hXfibQjEYeWKp6i0mblhiBmMtVewRn9xw33wfZ/VDJVYCCmubRKFUsAcV5aF/W2RaBQejYNo
Vu5KS/BHgv1Sox2xXnWPOzo1jMboS3JCWpfyV4DA6Dr9hXU/DlY7FcIl1cn/lMuFHxplJiY2hQ1C
zCtnb8WZ8+lytWGiGfvd+NRPXpfc5ChSZ2ZyqmXlMwCMWOblq7P/6E2l0wGcXg7WRYl8LLBiorGV
8FO7Wkb9Bqb5+qcePPQDjWfj5eQOGSpFX4OV2cdLCwyNpLauT9atcBmpmmQplupkfpcdbQaVar09
epZC+psh9/6Zw/OnDJQHK4dTkXnwFBbZTLk405fym28y7hsLN9dwqWkoLwIzGeXG2UyTmFhvhRoL
ah4Vb86kQ8K0fd6p984TCD5q9C8gFsUpqn6WwouQLJGTLst+QVKgljAXWhF1mzXFqp1R0UrfRmsQ
yon3bAXiNsFl5y3O7PvJwLH1YjRTA+BOkuxnwsH3QvL2Vstnn7i1Rs8rPWvdCTTuX/GQEPF+lNNa
Vqcg5O1zA5QJwTQt2bKnRex9acMR9dqnHgDCHfG3+UPrJa69+fiEqwWFnO/UeCXnfAi38Dwg5FeV
bUc54vShZo7jrFM6tMrVQRlYkwGtvHuJYVxUbGB/YX/OwBSFyXlH5q8NdauPv4gmP90BQbMj2SmJ
WerKJmZHCyHQcgkF2uzm0EmRruzEpCX7guZOFK1wkIyrajGdtpCYFqBUUd63KugElSU7YUz4amYv
xIQcEfoE+TGiEEYPzfavjgLlgge2NXio269ESqszJgwbUvISKhfCjKLmKrtuOPUddnyhtm6HCnL+
d8M1/ZAfLwdGHu9UKTliDf2OgnojFV35iRFh2lBXFyjeqEVOVqRiWuCDDKCaFOuHcoHSmVFS8B5l
Tivkzcu8iS4pVHyCwK/yM73UaJfBHqVECk0/RCn9IwfXhbgHkC4bImA33N3TTdd6GqmvX4bcqNry
CUKHuLOUjG0zvBIYE9mUVTlhXo6CIMlyMKsnnJQ9m+tB4QDKqvxX/tey44c70OSE1bP7owghLROj
7JRyeQ5aKOMvMl9iVQb6KBJFRI0DFQlLQBaCX3QDoV6CRAMRc8RLakXR/nrsrBFkwyI6Mt/R3R6L
MmbQtwwdJg8/IKJmk3EwGZiN0LnfePFKqLYsSgrlbp2zGmF3zqaXSHedA3uDQbqTL0u0TR7KZr9q
xTWHd9CminoiMyU7hfNNBG6//pkcqfbmV9NX312I6snQ1+k93aqxXrwJtubGkXQ1bSi8DExW5r10
zUbXqrdkdrJjcMv3Jq8y8ZViiXrnbps2IYZ0NyOtqCkkY3l6PNLo09idc9f98WE6qrcb4vptsnvt
HvQlg87gr2SDOyNZ+kbwbjI7IwlmcsWuNy2Yo48rYME2EF1Yh6AEyVXJEMjt6E/BWpfAdU5n6SCq
IivvvafehSW7uOVC2DkhjOAdEuXpHgZ7NkLPtyO9AFkZGIZwSnF8iMgTC5pOMx8jGM9WIHPao6Ho
twBlSrI6wUkHo+SbBU/C41deH9i4pjTL4xZd1R3JLJnHm0lt/WbEdOmQu1NmLGeVTa2IOldWmRr8
Cz9lpVkiZnDmvfYZ0SCecukuxK7OSDbqCGo4CR2fuK9L/eqVP9VahziAaDXtK8tIcKkdwxW/mW7r
rAXO6i2ic1817pMj0MyRRdVpwEZflO5Hx4GRWr3w6fnf0Me23K5fYVVlxwXjfgM4NGtDPQ6icO39
DsPvyYRgp8YJDQQT5EXpLI/x5W07l/PnwGasYX7+Q0nTvJm5nEwxwFKhfPbfc9b1cgE39y1UTZ9f
orZbE++po0YCnHqQ4IWwtU2VnfMhY/3xGO8MTdfqZCZgyEZXpGuVE426SMgQx5dn5sArJSPtrkDS
Uuo1udWFmcH0sTytSkPq4iEXqL170RdXv0s5I+v41yDNNbR5zCF1i3dT1H3+HnqUBR2vaAQv0YXv
/8w68jOfbf84FmqjfDbHveuivXBTMlVgtKAYTMwSoM0t72jz/3PlBJBlgEVDRNZ7TK+/IZ7jXGk/
mxiyQiKXE2RZJRuc7XqAKX2ElRkme5hjYd/PgC8ks9DvQ6wZOjTkICzhrh/ax6Sr9ncntZh57sFN
xRwSXRCrfNIGC5dyRzASx3HyiaXzLINW80EKlfo2hOthiXTLbT3RUQDm7/GTgKbBu06CBK37zcTi
TQ5qne749+KpIlG/Oxgfsq9rwzM8NjOLmk6KGs6aG11BAffP2wqChqRlseLURtHyM99ZnvcrnVHk
/1/j6n37vWvDebVr35jlpDJgKqpghO9zfuQshPo1lV7hspzjAheadIKUGjpDblSw1MrmsM6Kw22k
BRpYLg52zJozBaCaegHkRYX28cgwrdzSngGaVqz9J9DhylUAcbxfvuu1x2LNi/Kb6tYVxd142q9J
PMpuBwm2ANDcZ+JDPD5EUe8SCCNYePT+FgDvFoJHY//vjcdD59gbV0UoroGa4KGfU9U1XiQ+KhoF
0NTT8kRux5xgVFZxb+N0wqb01xkKzH7EzPqCIsUd7HEZI2fVTmzry9/HcMyc5l5sn5oMLHZKShGS
wxqCx/c6/2f5Ps/9VBshN/gzWwGvo8sieIM9+2om5Op5C7WBnQCNPUqKRal6WJWqbo8I3DdOs3FF
+llz9HulGYvQOInonz5nzZ5APGkmWgIv63qEnL+CuB8m/sEefJ2QGws/RuGmPCXvSKB78AfZ2Wct
r7O4ehn3Q3GhUFH7by9yxqrR0MnoFMSFFlC/cNpT2DE9yVgGNKOstAxSjdDQ9Y4zvDuazmMp2aCZ
tWrIxUOxt/YvBPmubKcukf4ox3eF86u893k6NaQxIJUvSKpUcFvYB1V5AzI9UV+O/ZIc8rRywzfX
qIG7Q008LJmzxX29SI6LyR9aAY/9VaJoPMdzMBUuCDLFSFA0X4dldU+22TWuHsgM8JNtNKhtymU5
L7qrYqyWNQ1pYByejPHPk/68nyijmJDKxLV0upUES20KcM+oIluGjY8U7lfttxupf2SUgKRHrvmU
d//qn6v2Y6mfy8foviY80DbiQ4mC6G0IkjzXFSdF2vN7iqfNzDk0BoFDUCn9/tXisgALfIe7LvwI
IdbuDLMpXOpgfmwvQPhkX34xbA/rsi4XYlIVdZ7b+o8P5G95oStjbS96GhFcxCXHmqQ5snShODi+
qL6yKwubFqFo8+KAZ54kOyMnMOmNSn5ig2Ri25LfHNlYuzLawG8TFaeJLazFmNwA6mYebddxbxvJ
Gq7qzQJ3ZCx1cRPRiF2m+ifra+UEGY7zVvxsX4zzGQVZ6l7UOjaez/atqawXLRKp5VsigQFiEjI8
SSBYNHBIPittgkUddciPyXklZCoT22Vfv2uEBXKfN1Li/55A7D5+ouSldA0L9s+f3DbHLTzz3TLq
WkhkKNivWN5yJ+rclv2VnBNO3rKjqq6ButPDBDckwDejoGqU3pV12/Q/sbaq69eNEjIra7v3YiAZ
oPEFb64g/qS8m7fm8ufGXApuERLCXb/6I5lY8U/LCGh4cav+RXQjmbXrO5v//A3fi7BfYuMf/JLW
UYtETETPQrZFue4xGgSpnMFa8KyUvdTqur+m+7D2jZYDNQUOixkRsCwRXAs3cJLACdXp/Yj+LtjC
HCtPj5Hbf3AAmBvgGM0Uj89rupFVl+BBWeKIbYlLTA9FctYPIeL72JASD1zgPCZ5tEzIQKYaStJ2
J2pHgwqPr/Fg01XfQHUtKEv2fIAvAeIWlJhD8ZT3rxoF+4xR1Dcm00fqoVHULwN+Ktr4aR/OQ+bG
KHQR6DkeF9fXij7NTLmL18XE8klZkBfrupyjdYtrw0r7CRSEa5iH4eAg1IxJb347h+g1pw4rAH1Y
nu0vM4U/iYy85oLEr8B9Zy3JRRKPm8h/IUUt8o+5rQpdmQbRDzuiuOQjovomAhhgd7b80eAhsHEn
R45Yv+DXa0a8JInaQ3A6yrii1pYBfyazw5xDvx18UdGtyfVUDDBJ8Kq78fRrENrdDK6P8Z+NUHaQ
yLOtFRNHBhxTDRbbOCkbtAo6jqEASzhlzpjx0l0tzOxEhnAKtlwfPAxZAFrE2oD0gI0wa5JzPXBR
VF+D5QuavUJMLUbYe0hCwCIy1qSyS6/hBgJ/6vMaTZoE7K7kwEdAY8M+gYJgBeXkIlEwRHMUOJCS
86npOU8VuYJOcS4gIaMeeSLV8/ungzMmcRsNVuahV9PsT6JhImknyPrVqikrAbksfLCuNEj0elRM
2DLV4CjIeGKTpxrrONTTn8xenzb4uYDWMc9NTXVnM/HMsDbJ/GCa9sNRpln+3pvHbCb64VKLRvhC
Qt889ozbZLcOJBdyIyjXkVovSBJC6KBbgmMS65EHUBwQnv1Hq+/jutbpXUVxlUZhzGOng+11pKp8
vrZALp7EPkdsvs5slRK9awwikibNjat4zBKrhbuiwGH/E0i1DtUEWmOhxnU3NqRJ9h2/n5Sq3Pif
sUumN2+APHpmG0+kE4x/gUQQX1bkyvFoQmsVfdrm1zbPnMqVJUtxNix896NR4V//dpWLKiKT6csE
HZw+lU4PAQU1xJEPkopa4Wv6NF9JLRtiJulmzav5cQ74vHt2K2dMx/cYEcxLaAJ/zRzpRCHB/uDb
OayQ+inqF15fVEMeaKVra3u/s0Z0XSzNn+4ELLMHk7531dYfVjM2ntAql/109F+cI61U3wxeHVfG
ud5FVKENYHemMlI1C7yyAnPpvqqdTpHJ0n91quPTFf6eZGRGxswuZA==
`pragma protect end_protected
