��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P_-�^t @)��>�{�<�M�Uj�2�0Jf^�7�_�A�;�fP}���Xnؠ�����S�)>z���f�PPE�:��	G|۷J@>Kf+�>��s<y�$���a�.��IѺf�J��2u'(P6��mz\�Z��H��iQ��5G�z(��6��'�!ur(���l���P�?'��EeB{�k��6��~�6d�Ҽ�-�g�̿�b�������H~w������=�q��)��rE�Y_R=��f`W:��9�%�+�V^s�j���0�ƫl�~��hЄ�cq�n�zG�� ��"�����y���ʰ!yX������ �U�aj�,�E
��:ziO� Mm�V�@0��{,�X���O��Nk�9��O�!E�Z8��
A	z4#�(9V��#��ͪJ_ #}���y-[�^��������*��~����&�	2��݆.���p� K��=�_,��m�^ɑ��`ѝPd�����2����c���xe�yN�z#p�%.{�c����X�@�+mXi��Vd�������җl`פ��1�H� E� N� �I����}E�,L��!�XZ��M�[+M���'�G
���N��;dO�q�X�s��������]G���+�	l�U��g棽�k�p�x���������hҤ����"3o��7�~�h��k/�W]D�����n����u�o����S���/��
�#�gרR�"��]o��8t��&_�ʽ
��ڬd?<�Ӱ�|]�>e^�G�8)� ʩidl ��%�G���-�ո��h��$�|O��p3��M��H�7U�C�սq-���֕�, ������2�>P�Ċ��[��[�7�Vl24���sC"��{�,ji�j"U����~L�!؝��G��1����ph�i�����@�����	d�h�Ŵ�
oc�
>5��e��Rs8�W��/'�cOWa�P@����62��e�${\Z��( Y�O��b'�w��A�[>|�ބ�6��r�c�Ɨ��Z#�:��s(�!�}�����'I�4��k[J��^E�� ����R��g�tm4�.�E0��NIY�;lJ}M/�	YY��M Ż����{��Eб�:��6����t��}d�L/�ڭ�N�,�D�Do�<�G��'���՜�����_X��]�X��4A���b,;�`bh=��Fp�5C�}�s��rlTZފAs�d�d�Q����sqK�_ q�l��;	o�I~��J{����Mh	(c���&�/��)`�R��� �m��~+�ݲ���
�N )k�T����z����]�W���'	9Ӵ<զ$CT�Mw��ih��󼿽ʐ��j��9L����]��H��@�\�_�Λ�+���D�x�ƨF��ÛG��� ���٪�P���?K95�[W���n����c��.j��a}>�VV���='��2�"��!������,�$�x�-/���g	g��/�l��!W�j	���d���I���k�g i �]hɥ^p6�e��DN�4�j�#Ĉ����%��P��0A��;v�D���T�v�/p�'��B5><Wf+�w�fqh3�O����i'<�6�/H��4�RȬ�=�DEw_9����J2�ƍD�b�EE���Z�SnwH8q�a|���X��;W��7{:���ZG�\�0�ҹ�s�=��IR��i��U-�'iw����,H��� �"� -kD�M��\�o�ˈ�S#<�W( ��KM���	@� > t�F=�	t��36�j���Nn��(��"�!�N�y`p#����_#�F��i��!������o͂��N~����ޱ�gi��E��ї��-*҂A-�~ˠ��O��NG԰�;=0#��=�M�Q�R2��.gbr�zu{*�g�&'��q�mֈ��'����Fl�߃ʥf��LŦ�_��܌�P@�����I}�h��x�i!y�Y�����E�q�>I^Dm��ApW:jd��}�s�}��gE��aI��I����T��Zv��!�b'%���sȼ�5(�i�~IܤSK0:�%��cY۳��a��@^-����(p�Q��DV,Ό<�����B�*���/�%�������s��$�R����3�}��=��霉3������sZ�ˆma\~Ʉ�4�_	Z��>~ǰ ޴�˛�Dn���P}�}`�64�fg��x�%��O�M@����y��7����c���18fq� ��%hVM��;G�?}LU���u��:�`�dYA(N�,1�? 4i��(pG��40ϖߓ��V8��`���w�s�U����}��e}f���|B��3��{8�e�`���f)b�J۷<�B`K>�C��g$	�Qw���.	��1S�iw��u�OXxf1�VvC�W3V2W��Nu@�|eʹ��<~AU��\���/��#�����<zN_��"E�����ѩ��9l��\���0�nL�0��;$ �0P�R	�K�y�nV�\k>rQ@��pt5�=T��d	|^��%�Ʀ�E��r���	�i:�	�J1��%$�G̛%�����h�ċNW#	�>{�{�vy�_�ԝ�鼗���⮟b�y�8n�v h�/��I���Mu�mII�43��Fת즎��{G�
���	�q3�4��h��.b�Cúc�e��:ぁa�`�:SO��%O�F�]l�s�Ojƻ]'w}�!3�h��jeI��C��?9c_yn�5�f�T[�)Ք�-�k���t»�OӦC��e��'�n��v��[a�Û]2Y#��%�godM��O	ֆ�-10��<�N	��,J�M���c}	�SLu���+Ю����"�'�x�/q���.�} ��#���r��vϐ2 *;�Sh��o���Oft������!���T^:��6��~
2��a�3���&�rs0�/w�]��>*p�ڸMί2�im�+��9w�E�$���A�?&8ګf�7(�bG`�?�A2��񂄟�d�wgs��e�iB���.�w��H%��R͆d�lj���Z/	�B ������!�ڋE��������d﷕z���W������K�X�����O�颐�?�9�&䪡Sg�ꡦA�|��Oի&�qB/Ö�>a.+���#1���쬈܌-)���,�n�$ݜ-Uk.&��������31͚��U�rgD$k�3�YBa V�ّ}1�22p��wr3;0���%��^�E��-S�V����%�H�?�
@[�����S�&SB�R����`@T�KI����I�M$kP=�$_e�F*��{A���V3�9�F[��f9��z�;�`�q�4�^AR�/�93�ih]����a�F��fRr��&�����=1ŏbm��<ub���WF��R�dD|�9�b�;���������Ki���d�ӵ���'9@�vR��q�b����qx��y���t��@F<�6\ ������4`)�o��@
cr�rx�D����5��;`c��{���WV�1a��`őPW���Ă�Sꪼ���H��GnENp�÷�C_W��U2_sD�g������*`�Ƶ�3I����<��cʣ�a�#kb�&f�L^��O� ��aP��+�б����Å��/�}(<���KK�&�.��qA�IY��E�E�>u(���]Q|��c������.H�́s5u#I��f��t���ƔPI:�����-�Po�g�OV�%����/��`��/�}Pg��)ev�8��sD�i�K��W�ed:���T��pTKF8��Vχ?#�d���ŐT���� )���`r[�����j?JډcO`�<N�ψxǳ��qa��E��a��*$������n�ՊVn
C�4�����A�R����g�w}+���\J���aL���
�r-��n�/55��+�vp_�j���}VG'��z�'W��ϒ��
�u���;mXYz�k�����#Ă���PB��+j��8S�Rh�` �,�l� G��x���u%��\���}��IA\r�*�?�M�Շ�c����$�%��.ߛ�-M�HBh5�A���h#N=�02�9Hf�~&V�^�/� ;���3�ƌH0_0�@� ;�9u�[�(��r>��jC5(�k�������T_��bJ!�\�Ļ��c��?���c�z������ҁ�f=�T����:�px����kw���)(Ţ�c�Ͱ�RE�Ӭ�el��"�9��\�K\�Ρ݂��[t��@�y�8��P�T��)m�Pk;�H�
n�K)�D������w�}!� El���_"�4��s�Ӝ�@�8?i�aF�b��PYӫ-(�@}L����\K[3����9��ʍ�h��� �\㗜iQz:�q�(�Qͷ����x��T��de�u,Ї��2�c���uQ���D ����ΰ�lL��S�
��� ��R��u!�c"׌l����G��WS�`�f̃9�:���<��+�,�$D�5��Y�8�!G���h#WE����}��j�*����fe�o�f��E�!�o�y��S@��q90"�z��ڸ]��G�qO�Ax
��Nܴ��g`ꭰZ�7#^�u�<��V� ��M�X����+�"��3��清"M��_7����\��(�YP���Lm�@���XE9�t`�q7�����F$-��U�!gڪ���R��;�ů���q4�|YM�B��H��m��'����Uy��GvHv��.�*
�%���9����w�Y��f�f��V�<#b�K�
j6��}���n�T/�C�΁�wNXݍ3Ad�r��L[�8|��~ign	�=`�R�'�� �6]G�x�cQ�=���`b�K� �*d�.D��6�!�έ�s6TԚ:B�)�pT*��F*�=�t�+I��Q|�Y�,1�Yl �V*	�� ��������<H�'Q��>^��4����|�7�5/$�����(s�Ә�y<$f0�¸��}�;]��Ffh0���ՋZP�t���u�}���s��Te���Ս@1����c�b�d� ���v]O-�td\�[A0��E�a�N��lhD*�Q�z"��3r�Ys���Ph[q���fJ���!{��O���^�[�Qk[�
rm%��O6��A�v���"�9r� F�M0�b�Mz���o�ʅ��z��	�[��Mn�&JS��$Y�,fӉ'�xy?!�mv��A�W��?��� _��i~-Ke�����XJ�����1��k�)l�ٺ�*�vrS�'_����Z��qĵ�l��	���}�*XD�M�d��J <�AUo�|��^�#�p�A�Cj	
�H����4	y
Tނ����פ�n�
qp��^)�l-�q��Mw[LX����pM�ڜ�J�f�����Y
 ��T�x��+-�'!*�-?qv�b����� �v�{eUj|��h��� L9F�C���f�&H��(��ɡ���
����y�xo�I���?���6��s`�A����e�w&�y�7�V����̖̚�������0��ve	�֔^sS��d�*;6���EA[K@p���HJA(KE#ae����TT�䟬�H�s촾���ô�A�6�g�M�����
�P�k�՟�|y*��	'��z��]��G�Ee|����� ���͜�EX��;���<oW�
'q<�����Ԁ�;>P�<�b�E���q���Q��"3��eC���V��L�H�3h��~�C��������{l"�ǎ,���4��[f��a��Dg�C�B��:�u���r�W����9���ow�zZ�P�x�sҤ�����(K�0\�<�Ľ1e��L�T�7 ��)��Ἠ;���ǵB�8�;�X���/@�_��?�.R`3{F}w�L;��U�'F~hiފb�����{hַ�a�|���.��`���&<-JC�y�GtC2������{���u���2�lyp�~l��y�;�r�����+����F[6ARs������>��{e=|�GS�;ʰ�zR��U?���<��ܪ�qM��w+�`2j`�{��Sn�S;#��j����3p�}�+� !?�'c4��[�W�iHz�=�f����XʹK8��j�c $��q�|p�Ã�e�+�-���z��؆�iK!S�]I���"/k�}p���O��|pmK�༄�P���,�b�pU�s�7�	�+�;�z7����z4059��z)`͡�G�����8]!��N�h$G<)w�DWB^��Ԑ�ٛ���7��1��W�8A��� m`������Z[FV|'��H�����=�����H�H[�IS^H��Z�U;>kE�'���i��e�\�I�J/��2K����jO	�oaO#р��	K`J;70���]��>�s!s�ĳ�u��$�,U&�>yq?��%O�h�neFt t���O^� �wD��l�v�>�M�)*eo�œƣ$|��rV	�X��pnh��ؔ��	��9�ъ�"�Ѷ���&��L�o�F���w��X��V������j���?N��l?��Eg׊7[��dM��,�g�kB{Y���Z�vF�A}8�Ve�pe�)bn<�;+W�-rmnxT��Xi�+��p�}fq&a��p<B��!�(<�	�B���>�j�� ��d����}򈀅���-�i%����x ����j��]ũ�!�H�l͂1&U�xOS�琏�a��kp�k��\J�j�-��@DFZ�Fw�2k;����9c9L+���W��7Z�u���a���f��9V�ڿ���JX��x�����4��/?[X�^!���ˍ���Kdp<W�򎫑�����J}�u�&���Hةm�4�Y�h�C����	*�e_�!��N�U|����O�HJ���:4���,]W�o��T|���=F�@c�47ϬB#��QkU\���4=����LS��ٯ^�w=
�'��bi5.�]���w4;�͠�<���VZ�;�!��Ў,ZB�� f;�w�wv�5��ёqR��9z��H�L_�Ȕu=
Yy�#���������i�����V /�XL�|�沟���$@��dA�	�3�ɟ2����Io�l.�W�bo'����d�V�� ��Xԅ����a���*��М_��:;nw}��ĺnM��;t�8F�񝫪Dg%M��D��\0:���L�T�N�ԓ`�:g_O2�r���,2��]z�90J}�?�S���<9H^w�w�
C�,S�,?ӓ+C�`��p��y��ׁ�PW�y�=ƱK؁ Xa�m(��3����n����E��3�R%H�2�mnyWe�<J�	C��r��uZ������(!F�w��jIP ��ni�� ��s}h��O���\�a��5��ցK
#Gt�����Geo>��g4��zsz ��E�.yE�9�b���}"���=��zE����P��+�\~O���6<��aN��Vf�.@�;F��XO3��2���ce[��c�#�j����@�AI��e�QP��!�*��\��8�뤕s��73u�N�c9,�2D����턋�.��0�Md��*����b�Җ��d�X��y���P$��
osuw|o1�-��u�v���S�hHJe?KB��f��uJ͒�*��K�WV#�>�C�?���ҷ��l���F팫��'�~�S�h|~�M�8xYt��<ئ��i!{;x��#v<���o5��E>������bj �\�|P��FE��7�H<�-��^�4�/�ю.�e=��2跐����=dD��X����E,��}ZY11"_���˻���vVj P>�e{�ϩ揷��3�H�l�s���xh��ս�>���{L�t&j-�,q�"RJr[ k�)�,s��Ӟt�ubB�����?F a���*� mz�yjW��jp�M�C��;�m��/�O� w�mq��
�*�4^4 ����m�͆%~��r{���
]0Ё�v�Z�[	/������b��� �&�rH�f_G�@�ސ�Dd��'DZ�������so���`�ٖ��)�l���+�+kOg"�Oq?b:�	(�X@��HZ(�#s������N{`��)����d<��N�u�D��7Od����_����
6�wlơ*�<�=Jɕ�ID�qDQ%����W��iO�%���K��i�(Q\o��Ь����B[�����N�cd�y�����n��
dQp��9��/_��*Ab�iJ����M��j�����З�9hiU�G��c���D�y���Ny%ا�8g��s�J{F)��Vrf��5$���X��o��'OVG_�jڗ�O��M�t�CL��7�A�d+B�6ҝ�nO����"�����0q񱺺|���f�
�ŷ���p�!��SG頋$l)��2�C�������f���������8E�7 Tڧ�VП�f���`��S֛:�@����o�A�9��ֶ��P#�gŋ�y�*��m��kJ�
-C>=L/.M'3� �o�	iw^O� �[< A������nf��l>��O
��5	xP��8`j�E�73��1k�ܼaq8qf~z����1��ry�L�mI1��=��������d�W<tD����	~f�6P̚�o@�|����"�zK����~�0v�W2m�j��ѯ��'�e�C�/�����8���1YD�&%Sp Z[ȱ��w�ހ�y;���T��	�ò�G����E�ݸ�)n�@ai��
Q��at^�����-{��t���pS�T�,��h �h֥����>y��Pp*�<�bP+��=���_���||Y�L�����ݱ��C��.)�,�����
�����/�e�&2>?��\vf̢�D�\H��M�R�u�����-�j��v�Q�x{㸏�¹�(4��龗��vW�Ak�<1g�ؤ*�N����_��H\��!���0�9�*=��S��T�G����M���y�C�x��ς��Zo� �t�-U��y�pc6'kIc����'*;���=������D�koX�"s�vTؚ6�U9x�,(H�(pJ��M�!u�pU���x����=~Q�<|�}@ n�i���)b�exd�,�;��68�F�q�r�xM
6Ȑ�#/�M��|)�w;�5�~)����rP)���G�G�M=�_�p<V*X2F�	Av�G��k1/'�/ZE��.�go�\����7��ok���c��0��~N�"�gE��bá���)���r���r�m�.{>(����GZ/�#Ḓ�x!֐�D}��� ��W��eUBl�o��!���`�n������k<2�E���L�f���("�Z.P�O-2��0���U��g�N�2eAL�����)Z���ɲ�Ya5�Z�\�M]���B�ufٲ��A��8�IP@ى��u����8�l����L�x��9YWf���0�$�i:ʢu�!��[��m�^&��掳hnHnyc�N{������b����3|�G�]��g#�ڼt[�ҷ�A���.�i
�0��k��	'��ך���:��`�MQ�m����?5� .�� ���diS��Zt!پ�D���,�):�*�[���d�֣KgTW;A����cS�Lז4��D��ZD���2k�l���uc�n�$7���Y�������LT8�� ��+Q϶(��|�]�$�p2qw���<�*��0θ�(��9Z-�;�ĉzi'��\M�������=���������JȟNքSB���AJ�m�V������h���":�?���5�ߘ�f�J����%0����1��J��q�����ܬBX=�{�܆��9x?#�����O�MR �$�'Yn&ABW��~�!X����U7�g~�Nn#!����L�kK ��jW׽&&0�O�$�uY�,�d�Ʉ <[�:����"<<c0�?���Pհ{g�EXaU]���(���}:�V0F�9�����D�i�S}_u
PC{��t�4JQ�����Ղ8\`�#:m����gy5ψ�U�3�Y���#H@����u���
K�T�m�!� 5��[`6�M���	�>�޶"u/�WzyG�v �x}��S�Wyo ��a�ƠK�/@7 �MB����D/h2����:t��m�]������3&��!�,�xX(#ى/�W���{��2@A�0cc���܂��5�h��ĮH���eMl��`�-Or�Q"�9t즪Zj+����������(���p�[U�����o��X�>�2ڐ�r˷�p|��C4�we�d�����Ɏ�ă� N��	�����.xxCV9;e�Z@H98����Q�#�"������﹆�$�$�K!�Zq �.g�R��2ˬJC^�]�0���j+ϐ�o�W6�(��@��M�f`�G7 �`�{���$`��m��O�M��]��4���IA<LHE]!�x5Sd��g3� 8�7���C�2�w�cгặ ��Ul6��$�'R;4[k�^�[�w����Ru����C�wWm���(l��vr=	���x�#�l������res5��O���m��α���B���.���$:
�E���!뀐��h�fB���X�i�4��V���8���Ǩ] ˷l�W\��R�Ws��z^��Bh��It �#�L�2��>#���g��󈶻X��
�[�� ~�l\ĺE��ZnY�!�hcd��!x�+Y<ۋ�'��4�k1)��Y�A!(����ӭB�ŁP������z	�>].�u�3��h��Q�"y�ъ����2Yƍ�;ţ2�!
v��3ޜ&����Z�!<_ iRG7����^�]���mQ�$H����:�7��)�h1����5��(c@e2��,^AX�P�~�to��h@���L"�Qh���P_xZVƢ�dێ3��G��4P�̱ݟ�g��K��l��� �H�Q�brtҌ9|�$&YЮ��X�Km�8d,�LL��Aߘ���h�~��FVQt���`��i���!Բ��M��t�w ~�Y��hM�L�Z��c�)1&+4wm:�	�
;큧q��7��"qgJ3���Ӕ��@[����ָ���-��b�`]���~!�×&���ӯ�h�/4��r�m��`q#P^R��]��&��A�n��=�C�/zk��7�'H�\���4�Ɉ)�r�g��~W��w4A�͛*�|�7r�^hcCd߁.��^�����_<��U����~�B�$*�&�SPzP�)�k҄
"��6{�3z�zP8��~e�fv��r����q#�wU=��6��e��`����p�^6�eW¦�VU�5T���]bAS�﹋h�X�@����x��a�پ��_��ppF&
����8	�Q$Xs	J��aѲ�2)�cO*��p~M�(B.�`7f�4E��
M�z��֊=z����Ʊ�ߐj*����-�S^6,�8�������g3���w�T�ǵ���g��󓬭s{R����Ⳇ���&e�u�$\�k53���溕j�'����v�e�_���Vﮏq\\�<O�S�����;��a��G*�Σ˛<�W5dw��$����kMZp/������x�Z
�?�}K捿����HP����ݽr&dÜ�֍߃���bw{���ծI�ҥ�vI��{+�M�t�2�ca.����Ely�>��Ǫ�Cf��� ����p-_�\��x3�i��ǣ=\9:���,�9=�۰��͆jױ$�a�4A�B�Ӗ8���s��ͤ@�Ɍh���@�b�%�����c�U�F沙`�g���@�T6��]�#�/�w�s��:��J��E�c���(�.w�FE�={gޝ�ߠ�e��c0T��nآs�l]���X��b�
'Q�g{X�#�.�,[*x�6=r
p�dϮNo�ˋpOR�����0�F7d� ���E�߿MQ���p +��Ɏ��+��GS�-ѵ\��N�;i���T	���y�2�~b<Ɇ��#s�I����zTl��J�S4�9=�q����0t�By�8lz�*qi��YIt��2.a��ѥ*����O^ֱ�Z䮺�-H�}1L�
Qk����3��S&�Y_����F��J�/��'�- cr��xSh����%,����|��8����$Ȃ{�:ld �2�mY2u0扪��_@�I?f%\9��#��돟�)�^^�t�|�g��^�p|D�΍�I�����Ղ���8IB���M�e!���;���D���f܎X_�[����;��������51�X�^S�q�P⧖}�����"#@ì��vG�ڶ0!�LT$�׏J�W#���9������9+��Ui��̿��k$S�����漃�����( 
�+�h���	U3��S~M�����	�N�[PX1`��bj��Y]m*���3�"�9�M�
W�ц�KFZF������>-	E�8���Ƨ�e
3�p�0!WӅw�b=�n3<�k�����Ve����6cv�Y����������%�MR!�^@��$ra���|&Q�	E�A�/*9(�K�" �5�ڱ{~W��+�Y��G8H�^W�[P��k8�Qa�� L�%=��~�	�����Pnj��W����}뇊Qk�S��%��GQzJ�ķ�hY7z8�s&5	ǎ�	&�2k;�h�������(��v?f>��影���M��.�6[:��9"����B�+��-ų,`(�%V�:ЫXq�X}ǐ��$ț�t�{�W%�}��e2��������5���q���7����fI�Ͼ�7̰0g.4�a�0׶���V�NۍZB�ݾ�[�GP.��"�2�z�o�J�Ҹ���~s�m����mT``�X�8Eˀkj���3��r��9\�f[=@�����7L�%:S��)�''�l�J�z���Qs���y,IۍL��9\��/@вк�'&�|����[w0贀R ��4`�����}��Jk��uY�CUb�2��n� Y2`�n��-+� <�݃vX��z��ϫ�����L�y=��"�HV8?:�5>�,'�%�ȃ��QeK�w��������%/��l�ǐ�*��G�\Ǉ��O�ˠ�!�ہ���H�$v�� 1�8�Q�#(���_��܍g���)n;��8ɵ�Q��v0��ix���zuL�b�W@Zo���"��?�W�ٙHP���(�崭����k1V|�IL�j!2�9��:�[����\��/Knj�Q�yv\(�?-�i�����% [..��L'�LVB�G>�a�y%&Z�[j��zx��|߆�W��Ij�n�S<�ڽN�l7���a'9N@��wq5���w��{l0'��5��Nq���[�����t�4����}?����"D*��4.!���xj��l�K+a�0�-��sXJ�9,?cy�-�Z8~�>K4��Yk@)��NXo8-.t��Y7A�'�J�����U��(����q�'s�}���J�YsL�*�R�J�=y/��o��W�:\0��[��D�^�R4�x�Ji��E&�a	�9���G^�H2�Q:����6Mb����'3e3r��8�����+�,po&����ǳ����v��
���l|!�k���>܉O�)Fq��I@��T��n2�x͈6�.�����9S=
~(W�=���I0Ha��Y���6�p;j���Q&�kv��+�n'�sk��pvk��p�*	{'������Ëd��b�����B�|`'Gc�>���Lݡ�Z^�Q^�5��I:��9�E>�k҄P��M���6u 2��:��Uwh<K����hbڔ��k���I�։d�f�o�e��_���ȁ�X���(��������Y{��z)��A�x2�:0p�̀�/�8��{�'��W@�l��X<�O����L�p`��'�yʽϘy��n� ����&�4:{�/芫���<�������^��������rȲ|@�ۃ;����6��+uxJ(�"�[�b�D�wbi����� �x�Q%d6��Vk[��C��5�OmC^`��C�&�j���ُ�7�ʬ��f�~x��v���1��>�4�d�oR
n#���� �S�aB�.�"�0����_�E��V�?��fU{���EgG<C���\�©��L��Z0����o�C$�R�Kn7��� cl���� )Q�fg�bSL���^�߯ƝH����+��/����ۃM-�y�	,P�r	�K��m9Ƹ��' ��n�g���q5�5)˲��A�s#p��0/`Uj�O������Ԓ_9��z<���շ��r�`�+:�ʖ5�Q�,wr? ��X��S���A�VG��הp$�!M#��X})2�w�lZ�s���`�!��e�'-N!�W�n ��ˊ-��zV�A&�"AS���h��W>�!�q���Y\������K�G@g�`2�G@&����|�-�l���Q�1��l����1�dH����<�_?;�Ϗ`������VЗ��~%>�?�32��&FlE9!���D���2�E'�B~�$$��ϴ�d���������`Zg�&[eU��&,lv��J�
iI�o?��dO�����9�~'�D�Ij�1�Z����Ql�rn�~�k)��}C� 4Yqw�_�N�����pፙ��^e��s�/?/�e�9� 8 ?Lu�,g�;�*,b��:��ď8��p=h�ߓ��	7���{�xv-���c��:���W.{�����$�[���"����e-�l���qS��LIF����3��*B T�,����/T��X��g��N��&�����w�b,�Zƅ%V���;�����2�%n?ǰ��"�ˀ��<�S��Y����PZ�|���	�X�q�d�A#���g��dkGBѶ��lŴ8���+Ю��z;|j��܄�����q�b��5��|]s�IJ�)�z�
�~u��3�����8����q<JMԕ�N�e��}�����b��Z��)��x>����O���w�6	�8y.!h[�Ҋ��i,<��p��ٓc)���(�D�c^�7vz��̊��,L�Vx{�;����$1���B�9v�Ǚ3-φb[�-C#�/?��j�ѽ2o�ok�Q��6��s�<���n�d�#���y�'�L,j�$����dR����b�̠�K�(�
��^���Rߥ��F�⏼W�an[�R'{g���cWPr=�唽�3D�&	�����Aj	���5�+U����� �::�{�c+ ��>Ƿ����Eࣨ~j���ZO�󸵕=Ez�t%8Q���-�x�;��B�<�~�F_��=wFԦ�4J:�y����$>���{J� '4���퉜���r��e���U���qy}�p����Yƅu8E�U�p�m^�EU{����M@xz,��KF�w��^�F�>e�*ɶ+o��3���v��e��߹����~��� ���.���U�;h��`̆��&@�˳�^/\��lB�)�(�N���&̔.Q��`���h)a��zF3�_%����A�����/������xu;��)��l|Vg� :�ў��H�X8�ϰ��I���Bׇ_jO��A���������ȣ;	�3Ö-q&BH+�%4���u�緬)�KA���jC{��a�Au��P��}���
�^w���g��֚_ڿ?����2����������Q�-#�,�N�,3�v����˞kO�������YQ_y�X��3
�ٜ�FS���<�3�Y\f�D�HC��6Ja�Yl^r�H�7;��]�����Cڴ���yn�����kW �3�� W��-�:����LK��G��i' ~�����JPy�:깔�,���ڧϔ�^�͵��#w�ڄc����Έyy�*~����T/��� VT�_�g	e��:u�DҚl����a�7zۼ�
�w5MM�c)��H�����r����=z[4h'���c`���1sm�>�!�F�^pʜh��
Ut��{���i�zrD��&�����U��^ST�u;lD�.�Op�������ZDTV<�ҬdB�*dW�Y�1���,T+�Y�7����"G���p��HBRزi�Dڈ���r%�&����{��r|�5��bh��h�3D,QK�f;	��0M��t2LЦC�d��)"hd��($~��H��>ݎ2����H�^(]�VO��>aJL��V,�%�R��C.�Q����cRʹP�U��9��]5{d�ܚ���j^�+���	w�N��d�p}����ͪ�3�&	��k45����N��Uϥ�R0��g"{�_t��x���ˊ�&����i6�.b ?E��/FS�wÀ�����ɢ�� GC�Y�h�	����8�WVz;"_tp8���E�v�=p/V�.l���'�3��<���}v�� R�_����L�������.�S0ː��SDMt@�쎺�*cS�Q�i�+p�b��?Nu�-�^®�v/x�`#���/�-D�u�9?,K�^�����p dߌN������)Β�
o�SlbA~׍���jxX������>�C|��g�v��]J�x�9�i�0c���xJ�t%���;u�5.����6�59{-- &z�{h	hR���3��̡��Bf���	���*|�נ{雃C����Us��f5/����|��C��E�����T�$b�M�r��Qz�sX��\��
ߗ��Jꉋ���ej\i�hz����{>RP��R�b��E����hq���bJ��
�p�=�%渰���b9E%ʷ���l��Dϓ`���K��w�O�Bi$!�D⇈�%�|�v�)�NFQ�A2�*�IC;��kUR8���*:�ZX�+H�`y^IP%ЀM��"���x��IG\�,���+�p�.���X]��ZUJ�깤��9�?����gh��.�Φ�Y��H�YC͓�Y�>�v�r*f����D��:�^�+�*o�0F��]$�zl3�<;�5V/�0d}v�)Yߜ��r��b�l�9g���\���9v������y��;;^�v&h�ܔ^W-�Gy%nj�ԙ�iO��e�]ʴJV�+d�~RW�ę9�����J^ަ�����6���SQ�ސ��q8�z]�[��d��A ��ֱ��I��"Ӆ}Թk��i���MX���ϲ�C��4������n���9��0r4�)e�����`؎�"�gg<O���i!��V8��O��j��"Ωkٹ)�ӆH����,˂�גl�����ց�A��e_qQ^Ozc��Xowj�w�RUl�&W�b"K,S�)q=cIu�������9n��~��i�'�w��_G�]��hOY���pe�UMTg�ܡLn��Dмa��7�(��6<�^p�`V�@�(2P�wέ5�~PV�O�T5/���(k��V2�u���,�F��!���41���g.ŝ��A�y���.���Ym
�P�$̑!��+ߕ��D��`�-)���f�4X�_5���o�ь��v�
�}#~]�UE��D�C�c��c<Lj62;6�.�ve�E��İ�̾��%L+XҢO��YK����M�w�~hW����`>Wܩ���aL9p$����
��/jʾ�[
�<�LV���d�w؊p�D�;[�:&Y&�z����>�*}��P��M������Sy���ߔI���9���'�1�k�U�伧�Z��w`(M�s�|��>W{�Gt�Y�_�iʈ\�d��3�ߦ����]l��:��X����h&*=��c]������ji���!�j�������A�<�|dXJTZ�Zs_��s�Ý�Z�?>tK��4�0���k�^���lq:��V*t����F�Y������q�5���t�ߖwW$��ƃuK1=z���Ԉ왪���Ś�V���Pti��[T{Vq ĔU-r��s0�#����4���r�	��K2f����S���wER߯�l�n�$ z��KP��L��<�^\�Ab��l�2yEW\G"�����u��[��	Jװ5;�yj�D��
<��/�З�.F{3����rЌt�u8q`����xw_6�⊍�v��J��<�b2����e��e�޲5a*&�B�d�+��<�j�ܝ/�R-yW\��МW�rb�9��Ǒ��*_����zr��5F��[׋t�8�T їT�Ʋ�O���\'#$^��6�N:�Ey��'^{�6��6��<�Aȳ��v(�����O�3���Ni�����5��p�qV��A��K/)(��>�J؇I;�%�z%�k�8
Z��09e���}�3��]���F>�H/�{��zn�����"�z`u�i-�XU,�
3f���c͸�����zP�2�軭`�=$<P��μ��Ճ���=�ȵ�)@	d$U4o'��%$]�W�_�v�`�ƛJ�h�I��XgW��,i!�c5��o�e��a��gT��#py$HB܂L���G��w�
R(�=���\Ԅ���u��>��?GW����:=D\���]�h�o�Psw��7��]�f�;I�5��}��5���6�!��A~u��}K��rֱX��9�rD�}��F-m,�ɾU�P�0���`g<��o�ȲE�fR���sLʍvj�F�Y�W|�mj&�vy$_�&�oi�\�qT4�ɗBս[�
I��ɮ�>�]�� �T��៩��۾���ݨ��g�9FHa�sk�Dx�ɴq$/uh��{��(U�yB���)�h{�Tk����ő�.�O��crf��=���ҹCj�7�Y��z �Ζ�*�~Th@&pc���ݽ�w�Oxb�dD�g�aH�2�W3q�LM$κL���T-Pm���=9��$�s&@g���0�H���ƿ&n �VSz��t:�B�lK��R�^F���ݑS�s�D�ĳ���d���Ѽ��
��y�q�F�f4aR��\��
_��b��yȣĖ�χ����`����yMڏ-��/�'�sw�,$�I����e�ɛm!��'�D��m�Щ���ղ���7\=�KBtQ�?Ł�����a)*��R0��lX+�N p�wo�)���ףCY�%q{f�5��xAk���&�W�ka�c/�%�}r)5����������%*�ɼղ(�_�>#����=v9%,/̵=��S9�$�ﮪ/�}�>�v�6�r%��E /!�� u��Cc!�;$e�//���SYgqdQ��JCf�.�u�t� ��C6#�LnêD����:�=G/��Pc<`P>&<6)�"���;TzSE	,���s2tJD�V,��Ϻlǝ��m�J�,��ƻ���!>%��;� ��E�o�z��]A�N�9���'wT �EO�Z�� �@%ӱj�p�_}�ڙ]3k\nj{��+�e��t~֊Fo0� 2 ��Vİ*	F�F�fؗhӲ3&�׀��;˿GL�ʽ�[��B��f�O��ӌh�B"�}�Y�*Їy�+��74Kڃ��$� �(}���F~m�:��#�ExZ�� {]�6�=�[��$4��(UW_��r���~'�{ا#�/M�w�tA��߆$D��)A5z�,��=#*�I�d
�L�v���Va���9��&E����r���CP�>=8�!ј����D��\MWU9��d48a�a-�>b�5ŭ@����3Y�
��b(��ʾ�`H�
�n4��Φ���C�����]0�}��e�.�;��r!�.-?�u3cGߝ�Z�~���"�4p�c�E�t����ݴT�_�JJ�?�l����Üxź'6?i�	)�o��pu6��$�MdC粦�fc,�!34�wh����?����X����ЩJ�O�!�Z���(��Ts�7y��-�˄��@�)Yq����c+�]AI�u9c��/�W��Q6;�R�u>�QI��t�V������_��v���B���Y�H�Ds���pHaG�`�f�����k�x�|]��.d����uj���˱�](��~��~]����8n�|��zȲ�;��p*vH�6�It���X�Tڽ1�E[������%Du`�n��rܯ�}�0	I���?� �����]ƕU�CA
�kћ�fÂ�~�(�m�Ϊk�E� ]բ���_�c�?\�6���gj��-��$�/������}�[�P+9�mfiw�} ��B���Q���4�� �|�Rz|S��TZV�#�L>�ϛ��O�F�����&�4��wi�AqI���B�P��F�m.����K�\������,�wޑ#�?O&�� �"��Vio���eh�@�I1Q����+���K�֟9	#���p�Y�68ʍ�V6Θ����P9=?o����` ?T8I��������_1�x���C���~N8#i�mI	��E]gz=_�5M�Þ&�.ts�#QS7o���s���F���ߙ��۰�LU޽x܈;q�Q}z0�4�_�a4\[Eh����Z��/�~p���嵎��Z���&�M^B�
8����p�������뭞�����+2�o�8��?��^co�ى����L�[`�*�P������{�~��xd�ݒ����X���~�U��q��b5,i�j�������.���YV��ŏ���uݽ#�!��`��� ���{�Vd`$���'���/6�/�Y����
/�څf�h?��̔u�#��(c_�Íܨ㗌t��q�Z��5�$v|s,��f�g�E�b��/�1S����fz������/��p��m^gt'���Biթ�K�h��չ�D�%jz�~'a�R
k���Z܁$Of�'^�M�1"���ӥhG���Y�>���������R�N�`=p�v���@xx�(}>�B�S�7~T��$x��a�2���G��Y�2��w��R�7+D � Ӊ%uhdq�zP�x�c%�=uׄۜO��K7m��0d��<.���U.��-�O=p�ЬҶ!�!�5�i.8���p��Z���ז��&+��=G�%�X��U"ԃ|hRJ�"j-[?6�H��1��
&l���V�k��s��T�0���:��:>i� ���d�q^
��<-�_.mto^����>9�ohJc$�l3	���'�g�
�L7Q*��!�A�5���x��h.w��h��4ᢇ���L��@�F!��� � �$>:�#�E���c�E�<\	 C��9��U7jm�g<ɜf�n�JG�D��C��g+�4������<�S���:W�!̒�^Pduϐ��=�Oʹ�F �{�UeL�����J$�����|�:F;1R}DZ?ظI����"/��8��PJ��v������&��^U/w�I�7�](�kTf�٥�E����8���2�1L���$M�~lH���L��V@I�s��1w� �h�NU��i��Cs܈��[�EI�e�� ��0�]��Ia�]���+�x�.���1��΁���{��77�:C@��-���J8d�&�����~B���'o�$vu����@�N��fr���U1�����ᦟ�����N7��, ���詘�C�W�?���&�հ���s�*,�c�'I��9QY�?���Ć�X��N�Ÿl�Ŷ�l��ӵf�=T�� ��t]��7㙱S"F�03 /jM�1�0k|�7DIa�?:�&�����|X��q�TX|��D,a8qD�-'�y�8��yC��қYƎϺ8?Gj��˹7qN���nۘ��vS���2åȯ���*�����&Կ���{+u�a�q}�ܩ���a���k��a'��9}�sF/ RK��?�ل�qwXO��~�>@yI<� ���{��ĢH
��S�����-��C寧��*�Ӛ��S�cB��+��h��T�?�C���
RHݿ�A�f�v2��w��qm��$~8c�l�b�vуvn�<�Č��I��@/{un��yQ��h��E�����
?"�M4▷N9QT���G%��[�+����Yޟ��;E��9ٔ/�y_��?J�h�=��ǖ/��l\:2x����*�>���%�B�{�@=�3�B���{)��}�+g�>؇ ���+�~Y���Kǉ�s�k�_R�Ѣ�=Ep�ӑ��r?���@��D�5�<�	��5���MP$e�ҏ�K��v���f����qx��?f6j6���#u˘;�?��S_Q�z2��}�!L�jd/_j�����
ݏ�o[@lAª]�a��� ��G�ݔ�qR��"G?������Db�s�����g��^BIR������5�B0`"�����ݰ_�Y˟�;Vi��	:�%�A-���^�F�ձf�l�k��1���W�17&�(����޹�}J�e���d�|O%�f��rl҃�#��خ�6I��X���_��+����Ub�t�v5��H���D71nJ��	
.�N��	f?���qe{�`[nDsc�0U�3��,҄�����gq��a����Mt����dB��N�9ث��q���4�?�D��/�a��_��g�Õl�L��nw?{X�'*9���\��bh3�T��BwpL�~�;X��y�?�,�ޜ/6�/Y�}���)��fK� 5Z*]�k�W���m�)0@�ޅ�$�	�����.��F\������r�L/�*6k�X E/z��r\�LY���fbt(�۝2���@��6�PeN��a�m��q���SA���7iURy�eL
��r~�%���A�Q�Hn	9��8���)�$�2���-��42��I���<Ά�p���#*s�V6+lw5��	�z�ws���Y_- L�$^�dS,*�#xշq�/��E8��)���L֪w�)5���ki~	���.�N�4�o�$q��g���P)���?Tج��Y ���}�#i*h�)*<��A%�"6�O�ޒ��v�7e&��
����[� �M��l�a�-�4UM~�h!��L��G�3�[��H���F�A������U�>�&_�fB+�T�������u
��nJ�E:�hc�*�F��㐉������j7��G��ڐ�M��%��F�ob�A�0.���,��ܶ����i*g�|�'1�>+S�_��FZ�=)@T1HI��(���E����$�%Wp�n0���d�-���	����]ٓ�F g�ԧxS�Jw&�k�@@.D5té�$�y"���?���KS�?|F�� f]Y��H~A^F$����=�*�#�#�x��(����heg9�W���5M�t�.ȩ� c� ��R�yx}��J�7Ͻ#0��j��_��`� �I�}s��vҶ^�Q�<Zf��S�	6B�Xy0ʔ�n�D9��ʓ��d?a�9�3~��O�d�>�Q\�1��G���ྴ�)�bt�UB|�j�cvB8B�5K���ۨ1�V��>B�<����������=,�Q(��`�5�4���6z��*��:QlvX��q�<0��?+f������U�\e��U��'��tj��YA[��i��B�����;F�u'b��\1��f]\ݿ4�EwD�.�u_�.��/g�o}�J_<���$�N�H0�g�����2:��W�R䬠󫡺��p�݌��&�E�{�`�6��$��C45� y<�\�"�J�y��㎛j68O��,���hV�둛�8�O���RH:�W���i`��T�6�[8�O�oA[`1i� G���lOcp�u���4K���T�Å�[��un���mG��2��V�"v��7v�2����R��yu������� Fٗ�xӳ���V�5�~��B��v/��>�oz�Ҍr�5s�Wg����ý=TbǢVJB�I�_�)�����CA4��͐�G#��,�'f<���Hx�>�3��Z�>��|?ɬ�7���E�p��e��Pd �̗Gl�<ύd}��Mɇ�/����rW}r̉!y����F��n%x��>e�E
*'j��%CjF�/�=��Z8Ξ3������E�i5��WqD!���Q���U����g�Ans�ws��+ �25o���Ө�]�z�g��
�+:k�vLb�c|��ʼgUfYacB;�Qu*�6׾�7�ysf}�aW�+��<�$pvnqu����z����N1�u�Cy��7��W[�����6)Bg�B^USO�r�}��g�?r>�YK���T�t��$K�V_,N�m	�JМ;�BuD�x��n$'�,��� �[#�:�b�C�u�с��)y4a/*�l�=]�d�F]�� B�xt��[]	9�t8���o������(��%�v�\ϕ����"�)���M:�rlGL�,zHU�ݞb�1Z#��5_U��� �(4cB|#mY�z�U��Q($*���<�����x@7����J5_�Ϧ|�/Uf�~�K�|���Դ���o̕�3#w�@,��,�� ���g�����=O��i4�K�d�l�/Gg9S�+-j)@��K։JP��W� ýY7���M��Fo}�W�AͬK��nsUͼ��3���y�
X��z ��1N��ݰ�F<Ö	$�p�hN�V@��Y,�~��c,H�o���7��)��@��hq4	�J$�XoU�b�76�BM���f'C<u�"3�?�D��$��6CY����:��B0; hbs1��%�G=t|���U[�z,?���O<`���?�|٭5}xb�;2��q�I^[J_�������:��+����3�)=!t�A�g�m���w��w��1�8�
�
9���o��K�bf��i��r&�u#���X/����n��~Я��f�8Zx��>A�t�X���]?�~��Z6�v�)�eZ3�f�[_,Y3�
�N�2l��q��f�#���#9��B��Q~��Б@ZFe�o���C���G�>q�b���G�V�,��yRӎ�@l-˂Ƙ�����Vh�i%5�1�B�B����~�F�N������/	dJ��Z�����'n��z�ִ��nW��"��;?؋�r�S���N$�/J�0��ak:fd�%�dp\ZL=�ʆ��qi�T�5i1��k��Q���{ �g�_��q�o�s�I����0��; %�?�������?6��YI��|cT�m�2go.�{�����Y���1��.�O��{�M�����\C�� �{�;���S��y]qy S�ś�wͧ��w��x�Sv �c�p��W>����֬~��ϸa��Ct1-K�h���{x��ڄ.6)�d�
w�[#��|��eAQ�Cu��ɽ"?w���?g��Dr. �\�$�ǵWd���g�:tq�<�O!�1�Os"�����xD4��K|L;[ѿ�@�6��T2A0���MYO�ېú//�אت�Xΐ��` P9���!�o�r��f�����\�ό� |����t%�S�Ī��D�8��p������@ wJBSθy)eYbb�	4l-�0����y��d�c�l2��M�/�Q�J#���7V�@IܭB���"�L$X���d6�s~ҳH�=\���%��ۖ�s�?�D/י��x��b��*l"��]�RH���6�-:�㑉P��p7��H�&�����/�]�$�mU"��MD��X�m�����L��2��(�b�M��bv���A�Z�t6h�#N��A���u^ʪVR��)\�#�U(��dw5ɩT����EM��>�������\�U?V�p�����&+B˖,g-��~����8�q�.X/n�dmX��O��<�uI&�m���4Ң�	y��#���7P�<�'���Hw��ߞ��BxJiy#&���>��7�6�I^�&���?W�{����ܩ��K�/��#�|�����s�g���0����UBm5Z^��l'��ԏ�`�k��[k�WF������n�1�<�pǞ1h�g�<M��3�D輵JDT8��%g�m�-^������3%�Җk� ]��"���1;V[�.	daH�Zus�OJR�@�C�\|C�M&��̇ �
�����=Y�1k�3<G��L���}��e(� ?hD�c�S}��v;��^�zƊ���x�gm�T��ݝ���p TM�U�T%�{�k�������=��q�H9Zgduv����#�����@�U�XY�d>Ur3~>u�.G�k���{��k�J\CnVRif)��6��-東r�Ѳ�F��${���|9��@3�s��D�����ɛ�[teźδF{�H�(ij�J��}���������aJ���9U
��q;��I�ZG��ç�YX�'7\Gŋ��qʭU���q:fm�If�u� K�:��=1�u?�@=l�[ ���ɔ�T�H�X���T�1L���o?��ԓ�a���`H�>�8�Ē	|J�ۊ�+j�,Q�� ��GM3��#�/��Fg��a�;֥�����e�Z�p�8�r��O����w��$�����B��k�[�ף�,zXY��x�л0��Qa�SS���x�S}g����f�4�V�L�w�Vz	�Q�.t��GU�Y��ӟ�1����6l��R� ��X���z�Sa�S��R���q_�s���[��S�E}�$EC�bM�{�r@(~d@�-G�۬���$'݈��I&.6x.b5�;��S�ce���I�%���U����<�����5�i�_�S8�-��4{o>�B���%ْr�s?@�l�,�W[v�E�>��vJ._�	n1,�q��	$���3/{��{|�X@����`�I���4���އ��ǛW�HiR���VD��>uG�&��x]�S�``뉃R1���>����9O|U
����bO��;���VB�dQ6���~+�Z�`� $�Ƃ#�hƼ���٧"���̦Kq��Mz��^w�Lb�]����Yz4�P��2�?�� .�8����_0	���������^�SF%���Ri�h�p�y�O�k�g�
����
"�h�[c��_F�mND��2��H�q� �3�@�_��o��o�T+xӗ��N5̦ҫ~7c�0T�AY��Dx%��/��~(�����E1�)�5"���B��K� �E0/_��w]W�i����@�@�z�<��5s�OnEi����j�N9!��:�
D��U�l�W�x�5�,�b$� 4ҏ��U�a�����=���'�m�s���,���Vui�l"�)����D�c��`F�N��SH�����l��x�w�d��(m!�FΌ�������_���k�2��)��>wc�-�g,�&�^�bs��F��\D�����%�
�(㎖�Ұ��(��b���L+���-�o�ʴ��BE�5����k�FL��A���B`I�5��pđ5��Gx8l9�0�/1,=fz�����$��@�0dJ U�E帝�D2���$GyB�q��,��p`)���+��܌� t���ks����i_�v���g#���v�z���3�F��GX wE3�G t���A�@�ڪ逦�Z�A+sk�Kr�4����T�j�Ԑz��j��	�=�By�2�JcɏyȊ4���q?]�T^f/�d7���d ��5�k�kdx"�E��7(p��Q��=�x=�g�5�U$��8�I�� A��y+a�2��Z���ٮ��(7AαJg'-|�_�<�7�#EG^h���B�+~Y�V�r����m����� �1il?,`��u�����gڥ��I������;��c�e��E�p���%�Z/�)�R3�Nh붞$��@A��<_, �&����Fp�A6\�i�\sa7�~����h�QR�c����e%��:�LT�����RѼ��H��jr<���3��{pH눋�4E㎧��	��>�H�I+����\,
�E��s���7^��(�ɸ��-!5� ��m�9�`�n��UU%����'#� �lZ���b���G���B3�]ǷKQ�U:Wظ)M��_����|b�<�����kM7��ԄO��ԻF�0v��i��:�f��������ː�5w���?Y�L���{�T��̬m3�y�FŹc��j
#µ��P�A,�h9�˦���	3>Uu� ���|��i���!_��=ڈ�^���?'����{}1 lc�&x0!�M[&=)Σ�)�R��#ޜ�r�e�&��#�� �&�V,���|;����V��c➩��,����GR˭�֮xGy�֥=|��xPY{�۩CW��˱�^ ؜%E���X���]�ŭ�B�ԑ�^��2o��ڎ��v����Oh|�7pFNJx u"P*b��qI�\5��,�!�,磝�a�0��i�8�b�V��{"���V�[�V)D�Q���39;���
�'��a@E\�Q�y��U�ę�|�	�q�d����4�-3�4d�@�i��n0K\�ܬ��A!P~} b*!�V.��R�AA����:���o.q���Y��X�-�U��EZ��G��qe.��4����!v������\�ɼ�jiw�(�(�B��R���xm�#�!mp��g�BŰ[�r�]���>|�(���^�qV S��!��3SR�!��Џ�H�+%Z�5�#�}Lg
ζ��4b1�B�$ʉ��	#"O$�UPu����8BA/�j���0��3��w]�K���JǍh@,ʔQ�Mr+�\R��C�+��X�ܳ��W�B�^ͲT'l>��u��l���́�ƻc���9��� G�^� �B�""���ȁ����[��RN��n��n��������\\�d�M��t��_w͑�;`%a>���p�Ps��,V�������Dq�~����<��	�]���&x�b�o�.��pܳ+���N7j���!�?_2�L�M&�!Ȅb����j�Efvg9�[B��^��`���;V ��f,�����+�V3�ƛM�*��l �>�����7�ƺ�%��U�Qk�a�4��\lo'����j�����R�=�}K��"mu{��8F]��>���`y�o%O�D�Ue%��FR��O�H�D0~�M�Hy6��Ӝ>��OL�3 ��i&{��Mߞ��f��2~�*���D�&gS��g�Ǌ�"nڒ���罶����,�m����h4�[��{?,�k�%9E`-r��*�ɹ�=Xk��ڹ�zE�g�gC)K���/�u��D���9bf���5{}5xr�`�RWt�R4`�o�I��؋Ǹ�DS��C���w�m�[N�)�C|�B+��m�ș0-� V�?�}�=��	�s�1�x�5��[
�.�u�o��v��TC,��������H>�o$wȈEn��
{��Y�E�X'��^��h ��qz��j�
>���G�Fc^��,�ҟA��I���4��-������=OA�o$�E��>p����s]��Y=�_�Y��{e��,du�\䓽 ���F��*u�����W��N�msˌb-�K��#�x<�5Bw�H�c���)��c�@��eL.6	���O��2���	�z�]���ɰ?���*�@UA�Y�tq�Li_\�fY 4���8 ݅��I��&�rav*U��f�ZN+��I+���
�2W�"x�#�x�q�l-��t���j�/s�����\����)rڱ��2�g��V>�����ɞ�N~�	�9�K|�u�+�j�}f�3��wm�E���w���ʱZ���m�Y�o#�_���ׂq2M*'���Q3=N��I�I���P�p���g�w2'
�op2�6�	Щ���1M�N$F4��o��$}�bl$��i�	��$���Q8��)5'����a�)���*h(W3�'���`;�e���!�l�}���AT��P�[��E���%;8���m�n���� �}���i����h bE�!&܍���IzbX.������b�u�c�%�N�&܊���O�B�̻�i�./�X��4�ɧ��GY��O>5+���U׮���kʃqLC r�W���a�u�����8x�k�7Y]]�##��iG������o�&�`yE���8�򺑜=J'�(֡��:���b"(�HG��IMI$u���:7����,9j�m���T�
-�a?�&<�>T������N�e�x����~��:͓?�X�G:����q�rC��mt�P�o�nҎ~4��r�ĵq�����;y�PM��@8)L\��N�]����qMC8�3!��؇<����ѷ���>^��"mi�#� �s�U_#��u83^�y�x݊2������&��y����җ�"6�lg�����a��U���J�
����a�i�����o��>N_j�#�yZ�x�NFΚ�l���&h��z[�m�o��s %H�-9�E���?95GZ�c�R����R�}�/�i[��R>k5�8�,QR�a?�2�} ɢ��!Y��͔������D$�-
���s'�T�U�'���vK.Ӛ.�)������ٌ�%�-71&����l�*���6�p\�M2��S2{!���4��),{G��ߟ夢���� x��S��`����J�{kϰ��է�@�����J@hl�)���նZ��N��@� ��+< h@`Whʢ�F#���s5�m*�0���m�b��Z���ۘ��@N��9�E�%�V��)�T�^���0>w0lmq=���H.}@��N��:��.v�kJ6��Uz9���.���}-�m�hM���!,���H�:E��I\JX����L  �:����<����C�#�e@,�`�9)O�g,)N��`A5��T;v�1"�M��煡x��1�����Z��rs2c]-��~�d����{54,61)HHB-��)����6�lƬ��ݛ����X��i�Z�O~�E��o�H�U��ǺH����5�L����R)�M�Q�����[�Il9S��G�H�IK0��#�O&2e��Zݽx���
��l<5���3�7t$k!r�kU��Øs3�m����F�)2�od�"%�3�����7-��~�I��Si\5{�u��/S'����y;^W�o,qsNS)J��4f���aE�l+JB��0�Y�̹�c��A�Nw>������n�m�d�{f�3�}Q�S�6Hz����ucCӽsE���ŝ�utMA���g��h�[�+�;��6!��2��)�+[�2�d��q�j'���Z�y�D��R���4.��X:Y���@ZO�)�kh*,GJ�
�1Ù��y�\Ŋ�q��h�)�K����6Ԙ�~"B��O��r���'����(m ~/�P�!��	Oq����vw�W�޻$W#�1ʦ��ΔW_l��n2¸�]�mo�z�nR�Š�����@���I�®�/���� �}ж�.���
�F7�˾�x5�q#��Ⱦ�/�E��5�*$��t�ny!	�&,�$	�N�~�t
���Ym@�N7q���b\�gq-����S��׺��mv�#+ �i�Oǐm�+��vf}�cK�5V?����Mj���i��Hl���Oe��
����>p���$ײ��0ڋ�����?��^*���J���ނ-�)ce�
^
?����c�I�.��;��� #���5�9�7�	p\�͋��Z+���mK� [!��qN��|��'�1ޖݽoº��6uo���ӫ4��|~��s�>D�ig��ٓ�J)s���f�75T�.D�n��'��n0�*�&���(���M-o������f�o�����;KJ�<xt�b����;�/��Ҽf�9y/�p|����,7'�r$zD�)C\Jb2
�(�AԞ��V8�(h��W�/��U�j$'����=��b �Ҳ͝OE#�O:�7����@Ǥ��](ON�	jFא��?D!E�
�M��F����>�0��	�oaKy#����;��tQ�!;q�{K}M572|����nz�6n�jgҽ����J��m�T�t��1���M��)���&N!�Ѽ�}C
yo&ɧ�:w]�J�$඿�lh�c�@%R�~���W2����\��7�+�lj�0ks��#%DM�D�#"]bO�c�V�X�s{����=�F��队�)�)5�gd�<:�R���N�|���D����i���&� ��C]�~4j�mzv�ag~�m`� �Xpy�I�=�(p`C}5��G)Q��k��๾>�qy��R	����J�ˋ�(�V��D��b��`��p�[�6\d~�*�b�Ʃl*䡜�
�%��z�~ޑ�Mi&c�}�����G��1�nh+)m����
8��a��U��h~�<*�VU��"��v��_�K��>�M%+���qY�6w��\Xz��VV�`BF�3)D��7&q����ֻ߰S��j��9���m�@׌�<i#b�s�ߟ�����3��8�m����G��e��6u��Τ{��p��y!��+�����m�0�E���o��-��ΐ��Hx�Z~��<lij.`xY��2l
��"X�L�LbA���zQJ������cVud�&�ǰ)άTx֝'~G/{0/c��� 1<�ߢ6F�w?�? ,~胄�A�v�*+�2z�e�������>�U��d�����XѰ�49��c�T�T^�H.}'x��H�RQ�x��!$�fn}ɺ$��B�X��n2�׏��yu#�� i�M�b��8��w�s���l���A������h�����]Ea=໑���xv3kB����:p4�r�]��%�t���{��oM�%D�Yo{|��h������cɖ�Cք��f })���saE�V]Zc����xИ��2o���XB����)4��di:������u�������m����}��֏�p��aێ�"�8[�(�E��Ӗ�w���Q6�2�d�=�/��0������N!�����Ɉ��Dn�[�i���B�ϔY�:�`J�4B�{�Ѻj��>o�A�¶� �F����{Or9�x��+���NP؎@ӭ'Ƌ���㒲𬇅e*2q�]����ol�y�V��]��V���v��a�`�֋���7=䈞�Hn=!g�2���+`��S��b��
ϔ��B_Vx�,�h0�-��v���2�Ic��%�g��([�S�4�K�{?�?=��s
EC/sq�n�gިNR�
!�1Ο#������mtV��B5i�b�s7$�	���`���� ���wY�f�������D��	�P� 6y�t�~��i����tW�v�9��@m&�/�Y�ې�x��L@�0u����C6���%J�t��G���{�k3���0��l�.��!�|��g��ktO��/؁���}H$�p��|	.1�����"�D�5�40��Ԥ,��WS{���䑔t��y���e�B��cm���-�A:��]S� �f�ΩlSr��߶��8��¶��j�h���Q&��k�,#$hs|�����QQ`����E������]o6	����W�����W�A�6U� �*�=|��8�gd ��|EʻE'Ƹ��P j4�aD��},(G*�1��i{u	2 &7e�|}� DPPA��o���)ҁ�QB��r����%�+���wus����o��&=n�y��~A�S8���&�͚F�75��d=��æ�2�Aq���Kk�ȵ����u��"6|`,Y��^�?1�g|�y5�`噡�,JJz� ���L�}���>��z���c%�8�9EO/|0���� ��CX5P
C���1�w�>�!D���{^�9��F�e������_`r���c�t��7s�$d�+��P!v.���Y[��l<�Ez�۱M��Ύv3���McT$���}�~B-І��d�6���	���J�3L��[����Vᷓ#��F^!6:�:���9�1/�ͱG�����?�1?�)3���]w	��t�� ����*P+���g�I2&�vW\N�͍�G��Ǽ�.Z���zf�"��r`��C��"�֥��p�����v�8uG�@9K*Z�y��I����5�e�B-u	7�P5�<d�.�+�U�ԧ��<��	��z~_������ߔ�$�\Ax"K�D��]�.�T�8��#H'yd�9w �?{�$\�DM	4�\}}^�,��A5P=,��!�� ބb� RF��8J��Jr ����QP[S'f"S�lll�^��CKj���� Q�BUK�E�~q�>)��*�զ��w|[�#��@�$B���8�Z���A�
�V��F���4劺�nf6�Ysي_NU� �n)�dq�{o!J���d�O���:�R��; b�4���@�FZ~�8_�Gn�,�b��;�'����;�b��Z���_��U��P3��#�e�4��/-�g��E�Q�C��A��ff����s�$n���X�2�Z�~�O��v�pj��N��{��f�e�r��B§���&�E1mQ�*�G�q��LƉ�%�Q�l��,��+�ҝ��3��å�e���Q0���wF}y�V�$K�a"`xP�j�΋@�O�!q7]�>z����+�`e^�o�Áa����>t�������".:���\T�lh�kHK�����������ʔ_.�%�\K�!0OEWĴ�c})����Pl`���z�Z��n���Y�tY� �̶0&a�t�����3��?�<Y���X��Wɢ�-�$h�eB���j�[�J���E��'йﰷ �;|"���-�5���-�~;v8��r*�E��Ꜷ>�ߒP�kxc�uk���VKi�J�혝ugeF�w����av3y��{�{��{�����H?���$�h4���[��;^2�ڮ�=î�E�Ș�3�Y階K�Y5ؖQD�I��Eh�����6�Ǥ���w��� �c3���3�E����>FĂ �6;nn�F����L��^����ܧ���S|#mN���A5�pgQSNa�TIh3Ո�h>���h�Ôj ���<�$��䰌Qz}�<8��ђ%o\^%�T!`,��t��MM�"\_u��'sss��Np�v^q'߈ׄ�HZ@�p߾@w�R������$�ai�HHgk���XЌ%.R�5N������W���9��
q�p]��qKU����t�����o�4�����a��Ab
2�aIv];2Pņ�❼�(���h���*����r��&�Ʋ���_���NɐC�ϕ"F!���<�+�ٟ��#�����m���1�g�Rhxǫr�E�ơ"Y�A�n.d�U�� ���+�C ��R�˨7%Sa<U�4�Q��Џ7���X�n��~�s�*j~F�����HuC
xl����yVXKQ�.�$mևҟ��Od�aӶ��VM��yF�@�_� V:v��J��f���q ���<̆��y9bl`ܦB;�ę�+��0?E��LprB��k��:%�F��Y�_�N�9�7%c|՘W8�_i�l	�����R%cܡ^�,TN����m��f ?%�U�����	��-��5��"��ǳ]���Ƹ�����8n�ʘI��N>g/�C4�c	OL�s��q��f��Dk"��%ִ9O�#�/��\�2��i�~�P���gW�n'~��3���E{E��XU�i���&���d���7G�\/P
�F�Np�P�Vx!��n�HKV�}�OI�E���I��'#�>p��s \�����1��LR1�h�����(CB�ƺ̿�ř+��1��<�	�a�ķ�S��:��ת�I�ʆ�-��P�x�源e�h��q	Y
P��`.C�����ɳ�#xw�t���j�t��������lEK�~o�O�#���;56�~`9����&?m��)[�.����5��3l�%��ȟ�C��<,Ҧ�i�5�w]�q]�d�u�l;e��,$�Thv�� �X�}/^�~�[tI�q�D����ٱ���Q�C��V}� ծB%�j�k
�UG9OhJn �+�
�����Q}�X!��G�-k�����'��Y���ו���
���Ȩ�r<�E���MD����|+�[���-�8��,�w�T�5;�u�rV<�aↀ0�V2X�&�!@x5�!��B�
DddRm��R�Ju�'�YSi���HXR�'װ���3]n�(mj����Hʋ��Dbش�� ��g�Z����99T�$�d#��.D*uSl��5�}�	�\
�IZt�����\�P3C�%<PL%m�zL���,7H#	�s/�o�{]�����g��NmM#��`M�6�~s����gg�t�9:�n��c��m�����T��I�j���������e��+t��������P��oȽ���l��W�Ò��K�k��5��4DP�۪{�1��D��hG|�+�Z�|���^W���l���]��w�e��(��(t����;�c(�@�"f5T���s7���yy�:����/8�;��ZR;��VA��]�9~�J�U�*���Ĳ���k�I#��C�,|�ex�A��qPڍ-�nNZ�z�4X+H��r�&�Ps�,آ����]�Ń��P�\[,�-�`�JF�O-�C�J�p�I��f�E���c]�m"*wfM%(�0_�ƏӉ�N���]#�c��f��G�<�Vs-ߍN�1��� 2��ۈ��v%��B]�6��ױh�9*K�b�*�N�+Q�qG���HA*�!0�0�')H k'P�M0b�/s�������}�Z?�￠�(�.S�R�_���@Ǖ�<����z�QI��;m-�߅�A
ym)/��&nU-*x@4x��6�{[��)`W�}�x����!�`�'���V��"riH3ē����X�{���ԙ9j�Ŏ�e�U�0�����[�zB�w�w�����C]U�/��4<�NR<�T"���%=�\��YϠ��;nCa~��hO8�\QC������	�>���c�~40���2��d���H�4��b�x�A��cv<��A\�E��L�B��ZP@�:tR�U�k�$�/>%�ՕSٽs�1���g���ˢ�Қ�'�<n�"H��Sع&%��L7i%˴ ���t��	�!#���r���/s�2֕�v� �O^u�ُx�d�;�^"E����\�洫f�� !�fV�b�)�4:�6���'S���j)|���_`��m"I��@z�7��Md �,�䱄�̗�L��4
s
TZ�B	)�T���m�#5a�:��<�Ҹ��}�6�ebX�N��.��ѣ�y�t��F�D��(Q�f�\�bp��'u4Ǝ�b��o�I���궁��
%��G^�x:��ch��ھY�<`�{�9z$�a�z���Zo �a���<���.R{(�6���*=wc��/��7�OJ$��#O���e������@n�(Q!����&k�lu�Ò�t/%r����Hǫh}y�/CC2a�:���������ФVaI�F��OИ�(j�(*��2BBϧ���щ,����Av$�@���5�گ��h�Ē��^�l�Z-0�?�cK���
W}J��]���"!YSJP�*�vOT��*�'`�P
������X>�R��&@���c��"������'�m?��Dw��g�х�ykN�����F�C�X�2��O�ؑ�j��3�
@)�f,Ѹ�Ç�d�Y����%8���.�;ړ���|9P��{I�����\����5�� \�T��x1WA_�9IG��XZhq�~��0��zL�0K����9�z��zQ�'�3�������Din5�n�BZ�%�[o����t��5�[��.�H�T�v���IЅF�Fs�HV�)�i���Äϴ �C�1�11�S���.JaU.PܔpD�������ځa�9����E�i�|��ŧ���N�?��hA�e����8�%q����.��L2�]�8�؆�n���O�Yʹ�4������Rj9�d��a����3h���w9��]�����,�Y��P�TW�DJ��*��o\�F#������K�D�3�:9�t8(�X�m�~������m�̌9k�a��J\c*��8���4v��Z�H�:)P�f=﬈!�dذو����|�gt��U^����r��ɶ�U��E7���cR�Xb/Pd�\=w*怬��p����K_���cV2�3�p�4�OQ[�����ȿ;�֧E/��x�g���i�셼�|��~�uu?o�[R��w^G�p@j��:'x՚�l2�ri}!i�Yo`�� ��\cH�$q&DZ�0n#��կէ��J�~��kS{y�3���uf耶�[PW��4��$C��i��0��=-�8��Q@^�ET�Ŏ��19��`dp|���m3�{��Vw������sϛ4�@e�tm4���Zs{�y݌�Vnr
�bh��'��@R��@�k��ϻ��� ��xk~�k�)[)t�@u�PmZ�
}�Ƌ�oVJ���`��H�e��x��n���4<��<�Ԇ�E�x_��{&�{�4����B�4�c���i"�t�N����lt>\��Կ���#I��{��J��M�:�
KJĥs�VO�b���R�:�EJ�cV?۸�yk �"�} 6�
�Tֆ�'�h�{=*ħ��൳nQ�k�K�ʇ�˼/���o��P��S � wOo��C��X��dۡ�=	��ꎯ����gB�a�'��uʂ0ޭ�e�d�*��o|��Qx蝺�Q��ًs*�(Q6����,�-P�<I5Lj�V���(l ������ȓ�>�B%}/�U�T����,�h���gË��*M�\���-]kzW-Owt'�6�{=�&��"��95 y#���7	��B�e< +��%􎽈�A���jiߗ�'��7|C�X��f��[�Y����D.�5ln�Xv�� ��E2�x^�?�r�����C \����㻝bd*4fi�[s�%X�A����snp�H�bJ9d=�ZT������t���X��R|t�Hg'��Q{uaH�L�n��Xu|�m�V�$ 7R�b�sNb"�ߪb��%���@!�	=݊� �Yc<�P�3�Y#k��t(ߧ�2�[�yoԓy���z��~j��씑�$2:��C)�c���}Q���Ł��Ӥ}3��8/z��j�6Ʌ��s)�H������1�a��|�XT%�7f��|�$]HZ�>��g�Ҕ36�/h������R�^��6Eq����\��8a��6� m�4PAq5����^lQ7�w�$���{ȃu��ߔ�ɩP6�l�׬�̈́����Eؕ��6����hpy���ɥ1��Ϗ?m@�}��Փ�r��	Ŀ�e����/h�	�$/a�ƣ��9�+���������,#�Rty(掁���eR;Fg<�\f�uKz,%���ή5D�8v����J�*��N,�fC��w���j�0���e۷�򕝴hݮ��Le&�^AQb����Ͻ:d(��ڧ��8�0��n�)��*���!�@P�*{q��h	����@�;�H <#e��4����T���5GoaA�!���!Dאָ�5`?��M~�T��+>��ФV�p�}�����Pm���%�\���$!R(oeo`�}[�׉},C@�p�$�F62�o��D�ԩ��0eN��P����:cofm$�P��µF�y�O�緗C�3[T7�9 ̽���I�������64;�cs�e^n�gxǕ�>��KU�_�!o�������l�_2��"]P��gQ>�QV�g8���)'1|�m̸J*��~��5W����	-o��?R6�c��drN���?��p�A8�S{�&|�B��?�)-<�Ĕ׫O'#g�o��!�h;���(I|����E���}�"(h�:��V��uwY�R NDq��:�=�����S�Y���}� L������M�o�2a�<ə"K3�RЄ2�,���r$����'������<}��R��là����r��i[��!ǘ��0n�f�<�,V�D'
�z�tL��b~)M��k9b;7<+W'�ʫ��w
�碐�����)�f����[�cy��_����&gTU-q�⪻���u�0�ā���s��0�44�xE���}8��=�@l	j����L�X�H ���4��4����"&�a3����d���O��,,�d^�lʅ��Lr'�a��ϲ�\6`YN(��ڀNv��24�+Y/�LS%Z�O���y	��������,���}�E�QǐK]��!X�#���i:�D�	2z$�N �A֌�m=3�4|���2�%��PM۹d��őf���H"P��T��%�R6�W)qw� ~\x�]���3�@�~�F��3��&���r�/���� �2����qok�l@��b"K|�*�R