// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:56 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ejOIHWDhRJF/uZuKgfi15cZjrfKmxDtbc+KSwngGrzUhDlb+4RlyJR56Uc2GoHnE
QbUD8/r9q42qArLbVv2p2IVAmb6vO9yFdeAXBFlylFxgHgBpLBYczW95zfK0+6Ps
M/KQc/9wFJ3+Ib8RzIaznM4DgeQ0rGiEiWRCm7l38S4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2192)
/7fbXmu7hqTGNiwrVXbStVRH+h7vLFWs9eRjA5hj3cD57Ztntw09g2106uo8sx8Q
zz4jYH1lpzshk651kzolLrrUmTYCJMnFobRThRXHQY89OM37v1YiRGh1NNwUI7jT
KRnlCOlCwVjhkdWpvds8K5tMyQOAVbyihV2MFXh5bEfVuIJujDuJsqN8UaQ9xwEk
IMtwDmXcEmgBVssCP/sbCewevzRHnT4pK4dEgp91adZMQ204374QYKmQBdTS5JzV
4sqNmfjK/LvvXR8kN8Qd5w1I58BUJsKbH4xiQF4se6O3h8ML94D65PBZ8KvM6Oy5
4R9ELFGx7AJx4BaVHW8UaId5ekTPk75iMwY1immGXYubgunEQyU87i/v0qhvee2k
uHwsveRR2eguxrmDzIY0Eu56w3xNjGlvAvYz/UP1uSm1zubC+zjL8mUIXk3ilL++
mhxbUdBxe7xyjbR+irfpLEIHGcYtGkj+Ae/9OVjoTecInk/Hl6AYOzaUaZU0nLaA
wG015l+nKIXefi8PhjjZ4GgZKVS2I2thgPXWV55QP19vrbNQEI9tU7PmSHIXOZ5o
2laKmovD2nH2hKNajDKZp63it99GVuwetckSSbMP7ai7FABl6D/Al1F/CHLuuERF
sxn12ySn80ThlYnI6VZ+KPScFNDJzRYH8CE90OIqsc3iR+FFtRGuVNgHH2bbWmuJ
iSa2LuRDP+zlhGVCbazaXo88iEQTgNCuwpMs+ClxJCfqqFZbMigAvWzOyQS/Gzkh
GB2L9CNyie34RLdGETrmCR3FMGU2vnsmKpIbjZ3a5HsNTXPjTKYvXePI1JKVeQjw
C6d4Nbq49tueOR+T1HodqPKguyFQp4pW67zxTa5gTzXDGD50fnht3LkNh7r/q9To
l08zed2Md9xhywZVvbuyuDSJNndUvSaWiFSgkAZCLWYmY5VA8SyyHHng9us8Ltrn
Dok3tEjtTfEncMNQ6kbsPZOYA1IqGBYf6hkQnI1R2LbTejLnVie3XRnWIonCIolM
cR0OYA4wmLe73bAHL4EJl0v9gwRAUmrptO0wQgheGLp5j9ZAoKtT3+a7ETY1xgV+
0UjvxMwZN3cuY+Y+6G4erKXHtkoX9bQqgCMJqqib0lgf9IH3NPfQpL9i0VhQ8cFM
CVqSNcCIgrlA2NcjRyaFAa+6c0a/zWGR3ptEQaht3goxu2YpJkVsToJS+zxQ7oqv
d6sXNFsPNGZQc8hw7tIkMS5zNHyR5XwUFAeD0Byxbl5HGrIH5pLkU5b9bHn0BM8w
KM1Tdl5d0zoVv3hA+hLVzIpXm5W2APxiEW/G1uf+Ch4gaV2BKGoJzB4RWJrWGnAE
24W8mSgDg2MO8ZUeucFayCCYKSQsTX5MV+k/lvBDZXuB8DsPx9co319AU/m4hUYq
+C+I/gSiMWnM8S6sPN6ejwR41k/6Mgw14VJw7qT/DIOayZpsZM3kvK+cazVsz/wb
4IUnR1SxktzesxOclLF6yyF56VUbS/+heMi4wbaDr4WKl1gHrQiTM+mGLBcGixas
hA2pTA1LSkekTQfjPTofN94dvJrb2pDLe3FABj57N55r3HNUdHCHdR8DDNNdzpcQ
Z48aulOkARLK1HRFefk/noo5+lxW8go5z/Fcv3vOiqpTmx0SXBz7uqVtW3OzMpeZ
+/hvI3KXBn6Yf0kXluA8YDSXBRXWVk33gTi4yA/pJQAkpmeCl9SkuPZlTNk0lvhV
CyNrzXh9xLTCxV/Yh+8CbjDJMctHeaOEB5Z1ZMNgrS8Nh7xtnM7gSIIC/m4uFdV6
0SUOIdtKl6O0Vl0QctTB3RutTSuJ8xGHdxecGWw5Fyl3jkqPE0dLe+2xSIWybvhY
ggBAstFh5yz4xm1n/ES2PqZW1cLRAgL/3Gm3TuPBzryu1fynsuEH/wUpuMff38dM
HEiezlsJRTdiorgdbmTsmgGP/laelkndjE18vUq2LwVN3VVFA/VfY85rxGacCd6A
V8Pakj96CS5pFEvxH1nuBiTB92zaweIFLRxuyuwrFYZuLUXqX/c1OIALUCYBuE8C
ZqiHdhqppuhUTEYW+uPaNJqyzoxDOUeYEdDgxiDaBgwUn5wTKQNXaLtr9Ubfap8i
5DNoDlfeBRD4J5IgqUII63OoqlRV3sy3/QUBeQr+BihnHG09RTx1fiTF1N69ViQX
P4mQMgymk2MF9VLwPcAGabltsacmpCaj9g+OxoS/10gvLnU8ZkXBrfW8yN4BvQpi
ELUzOMfQEAeSpAvG24yjGekwpquq3SrNtzUIRj+nMb4N9rNSlhQ7D8uSuYcSxORl
d/stqkMfVvd2580RS8jG+3SSXtEMw/sGu4rlBp9Sw4PA2sYXnKKrYk6ASFLs5vM7
0QnSCvesjKRiijcbCZr8jxPV3L+ilTH2+kTrJqez3mkkiMGlFRMWyct2+TbeR2wQ
/NYzsdiNFh7nRbc3uT267s33a2PrDPk4yAhPoRQSamh/IZ2/zGD3NmLoeZIXNqKI
nwfKTOg/DKI3Ax2v342xRd3uwChTlKrMI2M92Xzi8j/vBQlCtLls0q4P5xYDhSkM
cQbz/nfKcpFU7UBN2zDIYXzSWzQX3V7KE2EjfRr94uMIhRDRoKXnsheY74iPVNJj
Trf0QTA+rrteFbf+de2gIIIwrKySLVEtSlYLjSMsbWMaO+enagfPiAR++0GyxWto
kyCZd6AldWU8wMXkIPDnhJ42YTW3t+4iCUrw7Qrw4vroCBb9wXkZv7YROpHFgAMw
SkV4XYxdRv9Abnn4mIvWBPc5ag/QD9Nx0TV5rrZOh35Mz4whHYNp4CUIj9LWTHsn
X/ejxsVPcvKRXJe7m89LmP/5ezOwllsKn5oDUbelICSME0Gy0524HmAYlhT/KNOH
Dv7epAG42QNdmHbiyGjfc/J4LhU9N3oVzGIid33WFag=
`pragma protect end_protected
