-- system_sdram_0.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system_sdram_0 is
	port (
		clk_clk             : in    std_logic                     := '0';             --   clk.clk
		reset_reset_n       : in    std_logic                     := '0';             -- reset.reset_n
		sdout_waitrequest   : out   std_logic;                                        -- sdout.waitrequest
		sdout_readdata      : out   std_logic_vector(31 downto 0);                    --      .readdata
		sdout_readdatavalid : out   std_logic;                                        --      .readdatavalid
		sdout_burstcount    : in    std_logic_vector(0 downto 0)  := (others => '0'); --      .burstcount
		sdout_writedata     : in    std_logic_vector(31 downto 0) := (others => '0'); --      .writedata
		sdout_address       : in    std_logic_vector(29 downto 0) := (others => '0'); --      .address
		sdout_write         : in    std_logic                     := '0';             --      .write
		sdout_read          : in    std_logic                     := '0';             --      .read
		sdout_byteenable    : in    std_logic_vector(3 downto 0)  := (others => '0'); --      .byteenable
		sdout_debugaccess   : in    std_logic                     := '0';             --      .debugaccess
		sdram_addr          : out   std_logic_vector(12 downto 0);                    -- sdram.addr
		sdram_ba            : out   std_logic_vector(1 downto 0);                     --      .ba
		sdram_cas_n         : out   std_logic;                                        --      .cas_n
		sdram_cke           : out   std_logic;                                        --      .cke
		sdram_cs_n          : out   std_logic;                                        --      .cs_n
		sdram_dq            : inout std_logic_vector(15 downto 0) := (others => '0'); --      .dq
		sdram_dqm           : out   std_logic_vector(1 downto 0);                     --      .dqm
		sdram_ras_n         : out   std_logic;                                        --      .ras_n
		sdram_we_n          : out   std_logic                                         --      .we_n
	);
end entity system_sdram_0;

architecture rtl of system_sdram_0 is
	component system_sdram_0_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component system_sdram_0_sdram;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(29 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(29 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component system_sdram_0_mm_interconnect_0 is
		port (
			clk_0_clk_clk                               : in  std_logic                     := 'X';             -- clk
			sdram_out_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			sdram_out_m0_address                        : in  std_logic_vector(29 downto 0) := (others => 'X'); -- address
			sdram_out_m0_waitrequest                    : out std_logic;                                        -- waitrequest
			sdram_out_m0_burstcount                     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			sdram_out_m0_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			sdram_out_m0_read                           : in  std_logic                     := 'X';             -- read
			sdram_out_m0_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			sdram_out_m0_readdatavalid                  : out std_logic;                                        -- readdatavalid
			sdram_out_m0_write                          : in  std_logic                     := 'X';             -- write
			sdram_out_m0_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sdram_out_m0_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			sdram_s1_address                            : out std_logic_vector(23 downto 0);                    -- address
			sdram_s1_write                              : out std_logic;                                        -- write
			sdram_s1_read                               : out std_logic;                                        -- read
			sdram_s1_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                         : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                      : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                         : out std_logic                                         -- chipselect
		);
	end component system_sdram_0_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal sdram_out_m0_waitrequest                        : std_logic;                     -- mm_interconnect_0:sdram_out_m0_waitrequest -> sdram_out:m0_waitrequest
	signal sdram_out_m0_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_out_m0_readdata -> sdram_out:m0_readdata
	signal sdram_out_m0_debugaccess                        : std_logic;                     -- sdram_out:m0_debugaccess -> mm_interconnect_0:sdram_out_m0_debugaccess
	signal sdram_out_m0_address                            : std_logic_vector(29 downto 0); -- sdram_out:m0_address -> mm_interconnect_0:sdram_out_m0_address
	signal sdram_out_m0_read                               : std_logic;                     -- sdram_out:m0_read -> mm_interconnect_0:sdram_out_m0_read
	signal sdram_out_m0_byteenable                         : std_logic_vector(3 downto 0);  -- sdram_out:m0_byteenable -> mm_interconnect_0:sdram_out_m0_byteenable
	signal sdram_out_m0_readdatavalid                      : std_logic;                     -- mm_interconnect_0:sdram_out_m0_readdatavalid -> sdram_out:m0_readdatavalid
	signal sdram_out_m0_writedata                          : std_logic_vector(31 downto 0); -- sdram_out:m0_writedata -> mm_interconnect_0:sdram_out_m0_writedata
	signal sdram_out_m0_write                              : std_logic;                     -- sdram_out:m0_write -> mm_interconnect_0:sdram_out_m0_write
	signal sdram_out_m0_burstcount                         : std_logic_vector(0 downto 0);  -- sdram_out:m0_burstcount -> mm_interconnect_0:sdram_out_m0_burstcount
	signal mm_interconnect_0_sdram_s1_chipselect           : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata             : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest          : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address              : std_logic_vector(23 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                 : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid        : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal rst_controller_reset_out_reset                  : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:sdram_out_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, sdram_out:reset]
	signal reset_reset_n_ports_inv                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_sdram_s1_read_ports_inv       : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv      : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv        : std_logic;                     -- rst_controller_reset_out_reset:inv -> sdram:reset_n

begin

	sdram : component system_sdram_0_sdram
		port map (
			clk            => clk_clk,                                         --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	sdram_out : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 30,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => clk_clk,                        --   clk.clk
			reset            => rst_controller_reset_out_reset, -- reset.reset
			s0_waitrequest   => sdout_waitrequest,              --    s0.waitrequest
			s0_readdata      => sdout_readdata,                 --      .readdata
			s0_readdatavalid => sdout_readdatavalid,            --      .readdatavalid
			s0_burstcount    => sdout_burstcount,               --      .burstcount
			s0_writedata     => sdout_writedata,                --      .writedata
			s0_address       => sdout_address,                  --      .address
			s0_write         => sdout_write,                    --      .write
			s0_read          => sdout_read,                     --      .read
			s0_byteenable    => sdout_byteenable,               --      .byteenable
			s0_debugaccess   => sdout_debugaccess,              --      .debugaccess
			m0_waitrequest   => sdram_out_m0_waitrequest,       --    m0.waitrequest
			m0_readdata      => sdram_out_m0_readdata,          --      .readdata
			m0_readdatavalid => sdram_out_m0_readdatavalid,     --      .readdatavalid
			m0_burstcount    => sdram_out_m0_burstcount,        --      .burstcount
			m0_writedata     => sdram_out_m0_writedata,         --      .writedata
			m0_address       => sdram_out_m0_address,           --      .address
			m0_write         => sdram_out_m0_write,             --      .write
			m0_read          => sdram_out_m0_read,              --      .read
			m0_byteenable    => sdram_out_m0_byteenable,        --      .byteenable
			m0_debugaccess   => sdram_out_m0_debugaccess,       --      .debugaccess
			s0_response      => open,                           -- (terminated)
			m0_response      => "00"                            -- (terminated)
		);

	mm_interconnect_0 : component system_sdram_0_mm_interconnect_0
		port map (
			clk_0_clk_clk                               => clk_clk,                                  --                             clk_0_clk.clk
			sdram_out_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,           -- sdram_out_reset_reset_bridge_in_reset.reset
			sdram_out_m0_address                        => sdram_out_m0_address,                     --                          sdram_out_m0.address
			sdram_out_m0_waitrequest                    => sdram_out_m0_waitrequest,                 --                                      .waitrequest
			sdram_out_m0_burstcount                     => sdram_out_m0_burstcount,                  --                                      .burstcount
			sdram_out_m0_byteenable                     => sdram_out_m0_byteenable,                  --                                      .byteenable
			sdram_out_m0_read                           => sdram_out_m0_read,                        --                                      .read
			sdram_out_m0_readdata                       => sdram_out_m0_readdata,                    --                                      .readdata
			sdram_out_m0_readdatavalid                  => sdram_out_m0_readdatavalid,               --                                      .readdatavalid
			sdram_out_m0_write                          => sdram_out_m0_write,                       --                                      .write
			sdram_out_m0_writedata                      => sdram_out_m0_writedata,                   --                                      .writedata
			sdram_out_m0_debugaccess                    => sdram_out_m0_debugaccess,                 --                                      .debugaccess
			sdram_s1_address                            => mm_interconnect_0_sdram_s1_address,       --                              sdram_s1.address
			sdram_s1_write                              => mm_interconnect_0_sdram_s1_write,         --                                      .write
			sdram_s1_read                               => mm_interconnect_0_sdram_s1_read,          --                                      .read
			sdram_s1_readdata                           => mm_interconnect_0_sdram_s1_readdata,      --                                      .readdata
			sdram_s1_writedata                          => mm_interconnect_0_sdram_s1_writedata,     --                                      .writedata
			sdram_s1_byteenable                         => mm_interconnect_0_sdram_s1_byteenable,    --                                      .byteenable
			sdram_s1_readdatavalid                      => mm_interconnect_0_sdram_s1_readdatavalid, --                                      .readdatavalid
			sdram_s1_waitrequest                        => mm_interconnect_0_sdram_s1_waitrequest,   --                                      .waitrequest
			sdram_s1_chipselect                         => mm_interconnect_0_sdram_s1_chipselect     --                                      .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of system_sdram_0
