// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:59 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iIlkG0sZ2LlU2Z4uh11mIRok9q80Z9AePzm6B+TZdNQINS/FePuBBjDQ+uP79db0
Ed+WEvaRyDvV4HEFmhIjws0IHBPj5KUyhMt4GgvnVAtk30QhEyCINoxqPgHpAw4s
moVxhn8xK05ERqTzr9TAGiy0S4K9rapxqsBwximTdz4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8256)
2rE6M4Zsm6ipJ1QrUtfWYYA+ulU/jB6aBaeDXg20yqTW4xa4B8CrmVdYkdK0Micb
dea5/tnPCcE9s3lQX3zF+OD65UAjJgAtPDlivYUnPrtJYG9tkUdocIMG4y5VnUDm
ri1raXm8P8PYbibjMdPsdoqAxYfJll+zoNu7+CrH8tnkRL2lJvwilTiu6WbWyJrp
C7RNkTLu1ZA0eRcmFkLFVcJ5/AF8jp0cCHc+xTCpganXmbO83iYFlAjgHJxgpx07
EWNEtx7iRqm6jLW/F77HsXiN24WoVNb83TobnwxOnPRYT9naJzV4XHoLgDdaP5JW
DVl5mCZwx6uTdvKCh04IqM2z5OIL688/30pgFiS8Uyi7K39NxDSF4xPXC5vfrk46
KaNspulUOoEspsFVSzl+yKX4vmPZHkSpo68hGw9i3S2EHV66SMD6oVqdSmY7tDrO
ZtFKrgYa5Wty4rtuvCxAVcb9afsX+9JtmjzPNsvSErnBYN5Ynj3LuIcsE/xUG2CC
TxxWZITerGpNNonPIXRHN7YvWR6a/q9uxkd4O/oZNznhRF6HzixIxb5fGt+6AX4A
jVVSgndxJckd5fIL1TMjOYYs9cMQEVkAIpdlTBOYc8e1OEfas64YNBMfmzeIQqll
/RvMB0poEty8ZF6co0u+Qjir/3zwvU7hNQAkwEPiqZUjRJl+cR16dEWIjgHfYFIg
PmjmtkPCfmuH1KFlMuQDSYuyqvTyS7oaIbhQqhKHai8z/LH/gaDZRmRU+AnMzmV5
8RvFw1j1aH9J9eseY3yU6+2eEYnpJZEXe2sxjqrA/CKD9LxqDWVQaVx9EjzBCp2S
hQ40HBemNRVmUAzq2ffeGVWFmm49kl8FiGWR/FDy03TToqQWAzjlfMyS8DhtyGF0
pJlu/QEJlItISFtxjmmae33dccWUqNKVWYofGVzdZGq6nDlZqSrBCwfMIEKtschH
krcZZAvL8+Vzww7xcpaGOkQMM1fAK4dYgzm+43KgwAGtZdJ3AimPf2jOHIfuYY93
98H+5ysX+A+t3oPPcmkI55jKyhzxBe/d3v8VhtkWBWZbNs/rGHGVbV8qSA6AHz0j
ulW81oX2UkytUSRb5bvIEcBY16J3zbLWWCrjPCMbOzovJD7uzB9UHNfAq7o9hp7Z
M8vzi/dc7fbLkzpRxHeVKKVbenRNlNc6hvPNNkgv1J0d3TzT1GeurMBdzEHvu9fc
rlITvWWaE94lq7wOab8qa7unTZKANb64IOLmxNnThGGJPw9ozaP2rt5Yzt+p7tB3
JuNThlhvz0nOhzMGgFDikDilJiiQIbTEcWhTxTHJ/j5NKz0SPW00Akn0ib0HKa3a
sX3zziYC4QgFQVlBUHcbEbpKNX8cCn0lncynEDN18KOMgj2XhOG9lu6ZhtEg9nEy
e4CZTEGIp6Hk14YfdPY5QrTK1e/4FbiJ91qBbcsNVySDrPWvLuBVe52+mBa+zd3J
ZbgWlGNLh3b/eYdryC62flVWnOLRBr5oy/SaYTbJ2Tqieo6R3e1gA6zRyuBGvi4F
CZAVCwmbwKwYB+4JoyDA+KS4TXqYayHS5JmjkK5BtjxBfbA2PFHszqJVULUJWGd8
a6GdEo0PPHOQPwSUUYXOZxdQ/3kgobfyPDu33IcYQcT3H35g1uS5dJyXpWbBrv2F
MwVZYlOCU/FpdNpLqwbS+zxkwJlGKKpsYc29UmTM0SDjY6NGsknClNQJSwOCJuxU
nc7f5caFtY02JybU0/Wy6i+qpsG9hkoAp6RmAmHaYdxqWXULDCvs9RqqlRSotieY
WEjxeLNZAWO+B/IKJsEZ5Vq7YzTa/rpxV18twgKdnP3JpOSy+pVxAnGUiAEiMqn0
Uxt9dQHM7xCad6c+RTBOITPwUYBfLgj5L6G6aJwKikJs3vBa4dXKIrac+ojwYeYR
0VjlSeGKqOWr+TnXZZuxqii1CPcfPDPzAttOvQMkUdw99s3iVvmTlrhbEF8Cog2k
5cYPHNxGjqK2VRU24SCx1AyKsWrwYKK/SZ9FF5o4e4mFrAHvbEDpBILIU7rSMv3q
ibQcQrn+QzJodYuOW0Wd7EMj/4EYR9eRyUCuWznW0m443Fnx346bceNLvOCuLxMa
i2h+JpUqhL6zGXL75pG+O7YNWOazxkWP//ofWF1hmtUdfvDq4ktBmuOxYAh6pGKb
36LW3kYl5xe6fGiQ5LFNmwOW1vHZKY/xJv4Nd8dk9HS4hMQh67rK1QpcC4rAZaqO
Aiy/FlQ/ow1FpC/03Vz0kJNFwVf8WqxG+lrTG3TBbe2o2tRAoGdAE0fLFR6eWDt/
50MCR5rQdzKlZNczGcSstjV3SdglOmY90swO8ch9Kco8kjBFTKLXFLwfC1fsgblO
kIF+eq6Hp6LwowQYntKayfsv+lHTiIjUdhZwLvULSmIyvkj2b3JsxLHPJKpxJtPu
GV8iVx7VdNa4dUVF90eoEnMsEL0Q5wLJKwIHtJNbvhEQQQqMhBVwFhcvSdOq1TH0
/MMGslLd0n4vmQ9oS2hSKBMeIbdQsL6XVWwDbm3PlVXj6CprvOUfhLp1j/f4Dg3F
OTDmhhNZLJ6sKa6+w1gA5vTGLlp7RkZJiYUhzzYiU7/kvtR9Ib9KjZ1Vy7psXziJ
CRX6UVt3Ab28Y0bU8qM6KhuRq1Eqr4bMHvHjiHT1YhOfN/48g7UFxQUxTDfTKtgr
y28QRP2XT2LRAIqH8STRnEAdgET8Fy5YM+itzq2PjuNcC+DBg3ImLoiJMbiUxABb
ZXMTE6rndO9Kr88ve1XQjwE536wPEoY94RLcBMm8r7RXiQvJZYPbMJbj2EdOSkAw
J38CUcmpiOsxSJxa7Fjz5P6oHLDs3VFcb1F2pgpZVryAH2nrHtqJPukuJjo9IFv2
QrBW9VXMf1Gkd/DZrQi4DNy7RrY4vIRF9vI/sh38cJhGp8Iegen/AmVQFy7PgDhP
uUYE8V5794CrZp65A2lV5vm4IjuHHvdGzzB1l+w3YqZ3W60Cwt8JrU7OYHROK9iQ
UCStZlM5+TDvoqJlIB847pSDQlAw6yqXzOJSRnXswZkPx0WcUiOw8Pd+AEx4O50w
Ia161VTe/+i5DEcm46XmEsF9ZKqcHStjiZiO2VLqK5siKG6JOSAKbeKdXDhdJ9G7
gU9FSjXyCEDbWteK3tjTC0WPvPg0c9TCoKarhnht/q484wkNX10IdcK8ceuR2k68
3dARH/GfDbFLx626/g4YZBqXGUnUDJPsik7e5kpaHuP+YnMQ5D9WmBqSmcDQL/Qn
ozCF6uU8CEwBTqHUrq8lcOdwnkzlIe2yJp6phCxMQAspntXZhj+4WGLj+lx5eq08
v/VsMH7cEJFohJOcDhjb6noR7TleAxK67YPqX3xp2yLRE+Lov5iwpQBhJ0T3WwjH
Y2SmGzX01UeyDtCbvvw+l5naZzQLrD9Y1On/6Los99qIxTA+nFnGiCuWk5dYOJ+1
87aIoFhcZw8AfOkiMHyjJu8mhRAUwAoODLYyFB1uhBWDglaOPxxm9srxDAA7Hyrl
UZF0K12ojHA7ohhgLAtGmKsv1mEto3i1LqPpDJ2SyDXU4n6tF/G+zJe2IebQ+WEu
zZFBu69DyHrqz+uA831CTaPGUQax9mgY53peWd6amWGVY5LjEsqPTFU1UfXBQ56t
e4ZICJGj0UI68vCRVoixhciZjnVj6Ki/0fSTMkxklLQy5Fno6KeumTD8jkdEAlzg
kzOH+ur0NEgM1BcTAe8xa72FuiqaBkLbAZKW4RwFp/oQkB3eRY38WyJD3XFVK/Wc
xcc7ZUQPnaJK7A7lW3mIXW6kLS7Kgh1t3xqzMGoAvfZhZaz/XDfSxv7H+WfkB3BF
1rEiHYlyoQ+H0Okh+vbWHjTI9Rw9wPRde45fMQ4psDkCZmZN3lHv2yan7uNZwmFM
AbWV69yC6NnscJnYDWaTsECt8Y/NqtXLXka3X0k64W5SYoOkDzF2Qs7S44+4TI3e
zy7CIAXlR3eLllTJX/XVYIbqV7vi6zIm1vINstYyENCjyp9YmEhIYavviRuSJiwM
6E1tzEr3dMeMLbql/tJX3EzkyR5q/HiN0ep7iOGpCedFBraTa4GG50kAZxNL6I+z
Rh+JM3qOYKTjId5vihl4reMM8tuNrKl3lL4u4tabESKP2tZwrdjcqhehj9bcEpTz
4tUvXY562LNKCzBISqiWONThDDSc/LD8DmjVMQ9raAqHq6Y59T3UKLJCXcDEGOk5
PCnvwqxDeyk00yFe5wxyj3UGxT0fMcXFc0MKGtgZXL3S1FNDexhu7n3VtCStPD/5
geTdTK0b+OIxpTDteAuhpv/uKTFk/bcNq8EH0onoUAKng5SZW/lyHB4Z+2uEHq3B
QcrG5IRCmYTBKj4e/hX2hvL62JJqzn0zEjeDVqMOLrykwFWKB6e4aAYPzT8aPT7b
KmlfTsi21nkCeMA6JqVuGovRtMQ2DoX73bF27c7mdFLAfYoLjU0qAxeJmUDDo2n1
mNOCGUCPyn7AK2I6iQXJUeOhoiB8/8SgmleBbqa7qIl+chIGZazDYDdS+LxlE63t
M4DCLaw3LkJmtaQKp38wyf0kkyuYpBvbZOyPLd7Ofdfb4r9LHd5dktNCDQsnOZWF
J9cT1VffgbuTcpqXmX4K+kO6cEV5IGnCMgs+tJHdqB1qna/soWboSUn7LDX1Ydn+
AmvTju/qR5SKHpDetphk8MKhtRJTzCMkYMd/YFb70ONp2LnGDQep9n3HsCkKvDvh
Ufjf1jvrfCEouZGAm+w3UoK3kZ0+CbZKVWQ6EISL0PI7v4Py4yJ8VisMlson0ZNn
qU4kEyyFjCVQ2K/rHOJC8AYrOqBN3+TxBFb5/5EBN7vBF6Kp7tB7U2IRT9vircxX
RCh3Gdw6lACwMpzaB7pf1hosXTI5BuJvELRZ2EVWUpNpt9WaJunwBTvkySBKAmzm
mWp2xUIcjTCaRp/jA0fYftauxfWCeYSjFf34JbdkFw/jUeGRZCfZ8tXZlP+ZMURV
V56QNyFq1czPopNOGqiJh5DjYz7tcOkDJaq0IowM1itF8np+xIRQUwJMkXzkJZob
2fY6wb6dQsKVGXtpl5Saca3h/xJClfhxCqD2O0OPnMmKovDNLIkmgUiSIYn3bp1X
4f9vxU1jD9tGIn0B2tEVUe+eJTiFtf1AFYZ4OzSJ2OOIK3s2hizACDN8Jz/Gg2bo
UgeO9RKW2ZAJ3v6xvPoYb7aUTVTlFHWGsM2X/ClE6aGivUoRxEtJIF2OhBaeJ+Xz
4rj55yIlhrkkG8YVpjW3x8/2lU19li47NcN3uNIAndF7kJVKF76tSfx6pi0Rw6qL
WQvo4OS760GcGHrJKPg/t8w28O1gOhSrubif8eWRwJsoXKds8rnQ3dTlti1NQc6Q
A6Si8deWzzNqndO33eCMGN28kGQfpQVhHZgXbY8Xtsh1cCtGpm6VT7WzyPZeoTGM
xcPDrOH86uJyTyiNYOPpHdGEmrps54mjGtDC8WKnqmcoOm8FHAQOYVum2Yi2QZGs
4RVif2JZYvx42WS3MFasZeoJJUYMc1kGYDyjtIxuu9lCneBNfdvX04GphG9d3Uqp
bFOZ5Aycj80o8eQDzZ461bssFI+zHKLCU0cHEfa0Qcj4WyeZVOoB7jd0v+qowWrx
iU5RxFATsHPUNUuOu22z52LfQQswXBscQuHJtWdf2lIlBGcCufLsY2MdJFhvOi85
mYgdCFDDgAFJDJ1ZnS8xWZAvi+46GvzQkbMeEuCArgJTlzSL8DFY7b7mSR9TmoFR
FLBgUvzpA6JO11014PYA8ifMhe3c1bDgp5DuiH4NS5K5USKT5EaqJv9nLsC++/Al
2E+GLqHsr+qYD07oINWUBPQx4+8QZlSGlmtFrVmApR3d2zO7suZc3LB/dXfauJJm
nt8F+38dsVnZ9UQzjV5WLFY0sRu3ggMw2xea6mW8BBWw9CWpE4i9JrwJCkLVaLSz
3bxrNuAcxiW78SFic/RIXfkhYMRuCAHa/Xei7R5SOGEtinBrj2bnXM/2p1QGRWBI
duHG2ZzDjYPnBc7pnf3EAco3p325tJ/faKBQziIklYp+cUZILwi0FyoltjHrL5Es
2sbT0T3ChoYt8zqAGWyq3T5MqjxdI6Y9c7LjxM6ZKy8rTY/q0/Qb/om/qhvna5JN
DEC+v4haVEy1r3PyYxxGA9PNMidBcjabPfaHp2gDpcnPAA0xK2P3Mrh6C5m1eJcF
nQXKZMsmEAPXKiU9MskVwC4t6GhhRRZdV+AnBtSuALSkKErrl92Y2piwCLw7i1A1
WWqxMwTwaGSxGHZOVKB3f6gE6Rd+Dp0U+iBlHvdSdMYSrYQ3zm0THRZdCPwGLGBg
ThAFjtlnOvIUpDVeWooSS/1K1jATVxlqXonnzvn1mLvmhEyXwv0H5XZ7bCR+G8+g
5mdWmLuz1B4Wz335jKRafGEOxRuFJtYVt1PZqNi1WCwsSkLd0OwOOdnNMoJG6DdH
oqesjf6YziFrJ74xHczdNjgRSMu/dvlwInKg7p1JOUyBYFAsFVbej/8Eub+suiOb
+W0UqWVZI41MHKXC96HtP4nApgHK7YkohuRZWc1FbCfWb2r5Q61X2O9wJYCZr1Jr
dm4PIbEChJ6Gxsgfls6gimN/qSuiDEAZZpQkXra2TehZPsUz1VOTqkkJIjcJUey7
fOlH9ilsZpEkyBXUhDPE6pJGkns/0Vd9XeTLZ5rMWLW7DGxOMsJyscTwcMbYnzTy
2sABKowUI5cV+ZsLKwaMkUvqxNy8QBRmd5PlnO+yNROr0+yOjQ2Pxo0HgZKkLBRJ
EQEdWJkpIRIa69I9FEH+woskOUVWnSzsGBJLH+/SQiz/M4SsbfNnIl+V6x/dOhKQ
k/KwX+DQCjkMIV8DALY43ldE8ufAElszzP9dA2sqyudo34dr5D7gwLUlyXqFeWMh
txnv4i1nQ7NOJdPpfypjymMzJivHFB6wSkll0zjay8DFi8IfULYHXZ7f7FfL9uJS
1GzhDwRYgqT8re9ZMNNzNOfQeZl1jODBcwXk9qObTxth5nT7udLU/GcqLSfdjeuP
XHKNmhDBciOF+q0z0EtIV9UQCr2+LLRtk8hBfpu5apg8feY/438FAMYt2oZa0yQg
/gDYhl6TJbrV+F7Ouqj9YeF0uuQOr2IJcd8paCm2FU8IyGqiNDZ394Bi2XqNrkhY
g+ckmdE1ZdO6fysjs/ERDUm2JafC7Y48iBitJHTzz4TCFkoWFOkH4GlUXZ61pZAI
aCaB7JQEixSoePPEUefHr8IUVDwe3tdXq0ZlpSvw8NjZJKI9FaEWNztSf0uZLCVO
GIrczuVeOcd5YZ0SxOknJyjf8DRw2/vm/i46U0SFtUi0wB2aMkXzG19UpnDXw4EV
mdRoaujnWHY+G2LStifzp7XTkt0BY+0Nt/TGJpqX21M0+/YLWpb0Zr4hqteK1/0T
T/wgZN1AbwN1Hxd0ZlrS8RMziiwz/XCEtxRHEVmbCOPyar0ZylIGPKC7JRwKk8Er
9UWWsRarQG1BckRSNnxYMo0fNd+ilYQUX5DBhqsoR4KEA6ljEIxjspYMmS1O+WrG
cwRtbE4Gl99KyHzFzJgL+b40az4voBgeYIiPoZuVM0dR6zGamUtG1CFbaAshM9DK
lw4xmeDotaEE96E0I7rFSGPAKX583A08KMEOgRiNmVQM/NOx0kb9p+yY9Qy22OSW
n+udZzqhqLlcHx79qSzF6RksRdC58KXGSoReGzqZSrFg/gJNT9alPZHp/blRBJU9
feZS2gA3924aQ3GKFClQQvSIOfJJwDWXNZlQvyzHTrx4V/TqdNz6nSugwTSmLSy4
FbhqehiWFtd+cCDm6HjpBT10Kk87oD3wD0tb7kLy3wFSH9fVHF+nL58Y20lE6uGZ
5eTMHxwgE/hG/MK51Ud9MDiCEIqWj23wJAdkiOeJzgIozXbqGo2IihxvLk6mCD19
dlKUKf9Xk3QYBczZ9kcnceBwYYlrapeZDMctrYf15oN9JcsJqDTdpO3lVA+HuKIa
v2u4xTX3oCn6pLrJUSpjIf3g5HH9T+TaMZXR5mDnsbKTzAfgklfKVmldETyaM75s
0iAFqU//OQTQcjB2gNOwkwyT8hONR3DqCF74olGGcN/gWL02oxbfDxFYykrdgOlV
QhnDpAWyN4VcOOvEzEIrZRmYZj27p9xcm4mVcLQ1QovQyPFPHLxUOmn7ilMS3kgJ
PXqA45EHYYrCQtjLxPANY9eazWiKG2s0ekzQfu2VIuBpxcPFIbBMr5fJR/PgwjWs
mQA4w8t+eFUNZaZibaR5WIWrNcBrHVbVVPdD3cYnEbJxCTzZjQIqGBeZUGaKNUCX
old4iZqKn+pkE9eJW0AOj7xtHSBqKYSt9KTz/b3mXZZDos+qpLZqG/j5V/Idn8Ki
guHkeXp5wxUL5BCRNiIN/KVKXNpDlTxRf27eulgHxi9qSp6T5ycTw+gpPYVkWkZU
pHqi34rcz3aeAkEIxraC65jvSAWdRKE4a8r/jXwWgVdSByceOE0ADgMcOGt+RKnW
TllWg4K8yTcYhQoACWECCn37/oCxEV+EsPMo3cGBo+0cFzMFeYXDPM6V0NscILqn
5rUtD1cUnYAETTRkF6+9fuRBdax+1pr7EBrGtdKlKEswl/Lfn3FovanG9koeVME2
iIAs2PvyE6ApDggI828QCCn1gvBLQ/ZSWTCu32LYP4GCEdWJLoFK3UL9civWW8qm
wjri/pv9US/NR/3xNnG1kg0MZ4r4ao2eJAyt6dVv7v/3bQqReqPE9qBL5jfzPYkW
8Wra30ObkviknJdxa7/IsQ5dVTAGZlZL8smgg2n6zq+ZA4rkR2R61ejPOmy6HZ3m
5AYCld2KiaW9BsEkdivbsRaG7mToaZWEyVlBicfxxgkspuv/mGiuGXz+YToHSXkc
251nEPAnOm5K+M0xq+Ak+riMTsffE09TAVH6F4ndtlLAejgwIt6qSsPrlrO3aNLk
TuqrHWa4hSYWSaAA24lzlqLaDHrqQUx1loN+o59uHOBzHaXP928ceS9LGy58kPrD
uf83TLaugbWGFRejH9fAVDnfNQhC8Yow4+ikywPkKrMiwBY+ic0WzAURQp7HRT2G
Q83KhM9yzK9LgByrV1Dm1sqpdiOMYLPhFDAGxm+QgpVJG1eTbf2syOzLWUf5KXU6
XoNqdMX9YQAeQNDaESzBAgSKy2F5SnR3Npr4HNy4OpVdmJHZmL0tFyGEHlNFrV5H
xkkwF3APVusZ3UpARvAShJUP039mYFCTiCC/oXf0hmoWMNAkI5uh6mcKe1+WerlY
+IOY2kSPz29/eRsotfhSZlRigJyWC/WIbVP638bR0S86B24MYPJwtAQBYTv4kxen
k+rObhFDsR0XxQRcNVYvnAhkUoIVkIqM2EvYvmufpm8n/74iky3wjbPkGTHKKYWI
MwO+7cFILU/6VkvQrIcXSyJcUwsGN6mOpXyJsNtDx4OS8VDgLQ6Gzn8obmIgQq+E
3C3IQRqq8R6XFKYNnBflDs9QmM/oRM9/AjvRc/a84Ntf/+Tz+qeUt5f6VRLg0OxO
pa7zfiSqXM4LAjNdECbXGk+NfcvwuZuOYou9PGfAYhnkIo+6iNreeQCxfww2Xqgr
9NqvRs62RN3DiiOJksoJYbQtjRpWJmaafVmGk6bnb6X22V2y6acAM77+OwWj+7CN
4VmqO35FZYZiQZyf1tHYmtiJhV+DprIWLkXIXR3qXSvMYfdbiu3ttd+0MrmuddLJ
NJhjhigtSXmc8i6xsGU86fDWcU1cc95AsLS3OFa9PtMJ1FZPqgndIgY6JuLYKk3l
BwDur/eksD4q+BW8LgpgZ50pryWMuuc74a3l6ZuEMSZVaiOtHbgTVdHkQNqmgKEs
qhdDg3YLxTG1hOl5ZYq0J0GAYze6WgqSFifpE5Hhbv41x6fadV2zqdzCxjWYu8cA
LoPiam9iCvf3q17RoPTS8wywYP2IC9n5N2OZQxUD5gb11NWh35WhfG6ZDOhEjO1+
QyAq0++dwol9wOxCiDtVs0dMokp35MXp6Zn/YL3XzrCR9rwM61I2a3x0g7sPgGL5
0TIGe6iF9LC8JXlOQSnxg2pdDYMhtIpOA6f3jFx8d1LdOR50u6yH12ZnuwLCsWyd
YVqNHGh5hrm8oXz4WYIQjD/axDhh5vsSoqqkLWUrkS6tHsg3l3W6zC7y19yvrfp3
hFFr71T5ufr6bUINC2Joa098yURplYQkgEM1xijeoWbPQon+9UbrhwQl+vivRYji
QLsQRtEIxFzFL3KPYWf8ixVR25my6q1EVxUs4GqGyvrJJpmx7XeCQ2X44dmbSfmV
tvEUlN53gKck0BnVHa+tjoVn5fkBfkQSiPIFaLBylx75wmeT3/S47xK9OxUvkmv/
u5dzOWpdZJuGi1cRFtxE2BWzhvXZ+Ul+31q67xfJcsKvh3tUu3ydwYVW4V0/ed+1
BE7MDALr7o6got3n8GfwpBz3RCYTpsMPv30YxaYWNgTh8fqWP9GEYc8jZ/MuaO9+
zSd5enQdz81+Hh/s6Iw8vQittL9jE2R7oZ8DIIkN+dn8kwqXJ7Ny4Q7b6eC15Tzi
WzB0SLbljmXEvYNuKyIzHmkxG7BO3ww+//R57YUb2CN2aLiR0fpO0zRWweNAacC+
w7K6tU0x05hf0M8xvBJ1ZYCyvqGbLkfhWP94u0/DlsgeaR0m8ktl1TEz4fO0vop4
SXkG7KRWkrsoWCQPgwiWxnBCbZG0mw7Bb5Yqmeh0oArpviwYq9Nvd0eatu2dGWxL
b0umZP+8ze77i3bh6gQYtiogPn8Y5pGs7eB9FhCUP/xeG588kkcH4hk2hIs9OKzp
GFQ/1UYeC11Nq72f4YSnQRX9OS/6clLvbN/6kdLQOA8GbWSVz+Zzyv5PthB1JomS
EM7UfhAvlE+3N8jpM8fi1GWYXE3ViRx2iqofWkHAKX1GjjQaGJBL/2v+cBNHGBz5
t5RO2xdMUone09yz5VqmmJUTMnmrlNCQ+3Z5ElHRyzNv/WVUsr+2I01SOvEHyaYa
`pragma protect end_protected
