��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����Ղ�ɉ�%����r��? ���Vz�e�<j5�(�X��J�@Wu��f_<;�|'���� ��5�*$�����e²�堇��K���ѹRШ���ǽ1~�;�JV1Z��e��h�]�5���� T���f"���Bˊ������w���WV!�4+���VZr��U��3Hs���' �`]B�	����F�Q��#��;����nm����r��Q%�y���8(ZK^�������BN4V�W���`yS���	ÕF`�+�4T
��M���}е����(��&��	�rhy�Y-@@�d�@�z7S��1��{d	��Q��ʵ�P�P^7`�F�#�s��XkI�r6�usM}.�ЩB�˗�8Ȟg�zI��u�V��(�X\F���T����o�/��L���w��J�İ>un[���W�,�.�:Rzs�����T^�z��S~�4<��s���
oO��Ueȍ2���¦�I������ɕS�Uـ;�r�8��F>�%G�o2:J�6<&I2�����А���0O�h�f��nb�Y!�)��`/p��;}��E�9ғCe«#�X����h�����0�k�V�nQ���
`�3T$����� �l���x��u�j���@�&���dא[����� x�Lq	~/҂��^'�BP�x��z"/�.W����'�w�1u�������pgŒ-��,?���JS��pwP?|�2�V�Q�	����٩�K �ƅ΅�R@�����"$?�
N�͏�P��s��j����q��^ij	�v�*��C �sW��U��*Ǻ�d@��]d�S�SĚ�"���`^0������ŉ���LI5]����e����I|xl<�+y��G!u4Qd�:i�uRbM��� de6TJg�^�mCZ82~r|�HoU�ay���`�R��g��k�2�tz��4 &sP�#]̎28��X�W̥�g�s@rq�9���.�Z�L�8M�W-Y�x��s+���*h��T�1�ǌёh"��4����w?���#��$�~F�!�ыB��~�mKxQ7�!V�!��_�@���':m�/��t���9�u�"���ɶ����&��5��Q��� ���F1��Z�k�E����%'��}��Lx�pR��:2Ŵ&���A�C(�:4x`D�W&�2��k��+
=�Nkw��3�'��~
vlx�T/A�n�Zjh-+����Ȼ�s28\���C���SE��b��M�-�#�0_���3M��e��?��+����B�MV?Hak�oDk�g�c��w#�	(�v��э%ͧ�Z���Bɦ������2=#o����.�O�bx����Xk��3���Z|/ br�$ch�"��y����Fh��(1�Zl'�ˮ-�9��W	�F	�Õ�6��?�l�Xm*�J�s/�:p���v ʜ��B�-O��00�v�M;*J57�G��� r�K�(M��.u��m��o�Ye���C���u�9qri$_9� *�t�؃��QW��������^B$�e�?�%��uy���S��_�٭mo�S����gv�e�Ej�Y�gW`b�}Ir�(�FX�s��pɉ�{����vI3}{��pP&�F�' )��hUӈ��Y��^2'D�(W����Iq	���c��#/k�4\!못�8�$�&ޚ+�����[���м0�3��Od�<E��7A�����%O��܋��A�(�.�K(�;��`Cd ��� bݹ�/������ւal�����>�FmZ3�?�>�}�i��uL�K0��4�1\}?T�-�jjL�FF�e�0ߣ�P�����OI����>��lA�o�p0Yp�;�ƌV�{9ͷ �i��`�����T��8s,׻!��z���j|HP��f�򬀒�Օ~W���=��_GUMu�|a�Y�� �b�Лₜ|�k�X�o�1����8u��)��k[��߬���ζė>������H8`��V,�#¹�f�'ްH����9�B(��
�k��}ZGw(l�l�B=2&D�53nwN@�7C@�RPU��y�"�*[)��[NM�וń�tdcf��ۃO&�`����Ű���Z+�D_K�z�hx���8&
�:����h�Qn�����n�o��w\� �0�;�^9ʄ�kU{;s3\>o��o�`Ĺ�9��ԕd����d�ӝ;#��Zu���@(?��96�wZp��2(N*v�Rfv�z�Yx�o�HjUH�m=��(%��6#D�c`ׇ#5+abF`t��}��-�N�$3�s�X������g��\-�� t��Т�$���<���\�\ʀg����q �0��Z�{�������@���N���9�6VE�IZ)*ȵ$M��/`v�p�Kw�*��K`�t܉40�s^w�	�ڞ��|�y����|Mw�|�i��&�b�W��W����$���X��/�wP��t�� �(���U����!�M&z�F�1^G�%���
��/���L�M�{}-@\E�=}�ǡ���4�̳Gt������IO<M��#j��M��\�AY�~���z����Hs�^�9��X G#n4�'[m쩲f�$�z�e�";,StP8 Xx�s��1���b�wh6��|6&�/ߔ������'~��4�no�?��Y�`��tX򸕦��FF���5��������`N�~#�Kj`^��!�ԧ�^.0�U��q���q�n��롞��<���,2�!�!��вdt�wH�B>`���DW���8�,Sy�&���A*���殍��lm�Lu�YlK��I��86��_}�Ma猪ĭ�^t��|=����Ks�m�/������E��Y�{m7�w����5�Gb҈��IV���9���*���.�w.�S���"eL�.�N?��`�]x�Jd'��1��[�(V��M2㬒AK�"#�[�Ώ�a$+jĶ�@�91h�D��4{�$�Q����p�>�^�_�z�s�'���~�˯nn��=7E��M\��乘��=���!EWo��c�Z�{h�]�<k��%�9��B�]�E����B��Oh��pu֎0�TmmWP�r�gpG��d]f�\�J�y��l�̮�%&zk�`��@o_�ܨU�N��>RO��|'��N8���9<0���[��3�6�������_Y���Ǿ�0��B�Y&��J���u��ܯ�U.W�(��D�ޛ����Gz���&�A��I�0X�bo���cP�Gb˰�v�d���@D.�q�o�D+�_���rY�d쀓��[�S��z�&�Hw�3��0�G�b�<,�@�I/���k���|-��/F�:�*�t.x�I�D�R�\��)vsҪ��<��0r�����0��ҙ?L/ҁ�x�Z�6U9&y������ M<ۆ�2qK�X�ڎ_4�u`GM%��@�*���e:�Id�Y���_���H��R��lJd�@��h?�}�u�d�?*u;��t��B=%�p|?��#�|]��jo��e�_��d����M���3��!��#EG�H��7�A���F�-�]�x&���r$�>�fy[�m{.d���yr��h�d'yS����B�s �f�NZ³A�fX:(%i��tyZ^�o~�G��� �K.���;��v�P]�7���3kxZR���C�I���s��+fW`�rs�B�y!��B3�to�㷿�pIu{�~��f��'k�����X�:��zh{�-&����5��'�p �O}�3R�矖�=�Im���eP��`+g�,�n� :=�E�,�0��)��H�H�;��D)	;)0�	�!=��ǟʑb!��6f+lX�;��rn�b�e�mX�e�)?����J�,7�+D7;j��)�~�`XaQ9T1��ɫ�U����X�z�hIN
ۮ"��vײ���Y�^��H����uC�&���l���-�ֳO1��n<[�a��ٸO�����j1OL{�U�	�Ks@^X���V$��r��i�/����4"�e�CeX��6󀩃��e� дX����sQ�o~�iDZh��Nk�gd�_{�Dc+䭴Z����އ�'{�	(�3�<M[5��hy������7
�xU��L��˘2j �o{�dP?i*�͜�W�nA<�~�����B�0��9�����<=rh�l�\���cW�O�l������p���+�e�/H��z]S�P�����#�m2��o��M���Hd���K� �����%|�S��E RnI�y[%@qY܊
�8_�S��٫b��$KA
CeLĀn�t.mx���dƹ1�_��kn(*�Ƹ�������UU阂}|���qH#Xa����Q%��Pd׹#Җ���դ�8�Ҧ�P���`+�q�<d^�Ŗt��B��Y���[�����O�-�E9�;A�v��ɴ�'�Ջ�>}
	8e����3��Jz ���r%��!��|k����'�]��@jw����n$�z:�2�����;(--݁1Z�0S�C�2�0'߆O�k�=M�Ŋ��"��H�3��=T��֔�~d�s��2�ے� ��V�bR�s���f�f�; ��~Cmh��v'�Tx����d*p��%�V��>��q��Q�V����+y&３o���m��لi�Ph��>ڦ���������%>e�[(���$��TE�U�哽�*�#�����x�؍N.R�F��NF��+`�Q�ѐ��ךtR���5� �!  �8v;��x���ܓ3[-���_�p�h1AΙx>ɾ�
�<!r7��oݑT�����L�4��&�JQr٫����I�$! x�#�n���5��1�O]��mi�Ys0���r�U�#����~|*�A�]��b=/��P��(��ftf�����i~��T��Q�o�Sǟw��MTXN��!�<�����9�£�q�E�{J/���<�1Svu>�X/-�pr��kD5$"[��J}@Y�iBG����uYNF��A����S����cgle�({���4'\��_�P�[B��D�sH�Y���;�_h������׎S�6����Ş
r�cfթ���l�������3R����05?o�,��nh����(������۴�_i*�u��a�ޮ� �D�p��Х��yi���b#J.��ྴ-jW�K�QJ����wyz�[H3�O\0IW" 8<�7G���\0E��)`��f�Sim�巪l�2�4�i?`߸����M�l"p�(9�I`O�/��GH��ۖ)e&ZD���&z��:&w?�*������-T��2,+Xso�`����O�f�ւ��p�/��]�p��Z|�+�{|^Xm��G�j���zSۅ�]�k�$�m�(W�h�3Ĳ�G��ø�/��T�(bP����x�QR*�E4O��g
8;��2V1��3����<���OK���e�R~ٓ�Qs  [r!�:��aZ��(CC��>HSB�s�[�o�ޑ�N��Ex�����i���a;�)�����[򵈟�d���*�:~�G �������M���
��V�����pW�RD��7�$V�^����L������Ҧ�EL&H�_�����&��Z��y�9�^d?=���b��p�2�̂i�{\�I�^J��)>�k�kb�B(x�V�;P�9q�_�T�U�-��ʓ��~���/y������ݑd[�k,}e�F���$ڷ�^�
<7��:;Ō�[	����7����[�b��k��#���Ƥ/hu&/M��	�1�o���w$���X�)^x|b6cd�ϫ�6��ۣ�����[����;e��Zh�nwz�F�W%���=��(
�Y���������5t�hZ�y�ad�z\����Pw��=L�M��JD����oG`Z@n&/����>�֢f,�����M���̩U ƶ�m�t�Lb��^1������� �B�4���&\he��k�ٞ���ǘ�K�PXV���=u��H�����s���8R���d�s�CvǬ������S�?���nY՝$�G�~���h����H��(Fp���N�\V��o9@��\f��7�����~pl�"u�d��+)����Ir}��B�}�C��g��Mo�,7�>��@�M�D��`-����QpR��=�ac�½͈��Q�a)�X� 隤�u��Qѭ߮��^B>�;��(�毫�j�X��j0m��1f��Q`i�P:���h�".��oZ�?��d���I�_�H/+?���;2t�EJ�-�P����������I��O��š�¸	�̢Hl��X.���DϞO��#(|��`�V��-������;�#�����	�Y��2��.9~]V�?�`W�%t��Yû�����*����S#��
�c���Wk�d	�`���&O��d� ζ���5�.� 
��ׁ�4t��=-��fq;�Ӓ��~�(��cB�]�D��yi�*�}��xJ*&44<������7s�=�a0����ε@�"�R�w����m(�G\\�Tv["f �t��I��x_C��+N9H�f���:tF�����>�%d]��yT�栮�bGe�-	���1����r,�uu�I��]#�\.�=�������������/@< ��^q��}�m*W���^/�.Z�܄����t4��釞�lH#���"��$	h��$t�H���j!��6)�$}m�vA����9!=�Ly�G�6�u����Rw?�ueC�yR��
�Q��u��0);4�M�ڞ/[T]���pG�}�.�5�%�x�S�Y����C�L�P[y#!��ʆą�u!�_wv������S���*e�6g�k��mv{��X�/�v�배���1-��p;�)(���'���k��gkRJ9��ե�FIl�^v�Q��Po�?��9����ۃ�3V^��U��k��4�߹ё�Fh�K����(�>���&��g��yJ�x\hfc�)F��~�#�)Kk��npYp#b�=.sJ���tQ$x���I�[�d��T�}� C�ߟ���FB��sد�P6���+<;�cE�?��{�<*i±b�$zU@�Ȃ��av��21��皡c��,���T��&�ٝ1Qv#��X�O,�&q_��!�1bJ�ZO�RAF��F�"n|��v�8J��nE��A?��O��Q�!�X��hl.\�NZ�r]��ۨ1�kO
� �k/�<
��<�`�#<��ӿW��(��o���;�(*V���������f'c��KPrݔ��0�f�1" 3p풮�����y�YI#ׁB�e���KWh�a��~�R����ݪ��@�%#�2K�QZ3�nm*%و>ڽ�y�e�^��`�3�'�~�ǡݽ�i��8��>�����F��~� ����=a\�c��e�D9ο��������9�=,0GD /��gdL�&UD\.i�K��>x��e����VR쬮�����k7b8I����y����J�>����o��,��\��L�^1^z�h�ђm�x�.>�K-�O����"O���[�h��5Z��
� Wj��ꞗ��Ξkp[0�SE9��z�עvP�����[�TX���A �5�	u<W�;(bd�om�ݺ�4L��~�"'���s�8Ia�����
#K�z�d���B<�k�b�'��� �0�795�8	���[r��+�]��u�-��\�dAM���/ǲ��\���)%/�1.�}�H�L�2�؃��OP.�������MP��m|�{��V��_>,c�]c ��~���}��h/eZ�?��J�8�1��m��B�=�p61�2�5b%(Ǳ��TK+������CՉ$�9��͋�q7�e�lZ��Q_�"������^E{t3���ϸZ�|�K=��1r��U�Y�0`��:��,�fɒ,���og�����W���T[�� ?}W\�i�����(�Q���C��R�A��LԖt�p�(J�\�P��U�Y�VR�_����L/%�o�����Kj?,�˲4��	�*Y�\[k���d��|���Rć}O�]�_3��:b���=����f�&�C�w��<:��{�����/M���7��@���i\ƅ�pc�c7*a�r԰��*,��ض�pVG�(f@����̲�)�@=ڵ�Vr:��q��Ag䦲}+�4pfoQ�����Y�!w��ԹcФ/�N���2��Ń�o�8�؜�����r��R(���"N<V�6�TK"�;��'�Q3�>�]��L��A9� �Q���3�П�r�vS�I��J���CʗE#�8ߩ����N�. ޠM�_��|��HA�C�ǋH��^�S8eĺH�Fć'M�$��?��J���&$>��M��IG�G�����Ia&�iv�PN�>�N���\�QQP\{�"�1Mޅ�n���hB�^욘��lXx�.��MKt�!)�3���L���R�܆D�9`���Ha\e�;>GM�RV�B�LZ���&�p��Ȣ�؆CO�T9`.�oAц��A9�@���1O�q���X�\(������n��'���M����o"׍X+�����*�"�#�x�C�/�;�n����猓 (���k@��7ur��egF`cUO�,�5�D2A�ᚎ� ��h.��Z�!ԳoC�����f��H��<ж��.�Q�v
?"�(�}�u^g�S�#ݨ���K�TֺY9PTk��+�;Q	6����U!V�:� G��XV����܀%z����j
�.r:�W@�ytu��%g�%X�
	W�8f]�Lq�_�ˁC*�tRO���?�?A=;�����:ܫ�֗7A�9���v�0��σ2�C~ĳ�һx)��Kk��7�5�Z��o�L�)�?f,�
;2�j�·�f��d��	#J��� ��b�[�ބ�U�|}���>�?��Zh`����}	o�6��M�zI
����)�<��/��tͧ/��H�ȃq\�-&<����q���9Z���S�����>{֤���ܱ��EX(m�'��
�;_� 8G���o��V������p����clq��`�c���xe隼>ZjF�R��^u'����zGi�Ż�kp�_��:	m�
�ȴ �V)���h䆎%͒
vbI��o�����j��r���^���d��ƱG0<�H܌�O�}I����Ç�Mr!�OHbi�^:Z�>�EjO|(�Lm8�A�-���$AwQWS�`bP��h���(v#�e)�E��/B�����~&����ډ��)���(^"ő��x����{�ND��hqvJ�"^���ҹ��`2���#�X��q��T<�9��(��e����P/KU��Z���'{��ŧ������t';�(oߋ��C!{;J��@�n���97��P�[�5߻'���,��G���{��L՜A�Fݝ�:[���-����h�ye�t��ҕ$���]T
49�h!<�ڸT�j��yj'	ٸ_<�ar6!�+/䳴C�5"��A?O��K�AΠY�ȉ���^tc��c'G���)0��K|��R��2����g��$>�p��������*z���L1�-�K(_�N����A�t�Ruv*��P_�W���?L��y�vpkj�}uNd��'S,3$������̐�����[��:�(RI2p-�M��n�/3�a9��������N>�Ε��5��C�\}>a0��oʦȋ�ߕ��baR��ñUlB-����8m��(�� ҧ Ҷ�i
A:�e�i��d�7��Uvw�"|n�כh4�_7kiH�ڢ���Q�en��(�ǋA%�ҟ#��7~��O��m�X-H��Л����3߀�XM�1:���kUj�c�Q3)��
�nF]���Ά!{��Q~w ��F�y�+8��2��e�q��Q߬0����ת� �ӎ����_�	u�r�}���'���M��l���K�xW�QѶfi�����ƒ�W�$��VU,v.�I]�����D 6�� ��-H�.�������4������ x�#	�k�� �+ݻ^���KҔ�N��wBT�y�Q-�6f(w=���U?)d��N07��f��ɋ�C�� Pj_��&e�R{x)�+�('n�/����wduir�y!E0�t+�"�G���;�o��eC��e�>��-�4��u����x!sG:�Ǵ��F(T0�8F�^��aѴ��c�E:��o�@~���%(�������L�Z�߂��=�$��([�����DȲ+��{�/г7�~!����q�;���>>�ȹ����P*�a�����xQ�xӫqҗ(H}����1<6�� 6Y���׹��"h��坈=���o����1�_p�[o�iί����Y�BJ��O�$Tո
�Ƨ��½X�h1d�.u�ڦ�tU�_Ҏ��
W���Wp.��;Ӈ���h��尀)�IVF�N3��dk��Q �v�c�V�Y<&����Ѽv'��\E|g����'��������1
�`X�'�ۮ�l��w>�)ja���_��4��tB�z2�K)I|���mu����#�\]O�Ԝ�F3�n�Jul�ȶ4��-���__h�D����9A�Y��3���fn��O���E��ar����֨F!��{�'��&eƓ��g�,I������=/���5�����X�q��_+���=���9S_R��{b/eFth�W��c���ɘ��MyUt:S�t��3�.����ƔR:`�!K��H�%"䛮�3J��8$Gx� @�EA�ߋv�**�ʜ������2n�[�8�i�܅��݆b�`����YS�7�0v���gJ�Y�[C���B'Ŗl�ꏷC�T�iV�]�)$�n�E���>��!nĽA�̥-�#�7�/(�a�+��K�B���os]ܠ�%�HQ����?���w�ޞ~��*��9=S�	{Q�*�rJsU�g�#�lE�$�����Po���Q�TFA�`�<�q����(�V���k��Uh�v�|��	5R-�W�&���>��,�U��[\P)��X} 3d���3tj�q���	W$��|�L��IDVW���E�t��dTm����(�����9�G�zY���WC�,ߓ�e��tYcD�Z�=���eh��xW�QUx�3��r7����������(�u2�|�WW�<��z����RP���:�����ia����ԨC/��Vю���#��7s�[S��r~	���aL�f�)XsO�����y|+��;7-��a�0��9^����p��KΆ����9�
���(�$����=?�8�60f��kF��>zX��d�9��j��[y��1t�a͒�L<��5?���$�����7������w���i�C�юl@�"�0/�9a��d1�i��q�}}t�)ȩ��ڽ,^Q[��ݭ���sE͞��;Uߓ�PDީ�ǵ�n��ؔ�j�X�� k�,��5]�[�p,猣��{�H
1�i�m�O!��<�CUk�k>hoz=��H���ד����p���O���>�u�r��L��k���P��RJڰ�����)�����1�MUep����I�~�8���`LY�3_ѡ��G2H�}1�2�U:��ps_cY�����͹TE o�]1�[q�]����씐��4ˊ1��
Tu�]j\=�����j�G� g}���I�f��`�Ups�n����q��6�R �ƶ:���Qb�>�A�hnjs�����Z}4a����'��k����R���)E��.@����P������O��+0�7�a-O���w�;�������6d�K�4K��f:���{����5u��J��0�������Hª:�Ė�'��/��D��3�Ϣ�W��KW����|��`������E��ҭf7LcZD)?�ſN�Ao�m%+��,�d��k�j�ڙ=�:���"ml�0�cX���c]"In��}��	j7���	�����sȜ���B)�/�?pL+�;�P�1�YMeN-���t�m,�Fh��<
{�Jĉ�[V�K��a��W���"ך���K\k'x��}�n`y��W�{�/�D���~�в�s�;�o	�㹡�|Zj�@H�0���=V���U�� ˘\6=e�ʄ�!�sʃ�`�|���Oz�W4���IH ]����MB�xɷփ�T1����֣��3��"�[B�Z�t�ﱲ?Y�Z'/T~ՙ�П��D���7�T�;��!��1d*�!#�9��qf��TL��<P�Jk�||Ϩ.���:Z�C�	�k�I����j�{�W��^ϫ�Y���;��o��U�t���̴6S�g��2��8;>~ q�^_AK��`�z����uW*��D�o=���Q�L~�����Lk(^�]i�ӽ�Ĝ�0쇂{
�	0˻2��}���ߚ�OO���9K�2��.,�F\oūhR��j�21��7���ȹPN�O��\�(>B"��h��Og5w^��1,�g�k��%��SA{�i:����{�^��b�Z>���ʮk�����l*
1����g��2,�S����1�l�4�tɘ����\��ͨ�e]���5)Ƅ�_��y���kB�+.� s�s��5X��U�����V�{�h��y�Ǥ�p�ӷRh�؃Εs��]���1ƖC�ڜJ�p��jX�RF��Ϫ/wU�`�������6��:b�paai���,�P�(�<�(��X��%B����z�#�[2��A$ӟF�-=�[NL����������5���=��s-�0Ԉq�7��a0�0������K�$�9��"D��r!�(��'eH��+�N5F�è��"�.�����aI��"�-�p���E������)�lYj�{).'ar��M���1��U�� ��%�Z'�>���2�U8�u�����%"�Zϰqv���s|�����$�{j�f;�%�v�'���
6��S��SJ�����3�u��ɝ��xY���|k�4��C�;�&� pH%�[�����.��=��!����M��� ����E����W&v�@/rf�|��B+#���S��9�Ҋ��Y$Ȟ�T��B��<L��2�!z��sx1���²i^�^ Z���ㆲ�DzH�DG7�����t.!�KDɯ�
���[Cu,���;bq����Õ#Y�����q���+s����J�\��N^	��_��0�z9�=�=t�%h�!tX�e[��4�����4��&�c�?�'H��0�ͬP��� �M��Nr�o��������ZbÝ���9�*�L���M�����>�=��߮�ު(6�$5���[���$J����1L1�G/ۃ�?�T����Շ9�6uV�C�^W��$�k���/��X^6�+-�34(l1�p~�/ ZBs���*K>Os!.�y�eՏDd3���#�������{�ޢ�����*�ɝ�m�Pg��S5�<#�[S��L`����r:,k#g�LS~��XOJ @CX3���0�K�4c��LEϩ��w��r�}TQ�vV"�Ԉ>�p�AI	^E�.m^H8L�T^GՏ��~��w��X�Ȕ�<�;,"�c�����R~����̷*$���77\�
.���΄�������t�~��4��3N�N�vN�N���Æ�'�s�#�T.�fn� M����d�[L�Qk�T��Ĩ����Ւ��I�Q��\d���$���AZgA'�y#,��a��as���'�቟�"����~`~i�4eL&���8�b��]f�(d��EB��+soS�T\Sy�gԞ�}&O�������b�+|س5��8&]���&�$L<;1c�k�?[��R�G��j4G�4$�m�'_r���&LA\步�rۡ?-Z���7�� ����H��Am��QX��O��v�i�@�7��/�c� ��������VI������$@�#3Әms?Ò����U��p0��^˗�{��"ޤ�����T�z�|c��fpD?݆a��5@��"�DP��z��3#e�E}���#2K���I�� )0*!�$����1nUۅ����i�yITj�`����������M�(�����{RT�?W_�s��ϊ�a�,HN7W�': .���yߐ���%�;�H��i�"���q8M�Ad6!����O}3�t�r�s�LITy��1]�j ��=NB'�I��_ОmĪ�>r��,���@��"��H��<������aPG)��/��2Ă��U�u6��Hö6�H���4��<�������E%~���ָ����E���Ձ��D����\f��0&x����=�%�6��l#��`�D`���W<<t)̎�0�)X�:M�fx�r��p����8�n�O�U�k}���fg�BSņs+NB�N�t�0=N|�[��X.�}DX�o#%H'?�����.�_�Ӈ_��B�ƤJ���uHQ{�% �M"���t?gV�tXl�Km!-
8�:|�hy��;C�٢
�V�n =\�b�?��&���`^5��_|��jq� *�}��l�I��l��61��1mU�!�<' ʅ#�ƫ�!>�T�7~��_zV�����ĒuK��烝��w�HH{��"G�Xbq�_��5�x{�I��: �]�w?栥�@��|��2Uf��岶6n���xX���E�$,24O�A4��2C�����9�7[<�2�������)x#)�=�'�l�+�b^�6[�{�=g.0}m�˹'p�z�Rw��){@
�z����hՑh�d�d�nՐ��f����".Sun�&��醳��{��$
80���5�p	����&�G��!��7rb��1����zܴ�c��l	5G��XdP	M��i�BT(�p v��w��,��e�%J���@%��)��<w����ri}�g�m�1�Y��r���LY����c$,>��pX'���QY�a�%��o��qd�|fc�{���5A�'J��=/�ru|愴@� c���1�Qzd�Z��js��3�;��� riۡ�_}o��f������[��VD������q�O�-˓�$�ROy��k�������^��暰��G�� s˺��8ŀe;�D����0�8����r�W�e��6�y��k_ŪL[��������GL]��p.}BU�C�ѵ1yl�>������%���^
�v�и�vř�9|
46�)�j�7&��\<(8 |W7��S���V*��I�6v�
�Z�6�����NP R���_��c�ȃ?�i���mC ��?����nFXW|*�S��ix<(qڒ�q�����3�*�j��~�2�T��&�N.�Zi��U:�.���@��KYl��9����d{%�� q��r���'�۹<�Ww��T�7 �Y��w�T._�'#�G:{���إ�j�W�0�'�쬌d���c��nV0S)���{��7`���*dG��E���VU�0lS9^Yǆ����g�uid��R�\��>겖� �Kp4+l
�	
V�:W���#��t��Ã�r�ux.#����7hx�~��_	;�3�
-��?i����^����T�L݇}��2Q����aSe�8K;�^#.��Qtx;\ �y
YP0r-X�R�`U��A�����1
�!�xi�Tm�S�h�H�j{Òy;6%�.#��5��u] Qk2��Z.V�N���Fp�:p�Ʌa�e�M#�)�Zz�lvS<2[#��m ���`��H*�7'`B��ך@	s5��;9Vts<Z_�XkP9�#3������U`��� J��_~���6�1rw�8��3F80L��-�(�o����-���	��������M���_��a��Ñ(h|�M?������g��z\1��:V�q���%�ĺ�+ E��pEZ���!3Rw���4�.�~Nl�*'48u#��\�l�Q�5�ҽT8�}D�Y� ��Jy�^M�5u�&O��PI_�����)lf6Pt��}�+�����9&I�O�t�5�`��Z�a��22A�CRӻ��(�������&�B"!"�_H��s��8��{���֗#�r/[��V����9%GH#�yjir��2��@Ieə�0�Qo~��6����J@O7B
���xø�\UQ���yh*�)�*W�� �ņ������ҽQ�n�$kB��ʨ�Tc��Gd#6��m=�H��$b}|oDR�)����`u��s�H�L����u�HZ�ri�s��a�E�sԹ�\n����6%�<9��ZJx��H1�g���q6�,(�$�@e��NW����(�wt�����Z/U��J�_�b���.qM�ホ�U�/Vt��?��˺���N��w�'ϓce�ht���K=J8kVD4��� �k%�v�%%���[�f���[�;z#��d�E�y`���֢��a��cy��J�JK�^�V��˶j���7���+ɩ��. �}ΐ!�Lt�䰿r9��G �d� �8��.���WC u 3�`�����T!C�  ?�����.:ӆ(i�9�{(z�An��<�%�7��"k��؞�@̆�r�Ϙ�a3���A��j�#�`�Ą��$Mֈ@���a}�הXc��]��ʩ)Q�(^x�y;�b����0)�՝s���z'�����NY����x�1�B��~�g�B�x���N�)�7�2�3y��(�c��~�L8]�
���^�ߐ�P ����8U����<��(�����9-cB�����W�UW'�AF��v�V[��t��Ù���
{���e��C��s%�<�(M2a���������K�hڧ�MJx�xG-��ﾪyz�eM.�UzD��d;k�Ze��fcP]�`��t��ۍ�I�Di�3�?�k�qh'�lr�U�`T����YPB��R:T�A�3\f��_��3�Y�ߔ¬+M;�7� �.��<��
�ܞ�[���E�	�����[U(�b�Š>E���`.�mZ�q��
6���S
���{�D��˫���x��̅�W�1	F
� /���4���yѿ��
@��#R��+5�܄"��q�'�h^?	�kb��f[�1a^��zu{������ʕ^��Ϭ�eb�2����@-;�l�b�x�I����P�|��8?'w�Wi�}�vb��;�UӪz��b ���FK�;a���
�֫�c6���謪�x8�xv램&�@#5�(Fqn��Sv,D�M�̲�T\���T605��0��2�2�!��ų�JNtP��^>���0�Z��m��� Ռ�̹c����c.U�;@��.ߧyI-��ݥi��2��7x3A���%@�K�1�Ps�Wק������[�|@HfR�S�cד��#I/�d�*`�F���i#c'1Ҏ��X�$���;h��D�d>��zB�w�M����ǧ���WT��H��@�f�V���B=����u��	��]�u�{s���8o
K��#s�j�:�zV��8�@�0,�K�r���g�|���frBm5^�M@_�	؂��HbPt��6�}@� ���
e �nY���l�9�R۞�~Վ"��+Ԑ��Q��_�2�/VF��
�TuG�,�FXw�������E���`��♾�{L7a���������#�[���c� ϣ4���#�p6g��A�g����#�^�z�SՎR9NFWoɜM�=Gc$[���`�2z�t��a�ｿ�]4�BӹmI�&G�M�C,Tz4�t<�	�D;��x�@��=Z�o3��۽��������霦��)��F9�����!�tY9�������������A���?�s;ַ�c��F�E�A.�E\o���L	��8 h�&uvr��Y���,Ƚk���P_�9BJ�y
2����f���M_ē)J�lk��wd�����>�f��|>*!T\K��2�ͨ�>�#��H$���ṫ��"�1�5��,�w9n��5��_�m��Лy���k�F�J�B���Š���z*l6���R�n�W�gM*�����:uEK��Z���^����fKJ�P�V����XPBl�W�J+ު�MV�}l���n��p2u���%�kʰ��:?��_^v�};�^_"�U���w�1X��?rH޷Y���N�aa�B��s㸞�1 ���X8�*F�̴�p@铃�F�zGSo��nj�^�Qypc���R�Q�x��WT�w�v����3a!��N��A>��ed�#��%\r�6��F�%�M\}��'�P�,4���W�U�q��A�Ġ���$�X��^vv�ImIX]��䖁GEIVB>8L��j�����X�IO*�ʒw�R���' /9�˓���x47�G��g��͜W�-���j��|X�b&o���������}�n!����:S���^t���!݃������=6<0����5B0�G�Y�����������N@��^��	�)����
��'��1?��^ZH:�;�ta¬��v��jh8:T�P>h�WK<��3c�x�R����W!�q�Y����ӝ��
"%��#5�7%d�H4m(�-� �(������A�K����Ǉ����U��K����`���B���ӭo�(^�9i�����~�8r�����yR/-�V�8�z��9m\̋�W�t�� }��<UȀ\P)xmwW��QTir6ƫ�:�W�]����|��Zr�gG�򊫆<k\�FW}�����&�T����i# #cmǄ�!�	����X�=]�����8��Y�J��W����Ah*���h9�"G�S����Z���O����H���9-g����E��*���)2/�xn�Y�~�Zm;s��ʰ�&>�G5c�`KwJ��dk7 �9���0r˞*�K��Ix"�PS4��.�s����L���e����E�V�����M�))�<�>�i�N���������g��m�"f�@]��>��K�I�d
x���yo��R�����:_�s$�2s��Rz���s�$Y05v~�=i򦎴���2�hg�帄 <�����/1(p>��\�*NA+e��6B�GZ_�7|>}}i�.ݹ��~�*hz�ȯ�7�h�\�?�& ���j
5������N���R�+�o����{�3f���k���ї��f�&F�h2�2i&:��s
c�9+���M`��K���o����,_b��Ȥ*|�G7�@���G�s�J&,���^5�naT���"�!�b�K�
�2���MW��C��@�-L��Wf�]?\��Ih=���g�'K����٘�c"c���?_s=g���J�7��d~Q?�g��K��Pe?�]���kB��to��Ez�\�RA�UΨ������p��Q$������G�y�L�3�G
H���{�����(�U����"�x��K����x��`�qIu��3G�B���(>��%u��FuƟ��O�H4�NeJ��*���U��88����,�/g)\qoi�XY�����my �r�$�m��9������}�����˴\��!�͛�̩Y���!�]�p�O���%Y|x���<��~`�A$����<aβ�b��ڽغ���Hޚ:)B�!Z��p8$1�:�tԂ2!cw�_4L������T<�'������6Ԍ�=�F!U H���`+l���c�X��~����Ndj�$*�+�'�Tg���ȁ��ZUp���m)�����å�v�/b ���<�����h4� ���o��v6xQ��C����M d�J\~�x��"RV�T�>�ob��+zpQ��!xkM&�#�����Hi4|j)�������K��
�@��vQ+�ߓZE]eQb�[��%�� 7��=I���p�l�����juyD-O�C�2���Ӓ�f6JBϮ�B���hs�-��Kb=⍟��T�0�Żj���DsJ�|��"TS*���
vo�Zg��)^K�߈��9�y�63�P�
��Ʊk؊���p�mbȄdu�/ʊ�=��AWr�Suo4]�t�*��_��������(�H5U�@�nq�7v���S���CR�ǣ�����&<�L�j��mn���?�+r�`&A����nP���ƞ��Nf[��bQ�~K����]y�h��$:�K9�����ކj* �i?'���7�Oփ\��J���ݮW�X8��h�%��������ăeίEg�z���7X5K�Y��=u��D��MI\��D	��i6�S>����N�L�+��¶	�&��aɑb���!�Ѡ������E�A*��*��W^~��.«B�e:`�;�nf��~X{A�T<�vMOG0��lH��4hѻ��n�~��	���%*�,���r��5Hz3y��]U�Bx�����.053t��T����
��)�[%1�l/�fR�W�i*�H ꌧ�R�t��ݍ��8��ihè>�%h�j ���7-��x�:_�7�,��u�mNCR ZRZx��,�4v�T$*�h���V��J��L��Y�M��D^X�����r�����"9�6�����5o�<����i+�|	a5�ʦ��DU_���!\5�ݷ$c�J��Ek�ҺW3n���R��
�t7��"	Ƹ$lmo^<�� �.J����ȳ��U�3�&������TKm�}���*8��o�ba��?)�����%d$#����Eׇ�[�Md2��՛��g }l�d^-E�qs��?�	���G�g���kWYY���U��W��]���Í)��d�q�G�r�u�ӗQ3�`�˷2d�� ��%�f0'�}a-����3/�Q�YR�� ùz�a&0�J�>���s�3nL��0������?��a��G�:+8 �BN�OԔM��* �lAN(#��)�X@Q*��'�R����3�C7Ԁ��yp�W,MM�_��'M�_���.�o��³�p��v�PZ��rr)�-PQ��_9��[�/�r~�	\M1��ϥ�R�Qo$����VO��V5��;��y}G�!�)U��3IŠ1��"���6'��U�����ҧ����!����ޱ��O��I�Fvx���l��bd�d��	9��8
�S����������s�	�'A���)6�`o����m��|{b���p��� rQ�m���o�s�\�g��V�GF���A�C�`��9�W���ږy Qخ�.9�!��B=�6� ������qQ+��\�JԨ�G�xW�i���nW�lT��4(^8䒂ެ]v�7�$AxfFM\��gO�����[k�ș��^�*�%2B�S\����r�^�8�hJȫ�u�eAݛW�$G�}y�a?����2��/�Y��==�ɒ��qwtS�������f@���Re??����Q�X�7�����i��1�g"Ǎ�C��!y1���.��Z��ٽv;�C V"K5<�Z�
��_��R��J��Ky�7G��x ������"v�ĉn��M_NPMY�~8s[����	� Q������O��p1o8���Y�49�!�t�{[��	����@�8�傚k���*����%g���Lz�d*�Ahn���>s�o]g!���aܼG��0o��h���Ea:�J�wae�E��x��A1
�0i����E�W 5z�==�I��p��(�{�grj0g�1��zΗ��@@�dX&��X��	�haO��8��I7c
��`�bD_/a�^m�|g���:80x�<4\%r���ZVD&����."6���.I�뎞�[��q����]a�_���ɴx�wGaa�3U:�C�i�_�-1M[j��dC��-�.4��>��\�������^\��?;jX{G�k�=��Ln��9��hs����;�]��t�a�#�<+a�a���C�s���]��,������=��������yK=��ӣtTy����mw�ۯ� ��l/u
P� 6�'6!Ԛ�!��8"�x�@;�˺�!_����X}�e���L>��e������9�WءZVO�����cnu,7�6�`�oC,�R�Dd�o7�T%C����C(�~R�by4i��X�s*�~F:��3J��B�f�iO���?*��k�>7"�괋KJ^^&Y��R�OgC����U�m&n�=�	�I�ыIl�KG��>�'!b\����8� ��3�w;���G����Z���ہ�z`��XVn1���&[pTR��ke�W��4�y�����]I���4���:��g�����r�
����zwsf,u�b>i���bC��k�	���(�m* mT�%��rk�j���AH ut�[DD$��(nO1`
����
c%�\Sh�I��`K���r�8�
��SЃR��=�/�q^�T���O�:����!ǩ�4�X&�%������4��9
�������7�1��1���"�0`9R����r���B������@V $�F���8�Ȗ�����܄�+�Ĭ)h��䨰Ә:c!��5�+��Y�(�YUo��2;�� j�E \�Vp�Q����ּ��ӧ6PD���ID !g�w�=�K��,���3ם	�v���Y���Ȃ�e�.�?⣠3��_��5܆�5�i���v��0�1�T�!Va����ZX�����99:�+<�恻 �d����D������H��$>��s<��>�IXt��x_W��¢T�Nj�-.~?~��N�{P(��w Zk�0�^5��\���b��ݑ��ږB:( r���kj��C���f����dp��-��la�T#Q������/cES��Y#�Ő���_jHb��V�J�&�8)YY��|�8���`��{˗M���	�O�_�\)�>�0O7��-�x�܀(�*�����h�ĉs��x�|����l`���ux�ZC��OS�P�jjv���������v�cU���9W�%u�,���"_���@#+*F�/V�K���*��<b��:��N-��إ#e�q�||�e%�7#���WĮ��k��0�tu"W��+��X8m�s�����*� �4���Ď�Sd�(��n���c��{Z������>�h���y��L#���mk��;IM_�_����oe	J���N0��Q��q�*����O?�0�ӂ�o�A�O�o��yk(�LC�G(4�����+�>G�@��$�2٩T\Vh��d��*��yw�Ӥ��0�i�fA���,^���.���wp�	�A.���԰ZY�}���![������4�i�o��DޖKB�5�G�cdYm������X�����K�
����~��1.%�.<��7����"��P�jlpu�Q}F�å�~�wF�5�_��m_0��t<(c<�2½�4j<BN~��n�
HGB�
�86zˠ��hD�N����L��4��+A��Q��}gW��5m%q��)�Tgҭ��lBSK+���Le�0�ªZ���;L�@�����B_���lLkdy�s���D�!�W�U�4�R[�X�Z��O\*�4x�MD������
����0@!�0��6����,��&��rƕ�t8�ˑ��{��3	@�A"�0؅(2��`�ļilD��lc)�:�Ň;��u�����ɮ���4�2`0wL;;ʴ���MQ1�G)P�����	��_�j��4�O͚���h���?�UG��^;+��)��s,��U���UT�[P���]�ׂ��8��W	�/��s�VC[�\��:��x�52��KM���_�ALD�`�b��ӌ>���XG��7Οu�b���X�_�mpd/D���uU(�jl9YrB���@6<Jo�}����LNG�R�ר��`�(Sn%�Y�) (ڒ� 3�|j֑�3��u�rؽ��hVf ������^��6�.�����݋Y+d��F� ��/Y�⬲��d�<]��	�wr�Q8A�="�12�u�KF:�����G�\	�{�/���X��A�9t��b^���X�=��؀QN��)WD"���'�[8lωY�_7ik�,�)��l�5���}�� �0���h�W�>n��<v���� �6â�[
D6�&����pl��Q�6��a�7���BL���=P#{��V9)�b�5�&�5��pe\-0�gTҏ0�_f������Ps��B����l�U�4��֝�n�$IE.��P���VY��.�j_ܪ�Rh����p��w�`��'�*68����>��,0�KA�z;q�L+�Ə�ZO�J>���2�c���e����~X���f����j�+ ��Baőr�D��[
��Z�QFgZ����@¬aA��c�rN5�޷�W��#!Q���-�dV�w ��٣	�č�6K���tY`�87;c�.Z.h�U�W�k�_(��$O��X ��*16��\�ft������V;*iq��!�!I�X����@����Nܥ���e��� C��W��b`��K˸��7�K\�(:S�h�(�k�V)AU�SjU�)����_�ñg��^��z�.k�������żXx�����Ird����v��N�43�f���:�$z�`B(rx�Ӿc�N(�~��຃PQ�o��s��Qn�H0�o!���c@����?0�cڃՉ�@�
D���j[@X�0�{�"�C��'�N<�|p�2-���J��Q�[��8֦};��_'�����G���U�����=vhʝ^<�?3�ؖf[;�.�z�a{
���=�_���O2O�C}��� K�;�&^�CX�m����N<�
��_[�@�ДeP�nY=b��y�[�Ep ����6#��f\��Q�$I��&M�ׂ�z{�WD�;[OD��.��4����U ]Rh�^��|����X��������|���(4je �v�M��AJ�\T�X);�T��6k!pCS'��� �]�߽����_���Wޘ$�R+H������l)�h��e�*��r:�e	��äQ�m������l�����w$t��3��܌򭡽u� [���h+�\��:G5
�;�F�^g�uϛ(��Lv�ÂS�IW�O(���7������L;�)[i�S�٭�<�	DM
pE�\E��_����G�� ��2���h9h!6dG:�Fl��x���Gv�@H��ވ�g��q�4؁��.����3W�Ƣ�K�Pŀ���g���{�#t��r����^��Su�X��׀�^�����HP7r�Hެ_����E+�s�cX�ۤ\�n$�*�Tc��gGj�bOh��c��׎��E�kn.�Qa����u������y�f{P��.1G��1y��7
H[J N��W���y���{I�?�	|�Hw�?��u���隔?��:!~�͛�a���us�?;�p��w�m�)P�ê_������0��V��P��1zq��G$��&zF��se���YHS�n�ë�Ah*���֣yc|
t4W�����_�s�a���:ӝL�1�����v��_�qw���v��3ԗ���a���Q���3����&T��FKb���Yژ }�sN�y��!R?v�=i���i{��X��K�D�e�c���2T�f
�1���,��]�U;���������hY�hо�gZk�
M#!ϕ��U߶��m�6I7W{5�4�P�,���}e/Vf����B��9��lM�����ǝ�u~�	�H��w���}��*���1�c��5�.���c�[��LI& wȇ/7A"Tt�D����-xs:��hp0ݛWi���:Y�)��MV�L��(P[+�
<��Ǽ6�d��j�,�(�#�O4��l�|b����p��qu��A}�K���2T�J���a��hL�v�
���ŖK��f�?��b/������x��vŔ�p����i�PM��/��~��JEs�t��7�P�U������?�G(�V�g ��JW�� �n/�1F������g�_�~�.�>��ѯwE�$�~K!�ѯd��Us!�U�!���B� ��t.���f�#�G�Ҋ?c�&�����ea��x�T���Y��E�N�����`�=�`�)��..n�������Y�iyC[yai�	�2:R�����.�+|b��%��Z0(U/:'Q3u�Y��F�+��Wp�KΨ2��?�hWr�~,���Qz���}qw�_k�;׎��%�]4��8A�@l8$B�Y�I:d�'��2n�j��y�Pb�����9�aG&�ܖb"�T_+�־]�O�b�)��Q���Z�� �Ր ��U�v��[����|�3f5��H�¦�`"�<X~��nI�� S��Q,��hõ���-6f��� �O-M�2���x�����~g�?��5(���&�K��@���i�z�����c(R�'��pmyJ����"���o�a����Z?�!���k�BjLJxk�;���_���qu�hζ���DIp��h����TZ��8z	�<�l�"�g�	C���a�>�`�æ����3�ꂛ�����`��7�f��������Qj��k����{@�2Т_@�P֎q���|�-%�g o����%�\�K���~NC�F�S'��d����2�4�U�����̴��@Ke�rԿ��v��`� ���
�
@)w/r��Y��z`�(����}~h��xV=�'Hk�+��H!X�T�-�:�Vƭ<��3z|��aY�ka�]5�̜H���v���A�VDL�'7-�I<��7����
��}�c5?��d0�:��J�K��e|>�S�AXq����R�����WR�����hgi�~��6�>�*���<؇V'��!���sP�Q�7�<l5�kV �P��^ƭ��#�fu����g���D��Q��V��2�X�>y_��S��֫Tyj�p���Dm���~O�%K.u��k��f���*� �F$ 0�0��������K�C��+��K�S�O�=TP�a�<N�8tO0baGE��gzn^Ov{���-�8(���{�z-�ю'��?�;㧱���9 zY8?-��ye�cd<�{e�v�nN�Z��MO�����#o����'D��a�h��n�����|���x�5VR�nhK�/�z��\��٠4��S}���0�TS׆�ȡ6?��$��?�:`6�#eY'��گ��Z<>ί`ֵE�,0�0ew�~�����@�q�����L_�a�b�F� ��a�`�L��F�A\;6���$(8\b��i]�y��-0w�b�Y[d&o�r`@�7���HJq�0`Rx9��,��W��)�|I;�p�6����Y�l����� W��\gK(Un놴<9#Bo�-��TkJE6>9!z�����m�ƦiK`�фӮ��Cṉ�I�Q�����˄Z��ކ�_.�^];a����:��E�Z�H���SW���9��l�W�GE�{������V���K^~I�<(�kT�^'�����P�^ ~�n���9�bn(=��W���mo:���.���rQ�0���uՍ�<w1��]���&��թ�i��H�����Ahn�)t�;��;���4R�@��V�����^���"�2%�x퇝t���fI�"�dAZY�	��͏�(u���5"���!�ɒ��a����g�d�B��(�5�@:
�)ɖ����]�����е8Įb�xй�䗧9N�?�����$9���+��i�^�j'�xׇT��Z���ݙH|��(���n�eӕZ�ǖ���y�n 'xQ/���E�L��Zc�Gs�OG�0?%�
����/��EuQ�3P�\��_b���5J�Lk�ךp%ը4?rwY1�?*u�<�`�1w��I��^X�}D��FU�82+d��U.s�H��ɑ*�]9|�>N�P��Pʋ��_pS�
�<�fe��f:x����a�K����	'���D��1��2}
�E4�;h��|�N�J�7#h#{��9+56�< ��m�PC'���*?AWv�^E��7��+�&U�А~���س�eD��f��A�g�2���\< k�V�w }OP��uo�K�����I�_̶ /#u
�@F\W�LǮ�{��#3u��b�9b�V�3�_��.s�ϗÔ�	�|�/{�۶I��W�A���3o��{����'5_�����w�Ag�x�SDi%�1�Hh�2%����DbDGR�q�Y'x��@c�������$eW1-b'�:��S㝪��17��{$������Ꝋ����&ɷ%I�}�����q'P!�����=�]��%��I;�S6<e̋�h\���������({��tIx�]���*�[� $��;KcO��3S�����%K]�P�gs.���yn�Q ���u�"�#�I�Z��Q�z�t��sъrӊvJDR��diD=������]}�w�f�a��4�}O���F_���;U$�|��+��l.�'1G�� FV��"�����2��P!���!�� �Ss��N ��L�M^��Y�xS��G��V	�q�n�Z��{N9�R$`٭$����ӲRd'.~�efĞ�G-���'d)��F�����C\���v�b���O�m![m�n|-�����,+$�1�j�v��$��d����r��߉�`qŃ�N 2�R�4��\�c����=�r��3MN�J*�����.���UކS4�j>���Y"�ȇ?��{�s���?���x��춏����]�>�$O��3�P���M�t��l���~��'�����=˯8�VN���lK}����Оbh��H�m�Iȵ�ά�z�A@�8�:�����o��j��5zt��sm�o1"�-�G|���%��f�,�K^�d������x�no���s��t��3vL5_�DaQ��FyHKH�"�qm�܏hM�g�c�/�xPpЂh�F?�����(�W'Z�O�`�±W�&���5��~�y��t_{�8F�I.XP���eJ����:l!=֝�u���>l"a�s���g[�!f{�lE~�+R��huO�<�о0&�T{,=��ߤ5�q��������V�AP�L��Y2��b�#���K6�M*@��R��g���}� 3�J̹3j���*��p��F��es�������<U�I^f�i�Xe"85��Dȴ'2��f�G��h�:��I�Z����L+Y�z��)�nr]*���+��+iA���(
�K�&������iX��-�:��[?��^�ٞX������~�/HR�SG��� �aս��[8���o�/e���Ï�Kʩ�1�����l���Q~�M�����AQ����\ѻ2���0���B��n�h('ھ����82���1��|�۠[�j���è�L��b7o�.S� g�է�\4ٝ�����j�� a7�l�THv��q�T_�
�b��;��j�������]g��Ȇ�H����a+���8Rȵ6�o=�#�ӒH_QB�ba�E���%.�\�7�G��Ĥ����m#�$�^)�rx�CD ��A�zB]L����WT�{ݪX^�uR�s�����G]���LZ-��Ƥ���/ˎ_"�Z�9�R�e|�g�@[�X7r�~�R,D���Yeg*��g��p[� 4�*P��"�z���jz�+\��d}����Pn1x9�ǥ�A?<{Fs���K�+I�d�qE~g~�������
���r`��U&m��U�f/wkh�jo���Q���q~��  Ψ���E���Ĥ����PE!���;���_4��K&fXz)Z�@����/{���L4�k}l�����s����;�5����؜<ׅ�z�hHk�K( ��xe�8��62���Rh��5a�6|ڏf�P���Ap��`��ϤYa�AS�����G!09�FAt��'�q�ѕ��YR~3�h��7����=$��:P�DS�����Y���yd�nϱ�������̠��
��2����T�v�^�\2I�]�U���� ?.��lS7!���CR4����i��K�o-Bq�esH�\s@��Y�`,.����*6�Rvr�Hj�X4!���fli-�c��F�J�Hvx9�Ib�+��D�?�֞����ܦ�#���䥆%7
l�g��:���Or��SC}�)Q;�&��]p�?5$�|�I�ѯ!RqLz�����d���[���f�8j�T���<dj�]'s�^1�XkuH��Tt��m���}7�5mߖ��(�)A�ضd�c�����З�0<���;�Йm<�D�g�;_�W�ɱH��M(�s������k��a���7R�J�x�y�w|������e"�������.p[P�c�\�z�;*��p=�Ӧ��B)e��i��-��UL�y^E�x��md0HQ�}%vX4<��ғţ�K)\�T��x�6 �"����E��F�[Yw�y�� d��(_�SHi�O��Kn_jb��_�nO s�?��#V��~�0cg�9˦Fը��w����>)VL�&X�(�
;O?���b�v9^qv}�]0��+���rOŖ.j"����4�*&3ܺ>��G��jU�O��'�>X1`�v&�lfg�w���˅��+A�J4�K��^��G���w2͂�	b�_`���/���o/���+�K!':���M#�������rN������mj��Cvݬ�2��l�.��\����#m�B��"����5t�SE��Qh;���MQ��������/�����!W�Ѿ�ނ�H���K�\<�2���j\jZ�	\���H3��>`�{D�/�F:���ͅl�f\��u߅u��q���t����\���2s�
N��?>Xc�P�xu���3��t���"_}qu�T�&e�{�|��'�r
Ȧ2��p��o�%T�ׁ����&M�g8�E��a�%���m]����x�Ƽ@��OC�1m�k6Q�h�w�P��o���[&����n+{C&��2*Cq�I��x4me�!��% ��U���� ��)\J�k%�6����������綰�*�\�5�-J��Y��#��h'�X��B������C�4 a���Q!�N���-�>�߇Q�t�e��r�`).g�	�iex���~�+X.�D4�/̛�G�.s^�6� e�������FA�Ӗ���*:\?Ռ;)�uIC)K5�y�g�n���B�93Eϓ��n}�����_��\~¶����8$
����&Q��,*�,I�HPElv�S��=����u&������j���m�þ�8r�$���t�T�e������;i�7�.|l�d�/M�����U���їMҏ��3X'�-��&耂_��}�����z���H�[�ʖl"��퓃�'�C�֢d�P�%S��	51���r��")U"��Q(��y�U�U;������.�,���pI�֟�x�m��6�i`��ə{[�w:�h�p	)�]��@eV�k2�GL�7s�ֱ�Ф�o7�����
�����;��Ά�����<�ꄦ���\�~9��s@"V�uf���ǧxM��O�xX��]�p��K�L�kS�H?L��_Iw-@j+}�>bEX1͘�YƦ�{V.&��?���*sa+��qV4O��>�.����bu�~���
��U�J��	`XR,�׎}-�H�s���֛�l웱�l��]Z�!x���$I� O=�,����R�ܥ\r���fǼaNby�aa�{�i���y�Z5�;�6QB��r���<�3��5��SJ ���L���:m
���cO��6o�(��^m�{e!�&���9v��dr�D#�[����`��j��Ϻ�[q	}R~g����d���;S&��������$*��X��Rqip�7�T��������ɘV�����28�w����>�5�9P����l��I��m�T�,��B�}���,�J>��KC��2X�ƅ��}��#���`p�]0Tq��R:��%y[W&ܐD�s�6�l�{��6%�8�m.� k��*��j4(�;~8j�* *�SҡE2�.�6�������L��6�3/�(,�e��Sf�%�E�S���v�"��d�Xg�{��:*���^#l@�ς���UBC<q]|�*�D�[�VD��dw<<!��w59w�ZnW�Lm��6�tJ���fNBmggL�����Iא��?Wל.p�2� ����ZA�dY%È4���:Cs���S��Oa2O:��r5f���k�;F��1�QpD�N�,���5�Z�}Z�&?�%%��w2��R����V9���Q���ĵ��tǟo��`I�-�⽮�PA� �c�f��#���q|�M. �Vm<%l�dO"h*�$`�f����hPhE��YQG|��n���@�B:>1�g��������M�ުg��Ngl�74�K�ѿ�z��:�ć�u7k��~c\�[V��>Z�d���u;�M6��C�n�m�c�����Iǃ����|`�j3��T�K�F�8�U�`!��&�^���m�\����O��Q�eQi��]�y��ƊŞ�@��g$c�:p=S�����'D��qI⸺�����LP��J�L!sbv_]������}��~0ތ�`�U
�\�_n�
lЮ��x@�c����@@s�No����N��>ۥ]�ȴR��C�;�`���h�~�l���6k��%��GIb����P�wR��

0��N�i�؞[V�wu7+;��:,w��G�C�+�?#�awÍ�Y��\������{#��Q�[-�\|��Q��I`���@赂�Aw9�S5%;�I���g���	�3��8m�
}��O��[�rp
�[�.��n���A���%v��?�v	'M��t�Hד�ص���n�fF�i8-;7I�?������#��&<���Y��|�i����נ��!�6<��R�Z��v����)�E<�N ����#������̤��"�k�nR�������>ٱ~D}#QVߪ�π�ݒ��^ G���Pk�D�N��T@�\Y.+�6�![ݡא�>��SSft�U�g��zc_	F?�gw/�
���۸�κ��լ0�yi��/��'���KY�N��HS���|�j�ΘGq\4,�V��)�����?�RG7_	���'���\��M%�s�/��ͫg��fb����qn�#��Dr4u΃؋tq׎�z����>@eZ�\�f�;�z$;��$@�ּ����!�݀`��.���p������	ͼe�H��w�G�{L�Y$����[��/��{__�tԎK\�1�le�Pr�.x��]���V�]���VSq�ĆJ�x�$��ܙ�5��
�'YLu�#4�<mj4�+!P�"�C��"ߊ�I��ƴ]ǲNq����8�R��&2ŷ��T�������������'�FH����)��ln��<��v۰R�e՟+#���0����D�t��7����l��'}@�Tҽ\޵������/����J����� �-����Bs4�ۘ��k�}j�;GS�{��e\4���#p�5v<�k��0�F
�.�/�,��T�;��Xa��Nf����q�(4�ʅ��/����H&3������/���޾������x�����FO�L����	�G)j�wl@a�&��	�q��f֓xUF��߿�X�F���$�t���S�V{��vf��Vf���4n@��(�q�}��'�=�0����S�u���˟@���3��{������gHN��ō������������"�^ZF� �4�S#��A�eo���Ln�v�`Mb���K!C���i>IN~����g��M����
k��`E�� Pb\�sG!�
j�e0��q�))����m�'{�8�K�\�gw���H��I�s��)���kb�4Ny��~LO4'_�z�d`M����O��ߋ�/W���(������=�~����/�k��g�B$˾3�D H�Q����&$�wʡ���m63���s0�ńV���D�w'.�ZP'IP�(�;p��R���6���QQ�> m�y?�����f6\u)*�k�om�L����#Fs�n� �$����)��?Σ@~މ�-*o�S�>Q���5�V�"P����"J��.�Z���&u�B*&�o�m5Ty������l�����C��H��b�<Q�Ӏ���OG�"�%���������W�lc��(��T�=�n�!Kzl �/��l�q���z7犲Z�P�$�z�>^`�,�����*�C�1�ℱpOb/���Qj��-�g�98�nn�:f?��Չ�F��G���xr%�GG���[�T��7��+�@��M�����#=Rw�������Z
�p��%�O�ny�ے��==�6AW�v6w+���/FVX�`vkL�nu(;i�0�hk��GX�q(AVe�:�d!.�&
��vпc�вjZ?�`v�����y��I(��pv�Q`����1[\4������??�����G���G���C�|�~�%OB��"̈���b��>Kk�u8()����+b�z�3j�ӓ�����}��΁�2��b��F]j���5����/=U��Q�r�5j��d��I�F�!��Z.CDp��A��]wj����xǈ:��I�)B��2�`؞�*O
�]�$'�.n�+VG�"�1���(�f�����4Ʃ��Y,�� �G����Kw�h[�3sA�,(�$v-SH�;L�袽ʏnR�I��x+��x>1Y�]�R��Vpe�%`��ng �?�,�ue)�n��܄\�ڒr���M�=���й.�iV?��
�\u��9��!m���Fg\���Boߢ��z�x�^�����d�`!��N7�bt�&͌!�$�%�z@�_�!��NI��,aH5���j�J���* [~ēEz ��%��2t8��4��d��@�MPf��+=�S�*� g�>�l��'cB�{�~3H�������s6|��p'PI��$�NޯX`"H���X�|�6��(�h��Y{�޶G�~G~u��8�6��e:�RPb�6�OЧ(���0�� ���2^���
��Uh��g�l��S�t�ȓą<�ӠUk��±�q��4n�Ln���s�C;=6��m�|��KZ�W�2mpM�M�@�-�r���tl�zl?퍽q�x�� 8��x\C�`A	�ǎz�_V2p�ݹAdu�u�0�TQ(7�hC��l�([��Rm������u{N��q��o�/ۂ���<e�"X�]sG@[�#�5Qϋ�H7�z���=!��'H�I��(�~g�w�qUG�s�鯒��%B�\`VO�  ���z��ɼ�s&q���_XÃK�	ڎu�U3	���\pj���qU���-�rt�����wJ�l<��M�V���1h�\�Y�R�ߎR�l��wq �&g��ha]]ВM2������ˌ
��] �=����]��Ѵ�C�?b�U����彶�!�i���B�Gqba:#���z2�:�j��v�M�f�l	J|]��������n�q��Z�[����`�/�v�xY-߭j�R�G<~��4~�J_%y�����t��e(�]��?�q���l��c�/�T"{����1:g&�_X	�F�i/��mpϤ�z��9�J��'�>���v\0>}����D��%�� ũ8�������XU\��je8{>��z]倊Y���)��Yu�#5�{���G�G�m?���O�15��GԞ���	�'f�E�h���|q�����j`���g�՚���%j�i�"n�����6��4��i�o}W�@G ρ�V�����BR$�J�����j%��DP�� ���!$��s>н��_d�6�Cj��94�!�/���ً)\o��\;*�.#���) �6�DB�h���!��rЏk��l�p� � 1���Vg��S������Do��)�+_秃�~⩢�4r��Rk]��fꪭ)o����Ň�}���xޭ��<u�c�|nAG�x$����P�1ߝ���n
	�����ȅ���c�����v�<8+;��=\�$J[���@���:���������\�\E�]UBҗ��g��*�l�(ƥ����_-�>2�f���7�ư�)o��F���[�`�x++�N�(�<����� ����*5ZI�V�J��͏�2oOj%w�����L�*S�=*l��D��}�ø�+���%�[\w�ߜ�4}jѺ�w�D�T��/sK�J��GN�k�.1���j�y�֖�Nb�ܨZ�����\�>k	� ��+)�A��]W�1I�j�X��*
�9n(=
9���Ot�X����@�q�2)nڏcB��[�|�LU�A
�)�z1�u�|ʶ��!�i���#2�e!��=�ė#D�3jh��:yv��&{��sv�>�"��CӀ,�w
R����w�OT�|y��jEw��`��/�H�]UN�A��=+���~X!BϨ��΃��Y���
b�=�=dR�ۭ�"�I5�s߇~ vB�5����3����cP����\H%f��Z)�Z_�xY�0��o]�/�Cz:9
D��B�KJ��3������2m�EuA �[s�lɿw����wq����iʯ����������M��h��ż�^B� N�pg���.��z��qmjkS�_ϲ�ɡ] #�K�P*��e�W�G�ʗ����u����ɷ�$Ɋ�>>{�nƢ�lv� ��b۵�����w��4�f���NT��Rh�xBO�VH(���Ϻwo�w�l2%�u��r���Yd�k�ׄ'��a���@�j�֐��A)	��*���2e�f�	�D�|B'�1�%k袁�� ��L�l�b�]���S�h;���K�����C0U��v�:L�����"Ś�Y�����!��{]�
G2�W+�%?��ku@}�䂸sbiNճ�dP�A���f�q��3�d(j�4�iDhw�����T ��]���;^��H�H��׍�'����N�݇��H���_
���+��q�e����HܕO�iݥ��)f��"� 3���J\�}JjKAmø���%�D�8�)O���x�B����+���h�kXO�Eqi�S���_����{^#����Zijꪷ�D��]A �� ��r��,,�5	��&zW]9�&I
���#��k��R���w��-к��`�mbqX�6�CIrp����Ry�7+꺲 �}0���kJ���U�>s�t�P��V��n�0w�&g�4.<!�/v*�˙ഷ���": �BR�y��Q�n�\��d2�-C����������N7�Z�.e �$�nwoh�ۗ'1�����#�E�1}&�ji�W�a(дk:��(�Ħ5�pb���4@�z;P�P��S��c�B��ى�k�\;AUQ>9<���۵�H7��[9J���ܤ���%Xő�Ji=@�֫Ƽ�A��3�C��!�u�8��;��CpƑ��h����7],�/v��T�'}ڤ�ҫ'8�YrhY��u͢�U�Z��/�TXr1y��p+R�umM6\v|��)�;sF�	nj�t�����c֡��CY~�K�X�W!����O�r�B�m+ѹp4E���Z�^�q��*�Tj�֎�}�W-J;!�I����ȏ�D��} Q����Q���uN�/M'��+����_�v{�c���"9���\H�F�U^ �yxvySFv�[����H�w͝L�nz(a�Z��jYb��pN�i��*2~o�$Cǘ��0�B���i�dL�[�}�@]��0�Ľa$[����?#8��o�<�S�ogO8aɃѮnM"Qy+��|$�����%�^�����q�]�����(��3��J&x�}��/�dX#���F��o�Y��2|���F��An~S��8U����`���'��e��$ede~�Uo��Տ����z�Ԉ�n>�����"qy�����6�
��2s/�2:�i:�6���_�q�E�;?���4�'|��m[4�e~��BV�x�m~7�=�u��G�\t6����a�r�O;J�d-�yאEꕦ�ۄe#R��o�k�o�lO\p<FЉx������kJ�[��!�߁��B}���e>��.�_�Y�"}hꮍ�S�)��/�.u8���ߪ+�����+r����\��}�>�p�nr��a�fm��P.�d�w�#�C����i,����h���.A-k�-���Z򼍁=��Mh�>N09�)'o�Sqf�`ƚ�$Oz�͚��#dC&�	����T�sy��~�,n���a~,T&|�iБ���� ���m�2��q l3�ǂ�z�ϛs� =�a�jr���eϸ7�P��9����R���V����0��(Y��ۨ-y��s֕ƺ<���W�g���W�����;���W�ίoETxL�y/)#X�|v��4����X�2uvj8�s�8���tƬL��-8�k�C����h�Ƌ��I֮)�̪��3,�J�8���FR���YU
 *#�-�Q/!t�J�2
6��X��t��A�L��8@n�}ي�ŕ�����Kqq�lx���A�Q���W�И�q0�����;kv�pо��fP3�W	���x���9m��T	i+�fe��sv�2��ơ�������0H'�5��D@�bnL}χJZ���րvw����O@��{ڲt���V��&�ֽ/�i9��JTi��#����.ɾ��7�wV�1��F��\��P�W+��_�1���>'�xn���r�=$%�|9����愸�o4��T窟ڵ��T�`&�ю^�[{k!���D[hU�)tް�+O�E>%0�� �܂�9�ѧ?��'X`,=�k��u�EF�wH\𳹍ĳp�d���11R�
�ꂄj� �<1/��I�ySg}�0�ro��BV�$�ep�
� 
Y��+f:�x�ԡ��13����!tf7s�O�/47��Fe(��,z��-6�W�݁>�R���]����V��FdQ��O|�P�en�Á�c�ri�x�QH���]"7A�v#B(�zT�zh3�AMԳ��C�ڐ�%XA�k��YE��z�B�RaKv�y�pzb_��<gs�`f3��)�F�A�V*������sc$c/Wc3�:����7�N�������Ӥ;~�f�]�סS�0p�%8�P/\����j��pKل��6�b�=�4��������m�����P�T�3���w�I�� �Je�<ܺ�.��Q��m�i�c�����-!�{�<�cϋ��U��{/Gj�5�8۬��X��
�`M)-��wD&!-:�ݧ���j���j�;1	:�i&ʥ#m�2s�{g�_l#�+	\U'�����$L��o��D[�
�j>�З�4���{��
�c�.��Bn0��@옪ܳIeE����F�8f�N �v|��	�z����k [�`]9r=�/��f����RV��Ȳ~��ܝ��rlb�qK���,e/xX&\����H��k�{Ϗ�2�R�\CtSɬ��ъe�OL���1�s����U�*<����5�� �􄘓W9Tr ���#��(&x�'D��e�v`O�Aib*=�vG_=%��_O�����&a��[^�H�+����ٛs�8E��4x4#��o*E�)q'�C�@nRYW��ض"I��]�ǁB�(��>��J�e�9"�S�3YY\��wV�%:��+�QtL�5�`͊���#L���7���x�V�9��@\��o�4���'�F|�w��C�؛�Y�b�2�\�D�&M`V��7o���1PWg���Թ����+>�4-2,ж�I�P�	~Ċ���8 ��\��5NH��?�N�#+ˤ�W�~Ȋ��\T�����4w$cQ��BY��V���j�-��5������d���E�x�"ϳ$5G�8(B��x/U'~����O�Hq}U���g{�=~F�#�l?Q�y���U�c����y.
u�Uu���ؖ�#�`g���G��vN�)��ms�2�����^Ak�h7�9
x�<�ʍ�1-2II�A�~!���O�f�?����`�a�E�$Q��b�y���K�W���r���ܓ��^6�_�y~�B��J�~v��<�Ĭ.?g��e�\:���l�uU� Q���C�4nY�'�@\� tҌ8�6e^(�Wu��}�����)��#3}��(�_��y�bB�=z����3�<�r��?RmK��3snG�Z��#�W!����ը~��К��/!v-.|Q��
I�AYZ?��ZQ\�%�9���")��9�Q����/�˕������J̓m�2o!ׂ��	�3����H;[�Kh"�)s�_�0�A~�[��r��g�Y�*$��YtCc}:��|P�/���O3MZX�]EIn�x�se_9��=��]��ڎ��s�A��	s1 ��w�j7�^@fj{i��'`��_�og,_����M�?�:�#������%��
�-U}���N��xQ>���B�����o��`��(]ڽ�n�yo���:��8lCډb���lN�)��q[ל_����d�~e2���K������9@�ߍ;�]�{LI]�Wf�	8�<�Py������qZ���iU�G�#-��^��'s��\F�2�gT@vn�,�� �)yjM���f&;���,sF�,�(�6<�}����N�il��?� ]�#� �P�
, ��]#��Y5;��罹Pܔ M�{���5���Z��쀬�v��x98	�:�G�7�8����'�ǚJ;�t��_!�>oU~YVj�
!�Lh��AjG��B�A�c(�\������A4Qe��0nP�
�I��'<��ՀT���	
io02,��&��&��Y��ʹ�d���<��X")&���<?޼Ʀ�dZ��^��T��������Z9�����U��v�V6zY!o��N��Z_u�
�,h V��¶Ŭ�0!;§}������
�wͱ��ݣ�0� �N�x	��̛�i��e
uz� ΔPĔkD�W�^w��X���&|������Nk����H�x�j�p~׼�iJiz�����:vj�m��<į[��qW�����U4ܶ~���KZAq��6}�7����l��_0Z��da���t�e����JG�b���{	�+_z0�-ۏ��;6*�y�G��}48a�A����nK�Uc«����>܂�;�X�Y �.�|���$tJ�`�AuL�O��;e�P,������'�u�� �}��x�ce�݂�vt_�]_�c������6�ftx������+�2�T��B�H�,�Z?�Y��!Y���`m��ؓ��-�);���~zv��^�Ӭ\�&����ZYS�F��CJr�G��)����]|���um���7.��Nl���ޔ�F������vݛ����w�(��-�S]~3]�hH�Քa0|'U=*V�Z��H�7G7r�
~Ɏ[".��6�i�)�6 q��]b������Eq|�-�/FM�=6Q��)�5��h��G�J��s`���KWZ�UU����y٥'�@���y�e�"!�EmMX2,��U����`�8�g�x��ǆ/Ek��L��G�Aϴ����E��	=M�iU�n��Ft��J�Q��y�GBo�^T%��gްΒb[f��,=��t�,�i �DHb��\ʎ�ƫN��far�=|�ָ~�S�	�8j�{��