// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:56 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V5nm6MRvSwARLGK6+ZsW6jrIGgG3XJYa9L4k8kPLMMax9Mt20MMY7/4+7RZXJiLX
Ow/BHoRkh07+bG0+4QPYp41aKDNd+HQ/iM5Hds4KeCfbBI1sVNWUas9BSv3VgSBg
R4np2Sku+UBdTWdJKAzKm2Y96P23Sc3wxCo8tfKWrBk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17984)
BEkh6GFbmTUE6AVetXlWU452WwLwnKk5dJusq9t0vmUe1eI1kzQDZ3YvJYbE7OX4
mWdS6nnz5LGwxcKwqFCT46EGLd+f0T2ATuD3C+WqOBu5sMpJUqYjc46ocTI31XmY
8TiNoF8iEgI9C5vJvDowSVLQn4Y6fhp3XLzLgqJJSGVBHq+f245E458DTbTN484o
Ab6cE6qrVRyDJ21T1cBdSt0UBigpr5fZTs1Vz1ZnFwod6o91TZpvNMsBohwchsFb
JUBgBUAFMbkq7GG10TVzJ1fg+3Fb9HFtaNoAYIM5UzRfOBhI5dnsD70O4c4R1Gnr
ZCw9raVniwPNR3feee6D+FjGjPddjSo7dYITCfRqbbFBjcmnTkmmIZH963rwlvW9
N0l6QQ0AyB1PHy5LvhrE7sh50eKnO9mJ1NXu+PJp0DjAyROtPSMngSnQe6cW3WCp
TrtjvCDuKS9+xUxtb658X4pqU45HYieWQrvUUTltTExfL2u9R3L127O1CE6WOoWb
KxUobK7sUv4krhRGcmr/gau4Ix5C3WvIdO/pKT1x2icdgBn+SlHUqNylWdeFlSwc
6QzRZEC0pkcq4nd3jTZQQt55X9Pt9aTtM/gps/RPlyksfyv5urZwujq4YlHMy9fI
1uf7aJn3oEsFa3Wia6p+/iwjp9bAbPeQK6gOiCg0OR/EZ69HCPPjK6XJDEZ50GcU
VLAQc616sfjjDHl30EVbg7ggeFogxOddbti7LnWAJzBal31q0IcB0mGX6hn1d6fV
ThiTDvU1rwIahFr4ySXmu0mz3KiXueKLdmJhoeSzPwg60v6YCfdwzJwtnTbEkfbl
AuWYXy2skZ9tdYYDoB6+ACUGNdsvLdSuVU62O9vFymlz3iI+UPMIfMKH9Wjctu6W
4xtMWXunU5iNc/rVvYSPld4neSHDFB2ZVmdAMu7GdGB3cYjaGzZWfG+4M1ynK9JQ
nKTzwRzlLaPit6+q6a81lP1qRZGID0G4tOJfVjxH2/w+85+sqEGd2YdlZxMVPAB1
Cef8DA5dmlHmNK9y5Cbca1mv0EPWNFeI4cm8RJMcGcGQkV7sPQAZ+6TQNEQelmwb
3inwNfWW5qgoEVmxqMyxleONVBgDWJEG5avyL0N2i1afWaO/8DiMq+a4LyU1BWNm
vIurLhzbR90X29aOOfWWl8bUG2AwBq0xGIgKU6tweoBKbdAzhgfKyeCyw+y6zLX7
B74beU3zeCAJINM6mx0VD9cLe8VQ78GqAjAFzoD9yRq6k4zrR1s7tfKFydVwL0Gl
zDiiNPrTfMiYfwv53cNeUuciqNO0/LvncDU1CvetNHUBAD8hpj2KCtx9qUrxlU6t
CjfbCZ/GOvI7YGqvpNjnoL1MIp5OlhbNn9NgPfThYomEboNu9Yd8n6cA79Bqhuhg
u+X/F//3Mb3gAAjGznwyo59sPNsXViLLihMzOg4/89P2vO7bt2BpPOxVqTtSkT+X
JNc5IeRyB0hzu0OTcWftBNILcqgCfZZ3Ji+6OH2UPPvNvgSnK5b5reZLPniNndjM
xDAvbTJeaxL6fjo1QNE25iM8SXdyduGwtxCykyj3d7YrYCmTZnJldWeZ9/oG3WM4
wKIsJWZFVVLZyEEuyfEipDbn/z26bHd/JelN5OPtEYpL8f0pVg+P1biZgvVuizTI
rtNpB93CRibeACcE6foZcVidtDTNOJ9KoMsgAzR43mm/hFH7RC2SNwJDImeOoynu
Rjr0hVXCgbZU6leXokw+rZj9Fsy5bBaymODtrE6pl7Ct4wDB2Hyig3Az2vGWyk8C
N9mTJdwSp3hbOPh5LHS6aVQ/fcNWVtRKplnGW8ZHtd0wGd5STUWx8Ynrbl7RP7x9
dx30GA5eX7nbf300Jc5NxjUIgNzV6mSEZdn2XowsuQWziOgIbjiFjcZLdWONDYzH
Asg+Blg8dYrDkoJ50Q8ayhe4chjXQBhXFG9z4aDgv6vl5iFDeC6mv184qH+21WHX
W3nGuaXeFOEdjRgxkqzTIpotqBx/wGQ+uSTxk2GGTmmjJcb6pK5FlfiuIr1D7JRF
v9ZEG5TkO1cXOsDkbGD5ntEoyGccdUVdUjYsdsg+zLFLC3DYORZ9JJvoWCMVHbav
PcIe+KHFMqUPPC/uzajSP3tYuvsTnEWNwVX2TV88ZNwVKP4PwZjRj9Zlakc6ya9a
kbyzhksRPrjJf7DhItFT97wDl7jRn73/oL3KGkdw3Wk9Yxe4m7jCM1SlPAqnoqxo
aYh1xVntt6LJ3VPDcbYJ+m4WbcuVnVc5aLf9A5OWCzD4e4jjgVFmUDgyCPh7d10C
hD1++JTpD+cqyGC7pgnk//jEDcaS882M8kIERvreQ3MGVHqKmGVt+RFyc3k6sN7X
JBWZGQjNOcsckHiUntrRI4k4H7DZ4tRRVIbQTdPFp7bmRuNNtMsx4s/zJLOnijMX
UviXQ6GmD9z+WC10Jen1oGPivZlyMyr3/Omw9AQnZuw8xgZ+z6J8TIUxmvE8oZND
Z4VUXA2MCEzMvSlUztMYFYkvgfhiO4vKvu3WP5Mb7b8+9cIS6YFcnckM9Uo1Dc1e
T99rC4Fl3MSA2eIZqZYrqGz5r15LMyrHfE8C20Be58UIoZIpSr0o9ML/E7nzFygy
LqHfwUxVLMzE46WXNrklQh6yMWW/c8o0EEMRmw+/lM0ks48OEYOfhsgg1w2wgoIS
63qnp0WfLgAyqhcOrznQOlzWi+N2IvtoUNnmq8Ofwi6L8k/MyYe5oRdnFk2SkwKw
op1GBUrpQ2ZmEZ7P7duJngNqRcRks2KvHX6eKFhEBB19kSxcmWLgVbkUQleNweIA
VcMARutQ9U4DZJNlncuixdchxywf4ZUh0alotPAmPnwaZzc3KwPFakiGyHyc+8LR
BNCiowKZrujixq8w+jHSDHQtaCg+oKBD2Gzd0sTYN6mVeTpK9I6VAEd2RQZuUluo
HecUEXzVxzl5/84T+SZYEt6VLxsTlAelfCQ4nwUGWV1cC+ErrXp4uv2u/ACgp8b3
NHP19u5eNV68gpuKz+FzEpT8SDa1KrZe/CUvo8VShsBR9b/sDvyAtB3i/uW57zFL
bYvFSID48s0DGTghY8j97rfiV0UIzGAaTEgsQ7YXO+slL9WH64NrHAanKs7XVNnP
r+p57YNdlpvBYr25oZ0UEeLem8dY5IFGPs9uqFYoFJt4n060UhpzrZ4HJ13++Mhs
SXbUrgGnFvGbIXD6ClAGwmv9NTjALE6IHbpGEyXz5MJmPbJFm1Wb9oSkk67A+w61
rWAc2JUEbii6ZLspZz1ZGxqXEX3H79rGB7hUcIB5IWckEvnHM+fJntKBY/8h209M
SWEU00XcBEdzT9gpYDO06INUHSIlX7MN816MctnRiYJ3Wor63/qD4SSZXEQidVNR
6XbG61LGGmTOB4kf3trvw6Yq/Off5nIhO2ZOFBwi2fCRYl73kM2uF3shIBbdIlFD
4x1qJKcNQ5vpgZuNpVsSMnQaopNZA60vW9/GTzg6LQEIllKEj9pErOSR0iYOxLrR
Ygo3wEK2m04Hua9Ttwni4wBQ1OxjiqV5paMnMyAGR2eTkLdUXIPl27bdjiTcqbUO
sctH847H8PKSmt7okZkmTjln98lCn8+yyICNW2g/0tW2cJenNna6EC+OUmmXp/fJ
YsmaFx6iR70FjXE0lH/f94kDS4H1qJszYrYbzF0S2XAW6rH+wlqiih3HQ2ZvQCs9
Qs1aqy/KFgDEwt1T47zk3Ra/5S3vS7nI4QqLP9NyLZA1gNjauhMoBtTpoADXk2SC
Vs28QZ+b9nUaOQhVcmj7R/dOkRsoNIctn95ZZbtZuygiac9+pEXbqH3bcfG3mQpS
bwtYD8xdYqbOxZFBXEPELEq3xpQ5268eypVp7nV3baA4CIB/co2jBN0BXADOWYkk
9SiyqEONuzjb5CIHuhEAh8+R4Eh7RNcQUMXxzs5uXYZJvceVUC7rvUo6/ABiq4fU
fzgmyC+h/DUmIR0gk+9v9twx6gj/67AWyQttqnCqMHrTsW67/hb54dcn6aUoIK0l
t6fem4yakEyo4KX5rP8/QTRpBrBnheP3TrKILwT/PLYACyCo8P5tI1UHe1fzXsqm
udg0HsqZQZ9+wBcCkF9/C8msf6wVF9vuDD/hlGga8BT4lk8KvW9l69RdOkvVH+OY
72+oDSV+1nzs2o8jMs+PbB2n8mMAXg8Ld1Rcyv4F6gRs+gQgN+LPr0cb+OhX46e/
yrmmAotpAhwQ3TI8Yw3Fl0fNMSxY6iAJIZAuk9eyiUFo0oFS5DZGwVjtivZyDy/H
xCwNX740gJVVgU1qMdH6kX+TD5naJpu6VzZzPFnKaEhDOZLR01kVuH8EYqXi9gAK
VnFPxeJSMaDY8sJ/nInGe7lL0ICK8Lu82MOXk19AFQyndrFGnOQoDUrF2kx2+QHT
fljBWIFXZXv6FP31zPURDO366Ai5hTUyi2L5n2SOiVcuN9Bc8D+clNAsUDVGA5jZ
HnW2naGigWhSCsnfna3syuQqf4WRvR5DC9PVQzMb+UnpvUqQy5sStpEVl7YhZ1A6
ca2gxq92NKFU+jKfrbafN9eMxw1aFzdLT78rLLTIZrXbRuRCfznDPt/swIoNYriS
LtO6F+p+dbsJZrfxqgym4SQHZMSxepBD2JWQofrMVoPFjoypIFuheVoYZ8CpsSDZ
ALjQAA182f3bEbTlgU39rkDIqsYFCf2zYPTkExTTNRegIozy7ESuF0tdG2viCvHk
h1sb6HJlUuG0fiFVg5YUTrjnuJvokAEgeq9SrjAoV7kdStfGKVarONwnUWQ4m6GX
0X3rZfR2UBVuFnWtQz/l4AVoo5uq4ExQTaZoTF7RrX7d1eQgaOIIHV13jTsfg2xy
WLW2IKM3Wip37BmCsmeamx3Tyc0amuWHKNEbD3WEI31p1s+qsdUNpldUrqiAn0mW
7rT5qOUUjfgKM0z3/1koXed/cVa+rMLJmNjvQhOAyzvCLK5Aje6IeLrnirDR6/wD
H2pj0tLrQSk2cJdDpPY+OjB5mGnxk6+dOCilW6fM7rA1jpyLrHuxhE0Q/4numX9W
/PLu+M5L8gvkf/YcMX++dJuV58d1jgzp4anKodu+crunJb1LK/g+wk8R64PyEL4E
YZ8d+pv4wHPPMfx/5fq71P0sBmYlPQ4hRK7dDdu/0mFIEDDl965FG5A39WIx3GqZ
uu4uEMh7c2aQxFCfcalbYWqZ9OC/SOFpcCsP/aT3YKnckBrvtZ/FfpV6qwhuAyAo
zlTCYDTvRXIsiGrXckyc+BHUhv8VgAg6GYVXMLyQ/S0Qfq4fHllqhXGXQj29iOQb
fU9Nwaj979C/p1F5FPvBuzcDgn9tf6GsjDgmEyIu2ccTxjWzz6TH+KWOJB22aPBQ
bj7kjid3Hxinz9TGqCh2Ep7RuS73vGF9tC7SCr1Pjsb5QBg10OqIqsVCU5deeBZJ
hgQbx/xnxcf6riQiz1jnlp2Lo7ZZMAE7hCYpgKXmiuhGhX+/Zm7Pi6hSptthVSrZ
lajViLKbl86ufjfD04vRsvDphpBkYniEKsUHvT3YnadsuFHlUhQfmL90yJzb0Ia5
T4Lo+joic6TNgQXkr/NKWsWHFTt0U0mJOEc8TrAUzvKYWih1uMETiV2ExsHcZzy5
kd7AkWhdD8UCkiiqOuGOfev0VobLJTmOZ3pljc6uer0rnNdwRCCXYqkXmgcjWzX0
OAvTXt/HbpYMw/OSFudOnyghZIu70R7kkv/JovMd5+h3StudjcjBNWkZPk2rDY/7
wK28J+PIHOf4iuPLiDahTDbsLbhHkthK/knUaODE6erHZnoOvC9eOHAF5dIg99+Y
tG0/ku99bgGQW9/OQagPQAcisFjYRDhFXO5BRDUFr0XD2mcodgoKKqp9luEEZXXr
XNln5t94MTnaqf9OoUepQJyOs2kR08OOpKu5wPgu6X6PP+pK+mr8aj5xzxMGZSvH
c0p5TQ+Nw2Bm/BUJjqbewDo6YxUiVM5s2aAONJlZweiYIGrDzL4yHKJFaS2WoZGj
sSunAXQ/JxhCll8BEqFkgv6At1wFO/otpoz+1s0ZZEH/ePiPnCmU8v4oZuH5BnLc
jEc3boz1o9JPm7AEYJqb1vX47kxinR+gmsp3fAJYvW04ADQd6/0tHmmfRi1cxg3z
fifIqFFmJ/4BGDVi2lwFKyKNogU33Y5MMjjAY+hbks/pOrrzZJnzceC/rGg7Iwi/
Vs96TIQ/DG9xXgofy8aekeLKogP4qXazAkf7AdbsZWX0yvHDOswm6dYT86FNJtrU
UnHYOZZwQtz0nkSbJz/G5/umnBKkzL2R2vDB1S0g+ZJ501164Lzd5t9H54wZW+HY
XmPJkxponnveYnnRp+5xI+aU0iYxoHrB1aRQTZUgjAnnjM+iNwJpZg1/xPtv0E2i
fn4fKzWKpUmj6kZz8S5zTQhbhCNId7xVttIw+OxyOeJJyKCDkqsIFqDmB6+uYoC8
ZCBf94lBdJhxBmX7n2dZCK2V9QxLUbwIoIg43cXPjKjgyveNW8GxnEhFxDBFH8Ft
XK4ELALzP6bZr50wQuIP55MTNVxxbMKqi5V4AGVQwq14rA1xSoSW23rbognl/g1v
LaNUP2iC8gO7CdsnNgn0d5ACfNyM8dOb/NJweI5XTR1hQ/PCFtVQFhl4YCgLspXG
Bg965/BYU89+CAPjQyquWe10xLS+0VxhdE7EtdtfJY5y7ce2UqfZbiMNPbmY0prU
cCM3BmV2IQWTdHVwOkscJOeh0CL4ZUglw+VXHSYdnD5fML/GARsUq+fMebxooOPw
Iapohh+IGNbqwH8yH2aaoCQV6add9y1w0uQDDFTv/lzWOBW7h8UlhAc6IKRWfV64
PI0FXp/4bwV2fl3Wq16t3O6AgYoIpMBHB+IcpBs5ZsaKzMFIKtpvSgpKH9MmH3mn
YH6UT9TMcm1ug4yTGC8kJpikxF5QWHmBlOUlqUoZrSq3RfZ4t1RD7ZLoguzjtkv6
U3DHDhTn/JTz1uf6EpgJVzRYM82YkdHMPR3gPayCdklk56Yy853rR8iwY0z+nRAC
Prl/vR4w3aUtZF89LMwwmFDM9fb7TObM1L8GKfYkzlW7m3egjFQPdgExzhQhtspW
DgJ4S+s30jY7zCO6ITLkWr+PBqzI1wD0P+XBO0D5il7EQNVQ2Z9i0wSMS71xUeYM
/Xq8utnSjm6/nRRrFFoPvlgPiLMHGDlxOnVSP1/28Eo8FncIq8kaN/NtWmag0LR6
iA8hUSSXPp9oeIzI2hxncyoP0rapJ3aaPq/d0wHidt2xh98VAdVA2oCwsKzs60yJ
4QwzCzJcO40ZKaPRcbHxunzKPjqyM/EHAnBbXBDGVoFgORMDsJOYGJdMl6J+UyAs
/4OaeEVgzD0sMkeyOncxQp7wlQvaB6/pcKOCqrZfpyh+Pxm4u6iEgCO4CqODKJkS
789lWPYrbu2UrnoIIB4hAyyyWxdmKjQrBRMHjfbMJ/3q7MWgv+58B7d9ZHjuqaat
006IH+R2bGHsiI8uY5YIUzfv47xqyDfc50UOadfctJYlTIYe62xlftuvpYP6Yinq
T82puQReFspoNF1pG1nlfZlgm7xRHQeLbI4LMl314JGjQUfu+bfwMn4FDN46Faq7
rYylu8BaYfNymwqdJOYaLR7llqI/Qvm3qtL6FFmXSzgespU17oQKKXLHDK8GuKpK
+pITrbyOZKqPq5jAUOT4hvY5Kt7dwevJ8WzI/Ox3YlTrBeC1PhsNP3xydc9vMdX/
k+Aq/qPvvee8Qt4RQ5uRhGTthLoFjIKt0aLH7TFEInDLUel2zLS3p56XtLF7fTUL
mg5DV3HHXLL/PZO/ZXCeN2dKjLWFC1bh3WzlEOps053j8zqREOZFaa5PmMO08eAZ
ALuh06bW4Pp/uHPz+VGOQtkEcpyDOJgUsLvj/5dz8o5Utp6pLcFC3oPRXqRJ2jrW
zAo+xVIZtw1Ed2U4jU4T6j9sG5enVzmB0u7jLB8zYsz9wty+jn4WTu03IPawRZbk
0vE37Uit5NxwAv5ZozVIFX5J+X41cUYanp3Vba/rfHV432vsaUFwxNYknj/OaYIr
FEz8j5iETE8wnYmZmerMwyhEN4r4lk4h4OyGYTTgmyiD2erqhnVb1XrHMii8NCGW
FVeV9yTL08CzEs3iEu27lRcLMlAJn7rrEnnSZAkEfw4gOQqzIHz8j9rluYc+QlhW
DITp0rB1xb4KscZMMCeRXc/hFW8rDSmIEiw17wIFEpc4+gRljWO+3j85TOOwcjVB
cuKTF7DExjXm5V3+sTZ5rCd+lD4+tIp+icOqCUx+aEmFtdlr8843xrbqjTjJ286D
e1IxFQARzj4NYAsyR9K1rECQwKf0TYMPYXf3RSCzn0Ptnk1wCSKI7PF3OKZIhB16
oROXkdsbEWIkHkhDnxEXh6ciscogp1NscRzR1z/n8iJ8Q4xlX/9DTQ/S4croDwby
DZDWkUb7tJiQSYh/xUUf/D8pzyqQopvef5K3Z5EXqkhDnNU1mgvgDB4Luo56wJg/
znx5Mvpxn3lFNB7VRQpbD9WD3bESnTOm9txwnG8d2caCeRvBesQOVZx4xbS4E5Xd
tFNWZK9ceFWb9eqXz27BsQbBtOZrzhp2g8g2UQc3AARiPkqy5koW4GkMaIKukPGC
XZyQo1jmvSXejVpQy9aXl0bSX+5pNBGShxlLr8jcGJIS2F4AlqSaNRiRPDCHq7rL
lx0WxkIaYv8BFM798cpmALeHtea7x2em2It3aYHOf5pKeag1TpegzP7HoQ6Qj2cg
DzVgLqExOujSx8RBkIidsQUB89tDf6p6cdd2tYKI3+H/XIO6MvA5lxSIg3DbqIal
5oqavvoVJIXcRB1uBIyO7QGEyUTWHumSn/z76HZz9DeGvZR+qw9596dgF00t0DCE
GPk7weI+We1dttCYHY/AZz/7XjsTWVlKxacUFioEeRMf4eSgYiDflU2uVhwAzXr6
JOPk2OUAig1fzMe97+pZdFNQn3ZD0T4YK14txBQA3W3bNAK3xR8QquCDjZAwQHxR
fT4+l4QtUP4W/Vu3gkKZMkqGyMgNA20A62w3EazQmrlYnv3ztrLUSZEXdjQmfNPR
M8nk4Rl/jhKWNo2pggJSgnkNMn9E7gO1H1GYRBzyRWfDoEYZmqGTSBXrarXSi295
C93OKEcx/Sx2ijSsmByLRohiiHI/HK1Rhfqm5WL8yahWcNKm3jtqsseniOC9BaQy
O4Fj4MiuSssZ0ajX7/uSGldq7Btm1yFTogFpqSh5HCkU6eIdfkTScrfewLdLs+GM
kRu1meCB+2ceeUK3eoo7SURo+2zs89CVgMNtJuXO6TYZZq7UPfGncsbGS9ESrsrg
drGZ3Z2ZN7WXXFY0+aSR5qrdDLry/V06Gf6jYVK5zbNUFpQxhFxRXr1SDAiH0Lf7
IlEHoPTUTOzASlwvkKULjEcGSKrOvV/ydrlk0+cW6FhrBi1vXIpiG942btP3YMol
fZLrm14mtthvt5AlTj5z/IYDVP6IYRy1eYC1BED4wgdCPQ+qT8ZqFaGzT/5tayYi
u0ekC95L4k2JJPKeZHeqcWgIMCopnU4H8T+V6KOJ6qsZhPtlGMSP+Z4fo6HmOJ5u
0ASh8RA8tB7984tAUANulcK4I6+qa0uyhdUNacZdOBYUW4ULUgLUWgOjJON1YheC
jbF9WaAbHeJxCE6vRb+b98GM+vQ7pixVwSUdhYd9IAnB5Rhbv/F8j+t+0kWXVkNL
EfR6dTB6dgi9ZLZk9zoCaJyRjI0taXVStCXCXua0DobO2sQzHLt6WNoFgTLYenfK
xKa4BxsHdllz2xJ0wlO2tPcUqiDODAjNsBcCnHlGVvvTTotBQzoikM7Eg+ntbwu5
VMFYjYmWfo4AgQsy9MFOSEbR7ifUcTXXIPVdfaciFPD3VI/6981OizqDv+LQunZ2
E1XOQV1no+wHNpYgAinc+9BOF7MA4L2Yd++Dv+HKBOCY64+nTd1CddPd1WwiLHN2
kAWGRD8BbH0tUK0cElfhJJzSvb9ljRn+YNU7PoHQdIcxoHdgJgV9/3sCxakB1gwQ
fpE+lQb/2NTsGOwZrMljBwPKscnSmxM+TnJ4JLEwZzvzD9cPBvE49znC2nuwAfR/
s4P88WE9ZzXwsSfvRPeOaxPpqPa4kn0oQSuCFbxEFtQRkjkgmYvfLVAw6QkCpDdg
Ru/0yXQRtzEbkciygxnOIzq5RsSSpPUpu4r8QKenV9x5R/52zTO060oUHMfXJj95
fsIu84d15ni39LVjVuY/3F5mW5c+u7ceO+n0zm2r0E/LKqH7A++qepz4bSCG04aG
ALVQ/xubQfhdd9MydwUUeMmxpPUCSdK4vbQiu1LyzdUqRRg5FoVFu83EFiJnBJLL
lQDlB890y3kxGCQRnxYMo8iLU6TX9GxB1iZwW3jW1zQJ8kSEqNe30WfRnmOqqJ+/
nVfsYrAoBv6c6GmiMZsioRvs8Llu5cLFF9Wwlfw4WqP2WDJlfbgENBjfLxHLo1DV
G/UlNFBaBn1ioUR7U+0H6qCO03HFi3gHHu3xaIWplwh82gHr20BdGaG8geM4panm
y3zIPDNANOhJIpYesw5xduhz3U7waiM3u7O8Po0EpF3wHkhCG/jgram6JSp6KFTF
Wy6tuZ5MaYKfFFkX0RdHuGxzlTLu0aa4sDjcruTTDKLjaz1UOAteWGfNgJrvFPWu
xNqpqPkoR6KJL5x46GQ1J0PYuqvFk7lGBCu/cQsc89LQxE03l0e+OrDT81/5iiYN
cA7HggoUSpidxxY2m+e9THdhERrAdLVTR0y8UTafE+NNMm84SJxMaVouNAQrz7bM
zr2IMJ8BzbfK+A58/soREb1t32pXdspbyyrzNU+JqnVJyeVISySrwqLB5Ga94Pzj
p7U3iCeEpYQPVWmGIygRW+8ZRE1WOmP9AGkw4QJYKPTnUBYaO+W+tSJIA+CYk6nd
jUzgcOKcbQEGSl6gdE6x8CS1t056O8X8kISpwZpvnZ613DsV9pefEtzsIU7LPA1t
fK/IumDa6G4iXmxVoybaEwjAqDOPtQ5eYzq0DNUUNxE+ad48dujDuQ7pIeekbKPH
S45o7xs7XeVE4SgeX+A0v5wNTOI7CNmELvk4Er0OuUphuqrar+VblTNa+2V1nfay
PYlOqJVwbEmo/C5A2YUoFlpAdPezo2e1k6VOW1KNIdKS/IazLq0X353EsrYln/ja
jwCWlaj9oJuXHKcpJHIg0wK+SHfRWrabeZt73KYg8qJMDB8hq7pHJL5v31dxes2/
4MkmeTIDjofbAjmt2CBBqTJVHRQ0HMWdwugQM2apIg817wXH2t/w44+DeehjdZOK
ZVplyMQKGEIbkE4zit6Gd3iyoUrHvlEorREnHC5Ix9SMAZvkGjt+bN2lxdsyfraX
2HfWoq55o01IWu/PWSkbY4aHQ4eu0HPtXXzd+QkljYY9MEeRfKD9ljo/EkJ8w3eK
CItqtUzxmhR7Vx6s5PNc5Ud1I36hWLKxlu9pMlWM9V0kIK9wrNBOtn9L3QLqwxDx
LPR9Q+3FldptoL4xoG6TBxbY4X9td8bkQxpkBCkQcBOzJs8gnNWbOnmLWCDwpN0S
L3KJJJojlRmKNWt6nbTBIbZ9mCQccAfnmNIbd14lut5YPiBM/vPgYwM4kzaSrDVQ
WpcwMVidbY6rqub2AHtMVQOBlOPLgLptp+N54gLnCLT8QPe1etX04tylxVCkhwnf
XzumCU0u9qzHlYkrxbcQSNbtMOYRf9dSdEDVPc0WtIQ6IBhec3a3I1Zs/6Lblfsf
DnXhj/ko4wB9DgsfSQaqC3a/JUclIh7f7lDVukxAgqmhlc4CF/v3h81iQuHw0RHn
6Bz+VhLL7uqMtNxxLYUCQHUpsGMUQHpKKDionumQr3c885LrKzVqQC/0ZBjsrAnD
UdytI18eDYsKwsMFXeOKUmCeX1ZSwZst7k3RsoEYTsTwK6tuHLfkeYE6RtDQIVSm
ockyqBeV7+P+49T1ii9bHHCliRN2dU+wzW4y2a6JaEkWzHKweVn+tF54+3S8da4o
jBngJvJkTEBBJ8UCTqIgfHIKiTaGNkcZNx6rpddy+050LtgoRq6plWUt8d/MFUYe
QBNImjMUSi0ZzGsSXKOKgl3oBGFLO5y6s+R9+nU8gCmzIprLQ1Jy1r5CzjCUhN5L
Zm6+uTht02VQqO9VfgiYf/E+2GsmShKXzkPADnyQRFxTYXIQNu0g8TEk4wwbWoSJ
h24CQ5vaz9AMAcJDbxBagVadBtBUlmnesVTBJEnCtSzLCiZoNKYjyUojH2udaEwd
ghLHXf6nJ4DUcpqrKCXjTJ4NBLZixaG5fuX3rzjsL/RUN/5OmeiTBrq7z5qhvsjj
D/j/86Oxh5Da+ZDU+Ae5+WfK8P8yQqQqNK6o4G27UzU03WuxA2wbCT2389UdhZPY
OMvdyia6HHnXYFxYcu63QTfcyYGubVkVlYrQT1t7KK4/Hh+LawJIgZNCGziuAKGN
hjfvGqxOMYfKw+Hnizr+HkEQzLipDjmUcWaStWkoHdK/f0fuXOMHxkCe4Cx5bsjL
+Y3Zj5Wms6YQtuoZAVACNhbryICJ9gBfzgi6o1f1ZPdcTPfkGX5GLtkqG6j7R8m7
HvZNywM0Ko0ZrHUdBziv7at2K+8gHbeNB48xSLGeToFG2Lpl/aYY0bfFw3botxvE
fb8CdALzP79jCl3uWqaunvsAo3fZQ/eHtrqbBBM0hegzqwFWQAog9DMKw6Mbf3V9
x8VrpcHbyXIwz72KdJmU9Tfg0eJyNaXObfEKKmc5MFJYK2hHQVhVkDwEFBr3cwXQ
JT2jmg0WYlr8ww5DZZCG4lt/id39oHRHRlnk/z4xolea8HNEixvrDKAu+VY5V9Re
Dnxac9S9+nME3Jz9XEWG5W+uUSTwuEJxKBOIfnIbpyeiL4zs1Lo4QDIwBN1P41tJ
XiHeJyqZHOK2Bot+5nkJxLDfoC+yEEMTZcIsU0cOLJpIMWSdlG3YZajPTDC5eQ4s
ExtpujWbCR/SrDfVTUfYld0KU+AyHT6YeeADXckPzcj08HtlmMO/Fgq1DfHfJk0G
cmb5NrEvwKsgJrHQUX/QjreH3S7gzbat4hOqvsRkaylXxlfjqgK2iIMPuN33LFL5
UxTY3DBpoKVF7UVf/uzuN0/UTX3mD/hnbPuxIOdBZwkv65XRfTWuyqaV+lQEL8ML
lg8lZfqDi5OTfAKw0ZadjJxLd/P9UkKGQKpV4Ax1e3MfNVOtXP0CFjSj18YMjUNu
kfUrCxUyZq7F3M16PytRg17/M4Wsv+pZU2T9Hs+MKHVZK93HV2WT5KzxfqMHRdzP
5pr0hbkNlr94jk5FZ5SxbivlT1N/wWRLZgSSM7E9S9kYQYwlZwK8Z8ICaAa1/lAi
EcXyTMvmlwxbLQOjdOtq1BKysn1hAx5WNHCWY3MLEf7MpKScPL5HEjr1l0z0hLyR
WTcmP/UGLbJ3lP04wYAzglwU9D07pR8pwWjrxXbpt8o5GpodfPv4wUmCsEDlmZf3
kC8pqTZQTJh73g4CNa1Gucw2B4HCGxbztYri5PHX6xn12IS54v2qikTL1v/Qnov5
sPCzi9dWfZtRoZX4EkdaCJq6dfzrlpKotT1MFv7s+JlZ/fkDzCv1W0ucxkBVV77T
3nmAyZDBbQcIfyFidPV8WnUu6IFGhb27c2fBCc4lx0KHmuqrsqnXNsnsejK+Xmm1
zZ+3eTveVJaG4Lh+5/6BhEdfvTntu7NO2LH3UtHDwsaPuEmXBEan5L2xdygyqBX4
RdeOY+eX32qRpyt6n4KGiV8rUYmIOrmMC08IVLmXBVqVykR4UyidsPqsRiakwlpt
xROeFjTDMIWlLnbHeeU7QXt2F7Apv/fdwkjcz4soKh4/LkhHyOBdm1Dcc63zs7aP
l0eYTTVnBOfpxdU4fmC7IvyXGFMA1OhWrWbefUByWD9Utjn+YPUCDDkx81lMTDm8
VYwqiY5zBNEDwSHr+4u5FXNneZDjvTVoMfL5XKhY3E3+M38meShjfnT9Nm4xggJB
zSszjulRcBixrtjp3nbr2A8SVaIJn1AAJWoSFGSbF3T/ckKG4MD0gr+qzHdTEf0G
i/hC98/mDVpIN7A35wXUD3e20b3Fx4H0hbYK7hYmIXErHG0A6faLTBXfH8V6NWJ3
T9q9V9hsmNkpzyAhGtrCiH4pCoa/EEqasW2bxm0Braf5l25Y9NsVd+9a1ElWigR9
IgDo2fhJUhlj4lUZF+ZiLSrie+dqKvH0pFFAik2BgHLgD0N7gyYQcfQK/+mGpNF2
kxY38DU4zXx2eIrhuF9BabLN5h50w4ZFu5xCj6FHtDT4FQtJOjKpJt3wPP2id8w0
8xTThDRERDSfVZhKVP8dpmpFf8lJrLiwVCefsg7lF1zb5iXPkN1a/vHL08TBAG63
ioZrOp3Qps6FnOCH+LZ66WLCQhI7qYDOXyvj0wAiRLc6YnYvEP7g7fN6dIbHe5MI
ldakg+xTY3whqBrlSElkph+zQZHtBkY7EgaTJA8fGL5XA/ta8WrcmMxa/m93tz+s
J9mbaqoyWcV9SnRQNpeXUiTmr+HVwe8bZHTqSy7hV5wqZUgqKYAUSS+K2y12shwB
xTZv6RGwRsiTN25Pc9NI7bYlQMUgPoY+eUlmD83q7VeH254v9VSDNbNJpKzJETYb
5UYQdI8zPwUdyT5NLYojXqOnueRKsAoD233bAomOPvQvxXV/lkooZwse0C3x8ga3
hRSrvrcAnKfYDzkZD9LX6GGk+VWpaNg6xOiVm1nr0Mf8fWHkNp6u1YZOkWET5DUB
wLIcn0MwEUb6L0f9xbmQJn/l1Ps2OqviYfsOdfkBwrg7oOnsRJUcd1EFztxYU02A
s9Dshdpv0xSWSXrf8Ok6AuG2YFPGtAUEmCbiKI/6lf70hMRUF+8YMB1AYrhYbO7h
m+4IEfnpaa0/FZ2o3Kxk8bEx6+dZLBMPvnE6qCQuu8vd0ABzHAXW24r4KE5NZivd
+/WWlHp6nTWIjkV01jIlDEhtPBEkDLEW1fmwP+rfqgqS/BXJe5Th75YjJogFm/TV
1GKnqNZpdapN2BWu5p/E7L+YY6XQkZpxcFfUNn66WlN4qh1qkG6EuyltqcbscpQf
7UIk0MLB9CzeCE5z45yEAdFLGlkDsFZbKl+RBZxaphTKPAKEMMSLBxu4HGsS3I/y
IPefTIKx0VkH5UEZWPoSoDg14S9TvsD9I6kqIk75aisLYr2CADjdDXSuH60q+pAL
QNFFfS7UtOSOUlBm3AGuoYo8BmdpSraY55YGuyM9I2+at7y2iE1ZEtuJEtmNDs1X
8bwlKxsV5ECrh4XKa+zRVckNrMyZFi49meFm7oGxu+/JwNBcJydNLpW8+hThl2Ha
LCH/uPw8W7+GrS5lQaCNw4KpTSF41VC88lqNhUGfKK9r2B0L+CaBiDCrFD9G5bsW
ahfFCQJHi3n2mokPy2ceJh3+OcQXAdqC6wJjSPuIKryCEOooj4sHS+Kcj4hkBafO
TX5gZsVi5SSMY3tSnaBxlziQg+5Bwdrw3CkKKIfQeZ4AMjYUUeWZTzIa7tzjoPcM
MYEAXt58q0oXRHET/K7W+CQ+lMS1R9iB0Pb5vWsY26t9FNckkwVIu8vWgCcXuqy4
xrP/j3CdpjcmNMmIpwlObjWe3XFs0BfkeyOErergfD7BvbA2Up0euLlb3QShGYvx
3an5PiCzomx0DTUMxvCEuKTN1/7eWh0yYL4MjQ951yhIeO18ArUftWgjH8umvimm
YZ/DvULiCxwlnqW8ocsXvfUDiqYPQsTeqp6K3qI+Rqc1RdEtUkYY6+CFV7CTTrU/
YO1jBrRrmnN67OW4zIOIIZ7aCyB05VQm0KK2QtUFx68xZ8nbOc4pZmQnR3kuD5lR
ZNZFUN3uBxUiuSHtv9xFJ4WZYu8DhPa7s8hssotMpmpaLnkyDXwqMx6ReA9qV3VC
q3p4e2zmbItV2GyNRMf1G2JiKrr+HR43i+ySpOPRsA2HpCC2/MD/kMa0XJ8Z5MBX
Iy46yX1yzk1/hPjZx2cIzHvrqfjBCfXLJdcMEuOx0w3JZ6RjBxukB8nDaXx5jYGD
EsOtmKf3jMGV6B5JHGmKUOZj2xRhuiZJxulLLLvZWZYrdqEjAp4AaqA2zophKFJr
47clj3Y10+S+zxtwbcx+OTC+I+J3jY5D6eN85yx2rRYT/HdN80b/qi8uOSt5fhOF
zn3LJmwPX99EMJ7+Q7FpjDIaAWvS7a3lBGvngPxnCNQ5yT+cHvW5rjLwJ8ieB4aZ
VeguLia33K6qMcYPTlLAFZ40bNOQ1Y0ymBqgLEnuRSrU4DxfnMDfVh1PW8ADroR9
MUsv9l8R7BuSwVXTkrIUFh2GnXxp4pVNKCPbU6IDhS3/0IErjBlppnDOP6HSmMLy
1PVMT6r5KStZ+1X/u88YkTqS4nx3cF4ZO8PQ0LqvQtrCT0INjvAtFW70OKRVp9ps
YQJ2YIo7LjlBhkQEGJBfrX7reHx/JKUWu7rrzyILnR4FDjF+M/N//PNfYehhBapK
YM0hBoEnVyUKeIKERPXJHMtn8AIOq+/hiYU2/wgp/N8Qv+nQvLKu5cP2aZOwcEwM
WAOABBgM14275tbw3lakjg8X+ihf/QWLXzJ/+rcjBronOP9eMKvMQ44iqUH41hJl
vX6imZj0895E25Wqw7y9kNegOrOYRESXx8QGlSWX5R+BBDqTPh2EUoXrBxqkesO6
+UldHD1tj4O4X31GjWocRaBlR9PyY6woFtAdMt2q4dywNP7cjvx+w6hzzcRPNKVX
QvJvOE8pLfmTVDYzXn3zN+P4CHgav2hgHweL0jFQoiI/S2oNaUfXATrUxzoo0SBK
1THUkuR5O2rpFUYFct1BV53UHgr2DGaVjoos9kcES+l0L3+FcRXRY2i0XJjCezqx
a86PtgRrpWAOkxX+7e/o+iEtNV+LPRDCWQJWSbdopB1/LoxJFkyYUNvZh/2RoplV
kDRQU8idfzZFaJ0PLM8baRb761/6tPmth9aLdjUX0eDBRZwIYNkZ3GbZ4LJmcn9X
49X42oSoD+o779ozuV6+E7SvJmfWZBqLGhCjAj332gLUzJnyJUSElx54v1JOkdzh
Z7b7cNd3PVYJNxnLTPiz+atFYPCFCWnnKNf7+L6zfQ14u6lrJ3mm30S+vz+WivZs
K4GlaVjOS96Icsj+WIGCR0J+PpvF9SMxRwAbuIpI1MNN096Bypcd07ObNEc1cC8l
iN2zXkMR8hNxmIOv8OM6L4dIa04yb1dP00ohwAH9dNB1N+d83uLcr/mnkZfFe0Y8
Mcim0w3vpMZDEQpfSs32s33pCn3iUlykK5u/qzLp8KS3iq1PJsr+qNi3LTKzmkzr
UP46WtpF3o6UJwmpHA1B3Kiru3SI6xMqz5qQ/RLkzNxQW+VcDKbEtQ3aNHAX/lCZ
oKBfUOmLXUVeij/54dn0nZAjSQp4D+eT8/UIG2e3zdfcuu5zEVjZoRcMLd8eA6zl
O9LBhcHlW074jae/kfgx16sY7k1srgc5PQAR5M8k2fWeAGC0DOvgh43cyY1mUZNe
J95ItHTWxeAvB8CRgOefnUyodm4h1IUVpDcSTs/pDhXR2t5YCqDvFbDLeJNuuZeK
ylgA53ywjwENjeVq3p2ga1LLUK8+bSYv8w5AXYu/r+RqlRz/wSi/OkMZAAbrIGul
OnIqtjZ+wxZaIHa7nvaPUj1eNTJtNaYUKYqrQPyLk8oBN3iNHdrxqoEXX3OWvGPU
NThgaMLU7lDw6DAYb+JDJCklydhmHl3wcHWE2B7cWt/EtZGihHWxy2y79vH5LtOU
LcW20GuT2OV4pFi10d7usB2RIzlRYaGd60SEbdohmr8W0JfXZl/CQs2L21skcrO1
H7Q8WrX5Rk4XwJxiJCOdlwR1b83Hn0xvrdXHsYE+s/UkiyPyEP7bFhjCRrnHgE+x
Cj3ANn8Rd+e/deikenfmmhGy4nsyj5DtTLbLwPAnVCkOPVTzC57CYL0PqqvOOXvR
jABBvknEtdvzyE8+/xtO9NcAAbkSWUFvMua6BL2YpgZ4TZVHw1k7SMZgCpCj/Qh6
LzvCHM9M3wmcFlQqGCTPGMa3Ncn9St1yW7sBULXRSmPQYOaavBHXgQwDyMDQWi1j
Lx8BMliQNdkl/n6MR5NRIaPP+MQSbp+w2Vk8uHpv/TQ6EMgi9yBuK8xiDV99WCCe
0n015FPkhwEbjAutvXBy/CumrL4ovuSCmr9lNWP3dnsU+fhB8G1CWN3g962K9z5k
WpKSEpGKMX8y3vZWYY1eORqc4c57Koc1jfXzecQ2JNvBNkKF0vHP7KblKM1S1GNc
W+QQL46YHIVVChHMSSY3LKJXXarCj+O67yKLc19efe73IfYr0dvcMXMn8pqRqXRj
DSZtDmPNPYqQSexv7Zgh5ir8kHI3s3LbgKRwrN10ljuer7jDUzooyxUoj8SNm/2d
g+dSfG3dTb7a1Bz0cBJ7jyzVPTGEDkaK+7AqlMKekawRfoL3EGCPJHh3YTrUnVZW
oeFc3FFub8vEhcj/b9vlIfAoAnbM2A118oFbqbStm2IwQXp7Q34kQAhz5u/dtVYZ
VL0Ox5yoVTE8sfmuDDuEqv/iwvFmbT6R5UzXrM/ocMH+SErDryehAQRc+AhQApLe
cWi6s+I2tMX9X99LrWU++prs8Rq/fP4I+v9lsIaUuO1xchJC1Amw2EE2hmOMCD8Q
in6+cFOckHQlgfzPihjX+88lRom+xi/BPlhJIpuDQbzHG4hCvwT9EzINuaS602dx
U7yVS5eXWbc4LtlkOOfbKsz5uR03XYlqxgG0Y52MgeYcS16TV/S74Uwi1ALi763u
DjJLUHHWI9UivTbk9LTA2Yt25A7WEUaw3QDKdzFsAL5ALinYFxj6hWNqB7cgsG1/
flIFRCubmiBfwyrl6ji/hwo+/jDkwgIxRJF6WC1mD//0A7u5beudOsXrktObfkj+
iBo6FUh6mArh+x9iFh8lp3l58g8a83DLwzS3EKY6r3jPuXqPQ5k664gYdfluCPhp
W/112xrqZAMiwiGnbHwnRuPDafnJv6J35fqb/3AHORsRxAnzdiG69vJk9jQKzMuA
h49IMqwspQ5f1rCGbjtbbvl0RIIKflF4F04d74CnwfSOJo9/6rR6xsQyxSmgWL0K
m5xohqyiX1yBiEy9jY8h6At/0AzhaqNn2N4wGgNT/+qcWTKwEtGmW46bcbNgglYd
lWKa0POtHjNvy9KWhbBixTP9SZ1XmW1URVKO6ex4sMY+0BkYwt/0BSLnrgwrSes7
wALyfbXQKfuRTaqXNLj+5NhEqhp1g37tElEb7Cg9cgPjl5Bp/iErynMtDwax7WX3
imch5uw32BalPnihJC1PHa+99HFVq+1FLVRlnV9RxQekcFx2Cmi3pdfV3piqFGRP
aWDia7SUW0GBhgOrO4u2xjKAIm8QEJ1UhMTnWLjHeyC+ruBc+0A23ikIICp2Uwg3
yLaEyj8B8UGqasfqARjV0OHRBx5wc2dxu/eq35j8oODFR3DgMf17NXLAvKmkxRXk
6QVRxjBJFcHLnl0J2rywUbFy15MNCPfohHzMovxNY/8BP6/F/wWoXDf9jk2kP9+e
cdyIy3lD6PBXTEHpmu8MXswmlLFHmiWEOWek6lLlBYWAWkwuDaWkCsMIft+/0pQo
kQ4isLncOvApJouWH2yqs0lnZpIBGjfZWGLBfrp8BLCZ8HFaGbcBFJNTzTXJQ0Xc
BMHsf1Z83U+cPHCbGN0fIj1YDDyD6vEk4Bkd1tP9vvRSd032DMDTKK+RqXIUatcY
8d4oNbcvkspUJ6+/yQKW832syi/+Pj/WbOLpTwKBO3qT2rLD+nxdVtOdFU6fAbys
tjrEZYLe+tkke7lhFhY13/MWEtBZPzXy3QUr5rIDImVCNaehejH7j2VY++fQaeLv
aC3ybzGMw6LGXl5vnw/38G+/aIrIJu3xbyaLKn/+t6A/bGaGpzrYavKkq0PrCmxa
APJnIoxzbMU1hDd9Jf5fgNeee7dFUrODX+jkmudHE1vIfX2u+gJ58jIQz9QtUsuz
k1z/KTeOTtR84GmkuzfMG5wh6pIWPCKHElOvO89hrcFXYn0A6lb241B8NRQVvP30
WLVkas8Y1smINTgVWJY9emk7YW4nctSxqFAGGfdTAo82BWqm2aUi9RF70znN5D+Q
hFEn3aq3AvAfHK56LdWXAtKXq5QWeT6Gv9C57iRqoZpwDLlmOo4vlJyFKrLUJdJ+
cL83VZ1OqHVTHOi2Taa+P9xUpVR269kyfCmMTAKAHssGL9Dac6gmM3Mk4aXjq99U
LLLbhppWVOWYi5idHFjU+6ZDCgzTARaPr8sw1exfOJDBMH2sHrUBYVkvMYcqsdSb
epF8jn6D9vypDQOBxWJMXdS6ABjyvEjDZuHu/29zRsFQS05LUMoUnS8/O2mMURIH
yZmJw+8xZ6bXxAsceIaLxCcMV4bQ0DWXWm+hyoXdhHqDCLFY3BgWqfK1oMhtxNVN
4HFlm5FP0KWft0nDeuje79q9ctFjVb+30a+QPMZKiUQSyV/ufZBknV1zCPERHKqz
lNZn2Xuw83SdQEJBuro9c/zTO/UlIUR4sWXV/hUc8f1LOr9nCbOT7EdmNPnNb7kH
rWilU1BQlI82kgR9vvY5pimLrT5y/LlvcOSmrrhfqKpJW5RqVZhGNbQi19oOsxGU
7GptMR57qGOJppgXc8lO3EP+4MI7PWDZL4SawNzMnXWMqpPn7KNcym52wuOU4aHV
cN4UGVTGh+uRvkLV92koOJctkkKkrdwjM3ix5o2Iyc6rgYIZJtHCbb+j+Qj21+kO
LxysvgQpVrAnCKW2QEL/KuzgamL1omFgOOrbz74t73URb92xdF9GxsLmbnKIL+8R
xeSKpLUjmETzKcgcKaHxIfDsvnyiQpZDQratPKMUXxrvncAhdt7Fpv3E9c5K8EYL
vb3EdmI/fjTx99s+1XEcTnK+EEx1Z0qvX1g1Gep8wx+k8n8y7MuYTeQ2u5EGTBFA
ZpBapNBACLKPej33j2W6a16RDgCQpKM2diH6S8z6+N4BVOuQiYHvL6L8YCMFjqJS
0ZmEWK0hHQdOo37gI4AFure0tmlrMkZkWmxl87PskOX00vFydHmEy7Uo/GbjRX6G
p4gmAlM1gxB3GZXmtWZUyJ5IyNtv2POuWq3LUgHXM0q6lNG5YnAuVZeeml9fqVcT
2x2DTDYk9WcuseAF6QdIjTpDh9rfSnzRWfTIHSjvKz5aiZ+baiS45cqR3chRMG9G
yap1c47n9qAFfJ6pSlwWcxyYIfAmHwCZCxArKa3HGlH13SgWLI1hKRJM5ke5MrrK
vSQON8M3NPdf/OAS/dVGXQmOuX4gdFPXVUGNoLIxYTtirMT0fgjob9GJyK3lanP0
jZkZ4HVcW6BnyzPsDUQu/i3o+hRQJL4JpqWSZbosObT5VuKnJMUV3cuRB9YL3zrn
w7JvGPaFpiZNRxPIDOU9fq2P4eieBJofVtQMaWC780rSM8hqaubwY8sUTdrh1EQN
rjSFTkk98Z6xKDzy42nSPxrOm7LPjAAxus+vt2i/NP1pUflclsRW123WJv3QNIkz
FPp51tTadc9eIS6eIBGT2GjoJzJ/yIyyJJjhDsUvurZG95YrGZqfY6JneQv8wfEs
QvwQN4gRbj0Wdta7y67UYeJfhjLzi5SFAfMaQI3pVIjbrlw/EuXiPa5NszSEcjRH
MDPgiNQv7uxqi5WNbxwu3TQiZhgJjQgsr2cMEaxT5j4cGUKuwr/UVBt1bgWK/wI4
tGDJQfrI5VmunLupwWEOQd8Fks76nyjgGS3vi61Zh30jfXvzQ4XDGaiRQeASCsSd
30e/vejEQVxj1BtQ6AEYUYw3B7zKDVi+TB18yheowIHhgrE5t3r4IjoT1ZtXevE+
n5SIKzOZK+TowJ9Yet9cHi/6ozQc8bQtquQj1RCml9mZ6gkeyxoEtucXW2A4P2AP
7Vj7jSj+Li+CguSGAL7wGAYbcqyZMWQwwAeJuGHbA2NVgdnRRmbaHkj1mOAQu3GX
fAk+VzzK8YMjz0RRBPBN2hQ1xqLR0XxRNJLNR1VcZbfNmoxs8tvbWJm9r/RYuDTO
N/41OMFH2sMjAv+JBdxCm+3N1xvMluJggGwU2ilNSuGwmjzlZur87MOr7bW6eUKC
OM53FDl2m0rBptG00vUX/gFlmCEbjld5UJSdo8j4a40FWXSpzriw5kP75LWoXuE+
wcJpRxTqAlsIAP09Gy8JO6+rgjw/iOijcZiVH8GbMMuZRPR4WH2UGMBT1rPqHHrB
9RaHmpr4+CvnLsP7z3dGZA7MPNPpLz02A/7t7rfst1a3DBa8U3ym+ekzKprnwzEU
upobX9op3vrX8RBD/6P4lxcJ3NXqEATxwa9fottf0TPkztXjyUznz57ORYHal6jz
Jy3a0d8EIyfpoWCOYUVzH502sRy3ZH9PKlmXrM4LtdzX3jzm6PYSdh9TRrag/t8O
FtCoH7J6Kj9DoK4Gx/brQAkq+gMWIvTT3My8iy6837GcRn6DGzZaOzOD9j5OymMH
FLQxGQECQyw0GDIvfJRskdzaHasHivzbSPwunys02GGndeY0bKjoANxFQGKcQA3r
mwIwR9q7dr3HocaKjNfUm7K+tld4Zm/FhJbsnIwf75ogEGOIfxsbV4BbnVB9o1kq
qf31F+K+fEhgcDK72tdcoTudeXqN4pV773V/WfcZ1mrlJcmFAUtbn5sELh52+dBV
GuQjD/dB2m2q5dUFOAVW7ihiDZDn2DVIOq9isdNGJGR11kP+wmWyI3E6EV4F/o4O
n9fy/EMJprQ8/+HuzqBDxVjfJfAv8RiOP/xpUhfDJonKCYCo+/VU4VKxJuXHYqob
EcwQfsrgmdKu4U9gAWb5ULD/wdx/Bi0YltEpxEIOxHTmHrOiy9GT3qdl5mbQCc0p
VTygWNLZbwgsvLWyBLGoxjB263eIlP/MnzU4q6otDyPFXWtPM09un8xQroQISA+s
Fih8dVwNnz1+DeXn2ogVsKupfxXnfGeBV1KTVrbGEN8K+DKlO9z9yqRdvRAnIhhf
VtfVeyM3ThJ1xSyLSh34MgMoQBH4/3A0vh22ZHp7nNM4lnIooErZ9SnySiDmoAwP
b6MuwUgk8BWbKjJ8VDqrYlMX2pKi6MgMUpIGvQORCwWVSXO4JXpGwaGJ4iM1x/cS
iRF+rZ/rrZrnpf5WQoe+tQwIfn0UBr0zhJPXxGwCMrSfawWenA5KRTrv3emd9bxT
SEqKyUYJfgSKCTa+UlFKS5PRWqI6j6GPLcAe3F05v/V1feKzvILwOk7KFeQ0j8Lr
mR4oOc4L+qpSfJxgiwYtgMeGbh/vhQFTPneOVOYDiJ7Mo3g/rh1bTCq55JyNoQNn
hOJZv32zhyE2H2Alp2DS7A4PbrdGG2cPvzyCdZzKJ0g+rEWM1o/v4VQ9y9RyOmHY
0hH2/vz3aa9O02cXycSLKw+5Tnhh/gsxEiYQetNnmtWYM8HiVM3lCHy74/as95Eb
ov4XGpGMuAbraAA1NTPHQ7Eo6flq2BVvM1K/F071o1lqhuyJa1x4qDjGwcAOedIC
jWBhB0J78eJ+K5uKGwn7ZejKbDJpRT85nE5QMvydvHMNz8X5epN34NdSalCONzNp
o+nyb9z0Kczvvyc9MzT5cowZ6tUwy/l51zgTlBvuVZk+gbvO9zlvr69VpWkAIGPY
LPdWq+4gt0Zp5s/fyoAj/GMk1Lt3/vACG10U50bKcIfndSlecUFOvmPk7Q5gH30/
OIl+tiHS/XVnPG71U4AgjteqJLaIKV5pu6DtqHv53hUy3fb7Tu959XNWTtAuhdXx
7omanwtpfPnUYf0b0gK6bapD2xZcYk3qMpcSxB8OEmu8jsS6ivEmrU09xhwMY4VP
nD0A4+5d5ESHo5qXPLqtKHK8Na5P4ZtDPZbwPjq9lYMa7DNIsZXWz8bB+L+W6mfU
LhC7TxbahXPv0r/jPoHmCyGAR+yOo/LGQQN6FDfFQSA=
`pragma protect end_protected
