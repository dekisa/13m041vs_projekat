// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ilHzXN1igLGAKZHCH0dHzsJBI88S3DwIQQaHRqZDPxuT/gJDwEXoBmKqmww8MOs9sfUEHcciumUh
LqwLHFk0Nb2TdiPysQ5DHIhICjrAhWajdwjcbkjR4zwPZMMYJ+mCL4UQkv41zK0lvUeAH3FcbtXX
BQtAwGEW/cv2jnMc/tkJYCU7iNa77E+91i5FmbYJbnt8M6hvhCIbv1BXsuzW8VoErcLrFpK9Z3CT
bykOYBVKzOQT17sED7sTsumcCRsDNenYyRhLrc1DOQltZZlMnuYZNHYWyyrfcqjQK6vOgIDaeyLA
wt1oQKjCHxuTc96ni3NIi7EQGu91QvnNLQSCAA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6496)
P2eUtFnZr8QutW6xAk5N4WH6u0Y/xzPQjUct4N0uJzu25bp/s9nGr+2L5fIeOYXFPJQM09vlye/c
PqNo2/ZCKxK/nvrqL/pX+3RRwH2JcZxda0dScX/LEnZ50ppAel0LVr36XzR1ZiSXkdDX2Zjgcy5c
BgogkB44WLkEgvQOzNDDxiAcumnrbstb23kkiGdI2BGQgm/ME+TJSO8155AiuDSMXTe/TGgDr9n/
2nDtRcEWvXTh+iLA1I2ECX1o+/oMSeaXnS3FHPox8lazkkDHiJtgidZyqjH80vdTmCahL6zgnwFt
y3soSPNs/4uTfQ0LzULe5aFDP9x5epYLI4ZhJ9qRgxo+RzQTGFH2LBNdoh5yGXZ4ypNqSpFP9ZMm
nDblwr5yR98bh3m3mJVphSBZXFbWzuRDVsYLaMNlOTcs3LHTFNc+3+5lOc97K2B55uXSDSIiaumC
8oBVKl9Q4bNgOG40x89olMCgxyhyWGeUvRwgFx1phAYCLhsHnF9CdOYX+Yl66NbgrJIAUPq7ssJ3
EE9JTw3LWe5rOKPEFBrXvA/D98utg6Y9hgIaZ5lAQLWzezACiB6zcyFVSJLyv3qv9pIRvFalufCN
gZqucg2xnUihmbw5kyE+fVB9txgMo13+WCotDwzEA10Yt7p4AGT1FwG9+vPn5zr+DrKEbYsrxF/N
aD0p+pnhLs9GZtcxWhYLQSg3hRBvgBwRM95+ZYaZuxRp9FJ6CpTqc01CkBFqv17SFXdVFEBkMPgC
CvU/HuPwUuOQf/+338Zqi3PD6sPXLfP1EwNybFSIpo0ZVFBIiBPJHKkkSLKOfbKj7V6ykZ6oD6Uv
vfCOmqlk4Xma4fXNj6Ja1wWDZEM2sfodRC1QIbHCC4pYskBWuWh2zUHMXAWBukYRmqqswzQzweWh
kcPVhWSXdQuqeWH20jPUaEGnsAI802RyLzN0QBLtnZ+1UcWHG5Lpa+KWOFafvbgDHxOPwDWsKkZO
4xQcxALELRv4GxdhwC5lHeuYDwIpAuxUjWNMXWcZoa06b3FhyxugDOQM8wmVilkoMA5mbQSqHH6M
MD73J2XKnmF3JQl+DpRWgfSQ9YbcqNJYSjIUyDv1vNJJXh44csTm/CLyz1yEWrSods6OyRmLBZ15
nRr5IUmYlAxmb4Yn0Y/wI5HSs/PgME8MJY8CmaDeCGJm6d/dxZOSH3Psl1XcCLqLP8m/uxzqdJPg
dmuKxLH3Bli06repyd6b/o8LM7qLiiihk5J10BEs+PX4rKeL8d5VAsc7uRb6z7/96UcUGQupuyRm
FEHTaT/axPS7MgwRThsQ037645guuzIGnxYbhUu6XgUAcgx11DnjKH+fcBtwNGjk0V0/w2qLkTc0
tGiFUbhQmi0jkN5fJUbzdfYkSRdc1HYDEUW1S4+4qLt7zGFLRtQU5DzkEjdp+iVWx32MOmP5FFo7
FzCGdfEkanea8Xc0BwnTFntV65+b/o2/y+sPn7IutF9Qzk0kTBwXc6mdt7XsLckuUO7djJG22/9g
kfBoEWrzwaS1VwvRSk3ztr4ON33lvXB7MHV+o+xoxpQYD6eUMBU6H+uUbOWn5pl/CcdwdmyIZpTs
pPLCafdKPdZ6cR97uIWGKtNs0kV4FVYSEvLJItlGvCaz6eW2FsJmTZidDLE0J122ZInEHMZe8PYs
YY+QAGHODNlcUA29gmvkYa4OVXgNLhSTWZNiPhhrMFUwBxflJbotnMesjUVMtC/Unk8jP1UAxWVU
NAeu2tBMsBT+9Cma/eLFyH4TmMbpFVvQm8RPRnR2I92puviltYQ6Ok6+FeZV7lDbbs1asBqzpr87
HsaMLoH/yK/OfMCyY/3TO5/kcHvKPPWoNqnOj3LJWP91xg6GaTrV9jgmn1s+ILxMvBUVfKzk7dzy
zEx7VTMy03wPUxrgxWV3yntUCR1aR1tC3hWV5vu0RG+fYtP0yluLSyGvFylgtbRQlhM1CgG7myi3
lF/gXqSyGHP2UNLKvYNYdE5Rw+pgd9yUwO3b8XePd25R0GTernnUCV1xiS/fVvnudZF80uIegrHY
JRbZlQoC0Ce9HPTpUhGM8TytN+ifc5RuTKVND/FGIy25FgoEVyjzo3a/paHmrN/Q8q/mU0bEHoUV
M1mATcR9wlIiIdybD7sCRSE2KePcSk683Q4HIVkImA9jnF6Y3opiIWbz4wOv4Dg2BFLDqd/kLLvp
kQVcJGXBU4DqZ7odHUCXh0w4owQqhsFoLz4rsJQEUPe/GrSybEvW4v7FXjpCeDYI15Sr8tSPhKiA
KXMQuMf7O0Fhrs4KEqtIWSVb5iMzhEbr/YfPWxXDi0vaJ9Gw16tbpWSgdMwW/8nuDJckUJnWMkh7
4ut9fniRnytctsTXBOXLSFOH/AmP4+gZ6Iv1byLVZnwqe9p5KS1extHR1qdkHrc5K8xu9NGQ8yOl
FmHzMl8omXgiksskq34OC0pR1/7+a8k5LCExm26pHTq+cmKy/mTHdWF2znHEb1QgzkpHD3XTSpqU
NjO5Nn3IL4W/hrNCgFLIc/VFid2L8EaXDGoee4lo+jLstG4SVCZB23lyObM5i1LZSC0BHhUF3eeh
uOPeuXx9vodG2lF0y+07qkkS3yiti9eXYrSqmx7prm0fCDOzR22zye3l4Wuh5/DSX5Kd+SNh/53A
b1aUYLJPOVNUtpduf+Re28LU4tXvIq0W8NZ1MpZyRVQeH4Yo18kVi8J8v+7OEK3El+BYXZu2jeYF
CBUW8DRkp68B+j8FwbDpV3uLYad/UA0rtNuFw5MjdAYjc1eiXbuVYUScOy/6lBhBsoWzt7M8iebP
fnHRR9OD+55OPgN3EYRYxUNEFzItGhIi6VFI7bIvIv9fN8B+tK1StZf0Y0Pj1rk5ymclXZ+MsyUL
gX3zyXRhjlQmTEmUpVMxWbeTWbg38EBEw20IDgU5APCtmRyA7wWEbi8kdejL0TLJgvrdM2nBGPj5
hc/sLgEh+/iqtSEdQ53g3GDH6s7vMVI5J7Hc+6fxBPcj9+4tfYZ4D5/b9LgqwaqwmCWrzJ5MCFU5
XUXLFtbolqVzKf/cqnsAyKL6vXZSbG1B3mqUYGfO/orH/mpNEZ6siCVXxhfPuCz2UX9et5bmeZlS
wc0QSuPxYaLBX17YIJp2CcSUW6lY0hcLXODN42Cx6B6FrK/70Ba4dnYeWupXRRRfWfAG2RbigKy9
Pc2O+fLz3WETZ7w9fWm/nSOgbnCuc3gkz3yuuK7Mh7gkcwgO1w7wuNmkr11L1v6MM/f9IwCEDgVX
bVe51codbX50hjqdwr/wvkkN+6DEwcOtqqTR9Z99Ol9r/hd2GsNJLyaFYTjgzP2VxtzRNpP9d9y8
OPNi93CAnk8cS60r0ip5Tc4/jzyav0iVzIuCZE+46jmSC9sRFTkb+Q8JNCLikydL6mJ48vpcio3Z
8mL+BMVlnrlTW8jlh4+9o0w5OT8ajxPqJFj41XmStCFWHwj8Mbvk59r4jxpFqx6co0VDNlQXQcJr
9Dbg8UBHQ6gj1Nw1TSh3ADoDAZpTRNu1msJqYPlBHDID0FJCj0aH6n2Tt0o/uesWRUwjXn6jyCIM
SeTj+IdfufrNRleGth5at5MkR7J1isR4tMxrMaq2sY57/R+qSCLEy1ufF12z6uJmCD22XxuuINHK
40fciDp8OozrUmNkBg1UkcEe1BITmBySt/VhPjlVC50hTISGpCuI/PqRby79ZCo7iZY9laSL6jdp
TWII+SFyKnwyhsL51YVI+0SWHiQd9d4eBw5EHP1N1tSGY9JFCVwnaTnT+5dcdbxjNeC7eTkhL3Iu
4TVhPNxCr1ltYWJvvOjfcT8MesAXcxbTMMXkoTpxJaBx/FkAaxp79lwTmlxp3UzBFrVblrwmtmsD
JF5Q9qfD8pZycwd92tPOjy7cuVv2Xh0ygW6udxB1jMu+QP95uL0+wUB6bWghmqniHpag/4QikOC+
1YLAF1h3y0fEEbPu93104FzLN4IXmgQ1wvzC4XKMluzX5/C9d/zCBla6NWrmuDpgODTxmY7fETpF
0JK8KiOrfNnEDarxm/xGK6QVfg4Yt1J5XeOgNvZiJbpIUC+Jz1IA+vEL+3guiSW02QOSTUraP8/A
A9B3ezdBYPxfNCQO3AZ37ipmxyY71avL5y7WjoFrey2H936o3wjhWldEZut59OFmagTWBd5zSOqY
p8vH0Lix1c2xTsaAWopxh9jK+iv7SsAcuzu5hdXDNq0dTE4URizC58Zctufb3Iw8uxGrfyZXDubB
MfXU3aKqH6Fady5Rz5A/fGiBhqMooXl3zK40F2JOA3hmypGsATepjYMmO/SYIPhhi404E8CvMUSC
X2bAHgHRRpy7VOiML13NYs/orA3AB6tLtX0ZuF2lT+DlzptLkJ8ebgCJbF5qZhHsGjreFRYfmk1S
9ZyaSG4ezI/QoJNX+IRctyNisVF6153ngRx5eluBtN2jJPKD7KPmbTbV3c1Ijc3miiGDEHEFi9RH
yDseVkVNYApSh36u3E+yR6YvGzRLpknNGCBgf11BdMYHCoLrKzIUdbA2z3NSvpVWn0iAbs24xaHh
+jILXUenl0ulYVsLX46mrZg7KreoVoLi48G0itRWZq5RBrfIqtDu7gxI4y2CWAc85c6F7nZTY0GQ
d48yRjuOntF2NIhfjc59kLfB90vAZW/8skYN+NIx8bYjegqtHFEwo69weWFYFd1y7Rlsb57HEREM
rQ/v8LhmSBg8+HIfdAG1u2w4uYuPkHBt58NjprqiL/wh9WghyP8hEB9YOE+MpjPO4h9+uxUNonso
vaq/a/HjiD12XnVMsRlsXON0fwLGGrvGvqDbo+AZWtdMoCMZQrJAVXuAUexnbt1ZoSBXsSljDbGx
Oqg8HmI5FMDwsHl7Ch4Fbtty31PJDlact9floj272XbV8pzfa4gAZvQLjJ9ITVB4AJTf8B9bLKOk
rkj5hC1j6j2Ktuyd8Ws1uN0drYUoQnB2sdvfGPW9UeZlIR++2ODps4/eumADH5X/b4FVr8B0OaF9
D9oZERQy7uDapeAVID+7xMQ1E3dYeEHGY0RDAD5YGnAtEuHzUG8JKfujWHAqEc8yupGTFTf5vXIW
fUTE/eEc2Dk93lvymerMs5tOfaOT70G04iesU7kF4pkQCakVEc/w6hlcinWG0Jt5009VOQHhVAFK
B71RUaI1YCOJbSEyQ6on6IQFI/CXKRMP7ErmNJyrjTcjkJ0KpKp6eMPBc/STZEfZFZ8/yQ9sbpO8
B91Ztt09lszDFTsE+p0zAtVwaD9XyRbbrHjKpZfuFLu8izofVc4CQQpUX4lql/sGIyB3SCXYX6GN
Ytp9S4gTGYjhm5HWlANVWET8jj2QX8uM7X1W4rHk7i2TpMDK9E7QyI37bGKtJMG35Mm/73Z/Sse7
szU+U40LQzOJeBN15fmrQIrnIv9s148UqypEXh2tklfBa+NdktAt4wCZoqchjS/46ndld9qspTvL
vT812XIfSi407iQCT0l7I/3b/4HOU9tORKfRhruYiIWpOx+7uMweyvz9T3d0WyAtTowOTOyX9ujt
JMO84ZHYH09wyIV88FmHnZnemYvjFKPIx4vFFK2ZpHgyaudq6cq10M6qWfxF53CFa+6JgNuB8UMz
GzraKhcoUTFd0l4s1DGB0hkwFNd9HwiD7D7/VyD5x/VKe++VIG39yhiqzu9Td6SyTOyCOaf42r6y
goiq5AXUROYEq8cWEgb4gz9zpuVKN046wKxOsCYHs1MNcs66Wbgtd46pp2vjSiv0v1mZr2qkKK94
akWybqRcpfat+pv8NF1VUcSxJ+AnmboiIqCUCeNkgPzQIzJ8WJmFNTnxkitJhydMHDZWYQt+fbKi
rfDafNwwRfCQ1A5KZarqWGYkxDGPeoo7944n2WBo9o94L7j/hx+EV/BvdFQKNokY+Ipbg7bLipUd
eSa0zZQ9aIc0aDYHVeFfSWaMMUZlWZhO+1A6n1KwRSZE/P3RlUG6Dp8H6ucDG93A7Nuc0FYyBcab
a4ZjBP+JbK5MEhZ8CSfQ+4kLf+avG/7Bg7Sy4o0g9e6X/Pi0t8LiEGtAOBTA+tQQOgjugACkESIb
AFVkI12jWsRecJHwmM/A5iJI/qZON2eHoacKEG1V7w35P4KXNq09iwizSkhbBqvBbheuoD8IkAWV
5t+kXRCDEHtwGd65Q6KSb3JjoRUu1VmbR8/DoVeP/87Hi3BYb+V+rZ/g8OUBsreCyvSy+QFcbfvD
oO6bkM66tuz4RKm6vNyaCYgVhQGoIv5lYNfIiLY7826d7djQqbL5/12t7PpHdcft3pGT87T2xd5m
Y5xt8i4IALM1+lBY4X0DIMqw2rs0+52XXt4IdGICenMRBU3DgzvfzIIpulbjynYbbj5MBABF9Pau
yW+N2JxSIYGrMyJbihuXWPNoNZpefufbBM5Dt9+oQoMTEGllUy7se8TeAueA7Z6IAiOJ+mt3Mktw
xvmp22brtFod5WbvogVNVhudcQpWmA3TkxNmeGkvfY8nUBNpc9Xx2x7UW1nA6Vu2maE6XeEgyEhr
BwAtPi5umLGgoz6ockyV2+N83F+4kvk2TinMyTvOTvCSgqvilxVZetvfoE+rQX0asfvLxCsEGj2j
/7oMHBdpmc4A4HjH+2tEOTPQk5XuNu1Z5JHHpw/uucyImIllc1OII7+nIeQFKWeP1eI2imHe0VcH
EZGsjyE6bOT37w+Fdy6r/agwgPobaxoKtNUO1h7RJGsljg3oFwM0CVRPYTOwtNYIdqb2uZiG9xAt
1/EDkyHDgfHZMmFS0h7SQHxJtIoLWj9/8wtstKRCkzchCOLTQ4MT6KzQkajdgAKA75xnJ0xL5KF6
On/hEy6subiJ3ugAp9gy4Z+FfU/RX8po7k+GVg/fSnqKAgrvY4Aq2yh7yDuR5pSnr78F+HrtTlx1
JmvpxZRpSA09FX7EYouZ6I3LxlQ6aPNmx/Eubg84+YBooiKiewl9ZKFh9K803/rUCDCtS26PALf5
W9YG46aDoBWJ9yRV9ak5TyQWk4Os6VAy4kgKOlGT7JjchE0aTB4lbnPHRhTaROvvWj+xSDu8XvOZ
+9n1OpCbuOvsJHxjyyQ0zAGlDDslHm5InWwLQX1e3z9CeZ/C4sT5U7fMD5XUrB5tdUSFYa5LvJge
R1MDK7DkSSmCcm7CnBuyfmvfi/XsK04vHcSTlqeNhh4F+lrpyJFAEiY635hnWKmVuEbApfmSqe4i
GGV6HdS4h3I/LmC7t3S4dVbucXB7RGKryl0Ju0EmhKXZhdPjvdR7tc35t/g0LM+YHuRs3OCv0j3X
nBwm/E4Lc3OzYn57X/1F+mKVbTqRV4Q/6/xcueki8Oluhf8x6Lba5rOUG/wly4ayZ4z63rlrhlEJ
V/+jgCZGT5Op7sqwDc6MG8AMU2L6LgLYoD7rvYP/B+guVsFFTcQpv912FiD67gkUYQIfsdt53Msb
3LCuzscC/eszO0j48lDWBoMniEHS55VDHjt6HX/xpR1xevbLFbplRY2duujiMh3Pg2SrSHEAjhbL
ROstvH/S4KWspHBirSgw4s1LedWS3/JtJV+u+Utg8uKoI6n5v7RuAFaL23sGQYfPHXgc/a7mLPrg
vGLo7BJP1ri9rYHNUMOMfyt1qXrqXHJPiSQWvAlBDlPTCoFUeMtaUeaeeaUZ6r0UiYMVm+9+WkaM
RPNQi9liZrTWTBc0O+7RGAe5XN08vt7TpEHcm4/rKYHQ03FsiWUb4bjkZYzd9xPFbOoC+RX45oLO
/aI2PEF7Fm8nTj1IdL0NMXLFcQs8b057mIWklOBwzr/1R2D5U+jibenyJ1E5O5ozF3dGNwAwRM+P
P6/gxwRuQsKHqTGsIkCAkski83YZb9SRiQVCl0bBDkHI9XK0Oi5psQGJ1LNEds6T4BF40zfioh03
z8NvFX9OAQcdjA65rsTyCjDRrq8xXv761mhnWeMRo6OjMuIiUTcF/0L2uGtYdg2SMIYDGpmM/vz3
8+Udvegbz2bM66GVz/TO3N6REqXd0l9/z/dB3u3aI/71PokyAndnpGCFf08EIwPI7GnBTQEo6key
HL2G66omIRMOXJXWJlq5Df9if2IaUvFPLuXyfbfN0zMzbopPuApEtqJFUpe3dpmlJBPuZq7MjL4B
2bzM7bfDyaOKJ3g4nIisBnyzRPLGiTGMB7R/eyfzxaQhS2MJkr8Trf46auj7UGZp3ne2noNsENfW
Ek8W0lsHX6Un6hXFSXhaukG/R6Ch2viC9MYf9+TYaKirjJkp44SRbLXfabGwSugC9MELjuBHZDaW
Vqq+xe5gzT2R2hbpcTFq+dJz7se+ByTp7jTm1bsVgBQh+SM17dTNlPf2mDz0fjipI3ip/oL95BoW
CrBb6CcPLmzrGY7IYOKuvw21uKk+C1lHfR2Z7w9eB1AOsLX//LVabdQQLOzMAIFsyafJKNqL3V4S
G+bQ/mNb+GsyWaz7l1J42OjKA9Ctn3W5ZBx9CZEdUrnrhrrY7WjWJItmlUo2dE4x6RhrSDkIjxVy
9YUeeSFvafBfo2EDBVDShmlMJmwTELuiC6lbjrwvkWKbalPZ9WsHy0ZrryGUfmSQhm3cj8XLt2gl
4LFsNpPUyuA4l7Kj3bj5bd2A8AZi+aC1IaEDYLaBKb2MpLT1iCGBLOxDDseR62+ik4Ufsp42UA==
`pragma protect end_protected
