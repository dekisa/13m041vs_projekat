// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YXn7nP8cauz5cyou2vdxXEcHIZReWyox2+QfmWASh6lFExFi16GYFFGIb9gGAyef
vQvB9w4l+r0ulyBOLsNespgKycJQ7KnZwkgdxqC/4Smv9T7+eLdmH6trQH9vkzvy
oEzq17Ur6bHRnB/0PtxJi/KWr2YLUPEvOhBydWD79lo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 66768)
gm6VulNH+3v6v/Olf7IYcV/uLev5bhrDiX0E1KaiMXy+YvPD/mTO2zh+Z8Rd0d43
PQMsrhTLTsU6wk6cmBzP7OwpWHZH380f+3kgQpxAD9HxQbR5+lWU18ufbEpz6jhE
fX6YS6Stw1JOJHTJzwS0GkcglQve8EMjmxbMpCvaI+m2XnUTOHrcNfFl6whKke40
gd5WVOwi8HTPdOohR/cWYIZd3TmBcPGKZC/HKaxpgf7PrGPWGlIhTghro403uVxV
U9/c+akBeodxz+gr6t3rCVFI4iu5APRm4nRuB+HpKGWeeNCylCkbLLghO2od/5Gh
+htZOty4Ry343vJeBECieccEVXAe3+fVcKWvBGIzGHaG43ebz0xrgKMEIe8qHA44
zl2b2PUVZVy7H1vPkSaK6gFil08SPInsIX7cJu7srgLeh5VajY+qGq8pTsK0zo0y
RGmaQ1hPfGI91EDiLpiQeZa3j2ddw33Ks+x9YtQFxeWtnQXBucXyi0a38MHICzvn
/ZT3onoISsTTTdEbzUq0daXu0Up0M3WXHgznIZKbPgR43A3oIStwiVKYNG5y82yR
ObCJ1n/4dAutNTY8LpwiE2a1jEGlhaCYoIt81tc2yKZM8ODhZVd6rR5XqvJPJth8
Fn9laHk9UfTKFdUG++DH+SsSXOPLirlc/Io1hhqude2sc1DgHJiDXc7m9rlATfZ/
nATf69aAZl6kuXix/YlPvqdxU6ENlz1RmgwQ2oOOQ+iTqiXr2Vy2CPFm6hvHLUB+
RIwV2nG/Ggn3CqGpQD7LiiMBWiadqrvog2QpzBPrj8blwDGdL6stYfGdjdEK+ymp
RIglikLDL+goqzUlIQWUsD9onYWM8p/zeNnnKcg7x/LM4W7LiYkw4t/SkQWm3UZo
mPmSURYcidRsd6Z5hxRm2lqF195segDK1thvm2jZGVZJbk4eaYZUmzFY3/2QrLih
G0KKrg6nUTRfH979wTs2cdWw4mQBSrNrM5PdN2Iu9et8qsRs8WQNfwWS8MxCvMHJ
6Qkk0D5Ze4gDuohEqpADn0BYarNp3gzF7W++BUMlSvoHgx3seVpdYAXFHguhn0A5
w2Y4mBbNiePFTjKmAUZTjjr9q5ymyhBanyXC4a43jgBUIq+2tx7RXcAgaikT5q2C
EDBygavmzs1n3MYfjPBIQlJ2+UA2bvN0vVsjYGNqiCbKegWuddidXQsYYKFlOVBq
peQGW3zfTnBy2h4tjxaVvmlTfUgS+J3XDIOC0BynJ7isvCMUR341pXj0F1LWt0j4
FUA3r7Vi73EHdR+0OccognQUf3gLJp3/hsr3ap7KkqEK1fUP5ogXUlz2Dc3Crh0S
ZVLip91ou2vRcVQHT8b0PCKEB53kvgA/vbPkITtEwBjLQ4yQ83J6QSoY7wOh8rJf
pyeCqrO7tijinVlHxDkcgmrdVaRBONml9QD1B+nrVMnwXsx8IRXGBVFVx2mWYXtp
bZMH/QgpO+J+xdTjCTyRtOA/tkhA2k6EpHGlBWsaIBEL//5meiR7VQE8o7EVahTa
OxvMnT6YePbv6oyhU9IzJkW0B/YVCuLJ1I3JB9WUoLGXGmkSa62CP6PTgMDjfjAT
L0r1M3dvZJR3gMuofLBPrjvIqIjMU0XAAgfzAMkXwxCBTPkESbHf8q3dAxuxG0Cd
gut7q178AsrbSNL7zPuKGbIWnhAU+jXoZvD0vXdCghm2en5yUNY4fKGEgDR8ELrT
6pSrJuIA6N04d+b5x/LNwAbmO6D3T3g/XRnmSHKdTcdTlC3vfGfYzjmqSPnRmjCU
oqXfu+aL3sC3DUcuYlc5OOg5Rz/IYIf2hDc/uA4TEWum9X/o+uPMqYVVq/NRHT5s
5iD7rjYoxPAjdZys/tjhhcJSR++FPGx9uzG0SYG5IOt+zQ2tb+RE979pCAjhnqj4
OV5eG6fMnVn8m2iVCV8Ps+SgPvmlg52FegeCXV+fUqtoBjUL6LDNdCnq/UCIzGMZ
lrJUPglAPKiDNuA23d8uYN+0rLPQGmEkupOEzDlH7nxh84CqBif7tsJIRs8ObhhW
y4XBe2XW7GNOGu/x/ARrftYb4IJ9/84Pc6tM9sRZcYW2oTjpUnRT3BAqp4hr2USW
xrS28bdTl0NANJbBaCcttkB1pO2XaezYoYdcC/Wh4n+4vtqSUGugM0pbHRy/CgJP
lV6QOVHW5KyhpIHNUnlzg8jS1iO9D7K0It3H4NB1fbOvosyk4v1R1vhd6LUyHIul
nD5kZ98jl4xqEQdS/0vUZO/rzWQIRF5kbXi2EpzM64JnIw/rx4Bdqxh10Md+c8pL
38PjMTtMB4/48/nIIjAe8oLi0A4Gj0ZGPEo5RvMC58BBHf9+OeIRuHFy4tJV3btf
X8eJJXs/sAqg6S+20Ilc51WwZ5QY7DbQLQ+gxPSjdRVWhrMYsJoEXeY/W2++eCAL
XHb0mz0xXSxFVp2c5eA5R16i1x3YO32ruGFGQ/eaA6m7yBnedBCQSAvNgPrCWryu
RlypCmQP850ws/qnXeL35mA3HUod5EhTPHrTSE6tHN8jDCU7EqLUJQ1PlrsU2f9b
OAMp5ol77i13Ku61YmbGAuNYVXXG+vALKqF6f6L3TkJk8o5V7ue41trMDip17669
drk0bS7RZZnkJ167DDeanx8QGKQauyLYpGmZ4o3dhRfX4YY5yM6XXTWOOBv3YJvc
IqEGiYYFSyek1i0DQkhSxTTC45eJ6tk1x/nlL6N4mVF2OXDtHRx4P3zOZbJL9yTp
nYJCHWvbjhl5/y5gUzBT7IvfcdPFm+NFqoehvaLmE0cah65ysOSwZkbz2gLd4XpI
XnCVvpb/3Qoacjl2BN0t+RkxlzIsSJXuPSUtubhApmWjtmbNbH8cCzk/8KmBw44k
i/cB5gJJqWOB9Jw4/czCIxUL16SiNGmQuuVewIVcvZrYawlB7arP+mJzrqpxrv18
C30yzOcI2DUupkeymZyQxIO9vJmL7ZcsUNXkA9tccKfTY0yZey1mdHZiZFwaK9tH
+IG6RgGEBmZDAIiOnSUszMa5002Wurdkr+eELtmFkjse8mZavz8bsWTVtEArOXwF
egfJkZKKFuPJkxH0zB/NQI87dA+H8JrAXfBuwmF/SiHhJik6LCyn29ZqKuTUHhTl
vnTEJZ6X1GfWgPsFDkS9l7J9YyVU3OoCh+/wnSyzhjeeJJttHeYcQKcShsYkh2P3
652nrOPVIkQmQu1nDI8cZ2R02TrbVTPhEaAJuEY207odZ9sepgQZnLZmgwJPPyVs
aNwfmk1A2yDS6eWLTmwJprkaoHzZ8cJejmhGAtfybhEMeS4ymmw5sTcDVPHvxs8p
gIRTZ41w+ANoFx/vyGNDfGx87A7x7358vMx1wy6j08kO9uS5a4DwuUawEAFUpVCa
cpk7BDMVGHuHGby4d9nktsFrf8C27O+minAfYOFswiWpPMlAP13SsvIKa9ZNhQfd
PhtJp9vVUI+j/KXhrGeeolZY7l8j3nPOQqAfqDI5VQFOjBMAdqC+eA39YX7scWBG
zWczUC7Ec5Bl9Zshq0Czn35B+bWUTraO/wZXzyFlDt9Tp4zwcEhdhhhT7/D8TclK
WJVaYayB5yUXUaw1bVv6rNqQbkmda0uLeVFHtasilJYOTOBrzFkuZQTLR5Il9Mnp
wKaG1Rk+rQ/ge9tQ3Z0w0Thcza1bxyu6eDlWFpZ0CqowA68bqo0c4dBFGBAgb3cX
mbuTjnXEmQq0sQn2rgxkmBM25X/eItKmQT98ylbL+DM1PBYwSMPIj0yyvTH5h2BZ
Ql/tYLpPHhKUslhGq3YBhnuIqmrtN0ujG5BiSRaXS0eSK99JuD5zPyv6Y8z0FSMS
dZwOw8S5JEYuC1/fgonAWMoc6gr4XgntRltJ42mn57QPk23Vt4jaLSClvUoiSQXk
oq5A8qo15hHP/kDzZUaDp1xe289yneVj3F3E6T5CYIYhYAuYIms9JCytXl6HxOH9
szmr9nd22zHSD4Ny2+5TogHp4h7A7KzACg1uxKN4gJuHtwAlSRSBgmTuYhVJ0bBG
3CSuLvA/btArI+nt19XezGFxClxcO2PbJqo0VmBGCL7RkZDnAMTrgZzsNOSmR05s
D7tLQ2nBfbnmtlsQkjfr2jYSdJ6c1N9S5fcdShbFGkdmpX426M+2KT1l6iJK5nYb
bgvXSLffAO2gRsLF9ril7qkqbIqYKd1G3Nhp1OMyHGyD8gYyMD6bDsKSCurpF1Lu
mR9HtM8zfBkbylj/Pu0KdMClCudcPsmd+IV08r0n6YUUQPDrpKkTYNDHknBHmx3Z
yNgVx6ji+f2fz+Vky6Kx3WnvmgIlhxl71YljSt3KwRnCE6YxRVCDoUYkgqicqdAz
dbgaTBhjGEYr07cCOYeQBdypT/UVp+VwJUOL7BG3MJ0kEeP1SpnNh4Qbox4OBs+R
9F0ph3rXZCh8+UFBEeUjatLg+mCKANtyXqU0znjFH6/UIrxl+kCNulMkBfZOFOLq
hYq2pDhzcRcl6OyVdMHcyrisU1VIqyr3ZLQlgiAEQIrGLa4AeG31X+UzUZviaK5O
WsuMbtGMJXszguWVTXVoXRo7N45HRXpbeCd6WDXH6AfIRtw1up0BjLgX4Q7qgqGr
B0uWO6hcDitPY3X027GhiDmcQCmFpUvLoDrSxCtKv2TMfZAXtboEDNB9lRrQVO3H
qskzifm223VR60p8iczdMQn5CPXkxAN37OCjAuVL8IrkbsVPrQfJEOO0F3MlhaB9
vMuYY3+GxSCTHp2gofxI8ZyF9jZQMZA1BQdw8F6UpE77JMjhs4IeYWoN2puko9H9
VSEI9MrQqf1ARB3Ik0htt4X8mqDPA0l4b3QumiKnzW1bgHdYDw96K/jCKYvBayF8
Ps9tAvDoN73MWozSkr79oJK5RXJAFpF4r4rCEvWQRISvmumsKqi2c/WQB0ZV5Jj9
4qa83yItEbqNcDnedEb0BnI8uKJzAiUww33NQiOYnYiLBEqUqP08YjLnSn6wwiG9
yUKRFG8e0lNCcRi09hE3QPukApFXbXxMj19O8E1D4OvXfQfVZJ9ywJSPNBywWvYy
m67g4JcIZVv3T1ZX3gzBAQy2BS3zbKF+3FtVLPUi8GchNLRfZxEsEvJpnKCYKTAD
2q41i6WGCSF1iNW1d7uaBgMifDuH79H2VeWqlgrPmQta471mJgJojFDthCmJlccr
fCYSJcRetBaEN87D+HRXnF5/gmNUtxbfBVEgzhXx7YlvRSsRyU9uQrcfMekBPfI2
Jamxa5a2MZx/748txXBcauGN6TmVKa3qVDGYL28FfBuVGAvVkTtLMRGSieIMEPHs
q8tNdIxaECDj69jteoqPiXUFEicqbw5NsZfqoixwH4potPZJOHD/Ve0h7+/vGjgr
8/QrzyhhZ1mY+0XBEpDZVoldiYvTzdiFcq+BvVHWyQ1Rwrjc00Hsi/mUxo/MDuta
KHKu+uekJv/iGQGt95WX920dsPzu8ibeYt6h1+KZYWIIsmVkNbkzVyQt5I7Arrji
K00BddaBsCj01jItPsBvpDMScoAmjmmMlGUJfrNyuSk6mjdeI831LZZkt8S8AlZW
KdfWNfZG8MTpSpEto/WpKnUF0GRKKpo7w+mptpNtL6Pfwiokx0Juy75MNTceC38e
AO4k2IxtxK8GPUk3zWfJh0r362kx3Fn65+yiNeFgtmt+fHZgP52dSLmHpUNahQVq
csobROfHE/J9W90LyqhooBemAL8ROOD/O4muO4RGfUJ3aTh3agSfVz9CsRUkUJBr
1Aibxx/g81O0Dz8BYMvBjdCAvsBPSqgb820FRJI3tk7hCvl49UNYqTVkDnraLw83
Su/d80wTEqcv3+LCkWej72Ji23UvNZ8RAJj7YktZ6TlyQMejsV6DXVJfg8UFu38R
OcU/bFWLpzLevC8GuB07Mg41DLJYbRAfMtRajZi7QFXfwZK1u+KfgrTxTjckWROz
4M28Mujm0xp5t/ayfEWFPKeFpT8CrivCmNYjksQBVPCF9qqxoqt2qB+7tyHVtv0g
+JPaqQyOzW8/U+fzAUY8rLw0zdATUdndp2CobgdRCDB8hLgeY3IkFvp1upKjfBw6
EgbymSbw5Pr7vsunSbP4dXPPaseZggsEtKAQ7WgI4K6HyG8XGOHhfwr7k4Mt5QnI
mqIIZJZF45yIUpnfeZklNX2cTefgHGatZLDaRiDtox0HXimtqTSJ+mX4NgT8399A
GlG8XKuxk7VGzer1CHdQJ4D156zWMQ+IkI/kX+ynqWqL40aQLredMPv+2rWtDQP0
bQpiTZ3xkjYFlF1ObJ6REW5M6al6gpVICbQ9mfKvorLpmsTTQ7pEFCxSzmg/OQEn
Yz4/ZQGZ27BGlno32gB2FoGVHyJTv4k5pDjC74kDn0CGNoRspZLq+2RCLKFwCpSK
rvQtQRWqUDSvu7a2GUQsQiKNm1vr7JIYc5n5exwr01PHnPgVZNLxQq74SfM3puIu
UakUGfpwFS5rLGj3+c8jAqlYfONsNB4pwNp948mR9pEdh2RhuJ1lWsazvc694hF4
m3OBJMz5MalPYDagTzfGKjRT3ljmg95YGzSuezfyZQFMF6isWnpD1/qIt0M0qG1r
qp5D+ojm9lsWlTNMGnVNFZrnQJpghNk1Hy+0cWOiEVVoa55y5dWTFgnEJHRr2V7G
mR/Fqmpb40nahef2LiOJ7yEoemD1NbntLBWY5jB3icKHHwbQOyO6a+N+2NhH51Cn
LMjQ6aVYOxKHd3Ho2hukl1pDY8EBG8VcDajK+DHI0oLOnNJNQKJZ2Fjs65cN2tuN
e4H5u9chpQ89a73+yAbsWj8so5oddVFjFEPBGzvd0grEOReYbLJUdXAPnqDNe2Xj
qEUm8Bw2lFhkS1dBf+g5dZOABjcO/EVyYogZwmMwn8/DcyD3lJJAJpeeGstQ2Rqy
H9e/nWW3CJOahH7ATnR3Nfr/0nEW1yoRGXkmnrPIwkx6w4DNYncsjsBKJhnWTMNh
ms5tIrjo5VwA/ONW1+5o9SJd0wumQr8pZ4jkooPwXqiLmrTspxOxPI0s2txUYEdw
Cbr92ysX5ErkhJNzOMVwnvGwt6BbX/2AT+sZU0HSyq80z67NuPDiYidLpwHIxa5i
Q7peCTmTuEe4d0pe4jW7BGOxlBmB2avN/fG1ozFk/rnNk21+K/W1VegTYCHHgj1P
oiNbO24LCqoPbTuIugsuCu94qu/T0xP7z0ZALu2lqIBQhk5rxO55J+x+dDap5ypM
jiou02+pEEZGDT4PS03WgjWPdMjuH+abJ4PKyYuA3SqEGoVQKgDXFYNf0CrgsHib
+QqgqCck2VDQVLV7t8fzAB9X4I6myVHrQA9JJvIuOEBpV49GfzdqpAc8yesoT5Ho
E1+KFirVDBElr6n4bq142KBtWsj/FlBd5XEW6r+DSIMr84EOB8VgplCjEFUsDxlZ
fphTVbDO/6dsEKu+ovWhDEpWMttorE8gpXJ1AkIQtgH3/2+9m+99sWXz1i1G14eu
HBpWLIANuMzdchjjpt1scfAWBV7jMmfJrlBdMAPWwSWQiibI7j9Yd+e+zH1EwFV5
ptpJ8uDnb9Me4b5jVkfcydbTjtnEVh26q492N8PaXny4qkpLELPcH3jCEEm4ZB7g
s86M2yh9g/54cH7EDFJP7AFpFceaKpkjSWTVsc5dKmujOCQJv9Rr2Crqp11zrhz5
Ff1E1/5mjl63wEaw7r9sxopmU18fDFvRf9j7eHvVRQGaIX2+c0RuWeFJdQ92eAyt
UHkTZ5xPtPUqBqon/vTctOYLIFSHDywLZ21odcYRPhVmVMry+TZGkVqipZDMmWVr
R+un22JLEVgM0kPVLT7lpqykjgZ6wmSJIt+rmMVaSay9FrXwvCKz/nsPNYBBAa+d
+WXoYrpORy5GqROE6aL9Rxk5NDaPMYsiUQDKCS3MupvlyPSSEzgS+XrTH7a7TpWY
3w3klhoyJkpUV3BFfNPkwyDbCB7APZ2mWnTjTkcs4RzAthQjLfKaXlV6sb2MH39v
iqAu6k4MWKawt41Rwje3VdpKHtCcvNVUz/hyjn8soKUnOqLVYS9QAVe4weoqnStB
nOlDPGk8HcJ0f2yUiSKgxqtFpb0Pc7qk0hHDhzJHK7Yh+g7Sn+SNLv/c6ilu3P3g
Levv5HqsUWxdujhaCAQZRbqhuplPLikqRQNN0cCR2ClO5Ee9sQDR3HBRCG7KMdrp
UojiwpFo8sSBJvLMd8LMP6R4DEZzemjqp0lLUX6k5RQeP4d50hBZLrLG8t1B7aXE
vBL/17LSvTMWZADE2azI35+xkHdPY5vT6c0Y24nYUTwNd4bAVl0eJ2Pq8o/buNNp
lJJW8HUon3ZD6vZ4oCsRutvP+fQGGstrNt+KG+PLJrkMBG3386fLMYE+3BtWYfV8
ABIPMxLP+4dV9d4yaMgjRkxohtzTpOsKUnOrJYhnE/kCYM8LgVIcw4iqek1jBs4M
Fs9yKNcGI9vLJUvwmEai4RicTAjLWkqhT4hPKAXaJDiE28sgJffB6+4eAyaIA0PI
HDM2wHO6O0x/jneHh/njMwTdpK8Bd0pWL2moAnFXRAMXSV3U40dJwFlJ5K/2C1oD
3lxZ//r/xeNZgCZ4C/jVMg++/c7/XME6e7lvQv1mlxhyecMOtR92E4AdIW9pIrEh
f0uN1pJEYsbOruu7/ogjM6KqZea7rDtc/n5kC5BCIeKvPh//2588uCAm5numMVfN
Mv0ZNJ1yZgRjRja23DYszLqd3zfvIz5nKPABhlZ8zlYzyBXG2FuRAJ7mh1ONj2V1
24nI1xwKRireBRKUvhKxaCVm39Hq2jp1ZOuZjATNV+pn4I0m090aytqmsd+Ui84t
ORBpr0i+voebFu4y7Fs05uyDo3OhRGIigt+/hrShK8M2/16qS5eVVwpq5m+TxMQT
jOtsVaORln/yfTrXLjMyWYnayRd4EtchQJcuGFMPYcPxh3jIxZYWuWen2WA/PApj
WoVOl2Q/5bFb8rXHJJb4FJyYNNF7Kfy9LfJk3npHLKZHsMSJtDHqwAnK6GXNeVcL
lpCt0p6Xohfs79gtn/O9Xf/Zg8PzMcwzEP6LjRKdiAsqAWnyTBdfjdl5CFNB/SjT
XwP9dKJAlKmml6QFMZtBmYeXLwP/Oo90eR2yjK9fAAmZhuPImkO7Up0B1Olt4RFm
Vndyp0orLBH61zNk50j5R2OR/9n0yKZr6YjvSJjns+bWIIJu3X9sn98u9vhHa267
X4wq+ePm2V3mws1zOq38N3W99vZE+Oz1u65x5vZCx9/Li+PUWbRrm28twH0EmzXq
j4wHX6C5tdvgTl0NGNFo0p+rN2NxrofS8VL6jcfrJhjoOUjmZ/4fwN8NhjSKwNmV
/2z6mvSgvF13YleGXLC4OZh95E/YCn9qxkNnk5Q4HctKfP3gOHb9sl8FsG9DGk7j
TZAfNJ+OfL6TOCLoy6GjcVCdf704w0q1xbSec1Sl4FCnCTS1mwWjqn4UhMwZyXSv
kmC2kfk6kE27vCMmAF5g7OWU5CZ2jFjbkH1AS4tNIfTDuai7j0F+UIu2Y6peUy5h
Fuk1EqmN5xG220+ZHCw9Cku6P/rwhn9TkeXTXsZjSvg0HE6PyN/P9c+ElfguoLjn
ZOMKJBujSWC54547QVxCIc31JZLQnv/EnU1fyWpdzUSyO3ku0zkWNV4qlzLp8vXA
ktPL4a4Nhj0oxa7IH74+eK+b2+TPcrj+seQ3mraykJ8Vm51DolnV4MRJlXlJ0caI
l6JJYzS8WsB3ZGdIHj8jFXzSNalal/664G0RVm+MkW5Nvm9Ssp6RcR0Ol8J4IDV5
gTdVGOgVghJnHCGoqKDgrh94Ce8ILmPHlXnQuUPYVYjEAWO6cOAJM1A+hfLjg5MP
gJJVcwNEIo2MHtF5rrGinVDczBdVpAUnPLzP+dD7819VOWWm0zZYjN/JOgoDCF8A
RVB9sn33sEAn9LRiGtoKdc/z3NGBbfMylaJWKjELMrTsHMe4mEog83eyDG5dcoTt
QqSD6WcRfUdJTXPCh56A4kpXq65fR5LMpVD/VLQpasuyp17I44K+46+bTxr+R2v3
0305dRBGH2Nx5X13n23dLLdj3n4+qM2KcnyLltwHbAfgpZC4SqRmTs5CBc0EYYP/
YV85f0i64vFTYbcIXc7k5P/6zimvPCqAsZj4yB1Xw1Z3walrA3YKupSzuFunOO65
HCzqqsOvl+UiySLiU1aq1RvCX612Q8XM/ZOKajkzQs/w/+/gf4vQyiftHSrWBIpj
vLkAJVFCjiaM8shE1J5WZZtKAJx/4XQ8TqR+JwuKV1fQnuGLsr+yNXF0jmNx07i+
I7IqYRGd5HM60DQ1/pBAETb97av8D6YCM6dqAa25OVXBvOLvKN2CZM45jvo4+m7R
VTxcjkMrtwZVnths7DOWb6L/3GREb8cZP201XTHnfI5e66iEgCQuJ8TRAooHAmC1
rMh2yWMiAA90XE9xTASPvv3xVeOIGldNT5qBMZnaUWeOCWMSyo6E4Osg8k27W9vu
TFehOq4RfrCORiad5kUHSD+hJD2hpzCUX64c7oAJEFHQTAF7cFeMEppJNk0jYFTn
LqcKY9OLC5lDXU5ZWq7pxcNz/YCxW8wfKOPyjsQJKn1dbSLQU6UH3PFaPpL2FoYO
vflZ5AuQN1+Yu6KfX1ccsT6MaN4YynZ9V4eqxPmjNYbYJLnF/GLo/BsTY796aNe1
fC6ckPWFauS67mEZFgh8L/Vc1mAKjekL3xvexEI9DHqPjoBRV3yyqw/8PKAL5YcB
t40GEQ86fgxEQyvSG36hfp7gCoZNHaWk1AjdKNWUSqgFa03Wv77ZlDLYwlOVFUuZ
+laOAiOnTnaOpQR3CupFWQfbhiHmJylzXuidU6foEjFHRq+UH1veJrRTCRHftI/2
5vh9CHkBii28+2TQ+Y87OzzPuCDsCzEhwU1cmkDHh4rJD+twzu7NnU8pnoitKxHT
/187aO82TrwtJkAcXjOElq73K0w09voi3zcd4nXcwu25j4OjUZbMqXqATWseZw6u
tYlrRoIOI9BNQawkHTbuGwKQQD1cMFwpo7SVvJOS0f+iuE6gz3hQTNewqJPoaYv/
NQqAc8bmFumbjKY0asMw7yyhXZHfJVlKOy1Dv7HaESF04rK5Ev3PtH8xo8rX5D6f
1FnbaqOAxvbJCnq1J6paUG3eoWLIT+j17UdyflglJzLO3khPuAgWFxRv2pPgwAwX
BdugAhYrtbLsjrpdifeDn+a3TfWLTsERQRH/AA57jI84iW+TrsZfKnUIj/Nj19UO
Jmz9nYm39IThQMnUSpEmLidQXfed65t5zIeaq92Si+MJ5AfTgtmsYpAyYHQhI7TE
4u7RcvmwnnevhFjF9XEVy0eudX87v0GjQ9wmiOzRSYy/Gwys90fBGRTyFK7dYMlS
unuueF1tp5OFgHdvBV64H/IXw3PRO7Uf0Q/n/adaiDti2Ludu5pNRn+QBhyJrT/i
YUsSYqjdqfB8pb9ioYPMNtr2UpquIm2B+HhATrML/ynEBQrkkvuOEKTs031hkb5u
liL3c7o+aYUfxYb7IhvOMRWYKV+n7DMXcvImibPRv2RiX3Q1CsVOorIqiss9OR9R
BRymbFiJoILd0JqDv5hrlP/6ydzEP0NmAZQTGarEU8z2W7BctDgxG2FI9sDpVzIH
gSeUKLg5+xpTdBTkh/4vfP5Dn3YB6xjqw93DPVIJg9vvZ1btUJIbZoqzjGU3Ee25
VBtWSX53p4tuhIcAo9ItcmtGAWQs3ZEj91Q7i1Gadvv4cuE1EeGUGi6F8d1qqtBp
+eGmaL9GSMUhlrM8dw1D7fDiFCwarEtzXxAHQPSVV4g6L8MBueOJf1qd7cvhcHAl
mpPzZtohmfj7rxIKJuS2qwe7yifqrIM0l6Ap7tsq0kBnRFqU911Ai1To+n55g0Kt
tqxwRCDRRqI8holmPzzIOMB3ZXR5rzHNQ6k/EZVI2A2SLsgRaJXPFJ50pNGWvF9q
G4hvQVM5Au455PhiAAOFPr1ZhrQwVt/pis28M28AXwJxcR9QLriOLnPAujy6LQjm
Ntqt5MQ4NSEiF3pRLfqKy90c2iKU8i9ouCBYFnal9D6zAtowPyJDQezzeYeo+D0X
gJ+1RoT8HTIJwMxCsQbo1DxnQOPU5ob8wWD4+aQSeGrRjEffFzWQVKqE1Yy/8o2G
HGU0dlT1uZU/0lOBXjQQiDLLDKX/dkF4ycYf9cfgCDLNKVLKAJZ8KowlfaVLyin/
R7t9UoaXzXLIHAPm9Aow+MWNgXQFVg1Ac57WmWl9CVJSf0JWBV0a/pEn1mSXIpiQ
GhvYEb3Vod0+s2pZ9CcL0zWZDeyex6J0INsL188uOEpSao+QA/uFQxyY3dlhm/TM
JIpaQcxE0FB5WhVuZFTgtCFns5fekFIkhBirc0mOTRnE2StdqJgaBC16q6qnW/vw
USGglJO+aff8cWQOLruXw4uMdVBBpzX+NTvLFcDIRfuZUzpvIQny77cDupgh2P+j
9akGbry+RUAIzA22ecH1nYYsoJhWbbDYY1clKu5Du0SnuvpIM3YnUG4WL/5mKxfb
iM2kUoUGDIdjeCfZSnjEUh/lduo2r7wEeez1n1RnOhQUTXpkSfVnCPOMvmnVN+zW
KDO6qgnPzSpRdfm/5h4Pinat4vCzOmFhPJj1m6xZpexHfvMvF7638OQEK+xF+yGY
KAlSNcpuUgriG+EQBT1z2QZaVBdhlpDuuVzsaxvWk8wIOZv/7ucTAsWTFd2BxRXC
UoKnjIKzMMICLZa7Q4S/ohPQvWTIQLLVoF3/TTo0cizO94F2d9q38bkHFYnSpnIG
u2fL+xsPMr3iucgb7bX5NQPsYgAVoXX8E93Hw7q1YGGwXoahJ5FQqUeCy2bgA6Fp
QGlunTAAqZGbGPynudJZXodxhsOhTTStISExYrI1s89vNcMESn5VSla47DHLx/aA
6j1Za7qHlVtPE38SbRLnWj8j2uGZEHviYRkeD4/x1CfaeF/hLeFs346hF6+l6Opx
Tp0oWDOeTsCLWn70HEOIs8U3EQVVAlaWdz4om1fVZqpBMcSi97MrLdMEP6n44mHD
FA9BBB1e1HqOHZf6GakadzagK4ellZKT1cYBUMNvmRtflUTgiEKr5RvTaILFjfEG
+JYASfcufi9iJrvx9bNzNRQ26DUkkFI582E0CnAPR9+eVgmKOTQVArkfSwmDek2n
PK5t4In6d9nVnrxEeP/vy3WF63EqJeopwf+4CQDZwKhHJbF+dK81r+hXE92u79cA
9p9Dvr05+TZ4ys9+R5Cp63gGmG7noBil0GkGeQRyWOLpZEjvx13+eALTRi0XZl4A
fe9ZC1UgZ2NMlonuAdBgjh+DRki9VMcx4F80/ixcDU848/QeVhqZ3CNsHBJDp+QJ
/w6ENHgK5QbF9k6v1J7yaB8piOXPamU4Tfcdfh4QvcsMFljp12PEJfw2NWyhuNQM
WXP50wfp8pLE3gake+Og65vNFgRu9nEPqRRb8qmx6g8irMI+obiauYlm7JCUrgsw
GZPR4Y3WgV/Hthrs2vHUoOQD6zesLd8G4Ih2tyJ5qtVAk70qBcV8MKinKF/50BMh
tJhT9g5DjsF4Zga3zm4VTn3MAemGa5i26ozQSNz1i7On/MNxGXQfQAg0gqrmTmbW
Oeq2xTQ8FqY86uRQ0KdfzEjp0Uy2TfJ2BkQRXGGJAI2Gbws/Q3Oingcd662M6rCm
MHyfhql5DMfNPIWtnYlemzQPWDGX2r1liozn5f/88wlBb1rUavuHIr6VBuF86ffw
KsYg8G/WNDrKBNce/O9Tg3gbBUY5QAvEQdwmeq8bpsKjHapp0fEL7AKwHg3zPaqa
u26DaALZe4t2VD0XaeCT0llL7hhf/hat2pF/mJePxK/HBDzr364ZqF1VL3GJi003
cZ+4lvuMG/KpMxZ9qm+BFp7vJ9nmPERnK6l9kPcIwh0LHNna3GY4rhqpT1ZLpAi6
S6ldrWrj596AdmJNSJpoOsfetMey3xFIvY7gt60uV8bKZr5TGF1RqybdTII3GKEi
CsWYnJaEe4skB9IiWH4mhf1X1kehPT101fJSmTntl/istIHtqGdz0DxCDckgs2sK
Z8CcJSMvBIkDseQNGlCSpe0vZ4QNfWEx4znbFZ/5AbRc//VchN5oGaEsVXSU+SNs
mOQep38Tkyd1jBYoTp0Utw/prVUCER5Nf6LavvlAJuiyqs5T+fDzI5l1wcynVpxU
EkifguCY0elh/gTzB7jyaZGxjiwEprIyIsUvRBXkbuS8j3RyoVOoIUECslrf+jwY
2n+/53ktd+X09MXQrYCa31zt7hIxTwpEYamrPzEGl8cANG4ki3tRFTnvW9Cl1kqq
Eu7dYpf0p5K+9v813FJpS05HjOs7QXIvfBb4XqXQXPPBg0YG7jCsNZQxstPOMuYz
ktQQ1bxGSGWcdMLf8EjZEu5rDfPabi8wb7Jta71FjQaLKUvelKwpLmhbm9P0lxi/
fEJRMFMZI8+vEeOorpLqHAqaMfipHadRTR8sijnYkxsAr78Jc9UThWFmOHJG4Z3m
z8F4vjFMWephYgrLCHnNCzzIDu2NJFiAjFfTe/rHiFxlTRehqWaw2BQGKWmqjOV6
7JKFcItXIYgs8qSi/Q/7GsKVMJgKsusGieH6EUDFHRj/r/TGKZW2eRMVn8BCFTyD
KNr+/d4RFAmn3vuIfLDSWfMeofVK3xvPZIDcUMtnpHzz++spRO3LYHTGnUM818L6
SdJfZIHJNAl2tJd6LwR1mjC2rpUC6LLzMoTE0K+rO0gGfSKaqA31egVX9SQbUfp7
UF9AC252NPKFuRvK7YFm06iA5tqDJOtaqdXzHLrU0xDe14eFldrCDWK/8oSDhFUe
w0BiLo5QD80vWdb/SANHjsZ7UXiA10kIeBtydfSkSXnHkxSDxJX7E/3vbUFkqhGc
oFMfPDg+WZF7WijyhKlYyT1tZDZJp/B3+VnA/sbMpYKJG6BzFyNhZ7GkhyJKZmAI
Uxsious5O3kVOZJX2HbkrTR4faStYQzvohPseem1bgIcHN5Fy27L2AZ3eowSVVSY
u7jkvq69hYCiErWHZGBgIpkZBh2DlcSbMHEZmPNNOWO9XXXIv6zhhInBEsoCwf5Q
KdzMMsHDV70sAzKBM9Tk5G3Aki06sQbXjPtvMQhAsgZMqsmr73zLYCO2jkODNZr4
Ur1svUm0tS3hKJV97AzN/XZW/+uUSWELFSu+7HSHDUNTRx7mjndXcWOooXBVpT8o
VxwPaBRg4IAANr86DELHO7Bbd0TMdeZ/djbnPCTGEGFMsyxfzXP15IDl+uQpvIYX
7+KmNKKYxOe7e9qRh45ncXTyKMzh8HTiu3ATG7hQlGqq70qcHGaWECDgpEISx4z1
3uxUkDLaclewFBiyU6jwbMEvkIDc/20rAIxGpdXhT4G1hW7UevgaBBt+OOmWwuAe
DGV+K6UNvoBQsUJvwsTrh+p0AM7bO8tG+9EbZs32mjnvis9nI+d2ltUplFmV/MNN
E4AoMig75NZ26vM2z/cfp2BSYAG7VLJ0olGriTbmAgx5DG1Ms0RJpSy5dw99oezS
U9ljdvIfgdvMkiPmz78S03gOWDWG6ArtGkm0C23OBrPUM/WZOdM4HyfmFqzQssfe
J0J9ajmXcxNYOlVPTEchpesAuOE+2Clod2dJdVAR3DUDD5rOeiHlSh1CQPSxFEBn
2viYsHquyC5xFEvYBQthwW4JmanUkgOYM0ynItWBN4A31grdAOlIQuFDqFWUdpTM
rwFfKHT3Q4sIS8isEVKh05SgQSuY54uyrDtv3mlCXpismXGCnwEOEeE2pDMuyGy+
UBXuw8gf+JPq1jMzWSZyJvx/2gPanraWYvpDj+uZH0WfwgTD23AwZCobpHtIi18K
vtkHabS1vaGWQoryy2l38+S47t/lOh/9Y39h0kzvxhdfN6Mq2bORrC0ZgJ8v0Ber
/ZORfyP/ygBxBZ0K3nhOXaFZ+JRhgi1bpxmk/hW/7wjTqDeYmjzejZl7tUNWAV+/
mN+TM8U5XizSk1r36JfC3ln75IIat/1yhR050nnyD4hPN3+0KORxeeLLzHuFo3Vy
4MOwLIxaZLEilqKuo0CRGF2OPaOeeLj6LMron/GtMbTaHG4WIHYRCPvDfpcvLBRL
LUZ7gZAWAHM258dKmAh7AfDj1lUHEntpHXXhJKXKX791ifjYDNFL01N+qzU0B8RP
qbbCSr2rc97hyd+M4xGSv2GJHyG9+cDr3tDRIefQFIctmdd0TXhCsm8IF+N/4n7K
hj0Oww/pPHj4bLLlLujfrWWkfnWI44DBwROEqnt6f2a7Lon5/XwYuuLyWEVp/zFj
8QaYFOTWN8kNJU5tZLZFHEyp4k/zy4m2wRMV+DbQMddF0S/N8fmr2rltdP6ckSrC
Xq03yN7Lcbw7uIWYndjrRd4cN4a0ffviMfeeduwHkQnrjUSt1AfUolwDph5yjSee
uhDlOYMuqGLWhi2/pD/9TKNVM0bGNuVceWXDAlBoHuWYOTcs6X8ZZzrcq3YwDO6e
kXe74Advkxqfxg1rt15EYj7tGl9+SgiN4/bQ240Qu6P0DBWPm9Cm55S/FhhgampV
IKRAQvEtjIIJvaEwyUedoGNcZ6BSASdVJ0ZRFycZqNV5YfaW8juaMsGAGZWg8UIX
AmWkJgqVoWzlAABqtqSYs204IzNkwzi9rdlK4qT1FwxxL7UPxE00klDJahuXnJc5
egzw+s8EeoK1jpBzj71Skz+MBfPEte4TZZWz6Wnq7RcEMhUEsTNa+qdqDLDp0/cJ
xB1go3InuBfRcXxUN99SaI1UI9jbkAUPUJ6u20wb90QUQsh2HyEUfwCr9vea+vBU
gZBola49/YM642UMu2yNQYQ8DlBlvnYVaiuZhE4qYS/I189UPCuAgxnUPitS1E1f
TOnVq+821yDL2hE4IWhHjyBUHZ2XT9HOEdTzokWkJRhbkcETxGV1e1bjZm3fdTtu
2LKGYPmNhAJ1rCDoqPgT+llAlylwZ3aioZz0/T7q5spgNJeYIN88fvtEulwhl+yT
HjFYVHaYAJttBYw/5dZcc8UMgq+v11gTKWu/KdG0Ba3H1bkoJvQc/rf4nDdPx0Qh
lV0X4X9hWDByYLwnfMl43SlEoH5fx4afQ9nMP56W4esQ9S0Uc7c4KMCVWQ3JAU14
8IWNCwIJagvADIiBhz0LBwP/9wqFVsCc63A62KcoUhbbM3CnmA1HAPlB6PaVLH5g
mZ72xiusOK+QohbdXRe9iRrodpWrbrU+ekf3ZBFqxTEXbEF1sl+8ynttDhaAItjb
Az6i6ovYAMUbdKcDQgXBvyBi+jDdBdQrXU9HV5g5kfqjNwqbod5puB1TmVSatpji
44l8+EBZrqzSx7WTOTn6JEfg/rBPdt4B2detugzk5rsa8gEz2yETvpbXtkiO0f/g
0FZruNsop+T0nSPGGf/yYMTbpnu9FGDwKPrmpNyZY+T1ozsGiRvTfrPjnyy7Ilut
6GzvOypRUH/fTPJoUyh1Nz9KF1s0n6GXfkBKSiG1Y9utjA9SaQgNkqvqpgzS88yf
2vZXFPEyxZaICQvcmWOGVyHXUEz36/C3dzIrR+Kp8mPXXbA/Ht70SfQJFg0QVfMF
cy83i75IV6fVKkwaMD/HneR9Hgjol0GTAY1b71cpCYcM6hhRaP7ORqEbITcuhPkE
i+WfhUN3j+pRFb+NYhuNxLTT7yIvgHv2HC4zrZ1xhoD3atvuw1TVus9dq3jnLCjv
Lc57DuSHfxr144ykYqP8pa3P99lppqbwn2g0v7Al4Zg6r6MqDP9anVSFqln/6s8o
zs7cC4B/h5+BYm93TsVdWH3sduuLHQAiyNoPO4DGBoh1YjJoOMkxu5uYCuBkmbup
Y9zyvSFmOEMKqEhcILj0KuOFoEsuYXhWJ+1KprZ5BSd7ErUVW7B3sBDV2Gmml9e4
Th2627ed4tOLtZx9n2yT3VvuknpivhDmxXATca7vNbiIvSPzIQ+8AW5bixW3CHcl
1RndFfi86WjzGP8ohSPrcxdindPz4ySbJmJxrARDdbB1HwBUgllA+hPDrJ5+uc1n
jYWtUQE3xrun6r0MSMOZFznIcDRqPSk4CjoIlmGWvXPQCDjU6k2LYe/7/c6g2+HD
9Jxqc7pI+w2AE0TqaOXV6k0fzvzo82NKtNgkipHDWl/wjcCIDQ2zNfm830Hl110Z
Yv9BlVSbph71289ctQYkd4Xjs0U3jjOBDI8RqpMZWDnOdMRsGklltiWUyFjLSt3L
mVE6wuYWZNiMzPJK9Fza/bdN8iresEBx6q3X8gCuL5RhGqTaSEHVl+/ReSJZoTAM
PL+G+qlEKB6GWKujuzorheEngTqexJg8PpoVV3f9SI65tV7jhqQIQ+zlRIGac1rl
EmXPMa9qX4ZCfqSDS75UdCgl5n9EUY4chCFPBYQQB1xvyZ6uEVC0NnBiRpkhfk9A
xQQU+x+hXDORRKnLLQiSKq61SBiPPRSLS9/KLYRz1P1bbY/2x0TSa1oZzBNEFWJN
h3NMeLI9QMbSBKcsSOEYliqunfualn3qfuAwadjC3LhSU8mVIm45OuUuentIfGov
Yl5/O6hNgvKkJRQk/trKZEXDM9IC8qlwDV9mB6s7mpoEbVJSfZdNEWDzTf4k0dam
9zFsHC7aSXQpjGGbFnZ4w0IuURp1qn6nhG+pSUFXAJWTnYYj/mcznPFhOAmGw7ik
Kh0Vj3qLePY1M9p8DlT9RXlpY0S+qtJeERHUgB9j6ww1HUQobXiauci5L8oTOvDV
AQd5HlZxiwh9cslnJrO3YxKn2LqaeNhlSHljK/hrXfJgJRljyfnU51yc4SzBZ+fT
aLf1hORy2gFoGgzCpRzQagRP13Cv243ORFiHbUScuLkTdgG2PQm6d9pikxAeEfVF
PGmm6f+7gfW3acHBZlNESVvwH1ueZ+i05IX0QCwCPsbIshVejVd5lK8lI04uLLFL
bThyFC3EiAkyT+4aMXo9KTy3hxeaRr+99lSdZqEtkaI6yenfktU8lHWpgmaESBz0
IwOLkxNfCwgRB57D8Zuif+EA+1x/PRnTlTuFNe9RhPz0fIVUnBv5S4svBPr9+Ail
zj9J9OrHEFeF+yOk3YlHkcVLThU8wGL1mg5Nj85JdFy9P/dCy//XqJKXYQgXVkHJ
pyM7JimCCqC711SC9ivEeVCsRE9b+5m2C4zO5UswlPKyvlPnmuxOYSebV9piZboU
XXEraz6jbFEcGaPLLgVMnTqta61BESGdktIHhtL7cCQnSDrFPYoe0I90X4e99OBK
IC2aZFYvYsefeIH8fqIuSfiaw6jI8BvJjdYEa6Dc0EnlGj6yjv50BUOb4jAXJwEZ
iLPxvCDwk4gyopYcwXsepm4IyIa5mklA8j0gMhj8GTh4fkqCiS2p6mCg2BEVaBfr
77qTks9k/RQpvDeuJoSxr177slK6ot1VhGkvXEwa95SIv2vhmtvxGHLOB8AgJnBr
noMvmv6m30MvBPQ6o3QeCyMyPjyEHszBc4Bzt6PcKgSOHJmQJfQbI9aDd6bwZNf0
rLKSLodC9f0QgAGOupsoz3o3QgWJ9WKCE/KRjd8fdqvdUBC1VXY17D7vCm53i6By
uu50GFQsA6hxgADrYAMX7gBlrdsPcwCxLET+bJ0SAnMOUiTC+PREtH5+Bf9jzfYq
/LUl8uMEC1HN2Wpup4eoYX/rh2vF2c42ydNHDnzX5ft7IvzlglivqsXFHnkburZC
tyUeDvV2cpaiw9hG7A/oybNG18FjRCo3+54yx9+eiiWV1z3XWE2dMQ6SsKw/gg5A
9ARSF3UScT/776bywNNjAM2JhVe7dimDvOKb9S2itJoDYsPXw8dit/gFZ0IkSexk
vs6ZuWXcPkmH6w6F9qJv0ZPu+nqh2bLgxHQKzgWNmCPghCqaan1b9F0mKDMKGm3O
KL1G66IbZWWtumgFuE4LikBx31nL5eeo3PUjar1ofqYQ2YUGjZrVAHSEyAep7S6z
PWXdb6GpoZVbZiF3t7vYyFBYbBRAkonnzCp1io0PzCDNiaU1hskQaVoo4KntFbDg
lYSo2sXiYWhayHr673vorPterzR9hR+30DzX4QUQeJxe9PYAG5FjlO2mMJ2s7fSA
lM3mSj1FAMdTJadv1OfLauWdYoavasY/TRQRxK3gPx3raoatqzKUdTcd89UIJPIH
ob1hVO4taMnz23HsCg7o82YJ2JkcS5f/R047jJj3vl0vuBm+NrBBYPWMVUcEZIDI
qgWDtPoujJjsGbEt5RTeyFXp7zVP2/qfj9IV+HyzAT1WiZwIf986RRDKFps5oSZk
1KuNxiLLB0eqyumu7huehRd9Zr5TYYkED4E65fytvOLpR117qfNDdYBwn2Shyuea
Op/ABE965LhXM85MEDPX7NB6dAIC4Vfqu+HM+fFcLlYnRL7n6r9LqvVqsUUzwnNz
es3k5Nfzu5PPlJ5pbrL+mDB03//80utbN7XuUTPAdAbciuik9Mazmpq8/CnVb2gM
gDSi1KrWc0gfZzDzWb7N1VEDGQkERhrdCqlGnVjNZVDd72CpWRUDH3eLgf6gBZUw
DY5zRIzMJaD78ryv7Z9GRLT6Em6vPeouzL15Dqb+aKjfhEU3TdFpP1jrihL1vDku
Htn33woO6lkbeukbTQDPje4JhKavAYGxIPqwHhLc2JxFvj2A6AwS7NbgupAHfi0w
+lqN4D1/FCBfyAKUBiUU8lMU/kTiqXRRxizVzNqdJwlijGpwQ9BpZrfdAkBfi5UU
qd1jyDQ1O1UtjHNfQpvXJJsddj130ajEhQB/U4r6PsFcOJLBtTMECbycFaU+MQAx
jMaa/xUCbS2AtguzE4vkQ71H8umBOuF8HNLwp2VeVkSU2e058fhAtWZwpiXNmrtH
vPQBwt4SHudR8zHV/gLwXNuTtmMbmtSBvCO6MrzPdyvWjiOTvkYwfr1gsKcQ7TKt
WojNesCsssGCyGnYizPF3Lcv0JE2uTE+5L9nAAezBzTIB53WLxmmhCzJ93KUrddh
MEliYIMIGrwruUVdxz7isLq+OoACkY2TNwc2A8s0Mt3UJHaOxkz45p5harb7ScSY
YIrtNvA+foFVObZP0FjlaIuKXcvBktwWMFxOmTL7jLtJnNrT7UcHmEppVkNmQsDd
PPPQEt377Fs4iF5HTXvsmJEBsdA5DRc8OoOgeodTxw1ypqmiylBohBgfFvSOsDVJ
/dM88Mi+dCbgdpo5L2wABhBrsgEPcPS596vvj6db4zOQtpoUmS/Engnnrt8MpSxA
Tpk9UoT0I5NfZCigeNFLM6pZIS8M9Gb53SguOYjqc3LpSOjty1NkcXeIuS90qXb2
+r1IattsUFG/Y0LYy9I4EYxOqSLwPDKAjLnt99vi/27cw1ho29Ek2+y9IxGi2FEb
VpRyQhDNFt1Ri9AJADNW9N37UYw3B6eRqIcictg3gjBzGmgHHa4oIhAGYFg7LRjd
qG0fEtUtfcboQXwQx9S2GFWqIvf+l1Q3+o7nDJdYgZM5h9w2DNLgMfW91xvciiuR
hvWzdXzRGtoJwnZ7D38lv9SO6YnCxaB1cUC/6qxfVubEvfUa6jqb0DlxtE2zw2cx
5rYyXCw4wrbmEbVcIzbfDfqdQpF0ZhzAcaERvL/T/pTDEY9ZPWbuZf/Pz10G3QFp
lQvD0U+g5pPrw7HpH0+sB6OTimChdQ2z4gtw/e20obUwxeZU5UHMgZyH3zdTlu6P
PvOXfwq8vK+MAyNmB/FHA6Rim+Ar6QhKjdcGz6byWIByTI/roEQYT9RsV2mx1j0y
o5xWHQwdz9UP9Mt8HZEi/hzIjcuVA2GhESdy+e/q2mWxVlUI9H/XaM+15S53H+xy
U7/zrIPAN+xZbotAMzCKYeb4iDRs81xvhUdL5Ff5nSIKF4cI77DHQoLyezAN+H7b
irsRTsSX5gOKtKBO2A3p/0fb2j3fKB3XRnIjxR0hjYxQwDX7lGVn22JkcNbbvqU0
5D6u6uy367/pLaoVwo18MO9Xs5TBFURIZYtmIwt+KxSupaiF68Z17CR4BCPhzq1F
NupfbZpKBgQoAHOYNXx1MwcD1dlL19ogVUuxsCtVzXGXApv6f6QUBFdhP/6zHZGz
K8tG4JbNmhACobMuPrABVVFUbQu44s8aALX2JssIe2phjsnLfxi+QuPdUrUPHrC5
l+DI+xX7PEEXGjY4CizvuBPqFdWl6gnY2xwk5Pw3FKbiYQeW9OYXvCsLLtHVX29B
2pqkwjsx9C0//Yz36s2CYMGHHbiglc0fgOLz8KhExBhSy3zK3SHzz+THRifn3YmI
cvqRzNGyL1pyo3T3hzuwuOhY9rbqk0JLvYTAM0HbvsTa4Oqudyn1pQuRtQlGAGvC
OjrhoSkCoAHXpHuWVXC1aSGKU1yKB6H5+9Q/j5zYBJaoFqptrB+zQbOp0CGveslq
1PJQE5kwB6GD9pnkouXizEdDn/sbkC9EyTEUPBc+O43CIPweuUiKawqwf3E5EnR1
6vJH3Sm3szlSsPFM3g50ckY5joXz8P4xGZp9Qr1W2oWgl5nLFFmVoff41w5SxQDd
MZ+qjLyLp/I9vMJbYDN25KGHW/KIO0H2wZ95s/rcAPv/TTZHOLDHxU85rFaoUBwR
3G4UwUlzkzcOrfmzlmnIjoq01hRxofnJO4gk8QOpTdgYBoNTYplEK43Hh+lJ7hFg
0w4eA+aVjekPIqJrpox64AqFFtcDu4oACe8Bw4dwZhRB7Blfb40VSyO+/Tc/K3/u
jIWIR9qURZ0PqLkAZ4AZgQTGM6IX5O0c3krw3yt3BVz/1qY8wA+XFFfVN8U2TEFh
9SvR4bpSD6imlt0DQ7In9ZumO2+NLujo0sMHClAbsejnYg8Q7ah+WMh6q2NLff2f
1nPU+FH14sJws/WT1CaL2vknAXLQCJGgBxNdug+TBL5nE1X12pj5AeRjanruvipN
tk5p1hVZPFHz4ZlhPZUgVN72uiVvj9KV9A+6e/hYUlprPsXiN6TAqlDpxBA0PRzA
jT9iTehzSRldDg3bRx9J1vV8Y2lzFU82dWNes1W81GExkPN0ZoPD0lYK2TWlwCLr
/B0uN+koi+X3CiUBJspxIrnRIuOfTFYJsEnf2eUGFJCVIQk/MlLaZ0xhA0OH/5p4
FjDghYkCJ9m4pVCnlT3MTT0KHwoQB9vSa3WVVR6Zt3qKzWjGiv4jxB61JEql3HFp
ZgjvjHoX0jwxLe8es+3VL6CfuOynU5QJia85wHY0ZAmEoVKU0kDoQ2zkpYMaLDPy
kU9O5j5gnzH1fD9PEBni3+w3xEPgSK+RXeCdXBTQSZ2tv/C4JoMwG8p4DSiOSqwu
uSq+IJ/5gZc8EYgcaDD38kokNKUYCtWegbvzmYvyIXN1Iet8BbcmRTtcVryztN4f
/YpzZNYDQDYm5JSWXxqT/PF99g8dUCDtrBMRXDJg9Maer2XQQMiEJfQolHFh87GS
wd8e58JXrjXPdBtcRSS864M+t6tGVAqcH4MbVtDbKQwbQM4E6mCoraRjDQg0M0R+
UqivVroXk7t2uSrdtgb4VYlIFYao1BCnifTk5LbTuseTXAcGiPazRIJjyZ1PtqT2
D7k31XziLUxzILom2DzO0LlSOq4ZbBTLQAuNSxLDIkX5zcK6Sif48f7Z0XnbLxOT
E5Wz00n+TaKcBoXRjMvhnfZ4ntlBf1B8LAwBDUXuORxo/Ng5ANu6ctm+IAr9DZ74
8M8nqP5BfbVr3Xtl3AwRGmznAs1/MH7t7jvSGGUV84RZmUN0aKJQ6SY5tJHadfsI
Wdf5O44DCUDZfx2OQRYyM/PNy+r2KOMqqieSjtyZ8QSN9wqwFpXIWj7Vb9wWOHb9
tShrdNVPXFxehBzwnAczxyaAqp9n1V124EsIL78cFOC7vtqheo0lwnddOmHpt+bm
NENy+W5TIIuMYqg/6lmzngmYDdJmQDHnnY1K81CegKeASGlaQCYqyab25Bxe6FXq
HHoujsD4AlOwacXyjEcOd3c1KuOYoF1zxtMRh+r6KIVnY713Aq/JKIW/ss0TorJq
+9mahvGH903XmY4JwWRotYo6gqVjHOA1zLOuFPKttG3rrfTOuG2VTjfutQnm54ha
yzQkeinqReMACJObYFtbweErAE5WxiDZMEFeGadbDw7iBPDsN4M4J1QciL7VNjtg
LxiOQYh6dCvu1N0bmZI3vYksZYuvWEiJK72laSiIaDfV9fERI+WO4SKmren00pXM
taSrZb2zRpCbhlQ2piiUQ1GVRLUMqQylih1oJRat4YAX59c93/WWt7QIFmJDescg
T5kjANVJwuXDAI2DTBnLsRxTja+MIqFmB4FY6WH0wu9Vly3I/DLiYZXX+Hlhr3V1
m3SdyhjXioLhiNQBu87h897aTGjiUrWG9lGOvp412FTuV8lAu2p6zozZtFgWSlQh
cAMpvtrr8RWKfGzs2otDAxv3S2p9rQnrBodec0aCkhAkq3PwZdrE/6ZTQJSNxtpL
n6iRM5y+QOc7gM1FElwTBK0+uuHaKi9K4wzKc1q3kzG2x9WyfzSMmfCM8lt3Smn+
HN69YWpEZSsvuwCWUhb6NLi3aljVKDhK8reb9LYXAVjKqx3DT+MASgHaexSnzl+s
ecQpmBetYVkRipL7KXstOABNYa7fcokFzS21Fv1I3JB24WUNygM5dHYiirjHjHqg
icYZv603FLdK524IiVPQ+XmpXjLi9yECqkXEoX1OUtBJ/XySMs3mmEgHRAc/fWt+
nm3ANVsB+Svv+f62TULcucyHR1flXuU3WR/lvJMsCi5bcc4KzLEv3mX/ZSlGC76T
21s+UPZDcxrN5H3Bx22UIccuv+yaxgpLaOksNSzECFXEDPvGcup78IpriEzihYKr
XVZKfEOm6M+IpaCGOswWAjUkCip0M7JtWrTlJPgw7m8tnAMVcW7eMDXoB6OwsKR7
uAbPYv0dH/rmResEX9dJcaB1aF/wTQwZZNfeKh6ELH0a7oebrymRCteS3m2/Gou0
N60uMrPzEbo4V40tP3biZsPF7YUBSiWFhySXwWuX486+3jvS3MNNhUnkV0cKMXAV
bV0NrbdnYP2qYHzpYbrl0P/v0b/r+rIaZ5TE8IFJWTQjrw8zLRtAFuxlgS0/Mqe/
uNWWcpP9H4eS/d/zn5hvqK5AvN6AUuFUmv38rBZLDx9O67LF3J57z0Hsm7A7YqjW
ILfC/6bty184iIS03THca3gUAxqvPIv/fqDsVHex3nqGPwf/OOj+MR/gY4YlFtR6
OEE7rmgpoZ+70hqC0ym3rIy6DdoBpyh3kB5VCIIUGLBOsGf4iSyH5WwDT3W8D3jg
l3G1ig/z0EXA1P8OrqsH/UFimHWLxANFm3XkuqDewGj0vNxmfV6wqsj9JFLfj7Im
9pagapytFVW1vhd7UrOIEL4truFT64BjOlEoei5WYFGl2z89OHbFUE3jChfq2ud1
aswFdEK9COWWhq3T5HQ6p0E9RkW+Qm39KvPCtF10QDTCpFnjvzB7e+Oi64ej2AuE
+P+zihBZFAOma8K27CtQZbmOFzIsrI2apZWXEA0m6gt6S0UdsZCaqw+Wie3oqPyR
jL91Z072ox+iHYBZfSVlHNL4877dMXpUoDv+V0Q6hpuFe73AyPnhkuND7er7WqPW
Y1HWWTUdEs9NoNqR+8kjf58K+e8917aifb6gx1npEfj1Q7hCHwjjWkbKJoH6EvLR
xqUUeZ7YwLhMawfgflZ4I0pSTbTyroasotCKWXCVI89cUwTCB0cBBL9ih4yzKXf4
WbAGo2TljtUbJCPLOdFaFAOfgzPceVExkP97z/2mX3CaYD4pAmzmgYkdR0neetgf
ev34knwskytXgtt/EfBXW1ek0H1tyMq1REQFv9WZ4toTdLCaAmrbTrRj9U6vSfcQ
WiDv9wyYjdGdzvRHI4Zxy68+yQntgHW6o5CXxKDRhAXHiPZ34sD05MuOm6WCKBct
17IKnknXgRCni5tVJMCajFuYPcW9nMJ6urY30lbd43Hyjd92+9PwovGM5ZF3TVMx
Vv45mgpZsYLQ7a+G/bb+6oyoRR8hhK23ZneAgZHLf1MCIvYY9fuJ6mVjdDt/8omg
vEs1mC6pX74pFBqmYhJr203bsLFadYxtN8X3u5906JPY/xF6GY/J43UkrxRhWNhZ
SiJPGWUmB+m/kaJSaxYbqEXnx/46biKa4e66yTJKRQ0YDI62yX67r2a6KrKFgXdL
Hz10S37iLS3biW2vFyJ8Wuo17pwY+JWDZwXNjFgwe69djkckSvr0YzCI+hPi/VJq
LavoHDa3fWJ+apN1NcHwr6PZ5oDDVLKUYiL9jduyTlJUwgN/nyfG8lOeldlDSJoq
SN0yxzXPPnjD1hQ5QqZUc/8dCUe/xTdqJy8zu+sXjMRZnBxkEox5kqG/9BMhWQ4J
bnsNdV6U4rseRX7A1gvAM46TMYK5D/ZR/JcaXAw7ieROec0WxfhkOLE4V7ecC9k+
H/MAn4Tm2qsTDobs53bJYjtm+gT7xX5yztfYrmxaNqh3Vm01fhwmgtE79qnC5z+t
eMlMhILyhfQCtXMzT5ISdUef/Rax4r1WMS9g3GjXr2tpDT+u8MxSTsIc6omR89Sn
Wld3g7Oark/espl8T3vLH9/7Xd0fqDebHuym5U/SGF3MCY/IgsM+Bk/EOCOvSFGL
ht8MNiqrlYSB/6UZpLtvXjnF1StAG6Yxg97tRUQJ4lwL4WSbKwUsZbUbuQ3AMBEn
LnbeNYjm/kp85VHr4QcPzwRj7s1ZZRrwsQIbGnzFYNnxWn3/8GAn1kAFxMGqzZn6
h2xPWZSk18fC6cnamwN9P66SKy7H4C3MReFQhq+Vm5ePv3e+xDsm06SlndNdRmJu
fGfIrAzuShfsvUOWMjptt6oG3GlS51PxmKGkjkZ/O58MrRFDKEMrLq91GPOT6rMg
sEyk3fxZlyg8G5BvKqO0OWzy1QMul/sZYKRB/LgcY0KXINtCpTK8jfW+424xPRA8
50VEilgYueYa2/zEKxMO64/l6lONU4VzmjARfkvP2wMlf6YGdsx7ix/VkRHABrmE
1pB4P3eoDh3/mS941Fp8lOxa1FMUjOCJd/np1XCcTzBphyY54Q7DL73zyM0t0VJq
F89/IFxc1rav2IEE2rGdm26/0fLrd4VVzcDDlIOEMxCiBapbDW4xxRp2Is1m2Ge9
BOLz6kKeI3+J0nwFQcFyJEKZVt9NWMgCtsguIwYyqRSS2IkSWoQ1mSX26mgqbCwM
diAjxcxde84H2tnRa8LFCzUmY7piYIuw80xUayNY/fEGC2i1qpq5jzcG3mrnb5EB
nnFA1afGCQztZzbHRzVFGAvU4X8eiUqRuYcMfOplhKSTnfxDmX6Ngo6kE8pUcheu
OkhNjhZaGCbmjPR57t9rfPPyb0mnnplXWftLBRR+zApdThc0vWG/GqnmxbWeG42d
zGWHRLGS/DuuiYxh1j0CPIGNBVPVhITJLEZRHKMsz+CFdxIMPbfOoJPQ66bBEdhU
GLZCzn43hhlo37IL2t1b0BxBg8Yl5MKui18hDxLrYU0c1b/HPMhaJuTnxqeRkMDG
c0XBvXvcB4Q5Rq0UuxsNnt3ugjYhwrQaO2rwZqlGfxto+1FRBQbtvFIpgrxy9I00
z71qXwPy+vGygVsTv3phcBjtgQHzfqbBXPHwjdJqNsgonipb8BgE7Ftngdhd47X8
k8/UjpflfPLBrHr98TE0g1WemGbUqwnwO7duARM/c12tap+1OlilBFrKMCE2EBDg
tiF0UTQxSNPdzIQKvgiyA4R08aX0i63+pdsLh2fgVVAtFBbNs8Wudflfh87c2Gjg
IWzSB1QqWIfdRwDqzkh36tJYibT9Tj3oFI0z0YrEXXhrkCnmHYzpPm2gCQ1vCZ2X
BNQm8s05v91AVEs3+ntTfa+J8fcw4wJmW/bbEjrTL8goaxEw0aW8VyfeIMDD3tWH
zmNrHYyAj0ACEq4tXrW/6iYDwABhFsGCb+W4BKx+MqTc+BAsB0bNUHY315jgYdy0
qh/4ieqSv8y4RTGduoREh0x2QgtqOq2XLKDYTZ9vQrdI1YmCd976RCDb+Cnmv518
8udhAebWzidrc3gpWU2uUpGC458HiNHzgaLRUDQ063zwgPV30HceYIBNBUTi8Z4e
yY78vB1zPDTDKhQWVm+kNfKhVNcXoial64hGcH42HB+HrXHdOIdmoir/ppftSmOy
6oqAklXhJ99LPMhbUxzMEknDFw4sHfJ4HIyy1uRxHqHZOJO8JKabVGpiAhzA3Q/G
xDPDS57QJSv2R9ZHGj646FBPeJBVeE34Skn8mdUsgi8Wkf12ATnJA2J7mdYXJcw+
9AFaxMJA0RYR0jjAiWrpDLv5XIPKqlmkh2XYQQajQMuWiUHpBUI+IHGOuOosZXbE
hOjBTUj5N5Y2qcDmL9sfo4uA7nYEl1pi1OOLYaV7fxuqf3pMl1C5IVTZjpY4ha0d
2VcjOpAkeDo2yR4Q7jGvooQV7TmZ87TUK9AKX+PAzOfc94deZN+p1zlujykbRSM2
UXwYJRId8ZE/kTviUyFzwDWNqqXliPf4yq6cgnaTmWR2lmnJmwq1G2s59Sqat4AJ
RLXHt2BMMHpxUEzeOHlwPWPtte//gdTwt2OmNBbZDCeG/8PCPXh4E+jv9iJvU+bn
ivhNh2uc3+PgUloKjy6fSf7fvjcqA4sRj9afLEDx/0Cxhd0ZJZqUMQWrj50mxHBN
FD44mHrYeY8NHOeY/3AwoHz4QE9X71nKPW9+6olvkifmoO0bWm2LkkTmnuTGwOjM
f1Ob4Me1iLTUsfdOX0B46vjF9ChqZTrF2bULtfrF+9lWQYdtI/Kje1Cl6NNyVRnI
tAG99OLAPKHdnjQnN+/CKJJyupwtQbTOmQJ7UcSUFN2ZieLEPtm6WnYAiu2Cmcqo
/mg+id5XtBClPNe3OKQ40GQQU0vxnOTqaZIH7OVvBQy02evVaea8Nh7FpMdkOrbJ
hG1pYEm2q85l4hdqblJ1uF+sVOhcViIXLjR94nNapTmlpd7TGlrltlN0SCKcfQou
KHDxDsvdKS/T/2v9m78BKSoF9ArPp8T5yDdHHi+dNyAA5erem6yUPh5mXqNbnlqG
prmlveoj+GssTOn/uMqG+5i2HMbYXZInaJCvea2uyokOvj5c6+fK2PX7vNVL//je
5qFNRLGHSSv5LOg0eCX/+yFxvj8FLKX7xCU2P65Xi6nT74MWmfawFr4VSeFbL67y
O7MKBPjo0fTLlo7YkJTAfFZUmOx2seCAqFQ5vY/5FNs9/mByklkYUfvvLAcNDP/T
7172JCUe02h3Oh6/tM7P7a1u3BrwGbRnxrA5iORjCd59/P0dNp4V5vquHygxyr8L
YRPbEdnL3m0Qyc0CnzO4tD9KTbEglUQ6xZjlbcTU26IpePOJetiOUCZVcqfysSUi
hgkO2jwF2/QXC90eEllhtmt8jQPxtFxxaxdD9QsqFiHu+8jEZRhWlOEMWkryZM3c
b4u5wBjwoyzL9vLukSHUP0mwabCwuQjY34Bt0VYoRF3WMYgv2+80qm7JQo+kiZwT
Nh2xfRxkrpbF6cTxxNFIAMjz/xU4Nxjo1LPdwPCbInNjr4g2/vvbnP0UPrnas8B4
rwklJWFRb04QtbFCy1QZ2dy3F7osMrE+pYr1/k8hOnHVAo0HfP0VsLFS8kBnZInp
ZvYPUAK/9wdpiyPqXohzR4fgD66NE+gEYYECN8RkA5cebxVY1dnvyzQVwFSJKD1+
YO1CUNWdecldzd2qY+hQsK37/baVGdyAjAP0UaJQweKg7xQZ3CpCvibC2eloztnf
oe7YxxKx75N1QX5q/zpZ/gc/yYi4t2bAS0vZNrfYIBE1fLwL8oDmW/O2CbL/jzx0
lzopV6i1Ssdt9pxOMDdufCcZNaq9rVkeiasHRDhsTRhRgl17uWnJ3szSBCWdJEpX
uwW6FY6HqFkE4PVnNya1GqeQftYIunDGmOSCkHimLjjtMscalr9NjQIo5za116dZ
43sA7MAON0KXaT92pb4RNEWlIhOlybxoYw0rjCbH8KONYLJo0ybaYz57ZqvCHYsW
mQoUklVRsztEynsyKLq2luz059Q5nOCprQYw0fnTQpyu93EhXqhePbAggtVHa1au
vh099itjrtBd3zh4iUCmenlHifspzVPc/d/OQXHmI+Hv842O3vr2TGDUd5H6ZITk
4Lu6g1s2b2QANUa4C3PYCRjizbhhReJ74SywShzdlCthi/DlcnH7emZXdqwaRu63
jnN/ujyfG3+TCPY8CX1w0umNRy+FyRjgm6eTAwY4prVX0RcptJlXcuNzf7q4ojgo
qcJuOzQ/86+1jfSqgL97IITx74pfKQ+pJp4xReCw5K7p92vhVWm1Aq4nWUyPoPjZ
RrsXB+VGqTik5V0TcxPums+4sHALzqFb9q82lpBgzUt9OQbh94xTabAPbgyjw2Na
P4rwpvElZUmdhQqArZSIJ7xbUhCraz42Nmk9Rgp/hL9HwCft0oM66L5b/3/yTbW9
6mSR5QYh/0G6COyRtP1TAZcZKkaCfJC8KOdae5AUJX9MrUmxeqB3eE7EfuqQTldl
TcKsBsqFmK7qhfE2Gls++zkMRqD9/esNy8/JTAUxMA80OS4ds/a1BPoAZJt8mD5i
M5Vp/i9MCYo8khm71QEDVgy4VikNV0Icb7qMAXuHxlNUukfb6VYLSXDh2vR7/zgz
mTZPXy3+fNBEiN9lKwgIxhV7GwFH+U3rfQ7Z+vTIp+zN0J9Yf2+daTL8Fg5GA3tr
m8LfujJ7OV1xNlDKXI2m1m8BIvpemg3W4GNwjHtbjHEML3YgVzJtwoLfojvisyEB
DKLnTdCTOxzg0F86AqrGMoIl1s5NgyyTG4urGecBcng23XAMoBKJ5ZEXSJW7rdOJ
AfhAsopTtP/t4FVQinp4X7gJ3ETxYtSeS/ng8QZGjaTV3K4i3wRYxSjPjRSuSpDX
1u7c+qvgGy8iOltCc05mYSLhon4+IcqngZe0iUULV4JX8UTILWW2bzAxsXUBsfn5
4ZzL/+7LzGIU2Sh+UxbJTVIRPzPrFMY79hXYujOgjguWJpIC9ccVTKWpY2pjx7c5
p/yvoB1jUA2UcCP7hyUxxxHtUYeuCYCcSh6dmOvH73Dii/sy04nwAab2gNvfazT2
yCNOu3CIy9M7ss0nxwnMBAAJ7v4ZB1lCWRS/Th8BSAh6VUSHM6Ng3xNNsUJzaJy+
WDAmG14vd4KdSwzmivpBFODJcqowFfmXAEuETd3yDALKgRV9j+tXrG8BDBxz8tIt
+GSRuOXH3uaekUkcH3G83LuDY/LAMkfcwRLX/Z1T+i2g2faBDtWYJafM7zlush1d
/FTinev6Q6JpTtBfX41h0hduHL9NqaJtbCMd9Sl8+OCWQuAWKSYFYFMrPTZpBSkT
yIMMMACgrxPFGhYM+yOrRr1HLAfzwpMnSD+XZZRxNkM2i1iNtunEJMIbz9qNXrzO
DWVbvzYgJzUy8/Rd0pQFgVfBN2ALDQ4J/HOAp3VFdJiSwcVZz4YECfU+YgmBJYgd
GtjmIzMxj9SXwd9WFRfqMUllOJAGE1ADEkWqHZe1bMeIKfrnSefbtGNdnOnSIlvL
rtqrgn6Wh3nytPyJXuI6U8vb240DapMf2BEm7egJ7KxKntP4rT2Ix6H6NyBWp1jl
FujPAj06cXFb30NjdWQD0KDJ6uqdA2YQSx+1tV9M9voZSk9pDNE0x4Mtt4YowKBD
q4VYEuPInxGjGza0N8o4KHU9MVqW19uuyIVd9ZAu4svQhhxI5Yt1vQPPrdqnQ70G
a+kBlxo+gjFMYlL65vTPUzEerfQGSsQI7iGEfWE23H5Lqd2qlnfDYR8KK3ERgo/Z
poLKKMMoh5N9oyUrbNglYvhRWl8qFcVivZpx1rdSCDZSKD7MKKRQBkQ5WkoYbDky
Hk4/RyI1wshlfY45lqal+K4sigsxhL7zKny5CeHe6Q9Vt9d3/g7vvPDskMoAwnWB
ec7YCoDO5QwoduodArdL9lW0Bxc8Nk5h+0vzX1KQ3uD1dbN9v6Vr/Q98dKsmuFbV
2xfahrOzZG7kH4p9JUmWV1aL5rcFk/3VgOWht38tpyIaO/ZvA+/LlX6Fv4iKGBDw
RUh0sti37PLobntpwrhmqeL4Zs7UY04n3erFeraIJzvFn+cbfg67NLBX9S7rn8YA
Siy8k5T/x7Ae2E306ht3SBfQEjhAIUZOUro4slLjAyufVIYndVcXqVOdf3AZrAMy
AUuTzbRcn+/8AgpgGhjJWM1A9KiAIem5neJP8+VX0MFPwIkzgKLbOl5h3MlnXuOq
M+915t2eLxxMADjAAR5rGHWRTojDFGA6wuRFyLUNM2kYR6qbNtzHqIM6wYlhIxGt
LceLXbu/LAFgfF8q4XGKcTq5+hhAc9x4wyPsbDATP0+SjmZbL8LMyDRGAid47sYq
0RhE+A4Lk5XEE7DdCdOJYPs+LgbChI5V2mWaSgRIxxW66Njk6ez/ENSYsDh1Ra8N
c/bDnbNtHuEkgvcQ9AWAzSHYmQgCFJE3w7Gy5wl/xl+/kFySQVmw6/dKXBEumXs0
P8xol0F/81QYuwKSU/LjyB3Ymvc3F1leNVP3VkjHlZeoul0XYoek7tbbSR4ZlBgf
IVXYDwFpMVFr7hhf2vkN8BkDAntHPWI7b6jYh9TTeMplOhdmhNsD13ZuIck5DKoP
h614JETde+XwnJPULQL81zERzqK8Wh+K28KgAEtArGFxhJot/y1UDD3jb2DXfl+F
krpNe7d4u0XK2cFURdw1kbrVVSajvFdgZjGK6BWozEdUghrggTZcnE53ryXWXIlu
3pM5MJG7RtCEO7JhnWBp3dhH3unHBIbgn/lLzvSfewiE5EuwDIU7dRabQUs3ahdz
jMbxp05Rxmc+LZK3N9oLUxftAySu80XCCGboMyXwTuimGppwHYg1pxnitDEaepvZ
3kvwziP59UlHw+YemP4T1vaVn7ItQKTM+EDG62VELmr8M/2IIPHCPKlE6nrwvEC1
oWNkO4qUxWesGUa3FcPQ0uKxWgoNFdIGlgaWnV8CDjpNXdMAWrZL7rGiVpSfF3xE
1KMVIb3cyGR4eLsFYYM27U8zj/dchEtQ4O51ilPkNgQs4DDqWlwuHAb/C0pNELjE
TN3rYNvQdoVM0a9o2v0MIAn35HX6BIiH+W9RYk/egCB3KA8BLCqpbVW3lZ6JLjGl
7+pZ53XRuhLxkPjElIZO43tiK1ulMfbxEuRqqu3BoWxBjlI11yoxZNxL1dZu8a5O
AmsbxAyqzUQH8EZzFAZnTcdgiWMfroaYKbuT49QjvlEZI+pJqLZSBAwzlbHtsCUj
czsGZgCN63h7bwnsMM81ROIRoDverSb7RPh1hwdX9dHPrLtUp5PuXt70JmtrVhu8
ducAY51Kts9tx29N4srMATu4ub5/i54dW64b31/GIZIBmaPs/fFUr7wNImsL4A3N
3eGvZPKKZroWHlxIOFWWfSq4SupjzETCdwgWKlZnIN/G+/lsolmXOMDKq3cTRXdz
+LDuhkaClveZjJORoI2XrKwge47d2jtmrlU8FBPs3igEi/Wua0hevBd+bw7CpShp
5zIvq8PG+Bnfc18ToBif/7/JcopqdKPVDugZQqIWcpcKLo89FWGPZtRnM/nQ68lI
NujDpLLyagN/sJN9pTj6j+C1II969qW3f9VqA+IaCv2PipOt6x7YTyNkaWglJpxi
LpXsrSLdySFZ5dsVdeFUv3Qbz/SLF9l5RhPElCsY4lPIMTFrFdxFX3CR0D/tSDgm
QDcy17ELUO2UUKO9gwx3SnzguOJWT58n4ni+6xuFgDjr3OrkqdgSOUILdClr1qUh
BQpaVX966QakZtzslTXm3/SYl2IF0L4ndpEDy7xasW3Xa+UjGbqPj8jvCIWp1/3u
j7zI6Vl/yWq7tQfLWJEegji9vg2b4YTBbhdIelQXZEvgXi0WqyPs0wb8+qLOTY6c
uJKP7ZUAU8L0mp5PmdwnWB6GZ38yVlbazaMENyZMx47PlV++32BzJ7XWlA3YMwmw
h0+r6pXDxj6QD6e3Ze+1X1bK2RHqyCSQVAvTuJb5BQxoZA/TVPEMmZwotqbMPmbf
qBVHPzwsrnkmSVVnLSFhprUy2TB6b8xqsI624I+wjl7rtoJUBnpKJtcMO0WFLaeg
SqGd57wA8zYt3Ehuq0Wx4QngQadA3KPdGZfFilF/nhsSUVCb9ddHxmv3bHoqbbRF
U6OiAxtPw1Hiqnyl8qArUexW8IMvZj9OhFZhaGZLPWUHI6gS+T9sTqp7U0lOoqFQ
4PocADveuAwdxoYt/qt2mcS6Q94gzrKdCTROAgHty7RiZ5g8UsoTgFsxhdosSASc
RgfgRZZAIieRc5QjnVUGCe1SvOBHp1IlcsaLKWZXNtR0D2TCfu96o77DFBxGjfPj
OYPQ9m5TDp0MAOhibxjlyvr+0NkWWNFQw2oXq+Z1evTibqysVZXPcuvL+7u8OLsq
FfiRzFtXJbu7OP/Cbst9Bkt9/Rnc1nwk4S7VCPjduWRhy3j2nHkFvO8znVub7rx3
PLHvt24ZEnFMuZmthFSb5hqO/I+I2hR8SCTJ6xwcWhJZsu9ELqKCgjpLhhbhPluI
UUBoD7Is3ESNZqItKZfoX59pWVDjgB2mhk0iJFiBdCRPJGQvk5shwsi5OPVRU1+w
raU4DacgWXC0fvuj6WHxJCgvDcgk2Ei+Twz64cdw9GgAQ1/KgrFPskCbLE71jHcJ
tmFvZ9w/mmwcTDX5TqgWcmhAq9pCbzP6VqPGMMaeSz2fAbwXFWw89H6A748WzZ0Y
jaXsL20N12F0iKGRvw2mD/mynyjVeEold15DXMH77xGT26pHYHA1abvu6Bvj21Ue
Z6GQuIL5xph26pgcrT28DPy9B/eNUnusLD1wQNpkJnVjqLgCg906RVvFKu8dnfOU
WMsKupzgve1Kjt0tNmU4t1SH2ukJNmY2s7PTyCvNA2oP2QBnVBHUtyTXdm7KVvL3
wQhp3LeVC6wdogWvQMgJduGdmY99cQEQJ3zDzXNgbit0MeByh25Vsw4/6o4h6QOV
Jz6Vh+paSZP0cJ+uqv3+jtexVyEsEyOykd+BXvTqA6pwmdmj8O/F8ctrziWYvzKE
g5h+3J4H+yeB8mVDYXHW4HwJcBQDFJc3McuRyDx9Kkz5ztayQbw/IFwLxjyVJN/v
wBTygDqO69jLeGVt9s2/Jup58/Thg5Wi16Jj3QwuK9Byt9b4CMnUD1OIS4qEnUkr
OUMdgOdDjlsOagO92WxogkUmC2VWgC17JLjzM3hAQpXa2sNUBmylmYiinbaEU5mu
y4JnkhMK/bWje6QP18ZdK73M29yVD4h0GLh3cXYx554icNuivuoVBY9lqqVBHVtT
OnRj9QtxYKUPxSezD6FO8X/+dL5+JF7lUZNsMUvO8Bzt2De6SOnlhfEj9XlJWdki
7PW2+KhX9Jk8rgRhSAMGfc4/LQwGEei0jBOpwTO5SG6DKckS8leJlki6L7a9g6Jn
aUF9pd2HQWnnp7aMkGgpwPomVJymXj4aP8zvGXdMI1qA/pz4/c0yVLv7KUMcaUOB
s9IRBVekS79GcerKeXsEw3kZK3OMn8S6cbG2QcM9x0cIpWG64EZTIvdYM9FDQ9vN
ikjrJ/ZkzSD3vR4oCA1RDsnFNZVSufGL3UhBbZuX0A7zcKYKgXMd0KtuXwcnZMcs
p8Ox5BbtK0kfkl0UINN1Evxz/pUUlanS0NK/pGyL64Foa/9ucijT/elyNIInprKI
XtvTcvnNa/7S3+hon/YIzq6tzIanG56hEBY6mEMtK31TtgDaVaAhsPVFpbpVSNTT
otPbgwpNU1PQYVc/uNtW+q8VzXQ3sX1ufp6HZY1lgwpP2ADOk+5uw0VEtfH7W47y
dt3038BOKSvPPrqDrM/0yDwaIt1XQdf9LQ8LS/p7YIQID0JLpdnj83PF7tnuOiEK
jIk77IscLwqae0pJKNYGyD8nziVroUCbUL72+ZBoGXJnYgw/CzKIU5dOuhMyPVKk
B/xm1bmSntWNUijfhX2FL0R787nsKIh2i7LHTOo6CJ56QTzLeyrvXz5N7WLj4L43
BrEu1y55U8tnFgw/e9heXkE+9nzUVsLDNAHmZ4efTT0GjzF+1wO+3acLgQ8MtaIT
gtlrvo8cdlJaI+cmioCHYj5QQ3hlxryibfti3u41kFR28g/CeG0TP8w7mMf4TLVy
iC/4om3Fla76yChZfpVqo4sX9gggMQdaGO2X1+octOQuTkxrtTqvBe9YWm3ztO8X
HrDk4xNNlKDfR9Qa5jsr4E5D5Qn5cyDUZoG8134TYEbjpWj0Lwb//mcLfiFHRAi9
kzVO/qhlaYHeU2vPs90q6DMyQjNvnpOSxrx7Xc3ptlqN2yaQQCUhDkR0bLm7U+UD
1Ovn7omk3oKq4GSVhKuAgRi6HMBWr/yhFrwUSbTxpwxIOXe5wrsWaVjy7HBhYXvX
9LbzWi0Ld+RI5I4S1ThvACGokMLZ5Kph7YCRW8ltFvFzhMQlo920QRixFL5FOMxR
5LUvaj8jDfEIO0vytSumQu7R8d8uwQHxmGSNNWcMt7ofiqIhw30YvZmym5HZ7hDM
FbYgQQ2Vwyfc47xsr9GjB2JqV9AlOJHodVGJWaqEZ9RlLbnbV7scHZqiseXPnvnI
Kmr2eF9H0oj2fihY576e/MsAN25DFKR4zwg8tpKHnhdwFmn6Dtbsvnjg7Swt+dd3
01DqJi2Iva0g0u9YZfPQwCstCufVulHew853XxkBrT+K4MDrTrEzzSsjWWe9eAly
Htt2Cfwvu7osr54X3oheTZXFrWDEfthz/xZnXxaElDlpBTxiX9M0Na5Xb+GdFb1c
3X6a8XfzsJSrKybkvdUBECPvk+U3d5D6K4pMWm8oRee/uXy0oRWCZ3pUDzP5+I+D
LPHTIGR43dDDHpVd9M+8if5j/tK3OwGgsDvoXXX0JRhbo7YsjXGwmOAMOueAQTzD
hYDm4IbrVLW+1Cd8SGrPaw9zk+Q/4xqWZz6zp1EtulIZyhaQwfotKsm+YFxJW9mF
wcUqbsssrLb7aTsLGPADYNmIrueN2gPHuDoT1CNbwGUHqUnqfnoLSRuXvac55aM4
vgnww9FWT1nsvoa/H0LPSphWi7wMUS7AE3DF+LdsPqsJMbQjeiJoHdIKdjo6KOBy
dvk6CrBJmoLsSuxhx9ExzdWldLy+9bYCJBTKhaWVmjc6FvzdcBTgxEF7xRWWj1DF
8WwsxMlSmJFdauzRaWi/nyLRinwhNPGJRWVu/HgRc2eW44vlX+6A3yOHmECfFx5h
VLcw/G+fPyQd5CO0SXgJ0vtCtmfqDJaztG4D1dIPh9+pw5rHgukD83QVylB0va4I
VdnShOIt6wg53+zwe3DW3KpiwnbuM3q3j85sS+pcXIe+Ervs3vAdIIIxFOUWcLMU
2HJQhyZk5ozEWdEmIITW4ywZrkoa/3zx5HLqIudXvgMnHwe7NRcXlvN6nVwB4PuQ
unqrPogUsZhy2k0dx34avYABvXBB+/Uh3kIs4HNrBOT0nZ7mzMI7F3NkAhLc0Mrc
rqEfPeiNA5PZ2hJZgbZzhk9DqHNcfm8h3GbSSEo5YUn+ODwcSnSq3O/pL6WSeX1L
U5blVpRm+kSjtfBcIXrvcKjO6YKz3mxMC3bwmmSq50jf0X/Xiqf1NFytsu/spzyW
ORFQDdFpfCj7yR7dZIVdTvlOsBfJ8QBabNHDtLEgC3dIvn8qEHrfTL9i2I3EKyLi
wYh9+9BNXSZipyPVQNRtrjUgUx/rStsS1BafsUxPXbkSjgW6TDLYOUQZL3N6vqVM
wbWlncHbsgh9wDusBsBT8u7OEvgdjSvcEXGLbPIQ49XbcBhQmcvkpFPRWBP0dpAY
ZY8EWHSErmBWL4bDt2xbipY2U8swfD3Mgr2VzWV9nbnZuFklK8ReK2KIVmTRyVxr
Zvhj9YuO50AF5TRyk1I8bRu6MW84Z0T/F18EiLgtmv6msca/HG8Jv8MIuCRsz2FT
UTuK5RTvu08Kh3rdaiz3aFge/Fp047dJyaYBHWiE6dJE71kJi2L5Ge3NFyhWHJ89
bVT+fkoGDhYyE4WCYkVCJiQz3co6Y+C/y5ZPZk5qK4cHHom8vbTEUnut7mZjF5Nx
9TaWLfYAElqNGycLxKz5T5/u4GTZsZSwrcfAOHTbhzhR3yowTmMptPuQEit9+d8t
iP3qO3+HPgM31N4fyinGyKWxVH/t7pZZ5PG4JEY+c6/tL0JR5kG2NC9r53qEL+Vb
/R9JIMXx/BIx25TW0Xh2uoX5D7Ez5TGGf+3AN/F3PJinn2MQIwDV+MlYAgQvmYxK
bDeOh5ilL+8h8TgJMP0MtrRTphAoWafmjg1moptmBW1hbHXmzLx88wX08uARWKih
3OwgXpKaCJ05JCGpHng4DY6ogETpFHaRFKkGEeXHmb75gaNfByuEU4MKt3PGTCwu
dc+KJq95idlocyPKbY9ERncuDCfpUgVbKhxUzRBkwJmPhuYFwIQ9QIXelwdsor6k
8+YhXTkdN/dr3aO8sDk91Am5KEkUWBOo8+fvS4ZASaZSSbpprzGgOizWY7JfwHVm
Rg9tVDfMMoapL20fGJTzUK091E97jtsgsKXRnRgkI9q88fKzF2VSJcciKBbMhi3m
sALZYebmtNwqaQjwn3K16hhCzsvXmiu0zfeOPBppRzWEO4WytzzSotUljVOaxzL5
yY5NNTjEx/9rgg7Tpa/h4z6o5e0a2GK2txLmUNqT58YbgqljqlGo+hob4r25SOny
0Psbi2flFoiK3jlRVgD5HmrgnjMYdjaulXJH8iUJg9p3Acln0gbqhkgv/OU67CD8
9rKSSBCIUjaxGjaPC/fPQ+ZETQOl1cgkhEOs92TQRgz/3oy6WFNOan7XvOL8qRk1
YUURDhZrD993RJ55mUsN4PHAn+kqxOkzrkjvRpEVbou58sHWLcbRa8hkMZipdF7b
tvsCoT4PbCeOHBrWAYb/+BjrKZ0juq7X/HMGBIg00MqTDypT3J0PPNeM569cmtnh
6SNMNmXzsr+vm0Ws5GYiyG40nSOJ1Um3PvxLGdLvc1qNikUBwVbraVxd+vUwQdhM
WxWPlOvSq/bfrexocfIzgr2g/AntI3o+fBwDmazzk5PrJs0PS1+wjfnOBNWeYvcs
NuwW0kZ+2G1mM/iMMYvYZBrmJsfXmWuopZ8HJOl6Rmxv1q/VzIyD0RtiYRgywc7k
Lio8sLIu+JN8vRudTgU3pyaa3YIBQ2rZ1mNjjm5gSH1ev0PR8+ZlPHwMr/krddiV
r060GGnk2JlnIetUrBIir+AWpa/YEgyfULDBGUb9HAeiNg3gXel7SDDZADYS9MX2
GeIVBFh7s4CjJgvYeSKAvrV7uOaMjG2u2bchCPtE9fMiLXR9TJCQHnU89N0buSuU
9vzHsviocmb6IMRgJz2s2dcho1ik9RY9cpHJayMDuyq9bt0x6ufd8PdZQwUdsSbL
pmFOPtKFPrd6EQCNE9v6yyEUk1EEG9gwu6K05cnDM7smyRXB33JEiPDzSdtB8wZh
6NyKW9jTkj4qNkSYJtExO982gc5FoHeg0ZhAX+vBxB/lp8Okofbr+qw2UqV+hgou
PoN67excMvIxXdahLKzB2ZcoFLwIkzcPxJ0p9r+uF0QGvzGp7FyFkftrzQfmeavc
qRthrhD27u9ePIDGr2/1UiQz4J9QdRtl81dsLzUMTDx+tX0luuJBt9enD6mACnik
1B4X36HR9sXoV1qaWZI0V+4fO84E2v5jLF6RkT3d/phXNJ3Z3b2EDjWWKdZGvILp
9zzs+GW1dyMblyySe3aYYEe4xkcBLAKqndKrx70vZqXAlzo599D58OtJ2U5aujcM
E6Pgw+sJk0rZ5aLAn955vj07ILq6whuWQz+bmSsT8+n/vlvUqwrb5SII6vlQgmxQ
4Lqz4NyJx6enScVcMT0AvkYmRHJvHEbFKyLjK3sw99vyxymGDDNYnb1hg988DZ17
ZVwPzsUbY40W0KYzd5GuHVU3w/vKtKl1FO+0j+x8eLkzKBm6W3UeiHE5ukbQN+2+
nWELVVRCK4c3+zmtkn5xzvlqEjJCjPgRs6UQIZQG2tZgr2y749LOjDJ778wtLICf
0VboLzUUcWSEJCNSfOHW/oKBH5ziBiP737yhy+g6dpXA7LsxYjYKNyC9tlHiT19n
y9aoA8Kx3GeRN+F/UZHM6+HX6I87gZR6pcnUhLDbIGxyecvkmUBs14foIaEOSjrv
HayTZ3pKhFn4HmZq+CXpCGaQEdZwnhtRj+H2P8gEwPphBW8ktWfnRGdtLD5Ghz9O
X2BKO+VmZApz7FaQ9XqVIS67kbTX8mMAQPRgcB8WGdh0xl8kmZRm5kgb4S4nK4Pq
Mw5g9f/DyuF2TJ/22EqneSNGYVg9tpgjE9H3OSB/wQdH5fE/8WGxCRfE7IABiADj
VPIRDohAGPyrBHZr6HH1neZJKYi7dmPm8I8SZMy3xXhfLyBTz/jIhCDQDoGPCbK4
r0OWMLNtVLofYXp6HGEoqY8YYpUp1gro7lI05xEf+KsW7ncBDZ1IMYHmjW5iex6a
QbdbhPBHdrEITAQI1MeCtqipZbfOu9jJ5A49vPjxRIf7j7CmMx09jsFUxQYfxt0M
dPulPjQ0mJ0Q2OKKsBvXu3XEpeacV7mmwCIapoJeXuGPONuP0kmeZ6PYNO3VQA/w
tc5MFBeCg40+NzFD6cVlSeJiPqyq2iVSny+DkY3ShTOmIxa7q/8OdlQpCobinD41
TnnFPBPHpoYrgeE0XTGRcLRlF9xqxla/JbR/8YAV570Sn8vjYc9kQjpAIntSYxZ2
lktfmm3dRV4rXMZvXXUoHbNwLZADZOXfEDmtxYSWCW2be4OPBqOu80MaKT+GSS98
bQoOKB/4W1BgQRvE4KbmSUHsOTzH0r8iAxm6K0wrh4t/bwxIY4TZ9Dh47TbEdbPA
34LPUdJyLzI8dNLeWIN5UwtOF9jgyklAEBRI3APYQ8T4GG/AfJ6D1IVYPD/CkMIU
tRhw25hic07tt1mxS0SaOQdHSNjNsCH9ayuk96H/+fgdhq4sRrH8RJ599mrIDd1C
9bpgCcz4V7bGYY3sstI5fs5qHs6tI+kBNiDvl3V6DkCUjy8LRqjRpsVIicKor/7c
4BKmSmrKv+zkcL526X5lOlost80KqXnaNiy+kBJdit7ZdN7ibsWY1kt7l2MhgcJo
Bz38IZHhEmUpkSfqF9wBPzRg1VfGuaG/b1tfScEPReWfTJOt+ddGUrBx5lEqqDsS
Fhd7oPJ4hpe/u2DwZmu2nkiyl3hkLmLf/9C94Bf8Rt1evBpXibfkQTlf2wABme5T
rIAQe14wnKNdCcNV5GczNgIQOX7A40Y0QZ/Zd6NOMlzPeZ64NjnYK7rx2rDEmaY0
DI5SyRojWs5ogRPBY1umwLkrgdGhzGCJeuO9QOhjVNxyMiV5dH2J3I71aZLJ8Kdh
VflB5iQ4qQ2qUqlbBjTQVaPW6V8i5WgT6fVqcmFIOdUl0LDhT3FKRpfsmTB7CBgt
u7mO8AGIr98slqR/NWp7Fo5WWsHk13p5uEFuaMCqRdqNf6EIFz4xPpZGsGXPhl/A
BzN34E7YWwNIr5Aih9In7LZDXsVUmZJLC6aTRdxxQNKWG7GtDF6/CSemO6vBV9xx
hyrJeWEK5zIwtZXJLHHPDYFNk7HZ2kT9zNVzF0kFxBL3knp/SzU+oFm7ipVawRHU
xaSd5rE5+6K+AGBlTxNh+KkmGYycLXfqGweS6ZcKRUDJlqt9u9pLApXPnwM2cDEo
xQmgNFc9+JZ18oOAS2uh4LF4OSDYkC8Bz2DHPMoVijvg2J1q9T6cgCkbNuebITi7
uDOTCJ1HaydOT99EYCzvg5kqi4H44jTyJ1AIEroasovU/AMLEKbSoEF/iiwF5C5q
lrXFsWsBYoL44cJ9tFuxvhD3g8uPADaHQr/MXNi8dvZMHJ+T1JZoJAxIL7b2PzjP
b+bAFo7q+Ko01xoGBkCO9LgQ6tUMJo4mFsTXaP3GNiwhkY6Tw+EZOtYMfFvvaty2
wLuUeSyjXbn697I3cRaNTtODRI6J500vXpiUO5gFAp5citEqW6Y/xBiwAEApYw/V
RhAzY118d76Aq+3lYh1dmmIzdtqWYSDNbJgVuLd+tFG9neDpkSN3EFpBbliLAF2c
Ej3V8NX4nodHWx5TpESUEpJPUEtFtECJVDL0WwfFF5R+VvIBcDyy0678lokGVE3X
+dXBxUvxb+Mt6RNxRc5TwL5IhK+2WWQBCveMgrChm73SHEeClEvQp+lIZGogdQLW
eywgF3DOF3WzyLok2Fo2mTAhxikE69+ttnA1ZhsVTkbkPDSW34CZkTb0M+CeT/4h
X6R7nVko09j7XTEuMPtGVzT3TFHXbBvSY3SZppHsJbwi6DrHiamMGhyEN3Yp15cB
BpkyjocGJFjgLUKpl4ooMNWroxxTIDhQcWY9EepF0MHYN8wqhK7GrHR9oWmdIgKh
KcPn0aPHhbDr9++ZOq+1+L54yOw2TIDuJ221CvxiqsHGj1M38ERD9dhcvmigHxh8
EL4H5xI6nmP0IwuEzsB4zb0ZvizucYkbnOQTv4dXhBXJ7dICir0XngQ9OzFTx9JY
ivUBeuQ6rNwRiA0o1m41j2Nc5H+ERzw2oxCJ5NCbmsLhEFn4o39ZX7Ugdf2gH3yS
fykNnHjVTuhg5/CScUPEFoIDhDXtTOGMFJpamUPiuxeMHZAPGe/4DNKaHwV4Y+BD
nJmmkd2b0c4/mKu2pjxFe6ZaRC9bU3XONPDgIG7TZJMUIfd7MHBq2o0pyZ0oioRr
LkfCrXMG4+mkbWI4tqCJm6fQnVS66iHAUYLcYkNGiRRYNO0gqsyqSb9NbPkyyTh9
4HHIkHChnNuYX/SSjX+Jf28+9CEp2EQObbfZ51qLQqnk/FJ5yKvKTzoJ/F6WDTtI
lucQPnzLGeQjrTelDTBudkzXjPqAH7yXMX7b3VH4XUpDFhMwZ7LPWKxLTHJc6rkJ
OLy2V6qbP+nRTYftbAYRnPcppzij5om++kQ9QIk+IFVp2VSD8QI+aPxbiRnVZsVh
J103wI7wZX/sqx+FYvq9UrxE9okEVT31tKohQRROiO6sgh3bnPcGX0AHE3aFDZbZ
mlsEBHoBPn3dYljm6l37VuMf+ijYh1WM24cpXej6ktlXdcpXNPZ0EYoneM7szYaF
B2pApSSoFXRkwuH4waEU4a6Lq+yusa6/l3g5Y7mcxXJqtrnmn0IN+t2y5uJMgG74
Utxmfevvgq6IPqjyFlDtXgQrgxxKbp7gdKBsR0wpnQ9/D4n88IFFnANzHaO4VkEQ
hFtfjAShnHll/zVu7zhEcTrcJWP3TTEQHGZIWX22JbkuWH99liXzE9FBWHr+aKvJ
4bqXG3rbhZ7FLIAZEJQPm+sIWLxLIAxxBgCK0+XXyJxyttRDzB2HanRywc9ikzMf
2199/o7/+JxBs6mYkJqFvJGJRn9y5fNObUzCgdL9cZ78DZOceN1KftYSt0XSbUvv
TbjaJBCN/SRT389HSi2t703J6YuYX75WAdhrLytHjNAxQ9MrKIvz55ddLHLUpLD8
nv7TU4N1/iQCOe9/mCiLnajMY9ozkhocn4zt5ONOZez7DkwE35YY1taZ0UJoxwI7
QYU0WHOKN8TOMfksnrSR3+qZi1aTuj/108ntloQPSTluvW27PO/GfI+n0JDbjuV+
hS5RyrWLFqbXC5mnN05sQc825nFm1jCBBOITcn+AyKe3d8B8nfQawo8lV6oYnRC7
1GzoNobHOmMqKdNv64VsXUbjWid3Zju4stEVIpuM8XCB2zKL4R1nBqYaLwfY3AIw
Jtvw+XPtxUiEYoB5LO9xnmTfqibbiTw4SftjCG+B8iA1MvLgRFaDafL6nJ6ajQu9
QgoubeuxCXjnw2h2ak2o6iLSZru930s2V3hU9e0rKjYNTiXaglBXNfiA3ods4Zt4
UQwEAZxGYB4zjhzc1R70k63H17JQnynMQEiCVbJsmj756D63HZsAy8Sfx3lq3gh8
x+YxUWoGMWCQ5SZrecMLt0y/8HJwxedSBFOVNxS4K/TnHsUipZlZXVWRWVg3zJUj
2GJrJ5bZM4rh9Jg06ilY9kBeuZD7LxMdGYq/LDRAJ00ccOTXbA8T4gbnK9rfeSzl
pgFmFdbu2mAOVVkrUegJL/6RO5qj6pwLXnhHzgI9K31tzj5kXvgB2pw6OR3kF5rY
Tro6RQcH8I4Z/DdD/BLepfUGULguJ65tV96E/FPhgHXGGePL4AC0uD/mxA8n7A0V
G0eTSqf+YTyq/o55FOkkfkbk+/gNoBQh6ypTXjYZxRqOTdzZU3uNYPP/4+65IK8j
TzAfFXM5OOE9tds5XO0f4faVGKYgpwt2OyXhV5jI499s3Hut6IVN1mbUwK8XQKMj
Hip5yYLA7zxY6PwXxNTXiKz4/9LPz7I9VPe2aPmtQTzuSxJz7nK2oDS37uuOjS5f
p0hZQObwn4gVSKTHdlVwonccpj5QVWLGrFqXrtYMKQqFhG5G+L227/vTSiCGmU40
ue/52Xb7LKypNb73JU0EdMGqkuYJO2th6dszm2w2nfG8JnN77fv9PRmYl+JXKeYP
wtMxassaYiwdZLebFonxBOO/FVN8o4yuL7QCms1QUdlvBbhRuB/hNm8clVShoMfT
TVPCdVWz/ezlkT2z6cxu66tiZvs6gTbi9fmt76HBamSowkLFXYaVK1d5+gkqOdJM
xzJLkv2ym3R39UW23dxi4fYgYe4wgEmRizIVcjN9IOovd/xPX5Q9T5MUxjptHxoB
wYaw5ttTOZ9J8BXQLDCm8d3F48otDXTSyu3AQp4DbOOp6JGhOeiQ5BRMwxj8bkmi
GMNgANEFMprPzazFHaTAb6al79pAkjC/nzufLIQdTAzk0aC7BIdlGzNOvFuPcv+g
MB1M3dNvozoiBA9GJxNSO0GoegaL8bJUdnf1XeeXlXw6EtqYSERjWYzK5+ESB8n2
BBEVXRZgdj7mUpzUuXwZpWGl8eTXH2jWgdp4G4gEoXMd+CgP+KFB5criitwCeBxs
xj6fuwAGjJYfD6XLlUFNgGiuwUe6TnB1ojHH71KKP1E8nfozxqNpjbeWHG++O51z
z2ToNzxpm7Nba7BxCYXF6J0WWw85WFNJHcCuCPUm1ZXWI3lQrGk656eLPeofO9zt
NzdBSEc2LIDTA/i2SPc+80Z2CncFMIEdluDA8dJ236YBsiiQC36yO0ds7FloUCMJ
6HVkR6XBP/zDSim2sRnmBjIiobBasQcZ+HA2PSBIUE5ekfxX5ZkEYEhVALpVvJ+N
VDY3HchV/RfrqTavoekwE+v02mfIOKgDvcM3DJ6HtgAf0Si4pBO8Vq9WZ/qfA81A
nJYiWbmlhhGS5j+3bY4KPxJREU8/WUXdGObf9/wNJ8qvD7XyfVft8KUCECVfdUe8
jZeKgQWE3ZbCMLDEl6taRlq81t7J3r9gZJOd01gWI1Nhm47CQGqvOfpccssEbg90
TjqguEfg1at9dp/HIL8Lij2rCQ4kPPpRyqRWFJh9ZUIiCYxCrCHegbW6rD8t2FAw
iVwki1brsFnLpcCZRKyNznbPa7pt5mLyykUy3bI9FdkwyAxws60XIJwLv7T1k/iD
H9f5XF4Tn0cbyKrYsjp1PNM8cr5WhrQETgNeArie1SjFzzEVdDvo4xGJAI/XrgCV
X40/NLNYab6N4Riwvvz1FllpQVQ4WHvsUSf8lU1M/NovcQiGf36u34os06KPVABw
TS7gq8OmaQfYnyZTyWy9mIQzb6vgX8zY1b35KpaWDI4Fv0CNN2ZOTPDAO0XdrN/A
MOLk//LCjwXg2gf28swNjY1j9lNP8Xv73HfCseBZZq9faXboVsStST3breBM5+AU
80VTVSAQQdNV1bo5yMNsrqkD2Grvp2EDdF4fajMDFN/BLQyE9F7qnM9BH9kcMB9a
5NZK0+KaYJy1heG1YFvJRmu9YR3OS9xCU/3fV+GKiNqjrJcjumhpDL2pS23fduDZ
RSuBHcZi/WB1FDecIkSBE7fWB34M8e/k/r4dR4whYp2eIgjYM6pn8cW4uRRLQCLN
SxOPZnQEez0uZDpe694W9qUtTKkhtfrMmYyhS3tJRrtXvgKQcGeY3GSEE/kzPDkR
Sn6N78J15UNY9Lse3LOA4RHMZ09sOY7K3QkSTTGI9HQ/YeQ6ZGVEI+9cNf0wOe2+
uh2EquXk4mmwtmhynXx6ySEB0JR4l9QA4WRbxEwoc9onJtHOVEyedfd2bpRnWysH
gmopbFYEuNL4aOIaRzfsVn4zxHQmpTIRNx3Qlf3u7gDpw09cvIyFRlibk2C3IvwO
5rfdShwpwdhoC33BPsI0CZ90kfAt4j/XEMrGpBGV6r5NswUziH1xISx63G+eUxHU
YJ76NRE/paQ2RxgNCojy+AZjAeHSUvTgfZMuZo3OZznO5WCtQqr0O02s3F19h2lJ
oUgmoMx52kigmnTh5P/BXjZp0afWMYMvqoO5n8iQeWVQeaGO22nvbYl3ecOELe1z
nBvi+jHaiTLog3lVzJm3JRHpBkSw5EGSDznVtmZU88mc30PDRQOi+nyPPGVYUhyq
SS093if7LPQoOp77oyIjk3h3aV7JYB70E/Ya7q7XOmDGxndSHa3i51fB1yJLu4tx
ReXNB2o0upt5iU0sLR33JnFhNBaOdkzy38nr+eirYZXJHDs3U2cz/pCTEPlBTu9G
fbp0+LeNO+OlLbI09mzBYu3AHlEpaZHFgYE2E4U28dFfZ00Gae9IOjpF7GMz8deF
aHNTBLHEwgjngBlq0d551sz699TOqxmgbkPdy4X1GdnPYgMtKkhFSRUd8kVCUWD7
reyPfPROiSb+91hB94DRjHfvrWLB96UaKNqbqz8VOOfp5f+bMhpwnxNS+SESvf4T
rm7DNghAPaVRKpqJmrJGnrcX8w4zeREy42I3fvgoLGBneHQoQVOYByIdnbzAReDo
hACMp2PGQcRsfAfVWchz9Z/9pEFPJ4TEcYIfJHrkgeQ5eJZZJysHTWe2j24ujmbB
rminaH2x2yFZeEblP6EtmN39xXWvjIJkwVij9yoWeHZEAQ/TEIuHkbn2t004d3TR
i7JvY5C/YqiNSeoo40Q+jHN+UqiMSsvue8XmVcKFkL5F0nyTJoGdWkq6UT6Fj1yh
r9Yja3YJDpogAgq5EeUtmxvJkEc7NleRXDwNO6NhapXzO/MnQLTR+Ultezh1u4nA
2Y1gy9lAbyjcI3mNgzUk4EV+CcxlfWSH8EGgWF+Nu/UrPV6gS0Wr0JCL8CwAUT7s
DGDKR7DOnTOdQjwHrAW/qV4d4KC+3CosGGk4PORmWdXFP/oPaKhJ8dbsO91nZdLS
BtKZZX1J33O6X5LwG7+Z8qR8E9PUvjo5DUm0tN5trLm0Sw9gNO/7qQ9RnG1RTukA
+KAQsW5nbU9FZqBCa/duCht/rfY6LUBIcS/aMwIqPgwaNjg/VsqPcAyi+euQ4iAl
xzFpbOYPJ0Me40tYktMJ48V9ZOKxoIQCZl1iE7FuABqXpztsnX9O6XsPzjIF9xOk
ZCWLeeo2ynEmWclMn3C5lNWhSP8QzV4L5NAUoPgD6bu7Yj3Ccb05tivVcdSK+vD6
2YhgsiSy1a6KaGbvzRfTuUrUXpgpGiJuV769a58rAPYt7XLKOSAV8YngTs5pvRn6
OeCR5aGNMzvY/5DvSwckOD7owok3JeU4Scr6IeC9+UF7YJiwuOU7XIyK1AQBum2E
qP1q0fSQTLr4Jnr6sN1JO7hjCr1MDqOafXeNg317WrKUGIepMyNllogjSil4brs1
JpaAoe2UvA0V5X6fxdFQFJ9/Lse6XOD2KwSviHoTe9QYt7pPj9wNHJlLRU01n0S+
9vsgAO+jVbjVenn/x1JKgJd5GXecTvdI5i8UXtcmiv89JmCUrilXeved14dQWoBr
alHpIlFyrYqprFY50547uin8Co53+zAc05lhpW7TN+tgZcg8/XMGhvsK2NNTgnJB
NE8zMWqIViDHn5qMovCP2D8FidQ5WEouoCzZTolOL/gVtCexCjPMr3F4TETheusk
Kw2vaHlq2VhX0oTg3zBvcOtc2++x64UAfZ1ySDRrwZT62S6m8bZzzWblhG4OzgBf
z+fkwZkySN5GucruBHW58l+H7NlVcaffoxkh/SaBXywGUrbeSFFkjUML9Zop9/2h
Ym1yb19NmmjBtMO27//w4qH2KVAbbB0jHFeeBZnrK5H2r18aQMEdEPHQzF0uUDj/
3azauzXw2gEqiCYIovB9JWs2GpBnrLl0L2tC4jAe0fn1bi1NXLAW9xgn1s7XZic0
xMGdfGMYKgOiRAmZVJOPhsVrwa1R/S/zfBwuBWYeLyneGUS3V9MXufN8S0t/TMBw
QzbbUs+BvscjTQNwt8/yZHc/yqb2NLglwd3wvzOOXr6qSXjXsZxaFULUFq1eZOr+
xZBiktB+kiQUwazKBBUQfHF1ocQiDD7iae2JPE+MgsKvXPiqvP63+fSIByzZpP0v
IirRfThL/uVvMMKy5PBpK2sAdxukQs1WAmEzXjzYm+hK8jzDluO1hgr8etwHQfei
vpXwhhN3Q69R7NZBhHUp60pG7s3rp63fhRIuSkezHiefeVB6Xep+UjOO7zVpBfSU
HTUyIIqYaTDVBhCEcJRG6+rCLLboLBBxOhAMFpO5fUQBA3ILyN7++C4xiZOFM4g/
6qN2T23xsfTbMwhX7yslWf7FFd6oiTbWULTVtl6Y3DqmkNePgP+Jb7JPVW14zhZ1
z8exdCdLci3imFfboCUqaGyHCjhVBP9AT5vZQBTOoAZCfz3xtQEO3j2/el64kgQT
42u5bXthzwCVLOv8lUMTA710GPgGdp0hU+OueNtmSunEW/bWjPG/0BDHkiVs6NE6
8ExFFEX30NSer0lJJFV5pUOVYC/+VodrFv+ia16UbTmlAjjaBtX6Q5ejF6Jc9C9O
2dZu9SEwPSVcM81jrxPXK25LGmpAXAsxS8D3dehaabxufqKW1gJ+ow6M0XK0imGL
uqbYc0r92KG6vjaKHW88gbOOX3NK+yASeHuI+r0slDS4Lx+XQiLFe0CDLl8VmBTf
kBwkQvJqRZwYyUfVr7RjSryc41tMtgKtxuEUHTz2OMKwaSgYqBBH0GWVg4ehaF2R
U6Nx3nDPPbQsEP7RcIDItsRIvpIu3fK2bbDqjNcK9HGAM+PVl6o/Xv8jISydOG7/
0XZyP9PNMUXvYf9Pl9z1qnCZqBzXu3Obk924EjYZVf5CwQWjiXnXZHPJ3s4kS9BK
8730qDSW9lRdiJ3O3GDeA0vsU5Z/iDxISaBmaCs6U2xpAcaUHXJ6DjNWBjxeFjSA
cNnE/IZoeCFZYvrMeEfPR06WcFOw+yC/NBIxzq8UAYvyMHzu9MNMUbXCaQswT15C
YOYpYPW5v/yblpSuIF0d71MgYoVFFg6QLG7xhL93AZ3HenzomIVPtecPCtRRhSr8
qkj+x578mwUemJb4xffnc8/f+lLVChakTq1VjbGgvluV2AC1d80E3ydWbJmcEo0j
DvgYfZnEBzflvR3H2YBZZ/fl9u0a57SQfiUfrllDuAnJCde0Aw1pDhnrpNZCgl1c
E/XD4YuzeHLVLzQrLcfn5Wz5BGAIRopM+o3I6TkT+9CddrTtOE+fFfXPpLysecDJ
LMbb24/eIok0tZ0D8GCSojQqINklqB5CMcMLbX+9NUKw6T/u5Ds2dgq4n+jjJYhu
UMg87XjUhqC/Cyrs7/QgrNPo9g08PGk0xg8NLh42l0yX2vnegE0dAUKDwqsQ+hcU
jRje9Y5YnjoWiacdFskSUq16cwD8IAt9Zp4W8wIqaeyeeXqToMR5Xp9wk1RiTtll
ejeGgVh9jTInWS8oZesFhZp9zkU0oNYjvRedAQbG1aC3UKzUi+6vmG/XmRsJ6hIg
1tQ+/OCiOvWeJE5OVuujKaoq/uJYJgyeSqQ3/ma7s8btD2y+hWWPNHJ2Q3L9CGkr
s5nzdtPXdwT6T4kAXl3AC9d3KhdDIPH9B9tt/OD5Dy+x0/+Crhrv8CB+KfZkZB/0
v7S9kY/8DiOMyj5AfuJJdE9oend+8YcOdqcLHQoiIASrsWqyaGnnqGNBHTn/mFBx
sjAKksWuUCLEnkesmQ7PDLYvlYbJ/ykcjVDEgEGqzAQ13u8xdDurl6w0ok/Jjld7
bVmojaGWln9FMb7AMEhOgIevAmlIh5n7QiF7n25pGOTi4dbYqJffL9qJ9KPAFpe2
2K3+6mXOXiB5q3ksnsfA9v/Ui0moermIMYCGBAHcRGID8NrO3id7u/RKAXEnQfXF
UN5v6mpxaBpBRk/2qfbvjIX5OrYPuvPNF2dd86UZbI+lReEBHGZv3OqxZfCmP9pD
+u/muBPZ31iyuEilI0lAl0dT8QIgAlNBPgbhjRAGrTSSvI8R8ROGfY65t+Vk1BHW
V7oaW0bt9mizluH+0uPhsVMLHXIyz8eL5qtFHHtnZs5oAM/1zjP+H6014F23RT72
rp61c8elx1A7WAgOMNgu0ecZrLDl+RMTj8gXZM55PNTehl8sOoeslJUQboVZe4lW
cTAlRCHEgm0QY+bwZmhE7v7wUPo0nXri+w7pEI+qnN0JeH6Fn7GkE4DB0Q0T7Ctt
sM5c39qT6Ejd2sXjTaU3wFGS5hpb8C8DILwIAWavp/zgy9vU33+95KlCagjKCgWt
NbsSdcUDQL4AYgKj5Rt5rVF406R1HgPmaoKNpZDfdHuwrlapZNnwHnaWUyxUV9uJ
16FgLmWrIqx++7F7pUBYoSPJeWif7Dou/EB0tyKwj1u2AFo66/JiEdhw0TNYQ0fz
6jJ+Hhtm7nM6WtzxPoZLbnLDewxYfur7muZZk7X03T7uMrzF5T3ZzCqSk3V8m0JI
CCZ6ckBWvBNYBY49qW3U7bySxYA17yrK7Ei5T3qLuFfZMskxMYJ8zVDdhP+tRYyD
ZnLOPcy5Oq21h9VteLLXzwqYu/zZTmuNw8sVuNY8Hmsvk+xjDWMpJNg2hdYsVNf3
VIvwBAt7cRV5/rSL57KKFePdbHreoPs8QkEW/QXnslH/OuCd9PwFoewBHgqlYmNx
gxlAlGxLv7te3wrlNcJnr+HYgSqFv38rJ5k1W125EMN0pEQ1vXdYvRDx2TnPR28I
CQTVTPJcLf7PfggeGkrWk2XHgmPXZuCWSdMM7e/EVTARTzCWHvogl86VsU1U1cyR
/Qbv/BsjWEivKQkgTWf/KqnMTM+HxLAMa6ewWB+6PI2dIsxcjRrI79NC+MPk7KkR
q9jiGx+X8GZifaPFhCYvj5cSkRjx/A5g9NiOR8eX0kSgzH4+++gN91RsKL6pXPyI
pIZJA241h3mz9ch9Tdan1x386vX9wr3ctjh8r0f9VMdpsP2MZ+1BZVvVgLPf53k8
l5xPLMAcDZhfpRkpxVPShFEllAwOXiiLx0srYKxoBHfIMkhNtWS+7fuMIzzz6uG0
K3ZKd+f7zi774v1w0898V3xgrloP8/oFTtg5hbILqYsMBDiCbI7qrgwY+NR6BbRC
iGSLb4xL3Ziy9AwOViQB2JJc8UfV9RGROk6zL4pWyXBhmr+fWWBth0rDcHPA/Ndw
6AemfN3TsUGr1ZKpd96lTwefs72zP1lytdfhbJGLozNwI7fBRJrEf/7NkL6vsvcX
PCqJF5oP1vH/NXqNwt1BpXfsw00YzqFFZh5ATmZqR68uCVZI2wmb0G9j6Ep915+J
tIieDJFgq1Z+bQecuk5oRlJWHWPhsphVZw7raZlg0ma2Q9DKZsQ5VMitV/E1RtFQ
3cdQephkhVOw5EDyZlDS/JLAr9ynk9ghDYlTTsodkacjHa6IrpCtVSXx7qZR9+Ze
30n6yKwx1Bjae6A0wAIWWFZ1Ly+ZLRap964QS6jYtGbAuo5uZGcQlPVudxwsHChr
U6XCu7G8o66g/6aB3wRDKqZ/kAH0pNH7K9NVJ7Q4R4ORXQ2bfujVFjXo8oEG9duh
1zlhrp0bK3sCMcdmpqSUQ2dFzh51pzYDb8iyT6uMkX3Up/R9Rvzs/Aa5WLbYBKNO
k+g6MSFEDje0g6CG6W1LAaOFcgfQ5edHOJjHveX+g2AgKjGjHqjF7jwbvrNsahKn
GzTcxQgokJw1navWiGu9saSMd4CJNnfr2chJH2O6+T5+W4NJnsNfqjkTmYSpdfmB
8gcPcaR499LTTKaWZvMi2e8KNdpMIFuWTwgXCarSzaiLjJxbGhFO67oI81+xUIfL
DhXbuD2EwWCwFZM2wDaUJaPxS9+RCOi9OgPoa2ZprnO5Cpl/cSkJV5TJCMpaNRmk
1VDdjU4GP5TKrbelV2w7onhVsWhNtkW/cFISi9w/VTbNXC5/7v18KEqH+RX7ZlMz
GOdR+k2IShgiSYvBzmrqHJ7hmyd0A7D9SF6mx90FAXpASereDlFDMEnm1bHDlrnM
S+lFa639OTg9QSijkozOFlAM5yXtAw8HcKPbZOr/2PovcpbK5tNnIft5c3YUtt2J
hjgsJTmKnZ2Uc7lNGwsZG0uJh0koeACQveC2kfNkxQoxnxjFQISQi0keZ/ErNPYw
ejE3gpAn8EFicq9IfB9KuAdktJkYY1Jk6fIouRceZ7sCEXRYHQ4JRdF/ve46MlWE
5gK+FkUAWXeEXlADWLxa/HvMVw70PSufysxcCv5OEBdcpp8A+LMzCa/zge0fqWRu
6cUj0UIUeyRo5OlK2BRkmKJC6bqDxDSk+V5pKx3vnfI8OE+wHpc2PT1E3hwIonn0
N62Dw7l+zM1mlm6X2253e5gPVQbDED9RKHllA1XA761UFyZUUSgY9UC5C9kEQvh6
JsnLUxWaK6vM1XAOfkoNAitaVubVgiUZLWKtI/GYDyodMHUPrp6PK+9i8nVc4s9N
cwNk6bj5gBlMR0uPU5mU+yuHxN8Ehp6VFFZoEFFJWJ+dYl2twITRTPB9vWzbOB9K
U32A2RzasVqkVAIZywzL4nUTbIlwREFnSg6npVWbCOhmBS7yiepR0cXh+rkkIt+l
Ay3Om414j+NiAWb4KuSWwUPiHjmbAlvKLy3XEpRXEPRa3U47Os6xy6Riq1OmntGs
2YWhAIMnl6p1S9rlb4wO3H6pgwyrwWezPf6hfWdGDf0hq01QnZQHKHU12icXeLLX
5zlr4v9GJ/JDpZh8bPejFoBDrMQQY/njVIspxwkma+aRspQqqAlE5F7KsQ/FrXS5
BA8HPx+bSOHr+NGPtPQ3k5IwMTKVDPW1P53OowatUE5n9kKoukkxuAYrwq3ingZP
haeGu7Y1Mi98uZ85K1lhXUgS8YefRow10c/kkEIFWqkGiWol3GYPFxnAsW+9VNUg
WuVvZhiK7+I3tq/qo4vU8LghXEKlNRq1FUPCV0lK8EXFX/DU5ayXEUNIyEN2+Nxv
PrlnC4RbxJbPUVDTyqxqVKkGXu5ZbeocKs5ZB5T12xmWnAzLA8LblaGJ8wvJf44Y
7ZYL2BRT6ReDNLo6noRisXiinKKWUG2hFrH3OAzlQ1WubDLmp5x3Ve10hYkyaMBY
bJVI1L5zuupzUA+Re7zM1/oolLPZFLSeJ2Z8li9Zx8tz3/7Ne22Dyu379d6iHqIX
r7rFizdUAu8N0wBApQuNM3trZPUICJCyseCiiQxQItT70gHnrX+kvabzkbFsEd0f
K/fSS0gDatwdymWj5GKrRroXRvUa+dXcnMdWuuP+jtQV5Y+UXLiHdBTJeyGKWstK
RtEbUjb955xZTICdE2+UmIZKV9ClpHMd+62JNm2TpsD4PLN6zmKqtViV0RrkjYZ0
v5PRY5Bh33vSxNY36MgZmOJitl5OoIDSJXeShaIYZdFGwMB4jnXwuOcPmrDCZ/8d
04cOFXMH688f0EmbCFqlyG76DBcf5qNfgPGLQBnBQ/jqOgNZigWIaxYHu4ex+q+n
asgWstALhPj+4qc4UNJkBJ39bcDQ8D5W+FvzC3hJ/qcr6/iAKK3LVeK7l1GH99KS
i4qA3k8MCQvGjA3cv/rh4+z+dFAozUK+9A+Iy2/3gXYNqHBJXyBcPKjyKSotWMK5
ZJZ8vNkv3h30iT1kdqh+rmPzU4Kl8K/ezzs0gQTlg0b94IAyhE2kvliqI7rQJvBz
gph8qnALPhzEj0TKgyR0bUvVmXfAcVWPip7acwQzDUQNXvVja39yFtqug4tttAkh
QCQKjLe19HKqgYoKCCVYCmm9JQrzZd+tYxD3I/KIkONssgGkSSyCKs/Nh1Jzu7Tp
1rw8pupl2VKf+ozL2POs7L+BJdJ+Ce+fGzfIvlOQr1r5fXyjPw8wMD1csc8oXgRh
1GQkbFi3PBa5bIak85epbv5NrDDvG/fIBcS1eeVaxXre9y/RQf53IUKGRDVqiM+h
0Gv7HSkiu6UNJOjBhW1CNLAjNOPCBQRXhQ56hSHWjGKrRQslrDONishxm1gAJuY1
sYMTDaAXLQIkxfYurBfIfJ3jAGK/KjneojhZgiJIHiFU94TdC9JVI+ReKssfahVs
Sf8q7ajWOvPgyj3JJgSLhXYjY2zdyn0YMcdU2QksLM7Ra7P0AG4BZf3tt8las8OS
7pxuwNAV59eqJL9l2lUVJ/TieMvnVjOItJLaZL0YlKRXEB4gfI5FfjOureCGsGVX
qS8cAxbPpi0fxDOkTs4fx3iw24RvMSifD5S66G631IYcdlbayt9dR9mWhg7l9kJH
BuvIFyR5wrYf/jED7Atd5WT7eMWVnDK6Lv1OLOwFaEPgGPOEKHnfE1phVGwCqNpt
PyFeTRNCIOeo45BWcAYJJ0Fg58gy9E2czhAXaKpZWhQJQSXp2mLdWbe9AbDbQFlO
Cwawgl5yVrqaGkfnUzRI6ALOQhGYGU1tM31KEIN8sXGJs4ORrr+dfajlr8bEMAN2
b28e2Ijb75+WsAoQ9djQos+arpdgFdwa2o/XItj2Ie083RYJe9xj0RPH1QGEObHe
FDezV+HzXzvWVd4M2r22YS32wxJEkZgIg6NkB/d/5Viab7qvBboxU2w/JjIdO/1M
z3t3HvRWQbwTWAnEbrIXMENdJJZvmx6yP7noO3abYE1Z2L+5ACMP16m76uTwTtvI
9XtRq1y/+/Wepdu9Rv/wf1PUWE4k4SyUe89T1tEzwCZB63fMoxsPjHyodP0AfTbM
IOXuhu8DTQnu68ZkbdxLQGymEQGe0BaLmW7I1UzPIdCZi4tNjEMGSz03kTBnh0GR
Rhiq05SzYS1riyR5g51fAyKlCJy/NoLaSgRPnZDlkLi+h6Y0x6jPLhVFFmtfJVAw
4SQcfRWrGoyscw2EyYSA+h9NHilvKRIxwNoUMTedEYizMhVLqj0PEUJP9SySV7hr
FFSZ4c+LYkRYx1SG26DY31Z9GSxUe5y7HKDUWzMG5w6BT6JJwEeWpua+OoBDEchb
VDZKx7wDnd6LcSpcDQDOVm6k1v84QoG03qPPQhts9J1kANizPyM0fgo/n1G0xQDd
A74Y3RY/j6aOOJFNJmRp40gD8sewGAb6141jsOu3CqXrSvpi+rwtQzj3lwA9DFC1
VLos4mSRicNoHnEQnwvQfqsNRgQCE7T7leDNmLG9RbK7eryOtUkL1ABZJkGHMvEw
YnS0aYe3rQzYYID26GjpOOv4bg2B2n0xIGNC4XeXK2BczwRYU0m4Qqp3VR9IleCS
bt0Xz7G1fW7Y9YOLWbM/CsffvIrPLvYEt6UH18uWmPeRRtYdQI9+Mj7GHos2ntGs
t13hK8En5uBF3b5QS7XIZPYxkp6NDEXxjNfaIivke0FoSNtBi3g3/rys3vRC1utJ
5edLxht6ozkkQKYbA7zTJHUzNEPr+36WMe5iim5PUwjusvz1nJCWVfaLfibtMjZn
JEp7Ikw1YDtCuM4HEvNEBXJndCKoBvLx0toS3WHbZRJhz1n/tnR7nwIkW9RtNIUH
+6vXpCjMLOpjrMX2SAxUJuk3MIYLAIP1SbjEMRCBGJmnPvyBjfzGdDhfdQq7rmBe
EFw2hjPFKxwusXd4PbeNHv1Fxo3PrXT3B2r67FJNv5ArtZpBukR7qYgPuaF26qwY
+fXE7H2Go2LjKP6XRFNLbg3mHT3eBUWD3HnLcUR0LkzT7z/XdM/wqaHg6t+rc754
FS5ug+wjSFj1mqCZQh9qcGLiXvTMzLTtAdZQ3xulsKp+pyim52bufPHoVAIkPuB7
2KURajsEWB7039+MAbAwy6pzpbuz9l9m+oTkWg5WCwVkxXn3ldVRoO/eihaeObJc
xHoiIOU+1Ig9+g9DWTD4IA+2gmT0BH36PgL/zJDjf5O/Kb1nkWgcNOpQgsNMlGPR
gk4Jri4BOhqYAbpQSvBIx1/fAdMUUbWjhOcLNqWByfVagkmxDox6l3PCZWIHfmMF
MuxTxXeEzFdH9YHE4P5wsxPJmSgKSvl7dpsX+bJamak0BX40OadJNf6bixUj/ihV
qmjRbbn47eYPzyJ3f6Aai0Glu+zQ1MSHJUhemWQcRpxq8sCjukF+vvtW9XBRW6Yk
aE29JSN2j+x+HdBngRwXUenW6xioEa2mvsDBeZtg4uv4S8PqCwq5c4CQklGtAI+l
A7hwIDmJg24s93lk7KjqKH4Z9/TD/Z6A2QNU1l3NTHu5h1Ok/yb4JwbXibdbff3k
92tIpipc6IVA1x+QzV1GujQeOKUqE9K8URgkSf8mYGlSUEGL1H5y1Wx8U5R1v6Hh
ZwXmovi8bxMOIaCGE2Iid6gJltDDTctYU1da36suWBKJIR+vOH+NJrA4ciu7Nux0
hNRWX1MU2UxDLbobWPiQgwcYIz0GpJHr+KCMg+rJUsTVlv67/lOUnf+RY+jNRI5W
Wgv1Hlo2OjkpM8DRP+8IAhF0ktGzViSIicauHWTxdImt9jb2Vyi94GCdLtS0Oi+U
/p6q2C/ij1eAzR7J2BbK+7N6ZZgxn+XFrOwib9mnh3ExrcZnQQIkgAcscDNYTUNK
+ohotm5hRPVda0JC1TCjURlbAccjx5ZAlFs4Uj1QYO7yZZAUDuPt2tMMUaIRVmmu
nmHpII+ITa1ftvIqfATEqx5ub5o8BqyZoKKqvc5p6wW+e4FABm4fNLyJie/uI19/
fX0ATqoeU3mcFtcx/FsFzmRiUVIASeXbyO5HfWF/2f4bG29ZaB20AlqlhpE3xIe9
Rlaazwa+wCEI32INIddmKQeryWPyKQZJftglxHiF9G+owsNJc4gMzkoL2epfXtIE
/+l+wwQc7kyvszsLq6+sZJpMcQq5gmrNqwarBtmThyt5n+GAfqs25leMPTp6XzjE
KTaRat03SsZIULp9pgayreRzHRR6iR9/HNhw9ERPSdB9IqWpWME0Fu9ulIUi2i1L
T8+QzZW9wJ5sA/rFunJGccdBi9Me8v7YCgVUVtGewxz/RyMeFGUS7C2LRXPJcrc+
oseH4F+/BSJOBLo3mdVPXiiuVl5/LIx+8BDWiCFA0JjLlzN7K9XtxbIvTS1w5Ieb
qT/rDa+tCwZ/Xzjp2DQL2flWkq8fsFeempTSRcgLaPaMRNo9zvSn1JOCK+DjVBN4
pO7aVWxbs0RIPdyOCLuKemUinAWFuVIBi4956qASqMjft9nimGv+FayunIEQ6N4J
XSXwRZPpzPO7MSnTtcsyCYfmX4ID9WU3BiWq94UzZppBvZlN2BmuNa4R/88WnjP3
JHE+R6yrfctMwdBgkSUlYPK/4caMfxw3KptD7Cd2R0kDsU7mdXDIxexqxWXIpLrP
3b5oaIe6FvWz4A2G137RMGEegRTrK4BH5lVye5ONWxGwWfjbLU3Xn0ZZ21DJMsir
acj4iMVwKCRtnVV0Gun47Sv/H/6mt1np7pYC5YwoGFdx0MggZYRC2Es5xM0euhlL
KRYOOjLVHlL5N5HHkQIxGa4cRkgj0qOhujcqYRLf5ifeIjLYbw/qX/p6QH6w1NnN
/w14P0bRtwZwWqoTszxm0jnVHccBo0+Fi5UAsgdlsvOd+704dKjPlgnUjR5loZ07
BMVfcr7NBz0HCt2OpI68GY1GKc6v7Q5FhbH0YLVc8aKaHWI68YlQdDQxpXBzMzxk
sR1AjpcHq6aF8kg26jMmHnF4UD6dWLn2Nqxk2HlK4vv/WOfeRi+VEPp/kFV1VMk3
a275TpctCySUMGvSvzv+nZU+V5LdUjkKgogf3R3Qz/05Cv6mUe84EzZSnF0hwv9g
I3eMuerVR5oJDTUBUffgfXzn1wFxd4tuAfWYSn+Qh8jVOZHvCFF4iww1RTXjIrHn
2VERwGfH+6gLN0lsh7Jk1w1Xd2N8KpPATWVeRQ8F0FhJODIzs0h2eaRFvnuv5i00
6wY5r70EgU+32fMX5K+Kh0OdnoDyrFiuZte36Q5L3W636PtVDGsvr441SYch8j1W
VfPs0WeZrgolGpzCc1F09gp/w6WrULXlMGY5Ns+SfW5CoOQb+hg0cURhVG7jo+Hc
8RQwUG2G6KkI7xNBtGaiJ+LkuaJutJz/KnOY0ABwrPQwtZNeWS5Zppm/RLejKO5C
U8jRlQG3PQhJy465Z6xKSS63h3merp2U/uZcvQZ/hf8aTeSyI4XXpnow8I3XP65D
DCYCXvL0R7d8+d6dm/w2jwHfFjpT+LQP0l94pCILYVgaUs7oyHVyG3cyApQ/s41J
ZFySSgeNnPF1fKwXnuadNpC47pGJHUdUJQhe07ZrAAIfmCd05FVyexp4mMI4Czkv
Ps7rNwQot12iQpNFUwmaT1f9d0t8HqaUKYsBGisu76KD2rQtOyEKkhVn13AZd1tm
a74dDNzbEbqbVDXy54RJ3qTwrkgaUNMRAeXDCmpHr5BWKsWu2cgPhsClD+TsDq+A
jRrlUwevyPAqTnH1LSEuf8C0A8pK9nSBFt2kKmCd+y8d2dFkWem5H6ElOgBwlSXO
tWWqzUdCJQvOVQ8rUSwnVSBe6fF8BkukSYgpHAkaJeXku4l7TlLTycK68oPWWF7K
NaCnkwE7P1SztqKRA9YoJ2WC3ymhvSCyWd9CrDrIvaiIp6hULpoSLUi8vr88A1yf
mvg9UANRfzCkh+IX2XumtxymgLbYOsX0U1WO3nsQAkpqweUbfVobbQkQA5PnKOgt
OqpmcXC94sCO8EBd5tPbmybO7wCEdNXDpPvmxSlLI//z5KBLe9vIg5oYiUj3Jr4i
J/FX3yjV/sQs5ye2bRxXF5vOIun/GP76FuP9WUqIY6BJ2VbrGPj3S1ZVAZI1COW6
yDqU9GDJaQiadhYVp5zC7FPWGBFXOabgL6hEJQn2J9xQijK3u6KtwhMLJiiRMN79
xl2/xWdP+1x2ZMTkM2DgyJZZqD3FvDrDGpM1jFsE9JzfQ4X1FLR390jkVUgji5n4
tBDA4RYr65L9P6gKtnxc7d72ZMQsZzBMTx10X9jdAgKpHmZmBSX8jkFPkC1qdjTf
HssTIxnX0XLK3W/4qZ3oULibxqz5jYXdYjeqDn9z9xXrT4ELOdiq3lIRUFY4o3Ic
C/8N2vyadZu14cTZg9cyhneKrJ8uPt4NOH1iHRZLBX9I0/WKyC2F5gLrxWvOOZBd
JpjRfSmnxlG1NkDK+42eNAj5USZMHUlu8H7Xfra7v+gnK+BlH/Pb6I5rIe6Cmoo2
4iH7sD4MqUW6KJiHSTAvDjm0wvqeWdm8UdjIDTSJj1qugAjm+8fboQ6hnl3UCxSP
I6EXcv8NhZLo0Y8uXAEVc4hmcJAljX6Rl00mUFoijbL32n0Ko3wi0osX7pCkhWBJ
T9WOcCUsiYT1RIz7z38UfwROhfEA5UyNVESOTXQB8n5fFG1UH8+mCXWXsV3Fn+58
ruxvJhG2PFju4C55UnMdl4VhipkOi42OajvtFPTnXcXUdE3DrklvmE/1Ng2OsdXJ
GEOh0dQUBmOwM8wGq/PzmuwErJe/osQwuVcRIharG7g04wfvRUSFCPIgEU6tLOMx
y0fe7FcJlaPfRuqEq5ILJj+sUOHVMD9LtLLPxhp2pcqQEX6MzGmiW+RRRLRJO0Y2
oaCRzfI2G3T/waExPd7a5IAOFBkzmDJDfZftrj0Lo3cDesvwHMtt3QHzT5pmN2dI
MKlIO82O/fWpxAbwsNXOPTWzkMtnJF3hYYOroIsUAlUdMOa2KfxPOaJ6LgYfBUKO
kBXEvP8thSV0T//h21EZr5bA9n0XPJA1YUVzfWDGUeqZ5BQ9gG7AzHat2XNMNiM4
jgRHHghA1uoTANe2KEFgwnNwAlYMvJOb6ZtK1ZFrJ4uk5zWkRjO9FNJWnTYssFrL
3BUcbKmV9OebY/Se/eZpOfgQlVXz7iiTYLFLTHGcpNfKA8SqG/ULEhMNQZgy7spz
Js1NS+a3p1vuRh0zDL7nlt7cDGRMvnQNpkeqC3diiA2X2y3158LyK2nr/N6slCXQ
oQ0CBc7XPdosmz0D7MwAIh5s9CSyghs79ggQ8S4ueio/l60pJDZDhBLAwMvi4qkd
EG/lhjobFcI16v5EB9Ky/BiTirctfCS8wQowWGDQHGsSWXfDgNtXB28qRXxvASTT
Q4/nzP7mox4UUnGBEyqWvmqKyHkoxkjHDuIn2rnY0yoMBuzyOUAAAnhoSzfZpv8Y
fox8IRtxErBMFNhRz8+iz9IzG5B+QCmJ2+UCRzEiqUv8LRku961lGOJFtU+eKIBy
KY+3nELO9XuNyMrHnhGAixHzsoSJuSkXMe8yLUqEkL/X/SoewACSu8DMM5pgAdMQ
9Ed6eqnDXQHHZl+Gjcjzto9pYFIR0jLPHE3yEqxStTwrpelg9GRRKqkJSh5T7x88
szqy3Fug7FefEkhPp+nHLDoX/cpgXVGeiS+vz6asPxti2zsZzhbr/PsDm5CIcMjC
NnxDYcx2Z+N1tknUK/tW6hUSUaJmp793tCe+wlMNU9jmu38INQr6knaeqfKFBLNw
nYAqWeLNMAoFA+VoYF0ZFWgCpLykhvLvwQTvfYQgfl2i2OF+6wWH/j48nEOcHPmn
F6kWNHDdUPLuOLbXdnGkky+PT1wqcndzqvdgzoKwfkcf2tnvUJLv6qv+Lko1lSDC
v3ZIrhsJpArWTWFf91i+WA8FnnSJKYB1BuFLq3OvOtoZeFGa5V5KZ2MeGqLSGEoI
5slO9ZY/T1/r49P8ryo/gs9UyNMCSJD9zQL7HQgeqvi84yk75UGRNVvu0+M/iMN4
2+gohYmY9ouzFkhp1+G4tzA7Mg456gum/c1k/OZsuN7UF7rFbC/+sY2LOb5Rpbj+
FwUCOSw7EuYTi9w0hTYoNNjJ+YYPOiT+PXLqJnNzezn+wf4c2zdWukcxQAnBgsWo
yUGuotU9C0wkH7jSWAFMqWyDLku2PBDoLeGPgxYsgPZbH78tvvF+skXxdeoo5mR+
ffmJk5/em/mcb3/abVVLSJufqut5foLrd+UQD+q9iPGp2JBjU8s7MYKDvmkA/1ch
Oe5UTSvy5mf2sP5oCzfVuDIJrliHW6iEIPQZgdCnhFTZcwgg3YAshwr40CmnN8bZ
cIYlyVzEJlAsWBt7gvTfxF6AkHHkcZQ8QY37sYZ4ezsHFZZlB+vT2ArOTaW6pQbQ
8H8nooWgkLJGYWZhpaK4a9zYX7n0zQGegUImFBxSo3K1A23bukR1eexhFXooH8NE
FjupQ/1SZDo2m06RtReEdluVrPtFF3nxhWW/e+K+98Fj2aiQ8Vy080jHP1IdoxXq
4qmrW13LfUYCDQVOx6CMp5o2fcca4e3dd8pQPzqFx/FXKoPakm7AnAUNal7ogXbZ
B7mchvKh+NwT9SdC9saDkpZv0WNWvM7JQH2oRNTgcaqr3T513D3Ns2hSGZZXRGN4
C9Hg8jumCERvraqnKbaNWM3KhAAXoEicfHCsFwunFMQCh4uiVja57fA7LGztUbdy
M4kGrsY4xRqCnLQ7Powz7cQfc1Lf/zib6JjmE9ylhGykWFilu/GA3wKbaJpGCa1a
1SsycpXKqkfBjVXTP676h5IsGvwch5Lqcc4B4uQccuXLUHDTGyEr3YmWRFM0PZQo
joH7fmQ1ICYvy04GECnU+0U1ef65BB/75fj9FC9cDKRXMCgdQdCqqTJVFh0KtqS4
PywfN5/h74ciabh/a+Nl1lMQJUzeBhiyzWV0KUVYwM59GtCXHfjaSatQsHMaZB5g
e6A4fkkqYJXbwa1eiRn9ux+CjlsRNy6/sowaj3emOUYgNcRymbQAF8XLeqlgV0B2
6GhqnN8efeurFZCGLqEh5VKYGVmZ2jV2YEqwUjL0Oy5qtlsWLyvG79Fi4tm6R8mL
gpKrySIMVCwl8olfa9wTeXe6jzxlpbYXq8QfrcDTjizoD++pUUjcbNIAhcNfo2j2
Qh31ITZZ/z+RZXgQ9iBb4hv1+gMUHAYx41l1f4J8xH6hohlrwlZwFhUrsFQpINpA
h9XYxfmK6lPBIEg3VtmFdtF3K2KDHd+v1aFL5AYw4jZcROkzEdfh6xgGCOeaXQgt
DD5dGPx95WWpABj8de3QR5I/BvXZD2mBakChYOBoVCXqnD4gLuxiiDwNFvqTdskH
crcCkwxKTPGaNwUUfzmYF20vGgf3fFYqPGGCFQur/nG+w2cQNqZ0x51hzWMvL9BV
NwBR2tkelrcnWUaqfRiwlK0lqtTTO/BRp43BUtAAeG+ytjI+Rf9EZsQjHueN+7+A
o/WBP5zUGeDPrNDxWOpTp9Zdk8xC2MO7hY9y/53ShCIBT+44uKOBrU66CiSL5yJI
EXdSR6fkTgvqqzhHVNn5xn1F6/rceEZMys6StYtWXx6uVo1R7IeknMGCB0Cz9wVy
8Rb163F7MF7UJp0zH/3mmXH4XG8OFEosAVnFPGJHTmpTj7yMcdDhjfSipweGnqsG
192KTAENp9mc3wDPPet/E5/rRDFb48XZFJJVRPVVVqOsFOjpfHSMZEe53xR8VX8k
0Ub4Pm19l4DeoddlUbM0tI4iKfSfiYP3mb20SQFsIpl8Hrg3L58zPdQFmfE/DQff
H+xQGQNMPb4qD1B/zetMyNJl9kdE5Sfmz48pOaI0/gggWZbYU1K/46gV5biMThU8
sb3Dwj+WidtNZLvJhm76rVEpS/FjEPezLchpS8fx6OZJUGrN+/KPXukdT5lsYSe0
TdDVHzQ7k4UBdfEjVdyXWBvwa6I60MNbsyYtYucJ/3QcJ0rU5fZUif8Myv7uzOTC
/UUWod7CDKdh/pcV2RatDHWsRKbXTE2SlbxI+EF5f+LZKc8G/+/YhI6Pltzxe/Mu
rw4ZITj++OiKR+O6aeSOGV+NgXAMKsP1yJ0mQR/7OXXJJ3t/I6mJctnd77aRGE7e
oyYR3quWsqRHbThlGirBcW4De2RytCyYt4/J+gbOKuNe+dHxyMOmvMm9KT7Er0CF
nd46GXk8pHgaWd8AGnJIDaMTVgrKDujrIax53nlXsdcmoHXPcVxusIy+jFTZI3/Y
EqkkJuQt1vCMYuy10ziAlpN35/7KSYm2NmjKPYrWEQ+DRXMdPXReJqsWb4r0ha/7
jDzYMLXTpXleJ2u5vaG3xwQeA1MjkwWVnHySu38OY+R254DIaOrGjdH6SXPyu7rz
1PtR1+/4H+NsE465tRjSS2mvaxLYN3V2PPq3hqX61jasFBvNwm8med/8jomJ5DcQ
tIDNhCo9E0CuK5t7zOpeeCDPDFlGgghKuLyz8vk8JN3k5zksGGyLMteYkwzccC//
Ugj0proYh2Fkc43V9JJAOW8UVOAx4raXi3nniJ0RYrQVcBmkzm1XPT306xnMabRJ
EqaoSb3C+3SfDXX8gLJe62kn5OVATDaPFcw2fOiOuTc3N9awygJSbdyLnUZEL0xk
RtdlixrIlUrLCSDdRChnWDkwjlFgZuhgrP1fHXP2G0l/eEP6kOvxZkj9gI7N/brB
VE2JOG3LJZ/sf0XBouRhdj2dTnqWplto1j2mX+cGbWVTg22CmSginBOQn6BYE9Ie
B6bUuKshER/QsB4XkZKkFXnjCEeOq1tzrx8nNCHOieSAypKUqxpJikhDhAz/JYk5
7kbXT7NcIdnNwiO5mQ84yvjIA66tl+5JPuMy2qbd/aQ1cF4XvOtp+Zg6sEZzYOnN
dItgzm1NiaV1czmfA8cubcH4KBSs2ZFCpGViEbTSxopU2FZNLvHGNvoz8P9pCnbi
yjU+JlfrTKz8YkUIRt0GAgzc77ebCL0aI14r6BHW4npFt3j73XLTVAFF35o2N7gf
U83OAeU4WnKpGo3WVQv4Ixq3v8oIBCVKyznx1k6AqmjBlUMdrrA0RgC41PNHpCxt
ICMahmA7NjBbZkU4cGeJj7mIJIaX0Tgi81Q6NHUfTQKjbZKAuVkSI3nts0DGFZPm
tK4wdpJBHVAtC/AUWTLaDMZbBgAin+JaOC5AVo8WyVg8Vy+acT+ElCa9B2AcMxiF
aY+gsxyGSBCw9nha5/ZJqjRI8cmTKELXNFgm30KWn52KY0KsitA/aJmEleZx2ZN3
26KoddPbGEcV0vvu8WB8vJutwtwJIijWCXqtW2UfpLh3pE62E3c3fWhDtZG6MnBT
M5aP20H+Z1NxJZhLmr0Rhm/mY5nCnEEQkaK5ZT/241toJTZZocbHeATaTJN9QrTw
yh+Bb2hOe0gT8YKb/HqYi5hxdwoXnCmTrgCUV4I0g0QclOxzj9Gk52sp7LtT1dcs
5kXpEaaTa/Tmn/ipffuNwH0LG99/cTkrWdOCXH+8dhEXWZJRgmUz1qR5N8H3CQNR
iRD+Q7o/JWtRA6oqI7yG6UKr8QD+lHNRAirREW5jRf887VjmuL8bbV+gNQapWmXk
3I5kXO2RLMa/cphgw6Rrn1xkywpw9uS+g3WbVua8u5go8xjaJPMBRq1WQneiOttl
DNyWbd9z1mkSZxxiTCcxDp/uOqmdysSWR9BwDzhez4dgYDZ/6gDyGJ+kxwkZ0hAY
sUW2ZNnRnkfVpM4zeJIjStLVoM/bfx33Q7S84qQO50qgnycOiboM7w4MYwqZi0S+
k7mbXN2uDlTnr4lT7PZYzj/UvzTDP+8jZ9wsDRZfZgSgLCu0BffxxtT/9BbiOlVU
nh0zvAeExc0oM8r1Lqm0TV6UmEeXv2dP3YhJJT6K4isdViZaUU84qNUEYdZ3kAhF
PVuPoSrwTcNNSiZirBSFBsnyJrkWHMqXmvIhGhaEUh6SK6DmftDEW2MsOKRoGfNw
oUyU45XQgj22o1kz4VnNATzMWYYnuQyxs6yW19xGpOmD7voFSXh2af1RdC6DfXoD
cyq1ca/xVPXxuqxGvg363lcfw84utpaZqyYUHO9WfRip0vLCP8M/71LptfMo/4PI
2ZC/tkpc0iKwMyKjrAI7yY+4XDS0QUXO2zEB2XU8umUmFVYe/6ZpyQ5hNzZs8XqL
T+FCeNPGervLLQwNBtiu2PC/wwrwjQGHUKd+0qewHPSkwZmrREDXODe7cqNdNntz
JTiFG/J8UAHFuk2K/bnQdeaVnyJllFJQHeaHjgeE8aYhBMUUESBR13mFLs11e5Zx
tEEVEkmJeju4ZdTH144WxAwyjK+R53LJZTQW2BpvJHk0AJTs1312zgeWRoMXU+K3
JwfQNjW6ubgzYXYLdGcW6cSFcDzSMC7p9o5B6xcig+VfMJWpnQhW+SHRtgIsKSad
ZtVTTXobl3Ni96C4EMb4gOW8hz/IaTSWAgYNOn2e9V1C9tZofkDWP/Va8uyrzAsA
TJYYr+EFLaTZZlf/ESpjOzUJmcTsA88HBB/CAFkrPhobO1MwPQoTsIL2dEvyQR7b
SaZIHaC7u9lddwnlENJIGwutk2lh2i0++fVQeQqp3aBZ/YA3RmLa2UEs5nVdOibB
DxVOSJKHeoj4mcLhHjyrXSbu3qmiHpkFBSDjahk9MOeNifzJxtezbI1Rz7M5QKwq
1SCG2obiuKxAoxl5y0uGQLttNxbdd6FMwe4bVWcKdmJO2yOk+2Yv72GXc7EiHb5V
etRW8JqPF7+RCAUSXi+G218Mn9jZXKgB1oKypU1g7cOxRotckpPs8iE25zB5Jtrx
i1sRgQBTWZn7oNRJfSQDX9wiJPjTM5nQi0wpoMloHkQngEIy4efucc21fJ7crLns
GDIetFVuMl9w4V7eAUsIP5om0beSznBgMqJURDV1sHF3rdBObRrL/Eyd6w8TqRre
LxTOBMmGGJx6nhIp0/fLLw9j12FvAq9hkEwtrFkNihfNrk5EBjNxVhrCDsffL97J
z3oC8nWism8eWNKd/JgDZQaO/Q+bqsbjrPRQUpT1n2auKTu3LbPGJ9rDg0EXq9tm
RuhVYSL+mWNge2jbb07RQ12qvqCujxp9P7IFKpQrKks7MdMAoX1eA2VCnsE0wAQb
wSGiwbVkYaSz18rBooElM81Pj/+t2iU21U+zZutSNkL60n5JkB/YvZNyz8UX2nnD
1HI4FHdZIU4dLN56qOClrHY1FSDQ9hMgRmbPegmmJeRPGleWiHDV6xTSHUttyEh0
hbg+WZfopblzubvtTf+k68oVR8HZydNfvW2R0e5vPmr939BkpTOez3KPve9XAQJD
3AyNLw7fCxsXUCzeTN7FSb/0FDBUZN4ie7YOHz6BiG4WGVJrD7z+g4GjrJ1Bxx3L
tmFmL9OA+Btavhv0NQ33Q3H3tDG/S2x6BkddYt4UsOmkYeamxgYumnqya3ugawbE
vVYolY0IaLuSy6mydNvMlltXN4nkLHqZO5I3wINIflceT1qBkpxznCO/hNGOAHin
Wmt2mvt3h6RBhGlRD2CAtMAd07oL9zMMLw3PU8/hLRx3aXEapthdX46IZ0opbi6S
x3s6Vg9rA38hMtfa7wBX3O+ib5XjtbdHeLFrj+EEVo8T8SkBnA08PTlllEyFGmkI
yaUQnSL+H7r7KDwkgPlXvPvwSFYNm/k6w6g3rhzbdS3iOWNGU8wlCS5twJIYJkQP
SXwIrUUWXFG5jAsg9FOZBVhKSr19A+TLzkmuop1VyarLbNptlqaNCYm8YW4h2OCj
PXO3srv2+aHdUULAVAEmN0SJD1LSIQSmKjBDkABsD1TF8tZt68xR2kEAs12Za6A5
obj4ZO0qsHfBl7cLwgJxAB/QUXWz8DzGKjYwA/tZTYg2kt2kCBgR9LXVudwnLRra
oeKO6INaHUgdKKRIFlb5lvsM418tLLalD9gQ5ieg3CiIPFOh5MoNoxP7DeDUduZ3
X+0gtg2NgE6aMGX0CjxEXZzskcrbSy0RrsI0+nUJSRabflCBLCA1AIbIstjnzlSV
jS/imCuDy+Uz9qHpJFV/Zsd5cTKB5og+E9gWpyXJM71XeS7Z1NI8Ae/nn9tY0byQ
JNGuWRKsICdtsbVdhruowY5HF6d/zRtpksTEFMd4R9E32waYeQuFw4qAHgvWcXZK
fLbyzh3FNlXf2A8CWFhayYM3+YdzPQRZBcwMa5CkZrs/Pm1AymhYz5plk4BEVGc7
NJ6tapEGpwrP4v7MDCU+trAOBelCSlxD0jgXSZsUVQeDV8dXFFDz2e/WdykHdmWp
CkcXnuotMM14nAXaJ+lZJaEHWnWWxy+bPJrvxjXLe2RYloTwqod9KAneFsd9l+tF
80fytT/qOsqh483YFc4fZd+9UMlSNO342ziuqAIs2feWvEQXnyzRqrOP25qvNHds
gqvYJygQHhZIgO6rRbQH4PPje5Ml9oQ5oJgu5s40KJ147ythKMldaks0/tgVMXJA
HeR+1Q0HMNpX2vQ333mzfaQlee5BV1qTnDKXYZxiVyR+PdTFKS5jdd5pugcYVUcB
6V/kLw28jEhhPP4kV1G6vmBfvX2H+Fj1unmthstUHtfEgXGFlFEPpad6QqLR2/Li
jzlj1AHlMy7Ww9OzS2Rl8H3DgVr0TyvY7UurTv0Sh6oB0OS1W+Pqa5kzvkIiu8NK
6102svus7utGlNy1xXJQf8Yb0De9OLd/C+86aOuzDP8gQQIzKJyaIIUl2PjmspBh
Tc61R0MF/IJHmka3KWtKv7JDm2P7srGPH/Dtj+dd8fdERTqF6hI24yiyqJPTmB5A
xgMSCGkfAtEiFfbUX/LRRn7iyJ1qd922fiAfgNTYY6u/AeUGqdHWS/aZtiHL9GXI
KrL8aPQNFbgK2ojcsyTgihUXDarkLb2ENiGPHEWuxPC6ibOBH9FT0BFAKmNa3P0O
HajcaahricODxh7ZI0afn2O8tgm98JbERjhn+EbBnzWSsh6ZdGArx8QO/xo2zK9f
1tse/zwf/GF4Y7uoS0Duv9QzQTBJMNyiTWBxLqs0WD+aK4EvbxsEqqhyB9Q3OZp7
xTQDirkS8vkXK6dX5oj6+EtYMBGWcd/bxrh3ZcCOcZ3OlI2DwKpPnB2n/cTs8JWG
J3eG9404aEWTYWifd++OqkrkldeyPTnscam/6i/eVL6vNAhBAbU9WKa4XbdFPi+I
XMh2183hIo6bR7MG2hLPjHMK3BIdH37ZzAgye4MFYcvnnuAGZ6U5Wmo0bq5y8GbO
BdHZSIJqvbBch9Jf2PzL7CjIQcoHrSgp8+D3cdxE3ULIhTE4Uk3L2x/rxMM0z5yj
LXEQ1h60LMtsAxz99T4hY55z/7k3x0GeHO2q5q49f4H11jw+0V+SflJ6m38MnHUt
d5SEsKtWmgKTRVnrFmsLjcFPZLucHsVRXLWDd3oPips/myOY3eO2KMku4ibcIx1/
wg/JTiRLB30EphwmPu+x0lNmALdyJUz+iPYcd9z/Lf7Kc6waxHfzZn5eZfzaMv0G
mq2ylNqOnOI82GF9z3lx1Vm61zOzM91v5m7fnknPLtCjJLfYligOFaj58lLXtMbM
Yhc46zL+AtA+Cjtbfz7fL9+vNI5hUydMK93G1RJrKzaT9g5gNqxNp5nBvwaxbCqF
u7OGxBk8mi548jc+EBfywiF9LtltEOBMXgc6FiucrKlWIUsnFwFd3oqGyYVmxC5M
ErV35UuZwgw+K2z470a0WELmpUHa8bib2hiis1cutzptHCoKiUkp5x9ehFRyPvZl
mrMjwNXER9jMaUqpCL9Xyw0bczvxNoFud5tWgYIMrjfvPx+0mXTye10XOfF7knCP
sZC/W2dgWQUGL+eUQ0nnj3AQKXIQp9LGc/BdNCI9ukocBmH0gufxaaIaDzvRhRzg
/2b8EsnbFFo4Fa7dnOnRvxHZLdcH6BK0cQScASJtUflvAJkHfv+1nLsZapuAogDm
/+QJ0t3hH4g1i9DJk9McN5cinfnhm/7Rxh7E9yaaW1fNOXxJOtb0By4+bknMGEn4
wtFOnvFfdSMcKG/9fGXndJd99S0S5hCbKyzZ4+dOeyMnwLA4BXUCKgNxqrs/1uPA
1/Qcf7uF+46DqoGKGnJVHsr0DokZHFhELbQv5ReNqfoqvISMhNdMIAwWlBZx3f8e
JypNEQqUFNEmhzP3hf68S2SPmbPBOYxPDtUr/lkB3H3oGHlGllMdBtzU5vZ/Cz2G
lHv3F45FfDXhkxuZGKhaJVO6tn85hk2j1Z9tmXtAx8sq4nMSYqkRugJ4OHaSxDY3
S7bciSYvFEB14WZnifSiNtv+p7+L4Tf9blxOgbC61cOZmaq1n1SXlaWn4MfWn/0G
z0wU5MVrPy88vc3pjq+sx/Lk6j4rOaQzb2oaWbLXedlqogoaXnoV4PADydKwnNom
Q12SmOvtVuiaGH/tRu35IJWDwVRozj/hQ9OPqhX9W5+wGGkiBuxl+xHWwBKdgEAc
0YDAWDxDU9qA/nbZ63CQCKuZI21pGcHPnAWzUekQZO0SBlRWr2zdv4SfDVK9ryvC
GZhZ251BAUAEw4iCd02aTO55YXIIPUaISBU8YhHOWXsawQlkoJHUszY4/yfQCxuN
rNUvzTA7j2AMB4NJu9oYuEPY3R2yC8tYUOYQG1mlIQXssEapFDrHdS+o0UvxPd9w
yVs3DaibyS/LDZVhlTm9cVJvcfLt5zKOCP1pED9peQMjKTsQVjhfFFJ3jTibEhNQ
WU5ouUMuX0RU1nCmeltAvcUFjdLUsIlIhOXpcw/X1W6BJhA6Due89ggEMQUhEDxa
a38EigbnHccBTo35BvYgMlnUn6WpN2gH/YFWF0dbF2HhvG2C6aZaGsxSJbQJ/sFV
YGlGomfAAC31fXP/g+UiwWniyHw0sWWZKbuY6rovL3o+6K3vTECj6+mBDiQpgYyo
IuyB/w67Y4H75w4Ve7teQuVXLFBHQQpVUa5DJ3HP+4rV8bNSUgCdkUpvFzuDBCm9
PCr9UjQSsQL8nyp7f3e/r2ltvSEnn/xTUKhZSg4uH1IODTRYFTO1EE5sXaGaobqu
rgMF+9J60jqww6vhM0W1t74t0RiTZOHxKZyVycQzLvo0Vkfljcx/9Y8lDVG+JUDn
3pdxOVvbsIeBWeKyElrpYcvYDqEr7fjFLCNCT/RdAt4u6CDfCE8Ak4jVHNDC2YsM
ch/WdzbIy4J25ndUtRdXTAyd8xcUniJSm6Sk0Th4V7/70p020F00frkcK+EOXCun
LMr72eG6xEU+pFwwyK5xZBUE/6NjhMZ2xKAGnvP3R9Ja5jG35K9MRV1MDuLpKUqX
NJFrslZjERvYsF4tU06xng/R1lEuGrT8jSei3BNUESj2eM13LzITamTkzJKi38EM
bHmQOfiIRly4pU6j/360TjZPmoEARjE1QkIy18c2Kq+V/CeJvVv8DoYjRuQSaK/Z
nj5cXRKlEVGFyPyCQrG3TouXzYv+4KvM4Zg1MFW85uuX7amjcrgFMcLiyxfrypM1
Cu+Oyhq6cJCZ/3+FbG4Sgnh+TDsUgiTTochN7ZkGZlWbGUD3L5Ug5yL24RV5Aw9k
r0dt5lRRLTBF3Vo73+fIL4/MdYmLGfhaYyLJXkbVa3O+U7aQlU3N/E4u2dEB+2/6
umtBz1P3cWD9z+BCeueZxyYDrAQxxi6Y27qUd0vHY9O8S2WDU2f0tQQcwEVzeP9d
foeUy237CviD61di9EQo+T+9a85ssW2Kua3FCyB7aPfGJoXR4pUjc1NVtVZQgYG9
0KGbrK77aHvxFXZZWLMfbCiaIuxn0JqbVgQF00y9sa+C7+HcZ3WXxOj9r6I0on/A
8yWRK7EKEk2MIZYMrgT2TZ5+wZO0qxEV3DhYToSsJsSh4eau3RtCLzC50mNjVp9m
hPfehdMCpk9HR0uSXkrg6qg6uolGdqEBsSoRdSv71RQOUzsmR0nQ01PMT4MZ1rVN
/MAg3Bx0FR9LAcgUEWwKBR7yvHnqUCEpjDt5OZkovqeRPyiPrpJ/PEmZV4T/sA+w
S3mHpdfe+qfAcIGYYNz/ucR0VzF/5eUH9v85dlt9h0f5M1parjV7ixI5Xw/EZEm5
od56n1glzczf8RXu6FwxQIhCSkRndElXPaK2VInhTXRIX8l02+gD1wErG1su2zzv
/esCxM4o6vB227vDGrJFCVztivY6uAF6qCjotWzavaU+VX9hh5mPDbVsHFMBjJXt
uTRigYXyyly4b7ZtVpjJ2VqvPolew5fHKYZXGSrLyKf/4Uo66LBf9Ehno2Mo3tuT
wZQSrhQnw9R35Mvej0fEuC37yhJ1cFMNhcxujSyqLUNlQUs+0haZ+pbfUcC274wT
46HfbtIwqOYUNPnJVTtmGcRaIl4bIE1xLWU8TDwLyqr2Hy52LJuwVey0z6FxRYLa
pUuJPwFYTuObqejoE8d4VaeYeFrH9ipBAHAmpHJNFcebMhVXkWXiSqAgKMPFVVPC
oTZ6mkv2DbN6xanjKcEoMKZklufuVuLgshnjUEF5FMiiZz//5KdXoWo6XjBpba7q
IyCJrXbinLcshd8LqLgNutjjv41VAzeB94N7FFgDrl/5O4nORwRpBk/11ewuUikX
qEYvbC9hQzatPaZwNJE5A3hDW0nZBRoPhwMgkm3zuDfg7Vl1yxLvyBM5Rv4lO41V
5nz8OTer2La8+wehcSRH5qA1fUyZ6tX1gVskuB0CqAJEw6bR4iEDFmied4D0fSpw
bDURWkztnWPoUmG6ZsJTcglSJb1EbqagubFk8RvhcO1Ks9d3sceVtyGApgmo2xcs
VeL+qaqZScbnDKkAnZZLxb6LUTQj6vGtdJEBQ19ACikvebj3Jt7lgdFUUQoT1hWF
q8Jkrv2Vw9KGv03LlwSikGHECIdb6U91X+3qkMk0ZqyPAcQz3FKYPrC0DapwQVzg
180D/4LsCu7zY4txHTjIWN4ZbwoiUNug1B1AuTx5REmQBGQ7/2/P0FENjZUbK2mB
Mcx7o7tUO0zPTBgYzw+EHY4Y/qjiHzql4Fl+KQKU0UMZ7zAJH5GUZi1SkBF0kVaG
MhjwELF+skrCpn2/K/csa9WV6n1+grDv1Zgv1wnLpYJTe9mcH31aLhNftRXybpT4
t6Eu+yYstQj3BDi9uzl/dCjXSS3XXYXvZy5/+CXUkW0ohFx3wtmHiWhMJaOggIA9
/gOdq1FjhO2/sXyg67ANHjmRoDnCcRrpyNoza/W6jqC7JNEbXIeoMd+/N4eoWaU/
sINpEmpUrl89rpvvHkb0EzUV9kfHHNVt8qPA6jHc2wgnN0QSPg5KADA5dmivNEEc
e0cCKSi70mR2Vsb8WgIOzS9W2pHY7DUPrGYAe8ra2fAXD77x8A9e3OIHdHY7NBQQ
jYg7dglq2kCDPX6nul/9C1w4k5XC/n2ZRx9ltw/TTny+Yl0glh8WvhU9KOFr42re
3wRntDi8fTBrYmMEiTmNNh4AFWIwf6aJVtaCCaLBkZ48jQexfZZE8EV+8iaWRzXj
3zjW9Xd6YHDWCeS+JAfi/b9xiBfEmZMFRQhTMDFrw5N9OpsjBKpjXO2KEX1gRe42
siFCpA+j2ulWyw5TChHb8T9axwFlSVI3n3x7ABjLD9eacHcIL0NnuvPKRsgHKGxQ
KsTLLX5NgeO5Bib2YaRVofzmx83kZMmBFcQ7ZGIT54GZuXMpNF2XDd5eJDNI2+tU
XAIjyIFlzWOOeMBgRddCUkcWEUPp1F5UJXUi3IChcNDsqEtZ46IGxojj8hsNewbi
D402AZLTaQ1KGkXX+obohC68aBU6iy1Vy6pLOuWnvAOJentEGODphPyEjndIqQWx
9O47l1a62CIbrx3KO8Qay7s+ZgOu9G9l+lYwr8TYz3KfEonNMOIsiUNKd6tvIwGT
SrUkQc4E1eVZrAoxbrdn3KAwMuzbc2qveiYnkVZ7oZ6r2xqRffyLNeFWcWkNbQYd
uKcQheoP1BMDg8gzVikZBM1We1d4XAMrsuA1S1NgPTB0U4cFPrk7DEdfoxTMtMAM
3VKkkTPsYdctTf6dXeNskc0PHexSqgtEr83ljNLO+uVy2TIqOiA+OPDvKVPiyHlJ
am7ep/yf4s8GgAvo7zF6SNdsD8NkLU81sYCXRKMhd7yyFEvmESc4gDpFiJYVVqHj
hol8mq3f+RHDmQEe7gNH5BjGF8Av+jpR9SA9WP/682r94KLokaccNbVJXIw/gsD/
+h66NUy+eCzC8zVai086vYPcaf3J9TSA0qttv/XlmsXFWfMaIh9YIhANy/1s4C7a
WU1DruEnySW+I9tZxGj3SRmTw49PdnGoVaFzQUIKhz9Ob7k1OqXaq0fpigR1WmUb
X5e0QvhPI3oMgkWTuGSXb+TNEZOddAJXUe6fmFK9MvvtCumjCF2VBZwVS3tENGOu
Uj/MM9TZsB3/GUjl1s8FL1rnKRgiAFB1MbimLjy0U1HBG5eM/iZ6mKrgOG6yPYXS
Yk5k+rJ7xNJR/QpTjU+ZWeH0m6T7DxyqY9pOFG95O09r1UM4gl4fz7/lIEAEGS4D
UgdnzDtOXWY7g5HM2n7BZTVLJBjl8gK1KnM3Lhy85fOvhgFhmpsBzha0/EuIqn81
9tBTmx8k6z6BzgI+FHIv7uLem3yIuSR1xYnl/ICYFKv/XoS0unmiSWiqbGFZ6hrB
Fzwos+sQmnYDDEvAxPZc/FH34fCpwkG+eYEBYETbGY6/VnTuP38XeghDHghZMDdb
oNHlZ1uEpB7sNGkoKf0Q8+U1sX/0BBK7X/vQpzwU845P1aKjOaZr2yyqR27s0U/A
arBFInHss5altBqFD8+x7JTtfyi5D2EiEtgDNQIdIVerQlYByi5xElgp7WxvhhWC
8SvkYbDnyRjYLGVBxV0n0yt6WrSuH7UhLPLClEbwzlh1ij3JHbAzsPHH6FFaDUg+
/Tl26CciZNHSgIIDQ8MOPSUQWgQ9djdNChVCndGZAdJnQdy+tYEeYRXPbGAuW7jN
oXretA1LTf3QP8RvuqwjBb8RsgDbIyzHjJkq7LoMEsgGpEvu0XNkY3ro/tQvTSiu
hTJYXWccbPlaC24lGRzhVGQi4M/N+3zglrNvgTtEI7k+PoaZ0jeo8KWeXQfFfwcI
mvlPI41wK0wCB4cSpZAgxEv9BTM3C5maJ9TIvohnj/LcCnhngdgNW5DKvXmpYEQJ
SZI0INTiI6AokIUFwxmxEG/zjwS8p430iivyHqLyc2pcuVXn234WTMFrw/bmRCQg
Xqfo3jp+2J90awx6HBIh/Bb+v+wCrrvDqgfakpDSQUcWsUEFaqO14M3z9RFTyO3X
51sRAE6UIvZ/uFsc9aWr2m5aC5YoDotTYMqcv48iur2DKzxlZlpSN75bR6Pc5Zi9
jtJuRLkKeJDBdBZDS52oKYhtdFBZZwhW3OSgUC0N0TfCwjkmnOnbEOsDAFvEiEex
JKZQgp3NUT/lI5NjMQB5gRO0AUc0th12gqTtdXryq9K/7SD/3CyfVTQ2n0WlSH/z
uvhJ9R6DWnjtHS4vL0sc1TKqaVjGWRyqvg24azFYPZbDTsBtVa32blAk0rMGjDj/
7bx6/HdYtehn69BrXan6gEuZNJ1W9yep845PruKJ/Phgotwd3otfXAABIf/wrYCP
kU8JywTGfa1YWWMpXHrJkgeQejHEKFLVqtwL2VrBK8Tv/2LhQstnWpznT4ILIrNs
Tgb5emruwoMP2GX4ZKith/HjYCUe+LhVnmlCAuQFlD6uQbmG52ePZsBFx3xVMfBK
L5i45n7igMjQjuUJbBoUyxZhMCYEiVnp2xT2zCqqlKSbr5OmORsrbGoeVAoMeT0z
bQ6NczKM91JCWkEeQ+QFaRIZ26gjtJ5lkyJqDbvTzCJFY9y978nuBIeErulHqLWq
4x41/EYWuMlCG7B5NFElAyd/V+QtslJLU5z+1oiV3/I4Sxx7vhqp7xqvDtBVYUao
BLw9HvV7x+yGNhJJij9EhuJIDt9FAHuAI9n+C3jWvJ3e4KQv9DtYNLK0xtq6mJMy
SwdqhXv4mgfuokEFcGFwSCc1dmBnIpkAn+jDoS6sojtOZksPtOqRBIVKu4ILiW7U
HAqm8egpGqrBPmyWzoQopjv7U5erkl0vSwvGUY4117Ib1wiIE4ABdqiQX9phm5sW
sm0DS425fV8U8KYW7duVjCt5OI67BPoU6eLG3KEdIsVbWTRKG62SPUt1UKPnr8Q5
+1ZNsono3pAKi5UnDGqJPRUmnagoV4KZsZ2YnfYz9sBX6gPTbkZarHKI7al2hvwK
KwCNsDouDZJS09a9h7NxrdsHfRqik5ywa22dS8w9UWuSe0L3ukEavyu0mRYosGfn
QltYqFZjmFdAcpcVAdQ4BxQah4635kBF/xLlNaNHVCQKjNsPhOcjv6mzhdYJqCpq
51WSeiCEocR6yu1C55/gxx7j+K0InEHDuV+zJdDyThT9HGE/a1CG4hoKatRtTck6
yzNIU7/7jpIo5TPGD0M1kbO6pzrA1KFWF/hPUueHZuiKTVKwqH4TqP0NkB2tY470
LWLe5sKUsm84k5uz09OegC5Bm844vyGjgQVWFJIsxL1VV/CfSzRrbA7u1bAWzNsd
e2DoqY2JfnFqKmiQIRLDs5w6YDm4syIn7+6Ct0bVxfh9J3m1FOfbE7HPSXcDVDLE
3rVQI5vf8CHuXY/T2SiY7rd84KifP7UjprLKbFbQtyQ1EToQeoD1uXaX7dEu0gCK
HLY8TariSngUNFLRv3uvdAvad0GnDTjnsIb5v0bn7hTNjJRcXqkIYTUkhiFegiQA
kVctK41/RIGUeOASendpiVQkIDrgvFZhtQ3J1TK4W3vn6MRDNEMgI354gmB8voV3
giv17iwpEcZYyTRlwN2juepPEdjNLlyBLvBqBOmYYq17Ie5dPRvG8fs4ei1bmu//
HXlFiQq7+3lfEE5DPGpFIaYmZLDQ9q8wTkXxp0g0oQb349Kl9Scwn4v+OMl32g+R
BTu1dJd8yVt5UryQnCJ8et6lq09TtgnRh1hDwnxyTZ/KgtRgm4m8w7Om7lXDAEDP
yI9c1tDWGaahFOpyYvNSPwSoeRe2DdHqkrjta/cshNgRdSCH0qJ+V39fhgwMMJeH
b3EKc3DMEaK6VvfsFKlNB5bXklXLzYQfYHrKkJjEeKbuWgZSUC348vX67v2UT2oy
q6S46fyTtsV91ug3BQpM9chbrv47vDCPkbafBaocHMu0qqXH7pV3JYq66UoAvevE
1So6PWD1iBAl9luVyhw5aXAcTQIDIMyZIEnUcY65aKqkbzuBhX9Wwcp+QUZGobwX
0TsxANL/mLyW+w0Tl3Vwcc2Q8F0GY55Fg2LcM0Azf4Mhh0/9RPBB0jvzAC3dhJkx
pg5GVvj4BW3WV9P0tsLwNv4qD60wxbJ9ljA7UyvzpZ3grgfY9uTfpYGmIfnpt9kc
ktdJnQSwubM4ZZYH2DdwHASEmy32G/PThIaO+pKs9GmWv622v66IceBBp30Afb/7
Keyb3ZMBMDA2DupvzpWM8dRG8g0H/xxACq+VJNfx9V0zK1FJJKovbS6o6jmWPGBh
R6IDFlxde9jVauCsEooagopNwFZb0/LPXALLMhcHD5P5zc+SVvd9ph1hgTXsA6Nj
+KQGG3Hv8yfS463v+G8juJcWv4HctvXDgh071m/CKd4GcRTgxkhz2i6EHyVVWBVA
7vIQPqFNDiLa4avScrXFJpbmwiV95VVDkICn7gQAYx6FbHoqfENcqu1rXPbxCxVP
tQ5B8KnTjsg4m1fCE20ZhO3nIjkPbHsUafW1ae79hZHIiWVtrCRC15kFcso5fFPE
VUymYEigBv8CCJyY5Io90M0K4eIWL4hW2Q5WDXzgBkIlqylqA3hB+LB7bjQPgDx5
OLR2rH0Yc/w+BioTYexz7YiVIBRDsh4tnd/cz1WW5iswBFzIzMZ8YrercGMnsdCd
R/fH3Q/dFbfP3ZAx+pOHqLOjzGpsbg+XTcnogZ5vu6Q98rCxvQXJcikf81GrSpiT
wmTSpy/YrLtNraIweXHdUq5G+ZjiNlF1ZfYCLNdmPNeCbKS3uPC8Xkm4mlZfxcLL
XOMNH39f2QVT0ij7FJCApcapXHA9DgyAO6XyzW0AO5/Xmn8N9Yr1FjduFCaOo9lF
AIhzEdfRywkuLU1nhejI0NTE4LYN22jwHuDWajEqqPCA+d0pXMgVHWFFck4VBQA+
nb+pg/CoEi/lqRdZvM/yLB1Cul3nE4LaJA3gWpOC/MX+oKNIUw9+ZzEMKEjSCJqZ
iPLpkhV9VgH4As7sBl2xfCrji+ntA67ETM9b/AKndaM9+x5NRELbRgb2xwIyiQee
LQOl7sP43nIMZXZaqR8O8usNslP8waYLCLPLzs4MMtx2uEFSviWNGxJz558WVcFr
AQecbmoZzxGlUlccfW7vNTDcJtxRh8hi4ElpPsTsOy9w8U01wYJjNfkZUWhvwl1W
OGM1C26S5WXoPZpL4f2V1gywaY104CfUgHZYs8NjaE6AFj9BWJWYPNadvFYmwS9N
8Ttz20LkRIRYEpAVpK3SrulwyTVCp3TdH4IWhOW1AP3WAR0SvhAWbGTWfdFDdb6K
IQruz/mJw+k0BsmVCRhgbWM82rzQnyz7v0W+8Y+MpbCGZlyKBdw7WEJJQY168LMU
9A3KY6BZQApqP2CqVXl+yesrrC3c60KVxqBgr8kzk71lbBY8g+3EJd/ZuYcYpoNx
6NsHLD1R2q4pNhxcKRlq0e9ol04ZZpp34vI8Lw3YM7l2hRwkdL54tLcBW3ykmtHt
+pv0wIIn7gQb+F0PuB5PDYM9AiZ87slgrwH7PqBCOmJ2JTDwvMvDJKHD2qsFHaYF
L/6XJGl0AgUCeBKKNPkmm98gw5aUCZhgLBRLPtGRSiDVHCXGCw/t86II3ootnYtl
ar578atas7tJpnH4SU/APmMIeKjK4H2neK8N9QoFKmN/LXpPIE2eGIGs9/aTJta0
StdAdhaon2FAoCzW9EFMIS7G18Q72CZMcR020XZNay+Mkd19CYjjNfnlh2KMsE+g
bNWvIuFIZ5aRTHIVKmutT7fXUtgbecIjhj+lGttBfxugEMGvpCi/DXtcePc6c4bx
uvnX/b/jfcdo6MdLvkZ9qV48zKSqk4OuUpSg7zV7S7LpIUXjlFPuPyIVYXhteVtW
vHYFFNE49czVPxE6xsU8Mgztm8T2Eq+OZxQwAl2fhGXJrkUQ6i8zfSdKy4e+jFNY
/e+gK90MunDWja1lY+aYJiEJXuyHW5cuLh8ReMqxwen2LSYt6GOMwOsuRykl6zYY
nDXfDHPAj1LNmn2eM3haFebICFWgx+3aoMOO+Op7PxV0Fcu4dvnb72mRs8y9IY+I
fuh0CbVVNo/dJ0/5n3rR+deMpPH9HHH+02kQm6/qGJsGhumqjkgQPm/wSkin0jsa
adS1+PLJps4CmLBQm9+dGiEIvKztOo/zBvbC5J2K0veLV52zXMKJ0AhPx8xnxN5v
dnA0jJ+qGmA72nkZ0YPpZ+GP3vZ2qGaA6Sz2AFJZ/7Cqdw5QP6anmiJLQDbMuwIQ
eGWJlkNzp3ozrMvc1KynzKrV9GHKE309UlIlQ1AUicAdexPqbgph6yU75j3Xh1Gx
uGD2+3/3+Oieq4YxsiyiCX2DuEyV787xST7FhryjHTIVF54vAOThJMkzl31Bpetf
GthZkwYjqz5koHUbXhX4PWHLDwewr+2ZIThP6aYGsbsuJdE9ve0JpBlTKzUxXbQg
+KLLf3W3/7pI/OM4CwVYccaulwKhun/ab0KwKwtEiGabeOBcOWjWHPQ4O8lwpAQL
rBX3SzTBeHhtMUJMXl0SausqpumKNyfn/racO9uwYIXnz1yqjNRR8pFlQeDQfdeA
tk7I7KxtwwENxGk49SnqrNYd1IDQIj7WeauWk8EEY1cM15MIuKfrLYLgHBLffvtn
DdnHJgG3Xsvueg3Pa+f0TSuyU8+dIwKs9BxMZx4UhQE4xjIgTyF/Auo55Nq2m3fp
ydzC5xrggEeJHB8QlhMJeIOsYoZSRCybFfA4GKU248KY0r+STBj2wdjidRDODfid
DA1AcgyTM1H3/IB33PCp8BSKFwHbLA2xmz3WqZzdUJyu6lPcYtX/WXQsHogfejb4
G8kYTOpjec7TbvS0ptkeTqjhEBkdIoYYJrLT1Ovt5DpyEgB0MmxeAbBXcK0E6i3A
sx6rVQFMwvvcE+y/iitbIgrM4QsW5YiiRfphVMV4USQbPtYPsunQ4KxuUX/NbCtv
aYNmQr75Yop6A+wQuY9bVrU+Jbpe7YLTXPhBuQAv/a95ZAl2Bbfcs8T9/+i4Shm7
RuH/EZuOp7s1tg0jVZ17hFmGE/FKzd5p19862E1FsgkYy49HW4/9e9l5Ej11uG0r
Pe90zSmlHsipYOvtauc+6tXNDwA0MKzZLQHT9yk1fAxFeef4SIk+BrHptzSFUdNp
zxH2ICySNvFTfu/SJGPzTlR3Ro3IelFfQ1nZ1KJEx5vRdMozdDsWrsCxKTCIXppS
v+SZtUsLDX2QoYjbeAKA9OXZ0jzxZcYX+Y++5tciEj1seTJ2GCaIerl2ScpSbwMB
DGHMgLCQDsRqAVXlXrC9+qjDVFTp60drz6jXVUFS2lOeNa9dEA0V4TRzhpD4UH7i
Yb1HOOtP5hfgnOIPkswZgzu02owGMGkxVnO+e3GjQzrGcIbjW7pafaeueOyChgtI
N7kqD2N34fGDgvNFxnDYpkLsMROsaa9OPr8V/Uhqvj1TDNEhBzhuMxmsXcqWNkok
mKnqAGxLyYb4Tx/nkhkDnk4L0jQds17rL1gigJ5lhezHrJrATiao79XFxzRtjUFg
Nplfz/adxeRV1fDKZu/P3y7TgCWwcuIo9tP40AVZC8oO+lhUZ1fVd+GHIpE5JLTK
H8tG/2pP6hEJo/7kVYdEJtNFrHch0U3cP83n88V2yzCxmpoXQVdHEmQ7mRI+/VA1
T6Jm7AO9XJP+v3o9gp6n6WoqrIq/Zu75c8yWA2/1ECEkBIbbr8yB2UOQpQL6YZul
rcveANpUTrBMcBgp7IT177CrsDpJsPON5PN92Y971axK1RnUAorjP/4rqDCjJMc6
481wYaf/1vfMs4LvPvzvdRbxJ05h2B5CEJKJMz1gRWR7IC4qPmowR7NbI2odg4vy
rzyo24GbC9EyOxlX/metcNKo7kp+fJD+1uZl/P2XxrW8arapVn54pdaQAngYMDje
L4DDe94qOz+FU0uU6MQMO8Wn46OtgAnpp9wGMgVf0t4pUQH1AWY+dvngt2YfITLO
mvb4R3KoVR1OdQbk1cdjo3qVl09jpkx1YDMez3cvIYcTsmRmTs01SxdBhhegjn74
iv94xb9L3pN9MPG9xVIJt/8BmA2tku+9nkGX+AoGTh9FgkGV3vtIAV0AeU1El9hq
7ST/eWi1mgQ2LNrvYT6SI4tENy0k23/CRVHzz8QLwaT2AVdDaDTKHwB2lc8fKkqp
B4rGl7/ql/fl+utgkFBAA65SMRkUWmYR6wKsBuaNl1+u0RCrqgviQKDGaPOzBlw7
+dONWYeGJE4iNZlVb3byTgeMW6eqo0Vv77QxP2Hpv83AVqMo88qtS7U1F+y4RkaW
JQgUAABrCJaeRDEc95ZARSJt0CTXXn5r+4Z8TQY34hBEweJGEjrUjfSXdfuGEhXX
/OlVbLTFJgl3sEr2hWHRe39tAi8hEJGtlMK2RLEw/+mWhGcWg5CwosAIfDYxsHsn
+rZVFoB25uxlbuGsCr5Cu25lZNyN+H3bdOQWRZ3b0RFlCzw478OYH3o9GFZeM0H/
OkrehL1cnSfH1HfHFCoqozaJxd4EE9AdQKauwbVJYK4HumoI6fA6D2JvWHF33c8J
cs6iAd+ntAZONq6HVN05/zu2GoWGtOCsE0tjkoxMKh6VR8GZCC7lF+3QbnucuWnh
YGRLJeoCQ2tecLeYpsloE7c656Ps8GYqkzlYkFy5Ts4sR6xW6cHdx3h1QcjEuonI
otB9EA+QuV1FEZ9lUAw2/A3tLMFzea8LxN5rgY4vBGxy6cADxw+9EFy4vs9AyNnT
yfRFaiZRJ8W6SV2HbcjKCRzma6HxtPYgxi807t+nRYWHUbDfM2KJ8rKlRF1REx7F
1tCzwXcPBRoITriJlSDF4b9M4BMvCSq7mR67VUK8c8gcAc4M3tCweYwOEfy4onah
+T7bnGh3Ex9EfYZHYcYWkO7IlMr2U2yaZl0XFf2vFwrbzlyqotROiMWbeXFLh1G7
wp0QukcnaSEO+VvPObdKV6UvFXGKkqPmwObu3NAEkA1dxglBn4Ta70x5EyAyY7ii
8b90fqViwPXGut5RoEKcMsIO0XcCP7htnYniCm/dRVstFI2DYr+EdpN3HlmSBamI
lJe1McBncQ0W+BzQgEOsYxCEPLSEc5TnD+IsxLG/ybdajeWPU8MJH2O4RhTUI6qr
PBwYRoPnuMQbr96uodzVCoxlgUJZcC6K4mnXW4YcoaQKSP3KQgFafBnY44vZwjNr
EeUuqFFVLcLOo5dSHk4FTMQqIqG9ZAIh4+8agW8pK4ZJ5PBtPfw5/DA5gkel6WIG
0c/mlZS7hyZL11CIHAhAEAiseRPY2ZX52LNFajYwBr/EX3J5ZZRQvn4ec+EoS4QJ
l9mKlyns0kQ7x9rbTWoMZNjPcOHNZafM767j0DVVASAawy8T5OqYXE9yhMxseEdL
0OKmpJ/Tp30dFslASX7VEPyTJhOToQT1f9MaskcLCSMfIl1DrMCetzuFxh/L8hrS
i2Fz7BQDYL+2ICQ3NgomnyY1UwAmdSeYAUVUJiektnLVYuiUNgofo9mbyLzS4bT2
+QJzIIR85roTjZ6h/tV1Djm/KwWnO6rek0exs09MTc8stwzNBrk/ndFJ0v8pJfC2
OtamhTXPye/u1FeOwk9X6aqQt2Jf7VstQrl7UKI9If6Fwe52hmStz6UuNHj0PtNP
r/oqqL6m3E2mH2g6VFMCIIhRAE3SYTBoBFD8rPTk6Uyid1L4YqFi8XAA40xlabXu
gVGF7DQl4Rb/OfMPgt1ldrxT1b9gtuFaR1M0EmBr1Oaz6CVdGBaQkDCf/ts3a+B9
RBoqPNmp58s5bzQC1LAmRggb11inqxLEosZeobmIhwOYFS7+bn11OYRNB6qnli5c
ciEw1wEzwbHYXjvw0BOv0LVLbf1Ysu/5fCZ8NO2QrW3gyxoua5DWbSXGrU3iKDKw
5ewe64DwBGj8LtuC20TVu0OvgnKqaprlHMw0QPnc2jdAy3TVLN0N6574p0IXfS1a
gS1k4xx8XI7Bytrubd/5X5doKZartOFoBetFtgVBnb9kktpunz+s4coFhocaWWY6
9lpivzdOikwaTDVsvnlIN2G/L8drjiic20/0dEHEMtdICx/Emtf6DepQ1ldyrT7u
jEldvuFf4Nb7fY2pZaIhZkhQXmXPRUxVcSOqtcfZ+6TYlLuWP3gi2T4UgqKH9Z6V
9sj9+xz4XFvjt+cGf4Ue1mUJ1TJ/rmgyxc+d+Mb3ohhY2k402mvmsMlPJhNZkFxM
lQEOebKQO9j1KGaLFNEw/tsvhJhuuVE1EZ3a/F+cVuaA/I5yh4C9PxBjeqaJjP91
Ppnco1rIetDjwt0h4dE3r9INj4XpIQxekphtDs7Puk7/9iSgJWGMrrMIgPM9w3ZD
aQKDXvfdmAqIQlhkg9svh2Baxht0R99QAxt+aGTCw+Eif+aIrzRnDpttDPycgYxH
GlvuNx1fSG7IMrrqysDzlwNpB4mC3geWZ8Y0XvaUJqKG43RTNUvl4zYOozgVIIGm
FCdF9l7y5UWx13OKabsQG7n6vsaic4/DpV49sJbNTcfrZNmatXreH8Vt9HW5x8Tq
wTdRAmi7Q3uytL29vupUy4cIuEukHnaqUWj7FsyTwlsSAlbpdYPczcJlRyL/4mfU
BbZLjnRAA2RDflObfkcyIYfxL14PFH5qHTgo6EbIImC3EscMl3UoVvaMS6zSlRMC
7p2NKWvL8MKS/U0vRXBTl56ynAhUTzJ4fePyDJfHJYy/1xG+lMxVOnmbYEQ58+pW
kTkoTQelnxHaVN6V+LAlgRCtJpylWjKurHzGvKjjzCEI5CSSq+m+2pDtVuquPN/i
hLKiwrET8KxFrz3/pV1hG96KzJSiKj0Y3m+Nvg43nPxkakHKX0XqkN9LhsFwNt2P
9Iw5pO0bVn6+IZC5PTeYfwR7eGIaA99iQW3DhtmFNVLEGqcPWHrJxZ5q83JiA6fA
zc1GmW96bRxLPgeGcoWqP6pS2KSvQJtY9eW1Jc8jdstsWc2w9O2vRIlQxkuiiTpK
Go1Q1pOzWEm9U5rD3goKRsSC+5iLWFUtbibkM1KEXev9YUfRbXDr5RDjLIPmpGD1
ilB8ccSY12nk7kcLCe7fnDT5PTNPSAdLJJk3WvJQ6kehfa4JJYdHtzH5uLIK2nDJ
zWfxLOaiTTyk91cR+rG0M5sapnm5EMa3ALlMolexwYvYMvVZo0L22YRH+Er+rGeG
wlHKm5fli0qnmWy0KJ9rgENzxDzqfxFobHjJemJftlQm8qQwSGiMglWrbwMiLx/A
QIouCraOvXda09ZZK4ST1k1ct0NLzUFIfaw+79PRQUyVwcvUWbiogeap4gQEgN/T
h5VQgCqmQHmAsDDhSC6mGJj0EP2wNjcoT2s0x/pcm+aue3ekpG/PI7bS+kEqzDdd
QLb4VuhPNR8G5jKHpfECdbHLyDpMj8Lvs/ygSCro1oGyEbRGQHPb/Vzd6Y+b9oyS
m3Nsxr8cHf8O8U1L+psucguyXkZmsEMIDcYj/8eRYf9u+EIBKg//+ypWok2C+Z/X
GR/0+o5cButZbbIxzqgzlB377L7WtKcKxHg74pj7JQSIeY4qyjwyXqN9tR6wGt5p
B+KhDOTIFovFvwxgysNX/QwdmMOJfSn+/Roe/V29k/cHHm3hIRYH4QDL7thhxWGn
nhVy6ORgnc6c6y1TNFdLHmk0o0OS2xf6J8cJRMvyG+xl7DxAoQ8qAoJx2OYwztv2
FrTlQBn6yV+h9tQKhzYewCFzdzwWMROL/oyFxq/xIPbMje0Bi+UfiwAoNB05UGv6
lXfa4tWhTll75HzAD3Be+lo19T3k9Xg9SNYlld5Kf+WCMTGVbGXqJvW54e867c/O
J/uIFAQhfq3G6jXpTLOBJACKNGDSdHh8aEHfJ/6loEd8R0pAe/HAIxbSY0YvWfFW
7Hzl/N3fcCFW4o2b/hHh9shA3q4mEz4zMSF1F7OnDy/fJQxs2B/2yHu+gabxXIlf
R5qUAa6r8xwH1D0y0AepZIsELhBc/RbWPdynk0t8cw2Rv2kNohb8wRfcNfVMRGdT
8vC+VCLhnDK4HGt8PDEkEtPKfpiLYENQIRembvSxR6VS12d6uTHt7AdECFJR36Rs
iWpZEbbvWuJQ8u6j+hOeywMcDvfc8VveWhI4gCGpY99U+yB6KuzeVFjxd5CHqxBf
1jqO6oFaFUeifDvKLPWir0Enr9HWWzpi+fJlDgY/wYio62ckkrzBidpeGs8Sry3R
k2hto7FdmJPm5AWjYRPOwBOwverQb+55pOs/s9BplbA32i8LMmV8FIgX4mvk3DHj
sfoXYrgE8LXGxpbEthUcmbODhmdv4XBkTkzFKkfl6z5LuOGB9ubCxwMlyA0HpDzB
u/KWZAOImQANmmRg7lXuwtpMTv8ms0SWS6mipbig2GtpUsCQQcy29FeJ/Y4/h6QM
ZrDX21OxhvK3HGN/Rjm4mueYq8U+IFvqlway7Yj+YsZjJro45fNmO4tSA8yTjZJe
CK1/PW/ZkjpldcYXFbnd5mXJSiSRQLL1ItPZGuDXn5aoMTkoYeksBK8hc3M8TkWH
5rkkmZy4QKE40KuraTPIgT57WgLajRiOc+rPcJUEHoAkirdYiLVdocbuGMsNQuqD
uX48zKkdlXmhuHJBsBX/aVVFrsbHheUC1bWMvg4KV3ctQ5UINTjo/PREg+SzQnE0
VsZqedjn7jRMOS7RtS988lG+yhccRsGTM+Rc4ULOM6/N0qsZJXj0bbfnVVOjWfSq
90fKdltVVdAFSD/pwkrxa77ynCeMkcmMLUCQp3XMEm0Fxj/X5HQTFFSSWacq1J1u
yPz3MRNMVHOLdlemaJ4NVI29THFdFe3LEklnCZTdSjgqZ2ainFy6f1mLfIG4Aq8D
ffa+G7lxNBJOCSfrOpSyQLQihAYa6nRzWXZxU1OXH0HLmOEi3MKYfGaLFBKqRxCX
Sc46sIdp+Lk4nB96eborGF/qYqI8EOOSEiaKGY2CGtHkKGaBFMvO+NFwEbN1cZaI
+xejl63xsP/Hk3ldyyCxG7rPLz5ol9yKN1V19iYeBgVCdwN5aILtadtXRASRtt2r
P48RfMkVXRToh995ukdrg3h6ij5AXzuVIvNv0YYkHCEKPrK3v1lvXdTAdQueoSoX
OMgX3SmQcQcZK9b//Tpmk8iLl2Qu1yRJVWL3hXaH5Ml5N2aGkO7p44a2XqQWnO8h
EADPM0v5wlmoHpFMpJ0ceeOcsc952x8LhU3cw4s31+5vwgq5lGC4oQ1WgpHeGkpy
RtrgRILNmq8FoXmbbhFJDA3mFE1y2usjidKM20vcNkT0J5fTFA7c7H+zxxRUCiGu
XAjOF5LAsD+tSsRoPuU1ykDOB8Nj+Zp9rcHYheQ8Z5TtY3pUIn9HBol1YuV1vZhL
uTpMKNLTnikrqbwuD/e1B4hmDfc+mWuWddRpiNcSPcinhMLVVw7mfHzDrdvkANYr
ruBMVLeXI067qyZz2OQn5WhJtq9wy7SUH7fwc0drU6OWnzChNVgw7BEFD/YgyUc6
wSoxtXHn1W6WSjI1glHkLW3Z/0t4PJEmoUFOTEc0TEYswM7gRiIkX5oEIGaXCC3U
7tgx5FG4NBOqYgpeNMfh+D0dIbFEWSGMJBfIYr5HEQRkWN5RVA7XuthTyESmh9P6
ltFxA0vLezoTnKlpCqPHohPfsxUL882D/fZ59yqRXIG4DPh7T0+VnnQHPICu4OJR
QiwLzMunpFJM/Q5MTM5I1JzcYIzboAQPZFmDVUh02W9VwdoHepW3wm1AJVofdZ95
0xqPZUCJl0Jy09Le9JvNVq3dWfHLnDhuzwVJE2c3l5oOAP6DCLtdFqurpTgOBTUr
geWtJq+fe43PJP6P1FGJg6bXjc+ATK33gTXgwU1dSqBWk1DWWy7a0q/wpXLEtfub
Cvsd5ku5UKwJCb3JWhreSehXhwuOi+EglUi9uOSqLLahDqyM1jCNnxu7CIYmeeo5
eovtBdxyVpBsCLj8J63BE5kMfK8ysvGXt9KNRrO8BQXNtA9recL2UDziU562H7Yt
ChYDo1V9BLU1BPPIcB8H+0Q42vzOFZzThVNLf5DRROoCYE1okgjfC8SxwBK1bGgC
3VC//ZkjSSPtCi1ZNNarA+aGJNaXUD2QmDEKALCa3Bi0/RUqO9EGyPRxiSjO8HMn
HwX5tPHpOfM0nKTDUkn5dgE8ii62fH1r+g/s8ilIQ9u697+j0VPau2jEgrlktAQc
XHu3nnNKr+NArDfspl79FTRkWTmUhnsB3c57uGxXyFLshgQkDF/Uj0nWX5V89d7+
rqYqo/GTX08Zj3xn1Q9xp6C7qd2YJ5d28GJ/ThgTU6GDU3cKgnn7Dql4JBFOSmyP
4mw1I3Xuzy0tO4uuA0lnYOJqViGxJFa4sHL35iRldTyr1TT6u8dUoyBlqTYrG/r8
G0bcqkOLU0nTRGukuq92Y6NuFSZU8Oak+4Np1QRLLKvtHGwYBl4xH6P7uDsdRqLX
l+AFnfBpwnvYmJX63W6+5L2a2+QCIpVneYhzcYALyiwtP9fTxeMK/z7pNnGydca8
zLeacEE53xAJ4v9NXDvt6TgBzGVsh16u5k9+Hmk+mY25eBd4HsmTE7drh4sA/S2j
YSzYaSutc9x+tNRmxmKXFvNNJEuPL73RAo1ZY62GStmgICOjb14P1gVnXBAzCztp
cUKywifcFamflcXzVqOiDxlh+YQrd7qT3qFsMoxBCLmHjcIQqu/YxyzlyJmjEnd5
k69qPxdwyONIrrjcszWN4cFIjKGFT/nften1i/l8QGyR6cUwy8YlV5Mivl7mTFyq
6PEb5lau8XWGB/lpfHIu9kymECCnazafg1JY+6DqJe1/Hw6v1xb0kSy/fCwyJL6X
OWfQWOWAa7B6ub1LXxGObxUIKorpvkEdJi/R+hCIHWNPXvWcipzEjJ2hUqJCgt//
I7X43wpe8/rWNwGgOwWzBbmBfKk+rJZIzh1Xtm1LdnCXUBsKyOH16ZCBiUE5NhRL
dlqKmPLIWQ4jPP3DpeGMu1ToDLN0kdLNwkXWmALwU4Dv3NDVzeL+rv0OmzAOR1TI
XRwsv7puq4Qq4/auTqw4S7j7LeLoStZi0cml6JZO5hcDA89qNU1XrfaYQg0MXsUD
6JZjTTszK+bC95sXX/d01T0qAvWmpahtHpcmxQtxwrbU8J1pvbMRTZkzbzPQ2TrF
XlqEajO7n1/w52oJ9iXn0b9ZuhgneyUBU2Yw0vNaPLYMZwBP3GZ+3hIUCA2EBM9H
pNt8YGS5ibeobaVrj9gH/X0V9qRrLbTgT3GVM3ZPlC3hvkvL4kozwAaLhIueDc4p
J8Ns/14t4+zWQs0Z21cfWyvaPl14s10988VXLIIQyCZGXRQULVLau7f3B9EIACv1
j/lafLxHJsVMIq24AOKSq3SHxDHi9TCeFTyOwV5jqUwoV7TLJSgkjGzfxUYea4AZ
zamHro1kkwkVpHhVJqKXJiegZxEuoQlXa5jvEGIeJNnj7SsaG6oA9HdZg4fQott+
YiydKUE+4K3SsunBHt/KK7HOkbUI229/RFG+9O5cULjnMq8CMP4KRUJ3jPPrkvUb
KselZpgdtRJvhez9GVD+rvjmnpmUBFqNsS+ynOTD7Fy1AsKO/cPHJhm94kjEihbZ
OYD7YtBSRy1SDt8QHTD+/TQ/UOPSj0oquUgItMTDK877GFd2CarRd1eX1zg7PfQf
neJmSxC8rDo4AcpT2QZnh0NBQJaTVrhRpNtk2eJX5yg4pUwlv29MC7kQagW4mw2v
LvAevl3I/+8ldSFjIPIG6pLRNxMw9H0TYpdIkf+Ln62J5lJbVf10ejkmWmtd7L84
BHmOR1RfSNwD2CXFWNibSXIbgmgQN2ekp8fQOeqU+jMoKrknS2Ly3ML3KttUO7ua
O8f5tQXreRp2OhOdHNaoP4g8L4vmKkmtxR9O/oKEEU1uXzh4RzJx5AZ6Q+Ro4g9x
Au2E0fF6mF4FLxWBy+ZsBR3UqRo9P8dFzMr3gPaou6xKMD4EBzNl3rNTu36S6MLU
t706Acvs+d2SsrPphCFdDYhCUl+12rh0obZScYIcSjIPkuHX8Snka5g0wEwHYvvd
EmuJnQ35n/2B4pguzSCLKQVfp35S8yivTXPKwaGGYpyZulRBUA13OdiKRc/ze15S
8/pRB6wycqqQFkEmy0nYIuwMMTGnC/XBDNM9zRhCzA7hR9tVLeYJFHgz3pKJDR6x
lBWylX0vJxnyqAqAqUzeoEb7VgQIHj9fnjXdnHu7TwsE+u9uWc0QLusuu2bqcIbJ
sGm6TtpCPS3OIuZsQXyfZtndTx0befOx3s52F3hF6l9F3ZqEZOGa0Xv5k06YkwzU
rsDiNsc1mWyXmm+YNDJrX7r9wunyB2iQA35GMJiomCCBZRz8ZHKmx5uimjP8I+yt
oLkixJEXztZI34x+5hszft7DjKLOdujlTZR7Nuu5ryoY0C/2nNdmaHEVDQcm0GR8
JbLMAcLHZbFULt1H1NjFoiWuUuKsN/zmHQqd5NlZ49f84GkcHuTqmRkWNyY/Eh1a
fJ8C1JyKTHUgunoEB0dRQtjnf8lOv3pSTIFBg9drxwPTxYKg0O/TbG77lXS/SxF0
fSd2o0joJPYfAitT0oHX4qH74eYHO3VZLbQpUBS8Hop+IE2W7TJNbFBBus7Cja8+
FXY7VYfyuSgCQrXCNHUenoLQwOiT1GCdvcbhs4gT8At9IGGfWxS2qBgTrZhOg0Sk
f1/GNeMsxQHXOQUs4yk9Tl8OBSEyKjAsgbwS5LcKI7cTdAGQ7T+Ih7djnuXotslV
9QTZbeaGEqly0nEAYlP1lsZ/hz+CjButeoBLRSh3qquPycjsjT5ZOH2Yduol9LxQ
`pragma protect end_protected
