// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:01 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KUs5lyrt2NgopE6GEHwYq+nxXUQEj/Thuvk7kIW7ZPGvBYeakflK6XImqDZd6rIU
Le35kM1pkcscR7rzuscHtUBBPzqysX6D90W6ywfL7MXKbz4zG/Jt7zNEPshhGCV9
y4dKiXD1bpUjCbVJb5scNBGfPFqwvgwtxjkEKkBHBQ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16752)
BgZXmfEM8X6gw8Vkg80Ht2SiiZomk4cVT6B5rSQaSlo5ix9KQAncQ4zTx9ygnC7c
xMALh0U5JWFFRTRWnBaL1H7tLrn72vLcglC7vEH0j+mvrOGnRgtlFMvUbudiyYTX
cx+4INqhH/VM7ZCV4NRK3SXyktXeqoJrLU2T0SncGlez9bXPSXmWciF2gKR6Mnqc
q/wA5y9tDzxBytdSXQakgeSoyBeQHkd3Co45FrKNvs/PV15qApPyaB0g2MG6IKyY
sRHO61OvcxGCN0F5HUfLQB6WGyzbUOAIB9e90KjH/b2tKcFmJSMA9cOY6PNWyqMd
4V1K7Go913/1qFG5VwrulfGPZuTAVqRc60jg6JxGOkKbr9+DV8cM5qG99K0bkvGz
FuruVD40SK//nwgEm5Odj6XKN3O7NFpkK6Uv6kE6xORQtelN9A+dAUOPs+Z8ipd3
YO/vgNEU/sRhfuNTmawoa5GZhg9od/UOPz0JwhjoMD+3CVcR3DT+Eaz13dJllkjl
fKRViRnG4OeLPvKwE9Q5mU/2gAEuGvQbPsH3XogMpbGn3DO94/AKcL808TC2w+lc
2tSmBj5TbHuaqiB7unF6W4+SQ5GyH6kSilv7nVUVuxIoNSDgATv2M9hsgPm+SmDc
QljLjhwMXfjBR6RMNkK3i48FGndaMrjd2NdmLXqqYp9vgwSOrQq3rRoomu7S/Ixa
0I/JUXJoqnBrNqoJPvNzu83MiEyF7/L8UITdYv+fMWLagP2t5VHW9QEj3oiXvvnI
krt2QIBm1nlC2xtuJKxA3HJgWMD8v1JUQzsCAm90np8AQcvB0gnBBKkbTGYTdYek
loNkJMZw7O0llBc5moqhpPRua4cApNlvtRPezAvttee3ppEsqgXyn9R58CzgYXjU
q0AMVgoFXQx053kAQrmM3hzIjOonXaGrXOWvO6CLBvHEIWXh9xP7m7hC/o4705dc
rXXNCj7+2JA5oZY8u8pq1xKbegyaqMVtDuwxwATecH0tExC0/RY6y1VHfvwjgtpS
tJAH8L5CH/jnZVIYTBUmznfkKwms05Nb7oPEe5Wvmn4Lko4t3FR2wGLVs4cL2CEW
yS9PpnwIDBZHc63wsMVFYj89ZEXqavz/ZtvrIcL5LztxRBEum411W4G62q1TQFA/
9zp3OObekPPvho6p0gAIt0+uDt0OByCXDMgzG1KJbEFQgxcve1DiTP+gIXQbm+BJ
RzPMfLUtFR8aJnvqg4RmrdJo81F3X0CEVTAv3b6MzWARiwb9/BIFgEnsbQG7NH5D
r+868uM00O99pkRhntBwYUpWKEmn7MAMJvfJdLRT4U5NLbRZ45/XFW9gegpebLeO
33nZspMuF6A7KN6qdSrxHxO5dQEkCCHeucDZkgu1iTM+yNV61KkrLvOvoVPte+qw
8WDJgAJsrZ4Ws47LtrhJfM/bOlL4LiBHW7/adRzH49kcRoqxfWp3RziWZHHzmO6Y
X0dBWJVDZHfABPb7rIRUuBWGSEydLCr3c7wPmBAgQ6j17+1F3/NZ6Ykudusn265i
Rj56PpVr7JSwVquPgp4tY4hQMcEu27THtQXqUJCCE9Dzkcg9lj2OudZoZ9qC1Rk5
GCZFzZlfJ2Rbf6cKHZFk9q9c1BoY8TCe8FfYVBJb2D1HMLhuxoEfHnhq54Gn6rUY
EiLqhnRMlaOETmhVz4cN3bzCxWuAqBAQ3WO5ERIFOGMQugfhZsm2XHASBgWc+2HZ
+c+ZRyduJ9vnZXmhz8p5ov3JIaUAgZlt8JaCE48Po+1r2GbNadIUNRYUvN02oFdv
GLu1N4B8L9X0nmJtjIq1h8JN8oqmDey/nv88tqRcUkOztSIkrl/byvxSQM85aXZy
CglRGBqOj4nphbdvEDUnFJzg9bugKVSVoP3cgL3RQ1BIAx7/6EsgTtE7ERbkJXvm
SpkwBlOtrdhgOGJ1U8KlOiXHEHxA6vmyGGV9fTr626SNxpSASyeFCHoMZaHl9+s/
Magz16leXkOtutBJ26907UjJgml3xDEEuAW8v1OWfFakS9Q6T/miOZi7gm7MF/TI
NJ/Yj3wP0P/PUQSAvyUyAhr/aXI3FCTHlt4oGR+DwcAgvyhtc8lA9ljowew9ilzq
KjKkXPoNQ8vFWi5/LvyDAkmdyyUVetHcJVhofreGYmR2p1FiqYMkRvxXgDX50GqO
EwOfL1zh4KwPGIx7K/Pb4YdcdnFFgZmA915X8/doYSv6TeB3oTI/EftjS+KKg8K2
qjreVs+Smf8PKwZXz0Z1B+Z2FHbigg709JBhY/W2s8AjCm8G8nwQsS97LF6QNqBO
o4OTE0tAV76AndMsyrr4SplPysouXHQW2rp18z7bOysnFXwMckcJ2lLnygnvLklp
nA50ZSim3oI96kuUpKezFZ2whARtWPimvX/Fki+Inhps9SMaX9NekxrN45QwBXky
Nffp/31eewksEBuBb8yLdyQTbvo6JjWsobMVm85gK1XcLFmnTnjroDpvCFhrMwr7
OZ5e6rYtGkeOBFzOE7WEb6FjF4a9VwnUhV+0xkaGcsHJ88jhFe+nt0+wqvXZNmn1
HAczv5hJfwiUtAZURTJR5DQ0zqBmtIFT/FFX+LsU3J/yGGJZBFbOteFpF4Yjn9C/
XtnRi41cvkLsOgziOEslmCPal9LJPHqTIfJnHSy+3pfunrZA1Pj88aTT9jFH3Dmc
wqDguyOdbSgFSZIttRGjk/g1BsxO2o7191+OZB7sUG/HwNoTEfwOSn1eHFE4rwcn
82hwbfKQQpk9qwf42WZy4qLUM7oOzeBcWwNFBxtawOZnFBCTkca7Xd+lD/wCl36H
7ZMPvuW1AVZyHUIbbU1qbh7WoAy1auxMiQdmaGP8+lQQnCKTbQTmyekjqDqErVJe
2qQ9BFCdzb0pYJuTE+61yHi5fYhbBSIoQbg/IZazlZOdzPWQRVY3hBZ3xHSriERL
FZSWN4PxW5jsbUqhn/oYInJZNKn3kngBgvYk+2eWmnob+SeTdFpWRn2WO+uyaDDs
FjAlc+vK/ECYQVcMzBPPRZ0Jx4Om9JXjpQR5IgdElc49oJNFt4qIbJJXS4fuCphD
dgFZdETWX9p4jl0Iwm8iQKQdpL+3KAGYiLkvpagE2WULabbBxczEhFLBWbUpAqGS
wEFg0NUwbDfgi2kHZJe7FKOCOFiKvLLRdkhSbmNa0dkSt+FVhfacMpqu+ZDtAAsZ
pCnUYPzRE8iFtN0A6H/1Fpon/f3NCbfbmi3up2x9RplOe+HTqmV74IWWei+uF1la
PB6cDgWv0M2XctQHoDf1nSguvrxGgrP1eQB7082G/z1EDXulGoqD1TYl1su4Ip4L
XIofnCMZsfHv9l3VJoWugwLSnFlPxaR+xXniJZQusXXuvSnfZQ7qliZYyihDXWkq
1FuFt5jX59kqA8KCy+pJUHWEEjuSu0IihO0J269vXoJI9htFHlLFUZ4BSrJhUvMZ
Fz/Pva1xvbhetepOa/eEXimDjF+dhj29dGNs0TePXSufjX27zKqidjCF38x12d9Y
mNgcANkJ9e8D2tO/2Wml8vhiX/+vDytNoHGZrb2cAeGvtEQz5K4EYF6bAtccfi/V
+HchVVAoUrF248sHaRF1pMFwsFjfvPTwcDpbwNbd/GMjvwjJpWH1SgNdGDuq9lXh
4JxF3584w8F9OafLhmEC2S+N77G8sBXQ5o6d8crOzgJlGUN5jSb0Bysty3mr5ojR
MdRs4gjCU5XIH1nn3yyhbns9EB4emX0X1tsmzXRJQ5bZowAvXQv2TjNQ/jIS9zDJ
BSEKHVy00xyuJy0pdjghlGI/8p6TlzcmaDwZxW/DJSa9JXV6ErYg7fQtkgI6lO0u
AfuATUTSbxxuuMa2hHmfuA+k47kEJRKBirL4N7ebQct5ORH0xnZZO3YZtjzikJxS
dWhVUuOWtWZ14OXiHW2QN1Bc9pC5TjYep7lji9o4Tz82qBmZWpiQw88KBRgpYCU5
FL5Re7BApqOk56lfFkuLLS5xlQwDLGDq2YJre/YSn7o/2SkGJASWeiSGv8DsWrgf
6oklE1dpV6ggmIFEYMXLJrD7VE2d+M02MwTf6PuLlFHXW3vxB3OkYMsRZyrme58X
ZMYBCp6bfVGVhWnCW2UdIxmc82mVI5yIE2n/FK1pCpq0wU/YO8YuYKEWzfGg2PnX
S0QAm2hw4j72Fx7j3uoYvlmsF/XtX7OjPYz0RI4sE6MpT4UGH72bEjzd6LrsDQvE
vuc0B3hLzt0DrqS73ECCeCUQFPJp9Cwx89QQ7M1tlnnisf7t1Bnw7R1XkiBmGK0I
D9UCrPTh+TWyUV6YwurO/DpoTjJgVxNipCy3UYkXLuMVazCxWw4M76Z9KHWa//e+
ZBT9W8TSUL0AdFnlZeJ9GIMdohRkd2o9X65kg2p3nI4CSDVoNuX23v6OezxSX16r
QPGK4G0j7wM9C7EvDPZxhwMpJRNNpuizhkA5akiT4SqIM95i+/e2pfcEMb7fzmr3
ejuSkdRuT+MfFRucD5l5wWoKYDhcAFkj8in45tW4LF2gXHKaXFjWowGKzeQThW7j
s6o2/L0pyNswMivE5rppgkhbK34ODEWAoB8b1GhFKTG/hhLkApKX3YX8taW4vhdM
domrwG/f9pCk2yB8/WuGbkELspUaXMzG23J5LnW4ypIKIHoZ7VghHjmFUKqgNKIr
9riEyQZteO6epfPmcniSIUt7HHtwkUqmu+Z8me+FX2G4peryrhfZTHOlITtCNY+/
CgS15I1hY4gwmPLdQnjsFaqXwtG8WENZV5YIsv2MDsgozznDkm2Q7ms6DR1x5Q2v
JMk7DkxvFaD2J4bMWkKZy91FjxvvIjo1oVJS+LzCeyV70/cSU+XKM3ytB2N4tJdJ
s9TIgfv+tzOSdnPUfejv/yqDS925titQ09eZ4jyrz8wvD8S8ZmsyhKymBftet/La
GxVf/5QGgCug80OKPKfvER4QRAsnIsPcHAc5FtTEeZf4jp4za8AhcF/vE6Mv7ZpI
3MKfwl/cGus37Klj3GXhIRTzfQoFQkIgGCNNYQJAHBXLwPJO7m+lfIh39RmlYYxE
fROC2/BHfo5KmNxgryrjHmOiG58Yk57VoSvWQkm1sXqpv+WHRSLiczGbHMLtRSZW
o90HKn0h7jVtlTCx1IoYYtJTcOnlks05JIhYnTR5qmwSs4/Oy2TV3mKGvUXbLV/3
K1TSUp8t5DGo85UsIoZW6Up0QqrlmmngSLiLkXO1beh9wrHq43EKkUQQKxQxq6pA
CU9MAIlaEcDATiNmGxrBw5li06uxsAxOSPmvlYIjg2rIHEVooJ2hc8CTyCMFnmTO
rIzh6QV7cHH4kw8XBM2kKBUUX83wc3dH1C3HTutDgjmh8OOFkQjA3j1EBNdfjIB0
HtzRFdITa2gu8TaQ9xF0wtarxrqtSvTNWwtYPE0rRChyxG3fA+gmy/MoK2cFzhOB
sa0QAykB8JH611BNGtTqYXR58zvmw0P3dDKsbp6BY91BM/4Jdl8x4Ikm6McDLGEN
zJ9RDkOVipMHKOvJuOZEDPBtfjlzgXDf9rKlvh4ZD4He30NV7FLNTGUJEVddjAJ3
PrRyDOcQlWgMVovlKQ5aYUCd7cE+cfMArfyoUFqhcbWLR8LtSqKL2FPUONYhy8M4
qNJEcBpG4ioa9uft+ZYMF2XNZhENdW9KiPBX91GY46H9M0aARJjciV5lZu9SI29J
B/Ibt1acCuahiAik+sbvCQuf+Iv6QX9osqMe6NO7j3yMHbxIlVN3eBiJQPvQ8r/0
lkwd3F6PLmG3slox+TWqbrX+PzEhEyd7oc+sti/jABBmH+G6X7nA6hBr0uQT0+a4
koupUTHZzsJoKNosQJkmD6+JAa69fY3PLFB426yVmxXlJ/BPSV5JgIsTAbhkzieH
L3xCittzTWad/ZpWQfSDJqlxjdTojTyfQcMVDQXtIntnHoiEbwQVQ++NyEu2OIOg
mDOPEZI0/WLVV9VSMTu8vuHUyy63cqvSKTYlZBf0D70INhSuQILYMnl0T8mXkWuV
ztZL9d0I+K+vGTcvBiaroE5AWCSBYDNEO0EiMHsfPWjPjLSKcC8iDUBsiyCekCsq
c6+Z9CZ+TnRbJdCAO1eq/Jo6aWFN7melFk4EYTUNIYEieuhhOwcjYTqePwIlRJi1
Yxw5TwGtRKtLJGaTJv1G+tGCEc7HJF2Sh+F4YBtO03cKr6jpc1Fapks/Cy7gejX/
lZo9OnYJDzJ3BzWvdp7Mpf7BrXTMghFB+v86OAaJERnMHwS79zm6R1FFnts9U9VP
cRLNPOcEWVRTo8xMF/5UCTsIve8T2e9xsY7BvDKpRa2KOCnQ4K6ogYlbva5WZemo
NqnFtZVEyokqqK+17pzoVjpAfgzPCST/tvsGxbzhiwP+TKVt+Bn6JDW4KTflOOUJ
1LuUvMyNa6+qvbLs0+PkbyIa+jpTyOph3DRgxfZXn/+op2w6sQr/aGKOKlZyXywF
S47mpn0eLHAK7Eol+atZAU6hTluyjAqIxuD1yrEJh3oNhPCuLdeNtppryEs8YOe5
YABFrz7XtLRpt4QhNjS8miMVxoAdZvo9StDtZ8VUKLLb/QGPB31dfbjlk7yfzUc0
jWzkaeRz4Ex5JWxsEJ5xwSCzlLXeqzZFpSz/AdbsoeHCy0G4RkEpWDe7E1DacVYd
Xfj1rg7pO6zDRa5QKQaMmOm5N6s058LAt1zL5xXIMMcugukfW+IPyMR4X+mjZNP6
lbtk04WUq2M/b8e9v7Isz1d73yGnX+bTrdHC5h3nywSqHdbTjKmZHAx5m3mTsDFs
XZLSqAxFjVc1lJ+SH8wl+rh704teubbx6tEfPqaG5rTiLcMuemuo/mnaljPQjD0c
BudirvVmYtPl2GHL1OzUcP75IeiH44dhcSINYHobhaFXjtqm+UDFCRVn+7ALAkTf
Gx5jEzLA0irL9z6qixR1DkMxmqOntejmfF1Aw8BGawIexkk4RBMHeuzUjbyJEWdz
uVLl/RoV9ZdgAkviRkbVDdIiPDgPl6mXk/0nH7Qmw1GjsvUWQt/WVdl+2Xy+FhQJ
FbjynozQEYKoRiPDSkp9WmRIuZepBeWchjFS8PnRNFG/JU5FXzGQuiEnKhrJ6Rde
CsTYQzajT9N6pZn8aDnR4VOHHouC9VLc8uQNPw1aj1loVdnEIakeAmrnpyK8iQgd
pYGgWdiURddgx/zuntdEBljW+md+D0Ld+9tQm2LVupXO+rN4pkEBTOrLhh1F9nQ7
W9ZQIwAzD0A4E5QaVTxWEzTq2lRw9WxfMaFCWreQEgTsIpex6pGtY5pmj6XhUaXz
TpQdzKp2yNpdE452PjumJZ3xkTZ/Ug5qrCXhrmSIqBhSrOKcYql5/sQ+QRI36IdY
RJDNL9LwCN7yBcQUXJW5GSHgZu3ASqLXcAPW0X8ffB7fLE0fVUcgdyXyghuTiHA6
bAGDzippvwjuzzQ5OsJ+IdhBMp3bWxSi7RIJktHNTN/M8HzeEHA4vrAC5wu/GtLk
44mqSLz/wMNL9nI2G8Vw37isTXMA4VyrQ6BLEi+++Qzp7Z5KIzPiu2yYY9aWgui7
QQmkvP+/n+qoImBmCwG/x2Ei4lLY3TQtLPTCxB2nXVOEdx3+E64JCgpsrZ7EmYgN
GX574+UtBAvS0N2ynjWvQlrKQbGatNRo0R5RhkXdfsYA/bxksEg5Y37rPB2T7Uf5
OXiPNXuHSGxuuoyvEB9y1BwbRBcAxJBa4gXOW2ztcxr5jxnDEoqND07gBaVPQfl4
7XRuzC8aBL7CsaTKz1zq2572lT3oCDIv6yLCR9670+wFoZbcgImtRBBoP27SWp8A
KJV2defTQab2J/R111veXaCp8ZItAp3Zp/FYztTq+3vyKD2PN5hd8te8bPEeGLV8
TmkhRaW21LUtes5gr1y56qT/XiR2IlsE+AOqJ4kTQ/B4oDRu9tS9mB8Z3VCWAYvY
PH/WAaSmpuPFTGLraYC+3+n+VzXfFPe1VwiKdOO3m/HNcSau8DxJLHGe0McvQrpf
i5vJ4bZLbAdKwrkc/SyFmYSU+GAMC3Ps/ilSpSWaeGOzW4A6W0xQJWb8+B6u3d1Y
xt/ZnVB1l8kfcEJO4R1TOd+noEWihmSkt+XEJvU8x1TjFbSCqsx5GnT0OxgpCuCM
GqDZPfBfksE4CoYxkmNLBR+XT+s+35qDdxngQpnbwa1T3gE6CWgu1xDHHR9kz7OF
kt9fsaKiQuHfX2pQgfoIsP/N7K2UFPh9wnR+jRlL4aTJBjEuegBBnOCUJCfRMd8n
ojOWuYEeGVsqpAb17vcaM9+OnR0PXbQCEMLXsaHvd7OV6y78/c0qvB2LIt25YbNB
aX3KLja1my4CahOZylcWAIk9itJMyEEe22d0i6LdDvCrSZvzfGd6DA4kgTUFCS7r
Z9DzdlqPPfH63LiXyGGXFJ8xnC0+J/P+AqYXa47CMpN6fL9W/vhhU920dHrVl9zn
xaHX5inVcqo5Q1OD1xmViBRm2L3i/zrX3RAC8N0lpDzmQcWkeLz/lMEtQDQyQlHb
zUe76/sy2ntlExcIuCgeI69zLcn6UBkMR5BhiNicoQfFUbP5BZcOyl1pz4jCBei1
xsnUN2GXx8RQyl51LkxzzEN1a9ejawaPBZXqS18/gTL176lbqORMFPgW+M8zmqf8
Otmn11YDTSU9Kb/34BzpUpI9hvWw1AyEh3p75EKYYDKgrZ+0yYThglMOwdQBYFgw
j7Otpku0Du2tv0nQVMuKJ75b9Qe4Y8kY04Lkh0835GCm/1ZKxpigL9E5rGmTcxeQ
NEiQa0cg2E7cQR2ZuWgI24LrUu4lEe2uvtfxaY80wYgXCsLZDos4FBokcTIOqq0g
sw9twj0tJi3KxNJFpInh0AKvtQegaDMdBMwmyhBc4C0K/BEOCHK0R7rF9Rzw+8kV
00v1bL138hF4rsgx+tdBxAhhmITsvA1jk/q7MWscM4JJO1qf/XYXidGRu8eX5Z5/
YdVwBhbf3qR7wvYKbHDAI+iIyPUfR8veSGD7BIfQKINWdExxhIxW0J0NX3AtjWD2
hRi8x7CKMfzRoW/vkGGBNrZRh7nr7Kwje+3g2+7yJVqtFs+6aQlG4x9HKroPmpca
F8VTzd+0AyRtsq8uYYkRwtUb75FedPSS3PiG4KZUC96jV3g1EqsDtqyCPs7KcvTB
Bo51cAm1/CR/PlBgffY9Mw3hivinNUDQvgYdXdq63b+GtNXtiEDimuUtIWY/LnG+
ar5BnuNzCa1ICL/cimsO8Yl9z2NaDDwhnGABq+ff9Tjy+IIbPT4ckEAhc120Vg6n
r3PQv2Gn5RIDfDG5Q18ckAM4TmFSwtHBsE6yeoxU7tEk7O3h5hV+GyXMk+FYtjth
FDGGgYxtcOSD26orlgs2ADHCEx9Gmnpxc7tDqoKu6fnoSyxJP6kpygj+emReAoKm
t+/gwPoeq4ZB3oGtvCJeOQMQZ/rDBrnldoOu8hAcn/PDEdPVF8V9KQKW93QkgpdW
FfU+N5B2vqd21HOpUUuTWbqPAB+ZAifazIUOqd+NSgr8U1X4gXUejRuZPSHDgYB1
qCKI6s/TjsUPcDQ4ZCZdgTnF5ZkChZXHu/6KEiWOkPB/cEiMavGPu6lprsn8jFIF
JYNegOzzv+5wYmCdXASo7sMhOcHRvgmW0VSKEJ+q6jBM8ZxkVuthMbSTT8JJ09Jc
1ozgMHbAlMH6dr+BDYpK5tJlkFGMJIVPOcHFcSAJG82Hr8M5URnDsafZozgPdCpd
HvxYYnblPuDp/iRSrW4r6lJ354ff9ghKK2eUHr3uCsZNW/NCpOCO3DAFPs0njdn7
ze79wuoRRN9ePgLjfNplM8Phew5Va7Scfh5wZNMOxq3nUPnwzcT9WSDMl7G9JBww
rorZLiOS34mHLm4u4nYGaXogfyrnvcjD7tV7GQR8imBpXjmu9VJSH4ya9Tz7AuYc
39LNRw6kW+TIGAqM9eFscmzb/WanG76zFUdVGJ4dtd0mOnMuChlCy4jOSFsgkpdM
ZkbZ2Vz8IDpHq99f/5i9hLYLgLMJaMVMui7gU2OqCHxYWr/AFhRND/aQoyvfNCMS
JAJnrqM1CpqrtN2UwzVMFEsJuW84GeipOrgXIw5zL8yyQFYEEgpLWS3qlM+r50rl
5eK49SgQORARIqquOwbL/DhKDCaXG3baWLm5I23KhHuzeF3AyFiI+nWG1q/l3vjv
9Bl9AkGjcUVPq0f8WEDjIbnedSq1ZFevQzXyV1qOkMRw8YvK+L6dPUDtFofYrlVC
6l98QYXwwqKkB5MBdvCJQ8r9vX2ZlHlnHNLz7OyuZpWctv7qKHFB10exwmhTs7R9
aidGY7AoormmSW7JrQVVLDEeTWdIQ/ews4iTZZR+9FJ9qSPQcQHDqScB7/ddWXM3
Kpr0nRRr5qz8ubgpCjceSk2AvicqeXWCEK4uXFNeICDzhN0WdlhVO0kbyCP4gPNx
/CXjJ3n3nz8hO0oI+hdHOuJ2cm1YRpXH+qopER1easnMethmwJJRPJVOhHUKDInv
kD33jPPAb3LY15hCi1AwD1SJyA3g22xZ98uujv2Hn71Jx//G8v9Oor7ZhjXY5o/j
kf4B3oxzeXbpxmhlouCIFTvYXe/vgm/D5tn2w8xKa1R+mhdlRNOyllJ6hgbzJjTN
q9qflwUeeewr9+e+9oPGZafLu2Cdm0/6ZgaFg2rWatKStg6rnWltbhtiU5QVjZ0F
/hqSzSlFZtHQfc8WSSmaxut1cFiqv4YuSYqtFXC81s1u0GIX6IDTqiTfNI0Vh+3u
bjguXA6ieLumRBvZkCouYaotD9v8M7Qlplplut0PZu63wvYjQU9E+FMVATxoKoAx
JNq4dA3jNRp0H1gmAZMqu9pJxoYjU8vekyIuUeaAvngZT/aipITPujmN6+PsbdaW
tD1/3qR0LNtYLvojPSe3dy+FdvdDOGvIVCcCpDcPdsaJXAKs5BHGU3/IVAYFUDQn
8V1WjMamAgG9YzV4ttnbKyRhE2IW2i2Ua6QvXHa4S1Znj7L5ge5yMUFQntcwpCOn
saPQFBVFVP/EPAZ9GefQmqFvtyXOQePfyzKOSxHy5Xxc8FszMY/Zs5lASC7e5I50
AbA+rNdO2rknHqLojta9CC2U8HhQOhEyF5OyBeTE1eTolugFonB1P1gKrRoBAxKn
irNwN4XmvEKdPVvHXJ3Cqut+jEzkqVXmCNqvY11ERQAouwOr3i54t7GXZN1KhyB0
XSKzlUkna9O1HqG2lDyrJLXS2EnI6vTlb9UaPGYWOFM3wOwNeB1h1sdge3D8mwUl
WCc6q4SnfibvHt5d4co3XS7mLw43UtIA8v8oshiFQtoz0dGmcBqmvOisGtlSABoz
UZAk2lEdrGEJNe5zqZWbRfv4zGX19iWsZuFF0B+L6eUM1XTDaUwgpv61k96UoPgw
V55+m3+odrcBjPNrl7qkv4Scvc4zkW8iuYihsgjKkyvV2i198YOKj1Ou4KNIvY/2
deRgJjqTZwkUdO3Pn3EGDkZqwNR4Q38bs7BwxQ0mX9PvIje8Uk1L3yF6SdQG8H8r
3Jt0tbcLydT0sSwYc41VKT4McMB7Sl+uddardFCXLiJIZog2sreokHIUnmn0s4T9
BOP6pBtelttF5NBBySs1nO7Wke30oW3tLMeVtXEut63hE/qCDxYu0jDsnRvvUqHX
P//dKlbJ06nu53+aBYNnfn9EBx7t6xjrtBhVVl6tWLLdDoTCdWpZam75liNoELvx
qRiW+tQhdRaaeyM36Y3hTIU7692o+Up5Ucq8hLHZPkvIiFP5BmDVfoYNGFm5jwiA
M+XsVkSMABxdffahxTW5tfGN3RustpUj2+DjCQ/6wswYX7hZrpokf/V/XSOXRrWK
rH4Zv8yY7KRLYSyMB41kqOIz8BV8+5QkPslTh0t7HnBwriQ6voJUey2vlLwUlpxh
3QmXxQK3ILnl8IUu1oICuyPTMY+2a1umpNDcQDb7rurQTRAKfbIUhaFprsbXvn36
ndNLUm57odZE2A4+JZVqfO+tv8cceQiOfjHV5G2ZiJv1g6M1FIm77d9k3HCHOZHe
2PdgE3TXMTVkDmQX4e/69gYVBwfVNAnBPx9df0jv6FzPx9qVkLIfeYofvzGFImpH
lONDmf0IgskC2A0wXUP+8LZSCU1JlWeYwS/cWfGTIOnxv37iLTt+MAzftqBeqqhM
Vx8C5H2yusup6w19ouwfITZKq/Z1uSyGHG6SKjmTwPXp0g9JsXblwa8GChWi2VAf
K34vTNUpakmPX/cTEFxsxkeDVh4VJjAh58lAg7/2if6cLEOY4muvsc7JNyi76PoG
uLIO5/GDOy+d+373YrStj50IMcrVUiDr7HUYxM62jx6hD/jRSE1HltqZwjWq0GVN
EAuoHukro4VwVzbiatKIMC6yJySqPCIpq/gAxh+b86uanSaYtGpT5fxe5kRZRXqy
+ddXJQ7WVKw12l7gcW19ugD4dcnI7S1QovAS137sqJIcxsWeXz0U0d8VwgdFG0uP
4LTWcmhk42UuI7DZtBTj9XlZP1b1YTcuVy06SZSqxDevKobYOSt1DIPyQmLecMYH
d99/7FbJmJ58SLO+Blqo9A+XMvxkz5ic3F7SvWFK1DGb1H6vDpdmRVUa1K6gMNIo
ZadujKda0/fz9TdfAEljV/MMmFufZeou2RovL1G/5mhHr+qdNEe3cFtBw2cYadrT
YnYaAmgwz0MbRSiammUFhCJnOKnqzaZl/9uTqOKgXvL+NI9BoocKq70D31YBFxUN
MYdYwlHWIMfMUPTcAvtPyqHDrSO+j57sTViNkvMzXK7kj+kdZbRn5LZEOo77Tn7J
JrxhuhjMzVCibnfUKi/zWBG1/DLFtDJPNIp03Ldvemtp4VaA2ot4EwDvsjuw1IAJ
RHvBiU68I5fOsZlIzFkmqIP3IvUlfLwsk1E6/og8lvVypLAfeDzV5wVMK5SYNb9q
QOa37gPn64/RclgAm73Tvb5sbsm1CSk22+trATG29YlThupJsCaMPKN73CCxK1Nh
jj1fM1kR6oBKgIc+jyDltDvkW+a37Shh9HcdFS5z8/OKVpJ5yGnUdGcWdS+/hj1q
6mgnI9iwbQvcM46UujY0JlGsuPUQVroek9TY5VMjkv4AT/v3+/aRS7+nF/TM4Twa
mA7cnoRIbSifNTJY/EQYEjETO03zvTCJLCc9PhJaIZ5BnGTcH7tRgKQGVtVjQGN1
laHIanoFcQbe0wQj8fzYQ2FyZlZQVpc6Te3Lq1n+VdNg2CXqT7apWow7Uf88iwnv
AS6cMRzCb5jJtxKux3qFNj+CoH11nY5cprboXN3B3Nx7gameiWldqpEea97t/fAQ
tG9cxiKG4Ce088HSJWxszqBwCepxAQno7VIEJwm+SlNV/45UrbSfH9FpMoORFNYt
/mOjXxdtOPzodpVzwxFt8wyKEpdMcW5TyEHmKo0alZ2j2X2Sa4vXvGRBeS0QNqf+
vbKyRvH0QvqdaB5igHXrX3kQh5URpo6RNbDbUc/DNwpZCbdohhnqqXljjs2Rg7AQ
NYonGvZQfiJ+Y6Uw3l7cjep/Kscr72/LPTzsLxrdCqlCDWEWS3KPY0RM2AYMO2Ux
lWTq/cxVw4XsLXAJehNsYW+K3QSE/7mE9xkZrgjbhCZkIEItWxXmhlAJNF/Q1gPO
die/bgpQU7COXpBWZQJGrtw5YVUxIZW/f0sJ2IYPxfDhB2W2cCMPeAoin30mXoPG
BR+Xr/6rF4Xn1fkIFKnZCAJUHlbI2Ftzi6obGJeVMLJQG8KmvnPaEMdvrwbay5si
HDGA6Azw6dBkuFDpO1W7ARlMMv/W8bSuTreOOp9BOB2PWACvzems3xYBRabGC4MT
vKSUoCT0Y+SoVdfU72qMUg/Bqw2woOUBl5Ew4sSqGUOODSrFq0OyGGurQ1sWPIwN
6dckEQUmRnFhv1dmkbbwPOPhUnOi4/F7b+L2hZr1n1pkA6Bgjq2tOT00BvAJgggu
652E8L4SuJU4l1yszmTlGEXPOHb4ofCKLAq/7fIiyHRSI2DLzjhaOkymhQ9fLXX4
22FWN2/nGj8TKw1VGvN4b6VFDgvQtCEL/FYuPlSAB7OnB/sHI6THLuMQrrrLiC12
TEyROH7O5jEKQzF77bTqidTHdi8Bzc2DdnpBZqzyTlUvzGLwYaVU2P8kmLhwSAx9
LAJXc30fApZ9Z9rvq4awcqeKDdBwO609kTQchexHklWd9gtI1ODSqFwIG9Igx466
WSmdUDjrBs4WICHwzda0idi2GcXXQ26ssT83yspwTwH+n9NfYWqtJSvuecY8bj1g
CLjJ1gdOtlgIxIi6NKXFQcmz9mvskcgDwd+RDZMXCfTaI+0fSb+bzgbl9YxLTmmt
fS07V5/GkAE8La4YQP1amRksL0wsF3MFEIlKHzW2MFDrTIw9FC7Hz+DXSDPuzf6L
92XHEgpr9PTiKAnsTGQC4jXZoFiN/k88/NCgHhZ6GHRSfE/iMEhZptmDcjWqTVVY
teEtasmQto1/CnULEUfcqiaPGR8IL9gXKaHAy9RQH6AqH1oPAg62owMeI/6bCl6e
XtGxIDkgmNP1zwX6gEB3weOrh+tlgN4yNXoREqOZA7oDhWOp0qbX4bZEffnGfqgs
kvsGOguXpIAbgLcm22hr7GaHXFRRN9j7qWMxb5+vor23ccg8kphtcwxg+rJPQIc3
PBmDfmFZcnXPuwhydi/sw3u/P2UY3Y1JQaIPCK9hyKPPpP7rHIygTIoAeuUK9PGT
uc9Ro2oEiZ3ipc80YZhY9KBiTtPVWpBWORrUmf2iiizCHtF5/SWNw62A/KSUXr7I
RwK3I/X7+Get5hJbGCV3V1m3XOUvHYkXgRG98xFq8zAwa3oNAdvNJnBOzeVHanv+
Ao36kORwPy0MwKneA/0dfN8bkuHlccuHOLmjbsjNWULHIB6G7AH2z2QfecEZRnC/
JjTABCmXYhwXOVhBcRWtBNEHn+glP4A0Ozj4drR1dALZ1uumOBnvtjqt3rABwEPk
8voV2LWLfb2fBm3jdll19AzglFR79/9GDCQ63qvgS8sMmmJlcO5qKEw0hJMedt9o
Ose5n4VqVnu0P5lk8eezfubiXgL34ocbTDcCpWQb8dHkf9ffi37ZfpTejbCIruQ5
NX3pxJ0dLZtLaNvcPkEu8hVVF4csMRNsKBwBlfNkxnlOSdn3UZ+J9HWiw5QJAxyt
v8CURMrrK49cVu48aRNbgiUEypYfHXTeaNHfpNC1pxWMgV/405fcta7pITIh0d7s
Uabf14pEvPCzZCP3NttBo1GvqkfuMwD7ymW9UpN6619fln13aD1t6TkPUEQb1CFY
Uuu+jKwXGVXRW86xDGvr6B8rWVByZKCQvfYKIpZmTw6DnOvWwfl7G6hVflrze+Bi
OcnmWEtErWxUJ/LiMogEod+RmaS06Xaj9sNtSK3Xd6YwIkp0XTiPvDl/6vTKzZeO
kYmsF0PxCAKySRinVGczL6Im/bpSmkNLgtq+TjXDcFdzlwaTkCALsKDEX0QVXZkc
GDCIctC0+sDjRDb3tqesz8vuaxbthCJ6DmpKBfuFWVY7h4nd+Se0bUcUZkB3T+xW
SmqrARfOmMZQojwNtp0Tygh4qorij9/iEYvsLpGrpTZ3+x9b1oAlIPj1aLOT+O39
91pbi+O5E1Bkqoez1L+QjNOqDAWaMaCnlKCI7n68B1i48gNv8o3ai/5YxHwL8707
KlSY0R7VkhoK6oo5C8TVf93M5w6djyeptmlw4K8W/WLRt2OFlFbihYYwhDtXhj1h
3Br+FCHY++rPG34+RvmzRDhZCYAtY/RUBvH8ZHDvznTfb1UYo4I3lxAfXVctfww9
fSfcSK120LVk11LX7wSrvk1cGefTgW2BydQDrUT3XYuRNPnw+lN2BD3gK3Vj8IwI
JvqumJhSzADrUBjlLc+Q3FJ4mO8maLu9TOH53nKIpSagjzDy5eHNboOIkt9wkhG6
55Z/AxkYRzd9rYVOST/rFWZEuIviUp+6GlbnW11b9/BZrraG4ejhoIDeSY+aEjjS
usNF6cKuXw3dy45Ia+Pbwkir1CxVvArW9XOQSg6RXO+Ud/dNXq7kHuP3nda6aikr
lkbIKrrUdK373xKbe45+IhXky73Ej/TEZvAymLUG/YHZS5Xbqdkngy6Qm/mrJmqx
QrkV/mb0cj9eFRGmQd8L0aAfJR4Dy5KKSqTtxK7GDTaAIKkXw+c2WCIhuAfjdpPA
Mb3xGz8jyvxyWEQVrYfxM1RPylnNAoZ2gYoECVs5Gz44y3YYATUBQsH8L2sRnesZ
dWcgfu2rpEth7TBTQ/LtYABY/ATHLm7SGt3yzwzNm0BGV0DSyuEpCXHd156wK+Yp
AMDobK39GygWrW91PQt06T9jMA1Kva2Z+zHp5uhxbydFrDvDdovdfxf6BVtRm50r
/PhQhq2l3TJgAhTN2ohMRWD7uen0r5/Et3Ttm7px0iMAUmgiyxAJsbFFt08D+dJG
VuN/au0PTS7HzYNvbwo0vqL6AUirnZftTFSDWE+fLzEyFfTS5Ineyz6nE7bzVXEr
/85sLNX5RDHKrYjfDQ9FBUyl1LVv2jK1hEwvQIhNI7KFLw1IvUjLtFRVbHfTR5SS
XxbHJjxoG5ZJ0hNtdeLHXLUviXDpVzu00YM5898tHvXdFp2mFOcd+KjV9hBbgOyv
MlZ1U1QhhYoIQ0Ar2DY+r/T4sOBa9PWI6Dl7XMP7C/1cQSX/dPZN12AqmY6H44YF
NhJVSrSDXT8vfV1k2IziY3ydhpVf7J/YdCqwQsdLdGIr7zsXSCXJS2cirYKcWsuC
gJl7BtyFDY4tHnK5BZwiUvPUvoTmS3JUAYqMODlm11EVBN66dMWodxLD9ePsAk/y
IIatYNaCzMdpDxlcBtLDUHE+nqSCA5Ygx2sCD74mWWtliVznYmwXWwMtJla+UBtI
fHHK8lYR4eUhLdid6tk230GmJyWZBkuATJAfYjhruQU09FOMyZCUnaPUdqB62RYd
rp/mAJevcBjrglpNkiYLimAs/ExPkj8J2tv6fhTS1S/6Q5bOqeBE8U7nyKyHImHg
KwNdoUOo16DaFI2hiufWSviGj/j5HZ7J2Q8p7AQ4H6ckM2KxzgPrhIfmzx09h78U
h+JHvNbBQtzVEj1hMpjZnqQZsUJSjivegVSO1xJCYOUM7n25nvTUaVnNTpfklSgn
K/pqWaXxS8gQ6KYAqQyawBvAhGwJbClKed4NgVZOB15xt9ekvcvaoBPV9pgxnCwQ
7aovFqxU6ODG7FDjGtZKLLdHlDXVn1KhFQ5sohOIFrrs0wkmHjCydJh4jSWmQg2w
bbWvtibwoykf/urhr8DWXRaDMIXsHqnPkxu5IJXW00BPDZiPGYywbvfxOgcXCeiQ
ECbzbITV8vr27hVmnr+REv6vLHtq/JqXLUCyhyp27c/AG/u5N8xT9Kgx7vc8H8nV
9M2XWl4uEpcHsCN1t8dI7AHnEdJoSsijS5QZAFdJKCRp2ZhlhGzSHmeaVK0qjCeH
CsqpLgaXNoorfKCE3YaUqexT0XvDkCbwPFMKHpai/wG7kA8vFJN+iKI2Nrszld4k
jo22Kn74N3AXcgxRbu3JykEv+PqHqKMnzuCzRzIKtI8TYhhuCiaPa210AzoNTc9S
K0x8NlA7yM1vu45AYa4dU1/WvYZF1WY8khqVLyWVH11P+/qNasgpnchYgzyINxHB
808PvcUif+4OtCCZCLdlRMlhjGOF7NiBf2QYSl3Kb/tUleJTPS5WhSXaeZgao4PY
M186F1LhB8E0/iiuRFjnbFJCZS6v8dHOQHxRzqHPu4aljvzGyuiDQJ3QXJE15G5d
YhOBxAAwlLaKqkDQoqSAjcbroqB66Ji3SAhERLJzErusHGd0DxmmiypeQMpLVute
QGc4c1KiegSFumGcMLHCwsENVNpA5FJjP+VEHsqqpjMD499LdeeznXgl6YZFAY2W
8fVsptRFZ4xmHpfqNGqXawC38FQ/FDesagjNXhkv31tZW7h8xdgjLS/HkJge+n2O
wJ2peEN3WyovYInyH7YUJd7gUcNpH6rM7VUtWogPcFqJRo5L2BK8Hycxxyti27VX
PiM61eVeiderZ31MwttRVqtFalkYgIS8bbjpR0RlzvfaQH9Ir5hRlUXgNDWmKE80
cadAwvg59pY+Mfe8Lsv4tmyyXmoVwRuyP230JprUxabugnq7nGPub2H3uv+EMMdo
ByNHeqvLktKXq/4723NHNtTlGhodVr+FFeeTIv+utEqhwkrRQ3eToNodvER86e1S
HoK0sku1O2yF7MxSDnpnLlVkJ1GELKuyGMbUc6DyjAoLqJRh0urDVDVtyK1u5Arh
xoDw821VWBgXDhnT4xdhN37J9aq+bm9o3bIDnptMCZSwGL9y37KkcyAn+vxq41qw
YHZBAOEy4Y1r8EIv4IkTDTvRWywpDUgSkz6QnpdO/CroeP3XKC9j9dCK/MFInV5k
zK/g4QTSApImwMdwW7N0v11/7xs7fIpK2rv4N1jzJj5F4Ku3lX2DCzFXUrds2OHe
y8rKJ8XpOhRSAH/xZj4qvcAqTGGZ6+1Npz7/5hsLJlfL81NJ/aAlu5nYs5Qi86r9
166SxtchkzraUvA0BdEMeQFVshRKE7pHR3bh6NMfePhypeJeTxWIklcDD72MXmcu
oP4xJ/7AGH+ZBsA4JQ/M9yC76htUMvq9UeS+hvdKoydr7/VCiHNb3CbEtzHrf1MT
fWu6ir29xLl0ZSpvVe4Y7Zv85GtYJSbBsqDtebdwfpdOtj6G7Xddp290k2VlqNbC
d9NQVgMx2LhiVRlq8n7i/bKx8qM7RH99gnLF1GUGmnfoe1C2yNFyOTJHUhL/QWZO
rUZ0yF8QFFqG0uPf4LwnNXhNavjbkT65NaCl+GHoewrk32eqyxgtuv9QgsVuD7Ud
Fgao8AnaMguxgosWSh2ZBw64I22xN3Hq3LN39qRne1VKWvXtfLAXT2nHofupWP0I
E+HpWwY2Tm2ElyS0pYfYKDWAo+IxdQq+54kwaG25x3EpaECTbEYwjW6qF62vycZx
FRImBVwdo9ENEszrVg2lHKqflCRLBz6YEncKZ/JidgKafvV2RN0Slb5E61BIPC3W
JNOHg+3kk6N08mxXN74ScMTWl28tiDu3ZABrX3IcqegAslJ8rUKYmtf6ci9CUITW
we2MbzHqtUt4AyxnrBpm0XZ5f8cYzdRWgcNTLJ01Jbfu/M3VX07/7q15Sgip62Od
1iTzgXCs8tOBfGiCWFJlIYocyT7UIMIszzvklUm0GHi3718/1HH7Kp2PfWlNFkpd
Aj+fQl0I/W+4DZGDsq0y9cwxnvd/o3ybA7xC4atpgcZolym7XsnJFGjn8Y/sT+cG
yaNC2AzF4CNR6MnLVX97MjsUkIhQOYnDsV0M6dHqBJZfGlNtfTs385ogRfokw0vE
ppXVq2ejEFOUb3tszeXUBJQBpT6QlT2/EQ+KQ/JKWshQ+pZctWWK1HOHrSa6nPGn
h7cz+y3DsBhon80IW30RvSK1UBDmAchCX3fZoayX+CcPzTXwkuZG0tKISL5QNCV4
izAulo8KkS2PIlYIpWkENP9SxGZZP9LGvhs0f/UTZsMGuHlWhHIB3+C6SSCQjfJo
oBIvBcT9QO7Jj9wygFn73d6v2CoRnArsH/gks1uhuQfzw6e/kg9Xa+31u/SsJYlw
Vf94Wpej8YjXCQmRfz80COd4gRMvC8EPlOgL3CvQq/iGblER9lGayiA+D0aZzOE+
RbIpXJgdWQ+SgPduF53U2SceiLsK1pwar1XtMhjQNPXZtq7URyC6BMsisTh4pX7f
M3DwEnfZouY+sLGTFKZwxyM9x2oTlXYyCGKzrPD+LO175rRGhjlHihOxO2QjnLX8
k7+aJQZlrnlzu5slHXai5dFq+Iku4i03T4+jmTLDLeA1uKWNzfb22Qlcn6U2mdvx
mlgMJUCggA/y3+GF4pT9ziBPOCFel3/mPXSIf+qTAxWazf+Xt/APV/pdOWupdyhK
PzCk0QAuIcYjaAUNQsI4pGr2d3kLxmtxVMXhfswzplOmYyG//636So8dT2XPHKre
38fQpkgAWJ7VrTEjC9wj4lV5qGq98XjOcn2Jn3d+JMZMJuT4SDJwItsOvzHVoyzF
Kq5qBPfVxNTiSqFog2CjWfNPMQflxxSatr1D0LmkMBugR8T26vK1rgq1gViGGIoR
quDCjfW4Uth7X+ZiqAoJaN7+ecrp/H+juNR0IZoss1iy1fuyJx1CNyiVGC/MGPs7
NIofeHZOOmCNl3hLeOTWXsAMVgKs6/HRMShaM+PgNoYR9kuKhFf+B1Z08zs2R2U4
XuzZPD/xXBF/096NT66BlVv8eHC63zln7cUgtAZRqJL/yW9lNcBZ1YWUetBZZd/5
Y/3CmF/FYimU2DfC6kmCWWI3V42aL5Td8Hm1gQJdJBgZfp78B0ZzlfaoiTP/827p
aBEwmidZLJsV1hWP9DnOkjLk6WakZ4FWAu5f/Bbacq0e7Rdp/5QzEyAMSBJIGCCO
cTSvkm2TZW/eB0QWwtYxV35K7yTgdwYHSCGVG3iuqHxhF+fyNbfBpBQ+Fr1dIkcx
y4k/z3qVwmqV2jeeJ9P5wu9HhvGI0v9Jaq/GjbHX5azHb05yIcAGpWyUdsbzC3Qh
4leGkpnRDSB+EY2nh8iiDzoFYWNt+2Iy9dNRQyMZmyiSY/H2dpdRyDXfreHC8AtG
6FDezP908Ro4EoJeXwBPbiyBlhQlCsEujEdJdkisAml2kAkqxaKh1/mVnhVDSfgA
1AGPz3MFfO9RoBDlpDUZnzznnfUBchUhXgs47Dne4T+7eh9GzirXfzxEdzEht4J1
TNPhyM4fR+NJ8N333m6TvoUz2fo9OQxcQ9c6LPB2wz3IVlXbaptd36be0RvXCO79
59nNfO7xXydL1iwMXUArBEhJpEGqgOlK1x0S+mlGXGXB0qDYpV5MNcuMPfRji3F7
okLbteNQLHvghiDoKlwN8HGU51ObBOYC8HRnBvJqEosdS1jLriid+Te4d1a+Hxbn
Vnby5bX5FMcFCzVb6kkWeEzT3NhBBgQLucBJNyaiZFmXxEhO4qgpJhEW6B+mUu/C
pQ1vPUP1C7l0LultK9nQ9LXeU0YpZ0wkVS48mb8Rqylg2RYbiQ3wVtAU+YaGeVEo
VDeA8h/fiGXATnbCXy/7PT23YJ++D9g9B5fdivHd23pwKDTSsMdWc3GUzpL+tXO0
ecOs9rJ6cdn/giynAvfPztvgfFxhevZC1XA+DjY0c/xhJ6zrugRASVAwYoDWlti7
/NRSc7b6xr1zWQLKHrJTg3s1CFzyd4uxA2zzS8EtFHF6EGJbSi2iVMySaEI1SoNz
MS2FvM0/XPm8FXhqwybfbKGkfYuPiCBX5qVK4+Z5FnOMhGAxXV2/I/kWxIEzG2jF
bYsXlT1rioy+hBNShnRMMJk/zuycSYV2IbVry/9WBaCaKB7EDOuUuHjKkQApSUg4
HcZLqCpDKLFg68jgBrAj48aSfWQjHzbWwLTin+JfqxTvs2lytHpcUBfHYVYRTu0a
su3edMR6a8VN/NQ5Z/3R9vB1Zm5+ErIGhmRzXNQBph/ZbwSZNIruCWmmHHErucDO
wfuzaG+iFKAu9wBDAYRqmL71a+832W+iZHh95B+b952HsgBkEN1cEyqmiXl83Tys
pni+xVRzxzfFPEVJD2U7E6BCbRFTq/852nzm7H+BrxMLddWhTMX22fBiVqMIbY8F
nw1SJwHFWgP1IjNg5LV0uXZ0llBQaLPj1m2c+sgKFZm0ZzHvxvAxU6czrm7jsS9Q
mkNu9SVBWUeLqhS5sOvWqfYsiJKIN46tFU+Bj8GZAoz4FTy6SvPl/h6cpEgTnyHB
woPwzdnSQIs7461s3MRLbN6g1hDuw2l4bzyTc8Y4esEwnqxEWsR1sC6Ks8BmQ3rK
s9vJl2f5VDJAv1LTlUMocUXyOivQ/6jQt2RLTGBBRyXTS7LkCLiNiXemf6oQefrx
RnJYe1yZ0j6Exau7dS+yYhBgzjmSpBV/BsdmZ5ujAq/Yk9+PMoW4X91GvNbL2eKm
/s/8SI9BSHs+3kao4jHE3nhUUqirdKzlku4h2xaIdlDZgwolArAjBEInu36WCsjC
Zz10pCMpBNyoRa9Q6C52QIgZTZ1CKl2e7jybNuOnj3fWuhPEv9STJSkgt166DLpD
Nor5V/T/GYgEihkRjqKJ04UBFqkshascLMfrlxUx772CGDVuwKxE3qlHv5LH92EZ
mx5OVVElbllNmET6mJWuqm3oIhDUhROwogNXCSDrWcA1DDZtcUM68GNYcgripdWu
KQd7ME5U3/2kQWVXfqQXl0P/uUyMiToItirB7qbMso13+FNhzPA0vA0VH8P744Rh
`pragma protect end_protected
