��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����Ղ8�~��kD3~�bVwv'4�,�\w3-�P�^1G��8jH��|�Sq���� ��`�h�r�%1\��Tjk��qJ�T�"��]ۓ��P�Ҫ{�����`�w��c Mq�`CΦ<'c�>�"bxw]�؝ϳl�Yya�e�=���cq��oc~���25�ԭ���I����Dj��b`�V=�}�\�ڸ�E�y  ���N#w�������!������v���Yb>3������ō�c�Ҵ�	��C���g�y�B�W��0�WB=Ai���[Q�Y�q�.l��zDl�y���(�Ē"$��m�?-�i=�D�D&,>z�{g���觪sp�c�`X[�K�֤�M�]��ٲ�o���\ 	���Y�_�;J�LN!�Im@_�/oo�¨�m���O$w'�'i]��:0��9��^��b61�_N�!�f��-���4�f^���EI'`�[�nod�/�^��0�<��TT�����C��ɀ2x<kk��c�e�Y�@*�k�m�ݕ��w��C����}�^_��4"k���d�|��� ]�E��v>O�GP��	�:�a�v@X���{��.KTU2=�蓠�~0�w�"��e�V�y�;���lQ|�8�v�h�v�� �oh�ē���آ>���n+�o��IѪ	w����g���tTu�@���gtT�)�J�V�^_D���8�T}��ve�rT@�>�v�ϵ��K�{>ǎ'�GYބ���y~8�pn����P�����(�Os*��>1�㤪e8�+�1F�E�d��q*�Mp�x��h�6��H�Bs+�t�4<<�sn��<���¼a:��NB�ϣ	?F�	��|?��'5a��S󌼟�W��p?X!�kP�&ݱBġ�U��9v$��e�)�M �?��wh`+��b)�f%�ժ���Ǔi���m�+�J'�{�W��9��π�`��|&1($�cӢ�-��Ω5Z�Jɗ
սB��1-\��#6?ޅ\f�q>�pu�,qK�a�4���O"s��[L-��84��_RigٜML}�:9L�.�e�y�7E���C���F�9�]9�O�fG����cu��0$���j2�}��P1�%~aW�h�`�Z��cL�;��}����c�[����9�
�%��F��y B�]�Rkf�S���(?:�y�����B���R��C^-�b8^��٤�4��՝kC�����{e>]�	��X����Ue�;/P�"�1�]�����/Vp�&MqH8�F��O�cLb�?���?��f2^���4��7�#� 8���Q��JGG=����o�z7#ڵ�Lݨ���~8��:��kk�)�XC���.�"8H�R,0����_�R�F��#��=F��)�Ab�#�Sq=�*u��Ša��M��p��8>B�g�h��I�R���*Fg[qǝU��I���Xu���g~9�z�a��/Q!���_���"P���ao�b�A&�<q����Y{u�a��
�������[�_������
��ӟ�G����Q�f~�,�&�;7D���bL��ٲhF�L��cf9އ�(�.v�n�q���\*������'��ɦ̨�N�n�2Z}�`��e6�v�Q����O������]�Sӵb�9o���z�Q���7a�Lr�]�Wst��ę-lqć��c�&tP)�⏎C�c0��"
g�Z�T�\��I+Tn<�*�liE�ҭ�&㡆:C�+yբ��7e��I��A�tɿI�5�־�c�ޮ�e�&�i.��d@����秣��� Db�Z"l��_?�[����}�]�v�a��~��?B�&��å����\d������'�V=�@d)?���� 1�+� �Щ�dY2p8��"��2t��iŊ���t����R��ZutFf:�j�J҇��0��Y�t~N�5�7>;�0�.a��J��G���䴘D��]����P/_���9G�>�&�oJp�Ӕ�Y%����p܄Ǚ��	�A*�	=�I�[��c����a�Ӭ�b��s:��P:���0�P���1~Ŝ]+�ājKb�yNw��E��o�u��W��N܃���w%M���ߓ�z1)D�I�2�j&&H�j2�����Q&)#�@!h��0�|S�0,�g�b����1�0H�4����)WC���"�Z2k_�U�6<thN��[.�*����֒ʔ����w�)��,��\���c�;Yi�l:�9F����bl��F�Ӂ��	o�����R�]q5\������k?]�BC&*y�97Y��o�b0J<a����;�eq����8�0���	�ZyS��;Z��� �2��_�ƌ�4���[QZr؜}9o�	�ʥ�ˁ;$?���m���p�t���>	���Q۪|ǳ���в���Uط[{8�E�Nw(tM�����`�`W�d��``�E7	[��u���K �|����2�T���^e�������gE[���	�n��GU���~�a�L54���;�-	Ii�o��f�＂�Cv���v�y�K���I�w+��¾[3K�҂:/��$m�b0��b@YNE�l@�M��/fyZKJ{Z!����)f�f�"��O#��j4�w�I8���gg� D����QU�������
|.2���j�4����-ۡ�ν�� ��-ۜ"-�ͳ-�����7FJri�(�g�+����9�;�^�b�D�v���X���
��Es��<3�%�Z��m:W�H��|=d�p�$���?/+�,���c��Y���0)q�n�#MJ���Zu�>��t��YI���O2����2Tu����L�
y� �WFZ��$��U�&��(���sK_MO���q�^V���D������s,�.� �L��]B~����4!	θ;RV��d!8�#֭8ʮ-Q{P~�"�?%�VU%����cmPѯ�JF^a�W���vM�?�!�gv�Yt��7����"�=�.����NwB{�	�V�U���(�TP��Q���ٻ�� ʔ(L�]�"e�V�~e�z&&C,0g�=�H���*���&#�3U���k��	���R�8>)��/���9B��\N��ɷ�~�f��}ⳘPB��:�0_������J����,��6R`���j�,M�E���bЉg̟$v��D�c#��W��mk�Q�t�����>!GQQ����Z�H!#�:�f$�/������hE�AW?6'�5�˽K��~t��7y�/�4�#�x˸2���$4�����aHN4����yWv[Ƅ�א)E����ۣ(~[���"��ϒ1�3έAI�����#ݚ{\j�j_��J>QɹoC�S�X�t�6��W�4�]�zge�%�I}6��q+�E��0q�e��R�i���-�~���ڽ���8<�G�<]ł<��X���+��'-�)��df�ૡ�b~�H�0*5|@h��K��~��XX�6VL?��oDӠ�v;�4��x�ɔP�IDp�*U���~rh x��+4-2�w$��.�y�#�J/"0ȋȇ��0�Q����E��$�%6��U�pj_Pс���(H;%Q���\q�FD9�*��z4�?F� &��E�v������7baCF3Y^?�l1�MS�J|%!`��wNJ8�`�HB+Ƒ��*�}�k6u?I5��u�=�-S�a���X��t��iquih#p�^���w�()fc����E����������m�e��\I�.m%o��Q!���ʻ�'��޿S�-z'�Mǆq!�5��;�P�}���k�G��"2n���!�0��N�S������?��	I��i��b�B`����?��O(�H͉�"�]Q�n��m
�-��'�B�Ȥ/�_v���� �����$�;N�����Y J
=�:-3�7�y����_(~�b�kع��#�u.�K]j^|('���۩hyW�˖A�L^�G" (]幄6������4H:�"*[���*;3�� ��$L�$kE�"�/���|�^Ga�h���W'<Ii4�@u���ix�fhkU���Ҟ�T�ͧ~�(�E�o������P���Ն�95�+kz���W�AJ��[@�5�{tƛ��D���3���UG�"<��R=��uŦ�+��-��}z��w܋�y�w���G->�)"M;�R����@��99塞F,�x9���M:㟬���Û��Tޝf�q��"wg`���V�6�<�̨!1J��#���7EW�̷�#�M���?T]��Q�^��"UL�_4��áQ��J��l�yKu~ƵP���=���-��[R�  T��o%�Ki�x*İ��S8���ʱz[�ƨ͔_��֏t`�⻜�0�0:�&Jb��x#�Vd�1�S�a����d�_�k���Pk!���7�*�3�]�"K�{Ct�����Я]��39`d�u�@�.vM������@�"05By�+wƷ2t*�ka]�&H6ѷ�5�k� ��>�L�֟��}�ң N>=ˌȝ�ܸ��el�z£�t~zb��hK͚@��jR�b&h�R�K�i):�6s��B��H게���$̶��g
[���amZ7&� �'�p	e��4-_}�|�(���,[�
L���_�<�C��&tu۳�L���� �ڨ�n�8AM�J�uR�d(� �cn������D�����t�(�)x}���š��D>
��:~Evi)-t�A�a]89^�	һ������+z*�MDЬ�����k�Td`_k� �h��+đ�+�%N\YHt�����h8cA|�����dD뇖�*��x/�9,�h$�A�v!H'io��'Y���� �8]+b�Rĳ�.j��*[\�|?,��8��a=�!O��Ƌň5lߎՙ���,�O��h	M`�tvh�
0H��	���A~�d�̄q����߈���$&����0�"�{��K7vhV�W����baS�b��_s�eE�I��@*���f��� ��@�7_��|��Jt%#�GLҸ0P�K ��`�m2�U���*%��@t�ΉQH��T�CE��4�+�@�G.���$e�\v��mߦ*;�\>�m�-m��-Q�r�P�
꺋Ai��yuN��j/��.�.9�Toίm�K�R�@��]:��h���V�6������hu�2�$,�.�g,����Jԣ<�V�!{4��V��J
ON�x�sVݣ.*j�)_�̇�i���V����խ��}mY�++$�%�$��5ڑ��na���Xo\�����&솱j��BROdT1hN�����%}Ω�C輋��5<��
kp��U�o���T��'&eX�~�����T���_�D+>:5z�M���c��,�rW}����s�Lo�$�?�!��F��Yp<(�d�����*������Q��^<���v8Z�ͺ�TR(�H�B�����H�Z���^e�Z�;,�s�h���qx蛏g��>I�h̽��Wu7�h�έ4j��B�kr��Ю���<��1����$k���2�+
+��)�]j��`�u����t��L�M᳸;��o���#ݱ@p�&����q���&�i�Ɗ����r�n�=ɑ�����JN�p���3_�ٮ鑏��ޒ#�_6V�������9��y%@r���� �����
z��,x�Rf�/R��h:�R�+p�]p��d]S�*�L��[�ʙO���)�]��Pp�c�3�a�H=O��<�jsg�h;.��>���d�^�k<�ã�*����-w�u���4���U�@��Y�t��
N�@Շ8!bC���s����R?�ʄ1�ۖ�4��6QQ���W���F!�X����(�~��6��ˆ�\��R��-�!�ftY�����,;��6/~�������[�IA�bA�T|��b����d9�2�6�cof�2��ͦ��lkX�	�� ���WJ�3Ё�;�(�������|��4	Nl+���I�$�+��"�8��b3���D�ZӤ��@�7�B<���~��0:�&cw���)����kD#�����\|B5��>���ԥ1��u�A5|jl0ւ�:8,O�*C~f[/LѾW[D;�,D�Ѳ��V{`��Kr64������� �e�d܃�C5�9'����4׮K�<�Ӗ�����u4�Je��@�N��S	�1;�p���Ց�lZ"�a����km]��$�Ã*<T�O��l��+��q����OG��*���
˪��������=+���O�@p�LdO��йx�E�Щn�P)��0�RU#�v�^^����=?>%���d��cxf7��=����� ����C1
W��b���e�R��Vi�T����X*����F�i2����Z�s��G����Q�> ����n��"+���K��f�I|"����8v�e�SQ���o�>��*���]b�������ɾ��Ǖ�Ԏ��.k�mG1��h�b��m�g�l�ZdFED�~�B�����{Z,ou�T��T�B�nͼ�-l���Ǆ�a}楒�u��V���H��
G��@�5&�r����^�<>�����@}]*p�������o}%�8�%���[�|�B��%�4[�tr�`�c�#�a��l2�;���X}�d(���
�C-C}���Q�Yq �\L����~�P'O��G��z8s��r��^���o�}��7�oe��+���@-����Uf�XBj�P��G�7�.�u���ȭ�t� ���8��Rk%�M�t��nf��L���/��{Σ:�ϵ�(UE���@�j/9�i��"UkIĽ�2alU?�d?�r�E�`%`QM���9>�W��ǥ<v/R�����x��8�i��m�|sY�,�'yM�W��:�^A1��ʢ�)���)��M˴k��0x?D5W�7�����%�N�Vf�ln���5e�\�^K������ƞ���_@�c!C��_�bT�)0��,�Qu��MY�>vȒ��x�|ٰ�c���E�g�<�8�i�k��:$�8F�gb<��`�?��B+݃B+[c��1K�o\��[zOye�:�@�N̛�CC��Q/�%��c�{�C�"�������A�/ˌj��^��Q|�Dw���NA��WOQ>)�[X;�q�o䤦�ќ�`6�ӺK�* )o������@T��G2BUJ�x�$�7�	~r�=QUq�l��3����;L��'jZ�aLb����2U�c���]v�3�WD��r�"D�hՎ5�	�I�A~'���q�&A�� �bƍޑ�����߱K�I[��[�t#+�X�$K�R�b[��},8	������:�W��Č��Wqm}�3�s�����{�n��pnF�]�� �w�-�&9��/�iZ�{~O
*SOKU���Ry$1�!ݎ�Kq���t������)�9�zH���r&RXl�K�>8�M{�X�H�L"���W��&��Q�.jqch��KoF��x�����Q	8�Tm�ۚJ}��,��  �E_�n�0�r��GM��@��މ�
[�4���'éT�c�X<�\M�1Ŧ�|�ccgo���(��y��d7��?�8�;Ok��$ῢa6�~���\6�	��"L���|�8�T�
�>��<�����Ƹb��r�Y�&�Rc���s� �Z���>�F�7%���J�o֬f��r����~bs1q�s�ڥ�ҙ��#,~��ièmpv�,k��m��NT����h���gn&�a�@^bI��EZ�cM�z4��ѐx���Ǥ�I�H�(�pX; s�;�Ks�;/��].i��ta���n0z�F&d$��:�9�b���	�H�����H�|d��Y��0T?#	�o�vX��Z�Z
lq������ጆyI1�Uz���~��0��ZF�Ɂ��_�[;�Hco�5}��*�^��dl@;��
�,�
�+�6*����^�hp���W���3��N�K2vQ��(�G����Ĺ-,[TJ�XP���'s[B�r��Q�3�����$�ZH'c=���S�V H����K.JA$�Y�b�)����_艈!�A�![���"�p�=(�����0͏%���s n���������)h��*K��������uG��)����A2���!���D�EH�Q���(cue���{���H9U�����M9ƍ�vQ�|�G�aU��U�8�ɾ�����V��[l�
�߶�eN։�~�"���grv� ����ӅMN���L��p�&�+=%��k��׹X>��9,� ��Q��2�av'�����d��48����d�}�P�2bG��s2��(<w-�����,B�`B_�+b�xD�] �k7�y��PS^�Jَr+����Jy��& ���4ah�i7Ȓ �?Q��մ��o�@���L�Kf��;���$�؛����w2y>9~_mr�ӳ�Ä��G�W�8��T�Х��Xw=!�-HQ^3�Gx�L ��{��a������)������:��ZB�{�������T��S?���[&��ʘi^𠉺�`d6Q�k�20WcAO�7�F ^�@nȟ_�Lt9�K��ɶ�vd^�����p�*h ��(�Ó?��F�:\�ݟ�p�Á�§e�%�� ����&�[F��J
QAA�
K��j�����al��$t񕸋�8?��J�N�Wh��bZ����]А��m2����@�� unxrG��`�*d-��F+�fu�C���l����0Z�f���`���s !EΚ���A�)��zt�kN.�a�"VYk<�LL��^<�q�<�?|t	���G�� Y-�L�������cf+b������c�ZF�6]W�6����im�%�3��=�����NJ�S#_�/=_Ǆf���vw�ׅ��-A��ZO��;�Bt���f��*R25Z��"�N)D����x��\��Y\
��k���G71RK���1�a�v;V'/e?�][x�xT���z�L�v�F>׼<�������g8Bzt� � ڢF*�P�A�|s;?�ڜg�K||9[��}^���5\H�#N�a�+��q�Wj�h��_�Q�2��u!��+I���ow�o��|�@S&w�	��~<�]	�N�?�'D�h��W���G>�,J�!Q����O�@u�r��
COx*,�n��1
���ݧ��,)W�����&��&�O����=kGS�|�n%�^�}e���[�g:�v�,
N�Cz=gVqH�"`n�������E#��J P�W��M�,�.�V©�r�b�ZƔ�b���L�qo��'V� </w��qԹ� �)�x�(�u��g6�R����?�]c��~z4tD��e�9J^�5a��?�v�Փ�"�.=���������%vD;���+�#_���,B41� "] P�>��Y#S��z���� ��|D�/:���z���?�"c�X���Z��ѱ3�2��k���&��<1@�ˎ��܈�f�z��,�#���Z�TV���`2јK�I���D����)����_���u�*
��w;���(�Zu)��"?GV(Iz�62��Z+�������=���w�3>��(�%|�'��&�w��HCw�3c������E6[:�Q<�GvX��Q���qr�C��ꖃ�+Q�[��ʘ�$��2zm_.�$Ǳ�(`=̹�V�,���h��XI!�!��j��3��}���q���c'';�����ZU��$t�	��	�_Q���:�QD�V�KIU߳R���혥^�NH��'�D��_�Q>���hs˔����J���V��`��k�C��.L-6%c�$�J�g��b��Y�#��cTF�^N�s��r�si�Y���L��1V+"�dE�˭*S�$!N��g�����8Z�Y�|!��,&�6"�緆\���̥��8��Q�Ž�m*�A6,���!�GZ�\
=�@Jg��b1��B�3�1n��;�'ղrz֔<ܥо~���R_A1��8KTEu�(�g>�������"2�R�[#��b�'p��W#����?jow'߇5d�e�ށ��fٖ�sD�C���JdD\�&�����Ϧ\�0}3)(.����B.�~M���д�Q��C���
^����X���ì�1K��eEg�D�$>u>���@\�Qb,;pO�bpk��*D\�2�4�;�TQ�rM�/��#H�ni��}�y��z����	�h�E"9�� s���y5���:u����ѭĲ�c� �*7���_K��)'gj	�d��LB);t�k딤�Gա�10ݳ�)��+}���v�to��C16�j��P� `�pi>�w�OxI��H��xoZ���M�d_�PShj���}��4-�5�/ȹ2O79��ȃ��6{_<�e�&�G��XZ�?�>�_�Ȱ�_=�R�2m�_��m���F��H�[�S.�\�\@�.�)�h��L��7�Ti� �L�5u�����ؾ��i~��X��.��^�?��@�������N\J��*��6M��<��K��(s�Cj6�?��⮆⟴�ˬv"9����e��o��ݘ6�4MB]���[�v�"(����&K�a*��R�a��X��ʙ�W"��Lʔ(��	v~��I��9�rv�q��%�����M�}����<��7gB_5�,[�1��`e�<r�+�\ƳiЃ_qX}�<*�Tgr?�m�"FD="�{n�:�_�X|9,�3�$d��+���c8�����k6���]�F��n��2�c����@'�2�a��>�'/]<��Ш���K(X���əxݒ�������n\�܌��p&9E�ʫ
���0`������W��2�HgIKW�nbW�s����V����ނ��q��� ��Z}�RI���d�P��8�}WV�%F��ca뒏�MH���}�V�.��И���^�#=p0�@ӑ����R�7�k��Ų�/,¨Y��]���8���6�����;���K�r������vd�lˀ�-�;6Q�z�Z��S;�4���m�	�aʤDBA����q�J����HE���^ރn��QY,`z��c�l����Jf�
6��nV�V��h���'@���?�Иco�^��������nT�7�o�X���uY$�*7{�������S�E��s�=����
n��7~bX4��F�[fth�
y�Gl���G^o!3���7럡x!~��o�U ���hV��dE��&�kYG�~#� �V9V|C����>������(�e�ص/4�!������~"� /�@�,���.���'5�����*�+�.ݯ�� �!����^� �π#@Mh�[�c�QA-p���:������w��-E�r .�~�R�wY*������X߰Sp�t$ ��g��8��H���f�@�	9�Sx����||��c����E�A����`���+�Vj�1�%y�Kw��R/K[0"���{
gs��+	�^oi%a;��^vC�ۡ�����rL�|�om��g�<�&��( ����:A��p�N��$��V�r�#c���N��,��O�V!<��V�o��դ��Ϫ�&�^��4��"��K� z:gU~]g�Vl�o���I�a�j��+M�.�:x�&T����Jj\,��~(����;����O3���q�I���H��7�td=KF�C3��i
1ڽ�pd�Y񤼕g"�vl$o����$S�tv��"�Z�g�_O�1ʔc���<�.f�
"	��N�jW��@�3C警heh�lʹ�r+��٬w�0�T)kl��3:�{�����_����J-�Dm\�%�b,0uN����Pa�K@�j�;��DF���b�Vf�Ć��W���/�ZH�>�׿W�9 Z��?P�: ���^*��#�~�	|d��W<"~X���;r�`iY��D��~�9OʳWI�R��blh�,iWdy�+�&!Wb(䄈����?�� �&Z��ӛ�}w9Y�t`'	e߼�X�g�F���'�}����!ʇ�{�;�ͳA��d����k���Ϳ,���L�
/�R梈��ÔE�g�l��*�U���O��[x���j�+u�*�%t��P�L��cg���9qo��|ڡVNG��0r��J����pC����IN���ǆ�;3j�Ǹ�v(S=�,������d�"�sc��+9�r�oEi�tӖ=;M�_�k�iQI'!�Q���Ҧ��s���nZ���B����:�&�'.�[�z���t�'� Q�p�/�?�J�3�N��}0?N`+��ozK��_��p�޷�l�AG}W4��4a-�eg��n�U�p*�3Ư L�"2V�V���?y��\�]����Z�z��o�6�I%�R1}����$�تxg�d�9(Jf���G�&<�xp�U�n�:��D6��A��;�U�ߖ#�v��m��M�kݣ�΂�!���cw����/�`����kvM~i��8,i8����A�fZ���������H�g�����L�*�M�l�s'g<W"a7�6O��Cs�Y�&+U�y�{����5yn���Sm���i)t���k�ܔ��B�{U�ԣ+K�����|�cR�Vw�Y*j��mڠ� f�KZG���-�jR�1�����H�y��C�Sb�첰�`�R��gZP����9o�K1Nu*�KL�48J�H�ĖiT6PJ�+�D۟=h���+���/n� �2.�$pz9���_I���'�l��"����U���vbY1�5��g���\���1�#����0�|}r�G�Z�.?�����DG<�ȫ��2�n��dm	���5B�q�#�1?���m��J���3���և�^έhTQv��x[M��An�����x_W�22�����W��N�S(�L}>WF��y�P�V����?��O.:����,åW�v�٨J��1��Z�~>9���^b@B�*�Y�
��?�CYH1n�]�F[F�[��!ک�9>E�����1�o��d?b�X,SV��d��1�C�q�(�dS��:$���� �I�a� 'E��|b�CQs���T a��u�HZz���$`\�� ���.��8���e�s6��bx>
�Vt����]����Hv&��Wl�vO������ ��Ң�n����`��F�����<�E#j�%���Ij�D��Ų�E���9�����S_��!�_�����a�do]qC�U�y�ǥ��~��Y%��0=��9ɖ�ADӺ�}7��ʟ�\d�Ɓ46-����.&z�� s�W�����q^y�G��ѻ����\�sZ`Vه�&{�:�ag	7�m�6����W�w���oWJC��˯������{sC�уm��h�v��yc��W�O��Iy������/gGϾ���
�E#E��@5�e��/+��s������W�zB�l/�j���Դ�?r��8���7	���NS�#'f��=Z{�A���Ȼ�K��B����/���Y��Q
w������=������=auj��p�`��:Ѳ�.s�5zJv��WGo�?Ȓ���4͌��dс^��fSt���*s��������/��t�=B���Oj���~\3f�)
M;��#�����ǭ��M�y*[w�<��L�;>�DS�\?���RR��MX�؈�W�KX�tx���Wr�:~I�f��27��Y�b<O?hNީ%˕�T/�@�I�\QH�dd�E)mD�=ۀ�ȿ<B��Ȃf�]C�^b�zV� �B9x�k }�ݠ���d��N�Mz3�OQ`Ec�Q��^x3���2�t�2�)�����3���s��J��	(���߿-]2D���0��(�A2Kg��A�τ��#,_�k���$����%r8�%�U��W7o���2s챔m��*�E�9��`�đ�i���=�+"./�ǩ^�	�m�3���%M����>$��,���el���ș�袑�{����e�ɥ�B�5}�׭�2ނ�$ͻf���� )�\v��i;��1��P��m�OF�w*�"s&�|!���z��{����p�� ��ZI, �U%`]����Tbw�0�-��_@���J�=_(f�`JM�	@�X ܪ�̫�@�޹W�0���B�=6\�Ǳ��Z��r���gx�˭7��&0�AFY�wA���\MA�i���]��zn�k��̸0:�=���F�zjE��yX�8HDH�/��J�:����^!j̓�\Kx�]�$}RR��� �V]ܧ��t�%j	zX�`�Oo�ۤ>H���?~f�o�N�������ڿxe���=[Q���+uD�e99�L|EO$ya�9'h�IU�]��i]���wiy�UR5��=`�v�$<�J��55��d����}�x�?R\#`�!A���k��1Li<���!v�m�#5c��ܘ��T�n,a��I��u��g�g������ ��jQ�A�P�g˩ja��8Ŧ�%,���\���q�|���0	bw�j�	" ��6,<�l�^�/���c��K�?M��}��<�?�7?�
w��z��T���hϘ�zN5;u�'��\3������.���e�q�?������	� �@���6�t�y�]p#�j�ߎ��JV�l1,jv$�[���րN�.)�g�F�Q����Ȗ� �P�Dn ]Y�N��L��Y���
��SJ����nc�����*p����p�)2ək��Jq�#����	Ӏ0�&s�fC��w�U������9~� �r�J�vTn ���m8��<�u�J�zA ������d3%ǃ�nϰNt�L=QKvE:{%�iR�巶�sGK�`��!��mv/�y)���d��`s`)���f�����m���76q����&�鑹�3~�>ONF�DZY� ��������՜J�	�n��)\����U��c{R�j��rrs�s��L0�ګ�t+yD���s<��߷*	 %bwu�b�a��~f�����?f'owt�P0RS`�����/� ����X�L�+�T1�e-�~��70`}B�A2�� .���@E �Y��(�K��:׺O～��Ժ7�<��?CE}�K��ĭ��H�s��O��Ҝ}f��j�PW䕬=��~���d��"PYn#ށ�D�5=����k��`@+X��x��2�����@Q����yL�QLH�,��F�t���y;74J��a��GLu���b
{^٩՘:�ʫ-�e~�$�]L�&�:�1�E�i�|_����N1uKh��y�i��n�Xǒ,{��@������ݠ${V �F)5����/�����m���m�j�F��T��[���5%����[
|�%�����oD�Z+�I�_�o���
��U��ڠ�
��̿#� �2�y��D_U���F����B�o򵰬�rFQ|�	���
_ي���)�`��'�$����MMU~�n�i�����Ld2F������ǅ|1���Ջn���O�J��gJ/�L3�ֳh�wĊ�X�PD�1Y@ˣ�R� {m�����7�'F�y���;��/_EB�=���n�Q2�x�����#�P��fk����.յ��V�Mɷ�o<Ģ�E��͢��2��f����u@ƹ�<N�So�=P�����b x����t���cZ��bo��z[u,��o&Y�lt�[�<���ΫЫ,8�-R2�>4R�MdV������� X�B�A�qfS}�2����>�ⵊ���4�-���i����e�kb� h��M��9���Z�O�����p%��"�e�p�pэ	=!�|��ZV��� �T3��N9�Xy�</h�a��Q��T��|�_~�6���<A�8����2�����;X�>�;�H��܃�W�I�rj����HW�����:a�_��>Apg��P��z��P�\�U.���6(D��6���9�%\�6����晪t(LɗƔ�}[���������KBB����*�9�H?����uV�~2��P��)�Gy�^�)���.�� %*���C���e(V�}�y���eA�����������,�9��3D� �! Uj�#����)�;��!��v�2�(`��[��u�m(����f���-ucn�e���h�D[<+��5������i�^0O���;�TMLu ��)�6,x�[�g�n��Ⱥvą��ɀ��S�n^�?O$�rR�g,UlBm�E(�v�����*���5�.&�R���p�L%v24d9�m|c�ӡ��K��x2�N�@eq�m��EVp����$i5�p�����g�/u�1�M�����O�1�Q�,=f�(��#!�#�;Saw%(r�@�"j�j�ҳ>� _��2
{��`�JBi!��n&M��,m�)����}j�>i��h��g�q�"!�\�X��Ӣ��=Xg7�t�;+�ivG���w�Q�g��5y4��.f1�F͵
��q�xk3���:xqz)��J5'˭�Fh�Z��3�]�l��v����L�����}4�����~Q�e�%�"��Bۏ�sf�@����@������c�Fg����EA��a�� ���M���o��g��~>�(Yӗ�H+�)�i���O�T/n-�&Ҳ�o{<�S�W�b4�c�A�04�M���'U�H:�B���h�R�;O����j�)q�Е@�"ऱ��A~�5���`���x8:�g�U�j-��TQH�3��c�x�r��v�Ӣ�1���,�}��!�Y��#�����|��G���{~c#l���P�?�Kpt+���,ߣ�ܓ7Sm4k��;�?���y�!fa+�<�)��H6��A�x� �
��ov6F�d�$��e����4�"#�N
/��A�!�����=	S��TM���
8i���3v�!M�6��q��u� 1��Tӡ�j��Vz��ԺJjŝ��̉8zɢ~�� �nƂ� ���\�[͒L�:+R�u��5:���iu�B���(��F`���>��Z),���"��בF�mxP���y�Jz�D^큓�7.�Qm���MS`�Y�JF���y��ͱ���i y$�46�KI8�h��˹gE�V�F�Ch�P���b�~1b�CFoM0'��gI�$��*bXԞ�Њ���4�h���\ә���0�xH>�?.�f�!�2h���e��]]b�cG�<4ӓt\��@�[y}�]�(1?�B�bJ\�}�=��WV/��{��}�9H������d��/����b���iPO���-����o����P���=�(6�ƈ ��F�$y�K1x��jgz	�AZ���6}rP�y=�t!~!����/��A�qw>�4}��U8�+�z-;펈T��$�ܴ�?�i��l}����-У@+� Pi��	�*E����6��f\�eO��a�Y�E���N+��M�+���=�Ͽ�⦺�Y��9$x��쿎�#;���K�*�8��u����ʴ�'�$������p+sa�]��4*�TDk[���B��ޯ�h������3;MO�>�[������<�,�J���Z{������؃%I�����kEx^�j�b;�ڱ��Bu�w���[U�1����]�T�?�
���$�,���ո�p}��k"��T<?5`�8�?�U�[�ȼe!K��d�-`;b�I1Q����{��٩�ཕ���O���8��&>�\�_m%1�uo�h����q��⎨Ŗ]D��������V���?�I��p�$^f(>���Q�B��9��g^	a�ּ�q���utF�d��ǂP�W��L���r�U�	$�� �1Kw�������z: #Et
�Q�;���cUXZ>)eL�,�tak��q�2&_�Xoi���$dO�fM͗�`W;2�@�׽O�4W�ʥ5uiM{)��X<�Mݘ��4��T��c�4�5{��cԭ���:�
�ÑF�u��;M�I�^'p�R1�@P�����U�*	($�Tq�c����U~c�;��,�R\S8_�b�"��w��:����A�%M��Ì	,|h!C�'���j���Yb����-����y���r{+��	4ۊ,�
�ؑ�Խ#J�5��`QJI�P��\}���XiY�1��Pv���72��&���k�7���RW/�kZ��y��{X�YY\11�V�I�[.��=r�Z�la���1�NjŖcN��xuR�͛Jb��a#��^N�?o"����J���fG8�������ͻ�%�zN�����5�c�)����s��_;&�
AA�yl��6h�d������*�hk	�V�2"�/���٭�`���h��dMTǲbڻ$?�T��	�E��H�;�iaz�;s�W�ͽA1��-�-����?��<Fw��BP🀍���D gt��w��s�/��m�� ��&uO(,�"�?t�CK1���`,�T�吽���?�T�}�ŞgwJ?; `�x�F?^�D��4V���+���LY�[��J$"�>(��9�H�`�,������X%:7��d���O~��%wgD�� ���`d��6���e�[8h!��~�-�%����b��Fnt���� ��6�"�H��7�����"���N̉/�&65,�9� #T��o��<����Z*Ǥ��d�&�b�=t��*�m�����0�K���	EV��OJ�q���C�ɀ�Ws��3�a>����A����8�y�.^a�Z�"�&����>�n�oˎd+�pW���
�qS�J��4�ʪP�^>n #�v*��Mh�y0������ٳ~���~�U{Dn��\i��7ݰ���d��������5�������l2�F���>�mv�g���`:����e�����bLp�ܾ�b�S��Ԋ������-~Õ@�BBD�w�/�D�L���7k�wQuaC�� ��F��k���=��Ρr.�(⦤$����V��;�e��������������,o�N'e�����5(&V�,`	��zCXw��!Ylt�~����x���U�S%�ټ�P��;�,��߮���䟩i��5���8n�p�n0��8h���9F�11*R=j�N=t>ܙ��xG�}5�]{s� |�k�/����V���;�aP�>��ރ���'��ʥ�d�����e�@nu�h�V�pbh���̹x���j3g˓�6639]�>�6�E�˔�/�SܠJ�c�D���$}(b�:ř{�s݆WI^�ɣ|��Hă��y��!�D]�ԅ^jN�|b�����A"6<�����eQ�����x�'����6kCǕ$�� Kʣ���Y�E��}ja���y-�MpZ�y� em���������&;ν)���_ib��"5�|�r�@	/׮HW2����Q5�*N{{�m�4t���e렐���� ���I��Ol�>T�BK�ʚ+ſ���w7�Q~2y�ƧRs��c��$yN�5�D��	~4��Pz�.e�b���s����SE�E	LO_��#�F� ������q�N���o1I��B�ޗ��r�p8��j:����a��Ag3݇ �,�=�߹3�x�*Iث�� ������":"WX���J� ��?����4��U$�j=��R��>T�a�_�X��"��V���ףrG^+�B���{#��xYt<l/�y��$'Q֏b�L¸��i��������ʙ�%t�����d��2��Գ�g&�c���X�� ��4� �ݚf��\46"k'���%�������j{��t������{nQXHD
�������ξ+%�'5(���6?+x�w�P?=Q��_��>V���>m:��S��%��f��u�n��~,� ����¶�麂uB���>� ���I��/%K�Q�X�.jث�#�M
�R�`�3��R%��bg<k�v]M��L	{��lmRk����0���z�����$�T��[u����I��L#�@$��$���b��&l���]��=Ɩm��["��L�� gH�}5�� =�ݍ�:�<�#��ϊY�S�}p��ÈS�f�X�*�e�l�i�d��FX-ܷ �b�����o1�9�^๳j̥�:g;c��t�X����"���Ƈ�=�'3
���E|�Qx\v�Ƨb5�SON�GwŻ�Ԩ�5��oq�j�6*>�� ��O�Jħ�; ?��',�2�"t)馺nQ���G��0֣�����325���&��T��0��6�X}/e���E{��Σ�T�=׿
�_Vk��v��~� sF{	��3J�
�����<cl�A�<N����a�<�T���RT���D�
[Y�W���S��k;�w�"�̙	[�wY�k�I[��88�)���ޟ���j,��,y��*:���^^z	Y^x���Ô��Po����j��拝W-?���/���WA�������~�FM|e(*z��\xK���>���N�������4�{B%4^�x���	�s�{VhA�G��o�t)r�����:�����[	hX���2����Gs��XK�<.o�NBy�h+X�t��
��qq�r�F��,���.u�������/Vu���?�x�5�8i�r�����΄��u\͈�|ԭI\q�������5)Ҝ��f �I����+>�)8�s����GХ�P���u��T�&��~Z����F,�F.t]R���ڴ�֑b��6h�RI��dw/�gRkН���	s�,��:`\H�j�r�zgz�%Ld�56��ﴅx����q�i���/t�-on���%��B��d���~$7�ff2r����P���j�_+QG\����(���� ������/�Z:W	��}c/�{�(������%),�К�ˏ5�����x�����>����X�"'�k���QBκq���U����l۟����$��h��%����C{�%nsj[�v*���柃���_{K�*���@}��٥�~X8n ��qm�׹��u�2Z.����H��{�D�}��R�v�CR1�GП�r���K!j/_CΌ��'/-T5-	���Z�e���(���r�To�G�rً���ܷ"T*|��]ۑ���Y��f|[�X��- z��i�x�#�Э�y<�(��*3ȱu��̂7��ʦ���S�9o�ݬ�@QU�]�<�aj�/'A�)�c�U1Z��b>$<v@�&�B��+������Do��� ���^%O&e��[���	u;q4�,ɻ�-����z/=�������t���!>sg9 �Y���m޻Pr�r�#à�����J�R�6 ���ZOP�>��b��5Z��A:]$��[ҕ�P�E'sz�C\���E����ɨ��oN��M���{�� �q$����������\�i�g�o�Ls\H���!��,p���"�m<p�����12��?jdK�� *��`!��cA�!+�;�n���,���[�R����u��+����w?��W�J�* R�3N/i������'�{G�q�IA:��ζ�VMn@��>�V?�Vf�Й{��zLe���#�=�Z#~!k*�{d|ѪkOA1%b��	��VG��R���߄4�cjC0-�FKQ�>,�_����H�0���"��.T���:ѰU�/�T{�@&$i�_b�*�Q�L�L����ɚ���,7`"+��*ܫ���g��.;6��[���է�/z�},�ꎜ/o�����	I����1"�S:�����y�]��&lXh8S��u�S�h��V- �"?fS#O�+��ղ|>��F��'�5��Kݦ3��R�����_�y�j�!�a�u�q�LX��[hQ��[X��p�݋�,X���
����G{���D9_�c��U��6��8������
��J�d�'�m ���C��	]QK�&g��
�$��9!;l��b�0�Əc���.r8�1W�����}g�=�mj����+/���c�{�߽�0zj1C���[K?�G��*p~�:��F�^����1Hpkq��H�ո%���u��R!�0��iւ)�F�����g�I���z\��1r9���y�����6]�2.�-63�����cm��<
���|k�D
�F.����:���A��$��ٲ��(�I�����\]���<�Gr�����5���c�O�E��̏?DmT$�+&G���J۠~���<g�$p��<�~Lg���;�$E���{y��G��Ӛ����2{/��,�F �Wb���<��E
�Mr�F�b'����9�<�i�Y���Y)�'��ܧ��Չ^�Pa 7Mg�4Qnz�jx�N�ۍ��w&[ma�^���t�)̪M�Vg����@L�6 �j=~�|�[f;�KD��Ek��9��Z�P=������`O�L����=-��!�u&���xs�ݺT�`�F�z��97���o &�#�rmh|s���uy��H�2����
�![NKz�Ϧ�̠]D
rQ��:�n�p@1O���5Π5����ɒU�ކHK�G�]d&��s����:�YBk�p4����"��i�$Kc���@��|�����ru~�k�5�?+���~�D�x�D���� Sr��6���me�|��]������KltndH��|ݪ��L^ Js!f�,Ǵo1��<S�
J��*9���_����e���4�T�0�2	�(��f\oM�#Tntd1�;TұY�tx��u�=����h;����G�PmA�����ڔ��m���ʨ���(�4!(���u���)r�8�-M��`�qe�g�5j���8v�Hy�t�J�f������G���\��]5!�k��$�vmtY�ݜ8�?�T�����86��׏���f��gWK��Ї��(]�\���M���+Ć�F�U�q�C:��!z�/#}�/ [s�$"1ދؕ����8�!���#��|[�������>1�J���Nz�>sNE��B�Y\r���l�(���݂��?��8��?f����|A	����<~��'�AHO���J�^ϓ�A��=������f����.��4j������|�����:RW!��yi�ua6 ��![�@v�L-��5�~OX]9Z�9|�����|�g�͐S�:λhVC��ց�]8���%�����msU�<�i�C" ����} ف�:��~h�e��'��˙߲�㢷���I�i���N%wl-�]/x�2�|��S���J&�M  \�4�+8�O�5Q�|
�p���'^��AQ\3�H���ȅ��*�A9UO+��T6*�L������J�!�	 _!�,p��B�Z0����@a����e���5�<}�1�3�?�5�4N�|��rU���gF�_bS�y�Ǧ�T�_
�~�@�Ӹ0E���%Ȉ�(�@������ B,v񨗖������Ԇ�ʶ����Y֤ft�mO���KS:�r�D���c(M�@��d �i�B϶� v��@��e]��(�p�]���y��@�5�^|�����vg<R8Y��b Ye5������c>9��q�� �ܴzl{��H�|Z�T�Ph�,��~`�����v8i"��ͱ�_S�b�)���y���mمWe)q1��"�Ľ�����
���+��?l�L|��Z)�{�J���p/5��C'/��ø7�1ȋ�(Ee�S�%�h��5�T�q �� �[Йx�bE�e��
l�N�b�e�˪��h���MO a&�/l���H��NU=�hXL������Tz����RY��O3x�=�_�=$rs�^���2<�u%�p�J@�v��i��V��e������g<��U_���|%��Ĺ�L�v��N�Ǐ����ێv|��&��m�O׭$s�胞�
hD.��$y�w@���o)Lo�{���z����s�o�ˊ��F�2~�����7�Bê��"�0o�#��M�;2�9+z��兏9�Ǉ�����5����y����c��K��z��t��-t��J�P��Z?G+� uA<�{x�8����t��ɮa�cdpȱQjH<��&a�U�Rοc끻sݕ0�7e��Yt�e�L��^j�9*�2{v)��Vn1����Oa����~�Ha���u����Pu�� ���Pҍ���QHʴr�����Q�I�_�n!� �j��
]�ʻ0l�L�U�_@�nm�����Oj�X�>4�Qj+��l�-t��E^h+�:@[�CM=��#�F�ܖwG��+\t{�-�W!�)���~h�I����,ns|f��?�%�\|j�T���Q �t���7���ν#���?Xz�U���kn*�67,� S�	�s�����p�����̈���g:��7�G�wO��e�FC�귫�i�8��	R2�S}��{�S�K|FB�o�������e�1{�ԛ�p�A"UV���0ƙ�D��;5g��%�[E���.��0n�����������]9|,�ȳ75><S��䎏�Hʊt����E!`�L���@l�s	I���/�����B�ue���2xqӌP���/���T���Sk0�P	l3#�c�R+�D����Fܑ���xZJ~�����]��5";��_^��� ܟ��"j1cÅ���<NG]���攐U�-v3E�y,Ǳ^�'��JET!�O��h��_�qY:��{�N5�s����+�h��HrYG;u�4�������+�j���gP�n��C�	�&z�-݉G �ϋ)&�d�[K�����1U��Ӹ�P�|��$�m���6Lvp�3��p�$er�HI>�0����R��i�:k��Z�`tǓr�2F}�qĎ!$��Irm�{��%�.@��`�:ϗ�Mx��j���(
z��jY�̨����*?�#���A�r�Io8$����#��A����ߩ�)��d�2�|�X���z���0��`�9Tʲ�����S�����Y��7n�,Ɠ|2�f���@O�;6 +ebL�QU�<��w6/�G�Z�Z)���oQ͟�xHV� �Sa�
}ybLץ��q����!k��=Dͤ�����sF��a��x)ii�5��8��l���3(4k gb�e|x�ƫ2n��=�y�)(;�8���̈́P=��K!VW�a�|���5�}�gD+��L̪+I�H�����6���gO ��})Zq��B�(]^
��?JL%���NG����Ή�������v�Or��z���[**������\Q8�
�H���'����Щ��߫{Q�"���~��J� E^얘�Ӝj�P��<�$h���O��ؾ�'��v�mR.�)��ݢ�"�M������2� �2���3Vˁ��À-h�辐ވL�E^s&'�/?h�(�arA��q���:���&a������p�y��<��K`o1ӵ➥��n���X�$�����y�\�ty�.i� G���8�A}�3DC�4�}+D���h
��{��jq4c��nr�)�X� \4W ����D��� �������p�A9*�rKHd�f�]r`��7�<���(`���S����G����t�
�f�.�AXD	O�DY'=�ѐ��."~�ou�;�I<)��LS-v�YùP'�-�]ހ�I!���4�% L^�NO�dz�K�u����~��h�N����1_�����RT�9zT�kPtXE���V��2;x�l=
.1ì#饛��8J)�|ta]��4���t���b���'II�PK��c�ϙ���h���s��4n˦f��M�2��>����7��+\,�9&f��1|d�����K��LO�,ye���˙�w/.LԦ���t�9��w	D[o�l�ez��q*�u�i�ש#�w��Uu;����fh��}�zgC6����Nt�J�@
"c_ۀ�Ф<4i�Own[�w7!:��S�M�E���g@±���ļ_l�4�����Guo��$��M��"��������6 H^��T�vT�3���r�V���/�S4�4yu�ԍ���Ą���*@�x����Rz��ʉ{P[F�MO �d�jn4Pq<�_x����+\��T}v(��+��E�N�S�&�-,3�xRR-e�?��t�?)@�"�Q �Ws�$�	�;r�9S�@�ҵ�G�a*�	�(ư����p��t�=�	���M�^/L�(����]��n��D�_���	�Ї|��V$��mN�H�ab/�1���m�iR�'���|O�V��#W�t�M.X�ht뫆ł�L���a@<�N_h3Sĉj^\�<��s�����v����;؂3Y��\��</a�lY�����Lνa8���"l�s%��c}`k�g�4��m����PW�3ؖP-��]�D����靆_�~#8�Ã��ӫ`��Xm��6(V�EA�YQ���K�R�=7xܮ˲߅n9�^��<�K.�gQyBİq��'�59q�;�~��g5���h	�����Gl�-��������M�IA����j8�m�i���M<S?�8E:�N������1�5�h��_wX4���{��#,3V��W�hO$�L�&�f5�P����K���ϻ�V�ܭ�l(��}3,��Y7��ĵ�s(��L}q�+�M�����段t�yELT֕p5��������eX��ՓB�c�U�c���`
����@e�����(����9�ؖ�'��럊�J���	i0��;��^�<��#��`Vg�14�����o�
��-��3�p��+8����f*��h'v�b�+δ��+&��D�2y5�Wȏ��~\>+��ﮞO�SU#����K��(�
��M�Y���=q_��H(��ŠN�_�A?cR@�sAK�πL�*w�x��,�hF� 
���\Kn�2.c�	��ZmFq]<��`1{"4�8�X,q*��ؾ[�_|��+l��{�2DB����^D�Ui���ڨYr�~ȉ��T���;������fV���l�ɽ:=ʫ:"�F3��XTs��x���ց�d�b��mx��ϖ�@N,��r�^8�M���Q1p2�lw ��$�������!CA�`�|?�ս�;<ږ�$]�?�(�.������B�� ���C 9%����
r�Jf��U�G�G'S�<�@�MR?�F^���#�����#T��_�ilE�jN����D�8
��:�J��e�g�����̳
�-�H��]4�k��_��� ���͘�エd�[]q?Y�������e&����O�'�E��� 6��1A2A{j�d��WI�rӀ��t��b��$O�ъ�B>����r�Z�L/���~�E8��6#<���u'eAt
�[�M��8��:hQ!��O�cW,#��b�`�YS���*$���� j�O�R���l9�l��5"�`����wi[��sA��e4hg�^b����%��Kc��5'V�;f)"A�~��PIi�t�:����8�2Yϛp�XA-v���p��$K��'9�xQ�;a�{�J�T�_��n�j�?�ٛ��j�.򛹽6��)H!�l���"F�6���Y�����籎�Y�����<������$�h���Q[3@?uVwZ�3#�x�W�C��P�bȓJEؚ©�I�ެ@�n����܊��>��EV���������������FR�s4�$�{~��,�on7M�xʲ:� o)Y`������$V�<.��G+i��zw�,l9sp���j��ˍ��y��7�wr�\�E�,I�]���d�p���Ak��s��b��s;в�9��O(�$�/ܭ�M��t+���A�J���+����yt�S��#�k�1�Aeͺ�BZ/׼.�QN<�}T�4k�2ȾJ-V4������;�!��_��t�=��b Y�r�%�r� ��3vR��a4gP�&��4��/���9��q�(��1�w7a���Bѹ�*G����y�N l�I��e.����|���9��ڀBPj���سC�4��5HO����OwNA��	V)��(~��3�����1�r��%0�}�Z�����+��b�ۇ�R[!��&걟��C��"�e��7xWgC����
���Bp/FD�A��ŘO&�\���96Z$?��*bg.��y�lɬ�����Q|�����R3����P
&�C���:�D�����������I��H?�����>�3�8hq��@��ס_�0
.�aƾ	��{�|��ǵ�q4FΰT&�N�Hn�� v�V
���S�*G�fH���%f��Jsy�`�Y���b[�p�#����u[ѫ6Kn�o.�D��9���RK
�1����ú���Rf�F�>ݴ�#���!����8w�|$DSԆ�"Q]�2NM"��.v��^A+�����r���ܡk3a��)& �,!{z[Q0��#K��@�P��l^�0�p0~�W�9�JY3�~����ʰ7χR9)���ǒ�����ٻ/
�R�ҴH�=*�aP}=B�d�<���FX�J|������4�.\���:~��;	̙���l��V��ͅ�� �����$[��][�cJ�N��~/,�a^;H�
E;�y7eUp�ϩ� ���}^ylۮ��M"cƎ�*�<��npk�L�}A�a��M%c�_%&Zυ�!���
��H������텳z9��l,1�Ս{;���,��Q��ʹ���LG��� LH���=w;�e���	ߗq\|I�
@�.E+���\�f#�ڸg�
cf��8�#��K���C�����|��%����ĺZXK��� S���JN�P��v�F��Yҏ�uRA/��~�'�+dP�ai�5��u��?鶃4��MC(�r0�=p-2y-2�3�l�!@���559w�D8��͋�l
����=-�� ��(ˣ�����y\� 5i ��٬��{) qip f�����J��8�6����e/���_��y�k�F }���1,e�*p��8��hc��1�*#L�y/�_��J�;q��e>mY����ɷcc�K������������c"��<�x<*��>� !j�	MH����m8��*�h^9E��'o��-����'�	H z�[���42,�G��"���t�T�)��٘R9����]]�|pL"��6��I�����8�K��<�w���Ѐ�8����-i�3�l�PŴ��DúU���7rC�|l����7�఩���R�`8Ga�g^��=�e�W���ٵO�gBr�R�m˄j���t���x�=D�w���FN�4�CK�@�������9e�K���cKZv��6��.§.|K@�e�"�|���o|���6��6
K�����XPh��	�铺�x
[�]L~���ߪ+�H�y����[4�<� �M����c�eO��
4Axd{KK6ֶf�<�����:*�dq����\���� .p.���"2���/k�6�U튛Ѹ�3�z߰�N�ܼ[�i��9|7|�;�.��"YK@U2��1�:u�T-��ȣ���#�-u�X!@ƶt��v��C��O����������C&�� ���t�JSKQ�Y����l_�8�Ak��-խ)�p( iX��H����8�s�v�� �o�iRA(��S���ʃ��.:v�S�T*R9[	�UG=�\ǻ;�����k�B��u��[�-�ݷ��Y�T��>�Tڄ�r�W�� ����%���&$Q��H�El3S��R��aה�����X)2b�JuJ��+�U�L�����̵k�qYG�̠n����J!�V2�.�(m�dk�=��9Υ��iݼ'�pt����=�����*�׍�g�I�Q��zD=�����E�P��âk����*tk`��h�٧��H�U\Y�?~b����Gh�]Ȃ��1K4Oo�Y�ۢ�������a��̃u��5����w��R�	F�Bz"B}c�}wVWO�@V�*�(�_�J� ��ܟ�,��0�6w�\|��c��h�;�������P�l\1�m�J
���P�������DoW5����q#�@�:��H����]H?�
����9��t9z�YI�<׹���2��j�V}�o�yd���y̽&�-D-����LO����9���9��`0�}��`�cule�V�����4�#̞���㐀�Jw~�wx�d��D���́�N[��}Qn�u8q�)��(g�U��2��Pց����qdo8@�x�`<�JZ��܊�a�5��$����+\Y�B��4�j�[Zq�]��#��ڻ|l8�O�uC/��Ի�%��(��Lnj=$p������c�r����������'A0�����|pG	qK�� �rJL���;�6]��?"� >Bkd D��K�b�=�=t*o�P���M�N�O<Oxa��rOݜq��� �����;(jB �����B�d�\�;7I�����B\�)�m��<k\����R20�ȵ���0w.QR��)C�pt�E���VA��m�l�R���u�Kc/Qlܶ��{�������7+#kl.Un?�+_��r����nA�j3\_��2r峇�*�Z�c(q�uL��M�4���1��6�j��z̭ �ES���d�2�3WLԛ�pQ|+��pW�r��y�ּ�����Ξ62�,,�������e�ϼ�A��K�S�ą["��c!W�-C��Dɛ�~�)3$�wɑ�nuY�{�Ö�M�є�KB��;��G��eе_�+�uk`6l��߿�/�SiA�Z�{H�%���K&�]�s�nd������Bay(E�yt�s��U�/��k��O_ �E�tz�=��knG�L��便��ވ��.�B��G�y�D�lw�������؈�:��̤]U���M�^Ps4��"I��iq��N���^¿�Rsx����6���3��&	eOAp�G����n=�Ͽ�]��O,��9�f�p�4��y�m�o�ur�p"�Ε�Bh��|p�1;����\ˣ"����%P��c@X F�s��1�R_e���g��K��'��������׎�N��TS�*C�m�n*F�.��4���a+�n��[�].�e���RĜ�ߝ� �bw�s�$�>2������?�U�#��:�I���'�«'Z�-�b��plX���Q�-���Dћ+$7DT�nTk�6Zbb��F���1�f��$۲�ɛ����h���*���X�"�fs�}�U>�
��3��X�0�@* 4 �����}�>�Ҷap5���=n��/��%?͞pu�V�
m8G��9ɇ��yBL>ԧQ���re�	���/T������T�Q�GS�́�5Io���z�f=Ua�c�Er���x�dM<��`vt�e���hB�:���,��"����(����T��_G�$��!(5@��v:uNT��:�j���%��U��w�(��c\�T�&#�oF���P?ԋ%>hڮ$4�v{���͸B��Un��>~� A,�[#�@(1C�	�����Յ�y�)4x��0@����v�u���1clzr	�d��z
,�ڃ9�hGBw�f.r�	�	�x�H��^��A㷶�{M�*=��fQ =�Yc諾X,��<�Lʀ�X*�-�*���yT�Fn%�A������)\q�6�nAǋ���I�(ufƼS���EP�L�]]�׸�p�D)R�$�z�Yª�Y�6�@�v@Y�#�Fb�ҋ�C���^>m{G�E����z���Qpg�F���͂���K��ڷj�����3w�Ykڔ����R���bWҮ=bp���ҽ�{i��C�������^�TA���j�x;�.)׻}��;�m�Lfn�����u�|
��p��)k�A�Zf���2g�~��\���"������;2�6� �v_�6$��M�J�w�7��u��pP�}w䖿���G(43Y}r���!�2O;���=`4�>�Q�V ��$sQ�PW����:D	Rg�3.:R��.�%|_���b��+�������zD���5W��H��Ѝa�*u���ł��W�^��-�$�F������d�ܨ�H�p���os~�~h���X"$��6}I��TAo�b�W��t�
U��a���=�]��~F6��t_��$��yGD��ZU��A��%o��ZuU��a���G���8�I�?�@p5W�����<��.�5"�8�����?Q�x/I\�ʁ	��!�qi�;�s�H&MsxG�H�@�.��f�}m�'�mTtol�.~���+6/�2ک���E�֥�}je��1�Q�O��`��B:�!6z��e�m#_/>�BK�@o��Ă��X�T-�����
�n�����#k����$�XI���=ǣ�0��7{�ȋn:�.׹��O)!u�@-����'W��}�<��T'-��WO�рY��4P��M�b�^���)9��6X�4�es�\���`7�)	�~�g+��'���'(] ����Xͪ¯��8�����y�A��{�l�Ɍ�Hh�|�e���ǾO������H���"�5cՕ �G������bTb��i��}��n�exN��#�lʼ&)��|�0Re��xS��|{�+R��'_g�<��K�>r��HqjC��I�_U��D%��󜖕��z���	i�8�sU�tF�I��nP�VtJGUpr�T��u�QB�KLp~���g|���ԺE�������ǿ���W����$&�6���-|�0<�#�3*@n���ܾ&cƊ���� WB8dT�2`9�P#k&���	��=Ai9фKN�]In�N��'i/�?�X2y��*K 8�5 h���n�#�q�I1U�sؤT)�24����;����j�EIw��'���/�al���[�G��<z^+<~�|�{��l�R����Bk	VF,��2��@.}BTF갚�∟֙�{B=�Ӕl҉݌����>m�֎��[�i਱����4�1&h�r�mX��������F���ͤGpa��
-���:$sۂ*����W�%7����EA��
G#�_H�̧�U�S[����y�Lj,�(���n�:Uc���j���/E?
�S?:��9NC4W���^m;O�8�S��(�G�xT���8N�?e���Å���Z���q�`QVy��ş�h�l����]���f�ܽ�sћ g!��zs�'�����5{�V�d�Sw����/������"�r�%�1� �ӏ8��R!u�汷O#�s�����]^J>�l$=�P��Ml���LdiM6}�T�B�=�g`�ͪ���s�YqDf2����dV)��^O���}�k��H;�X=}�@`Bz8�@�@����gv�-f0n���IoM̕���S� �*���J�d�,ӹi�е�	u&z~�,1���$��3���M���.�|-��5dʕ���je��0�I$h���7�Q�޹��{վϒ�˵�)��|3����|��.��V���Gf���&��Z�)䔲�B]|ᢢG�p�#��O%#f�]i_���lL g�.���E����ڰ;9Ȏ�1�i����%Kً�_Ό�)D��b��M����g�$M>T{��p��9��>e�v��,�TG��BI|�A��Ė�.Z
�ŭ9��cZ0���a���T�ÎG��
���Vf�HrE�3a
���G��ĆR(~�Z1��8��fe�hs:K���������,UjE�O�ߐ�)�9A��MVQ�z����5k��?�9�� ����L�D�{ئ�ل�;Cܒ8il���C׌��'cnyv7��*�(�퀰�F0n@f�ˁh@6�ʚhsԌ���kS�m��]{/��3�x=8!ت]���wR�äֆj��Mn�̝$k��
�����j��Qz��
�U]�����z�S�6$K)���L����)}��(	3�k]���'��_{�#�W*��P8��9ڥZl�;��m��k1
t9��u��q.��O�m�AƵ�Yˋ(u�]��H�Ưwm1�w%�7�	TmN��b�R�o�A��vq�8�Uf���n�H����������X������/y+˻��x�E�kAN±9Ӟf;(��@[uT�9��/��eIZ�L'cC=Y^�����Zq`��j<𪗫	=&�Ac93�4~)���O�{�kR=[|C6M&�#�!��ĩ�m6E�7��v�z��X�^U[ jt��VT�ۓ�1>�9<a���y�F8��8�.��w}��2=Fk�
d�̷������h+;彯~fk�S��(	\99���~�+�tj�lmMgx�&΢�-e��z���E�ۥƔ��-�P n��1R�ேt����^��g�D>j%��	W��d Af2�0y�h��� r���	3�?+��b}Y
��dy���$[�6��7���<xTk�Mu�"�Im1�j���<��Im�SI�C���1����ۦT���{t�o��>S_���`�$^��>��Y����6� {�u�P����x̥&0��k�]Gտ����.Zy�<4���^�.tf�5E4E}����2�35�8Q8^��6�BJ���5|t6���@��2
u��j0�uvֆa��7�~�n`O�����]J�����85�u�k��X˅�F�w�a� V�h�ȃ{�\?ѧ���@c� j�L�y�]��-R:�N�{6J�ig�=���L�֒Kz�'CW�����.��7
%��nZ$DSF/��r�ց���&t�i�}�Iy_��A��)�,ҵ���#D(i�
)��x>m�<P��̕G�Ӫv�*��&h�����)H�}��nx|<%���c�E_��.�5����)��^4X,�8DD��2VV7�θ�����������E�DS.B�'4T��+�0Ec�Ji�Jp!��o�W�����a���Ç$��Oa�r�YL~�=ʡպ�J�"Ջ��)��a���]�S{ʾ4��ִ�`��C�6�y��/+���A:�qT��$�z�z�L�A>[�!�K/��qj�Z1��:�$��������7�I|�|��*����|C�	U$�s���'_Rj��Q f��緥=盫Lպ	j�Z��1�5��R5��3ȑ����4;;��Ķ����)��vOrQ-�m���\7��μG)6t��7<�"_�^����:�v�{��w�zL��E>\�k.s�?�0����X�C~�x朆��G�ci��U���[֞In�']��8�v���w�c�N���܃������ؘ�}��R��֦�K֦18m z�6��h�z4�	f\�M��'	u���|*�w�7 �'u��D�	�
ӐF���e�/É�,�X�'K��W�2���� �YT�݉�BR���^n�q���T�ٵ1h�4�������x�6L��L~R�{:s��e1�<ro�TD5�k�6-�����C|�%�����}e����g+<���w+R��~/�7���{�+�O�Q��0�H���>f�~�I�4~��}7V�Y$��`������)K�!U0]s��qf�/'޵}��9�ۛnw�PT�F����&�A����΁��k�5n�G'pSk����gQ�w��#3�����ў��,�(C��J��'�D4�cM���^L^b���Wh������3w&!zotW��q��E��S��U��9&nP�zo0I���n�+��H��������5�^3I�A�� ��W���,i=��4�[�7��/��UJ2�%��t������^k�P���y��D�����FJ؂��{��K��k��>B�v���]���c���)��=aI?e�H���~C�[�z�s�b7�KI��z'�-���Q��	�Q��&HA���Q�"ՅÃ�	�G��~:�i!�F�-d�Ly
'�$�6E�rǲ,X�ne�3NP��JڭНE
��/|K��M�9�\-�=�j�H�/BZpfz�� eR@S�E���+ID�
�/
��0 ��A���������+]߶O��UC\�D�ay��ֵ&j������s��5Ⱦ
�Ch7��Sf�N��s��p,��̓��J�i�"9w����G�fʎ�8r�SD�@�[����bw�$?˰�,��,#���û�oŃ���e
ΦS	����ʬ ^ݤ�9�o�ÏUN�di��C�N�X��d����}�G	�R�����1~25Rn�������C?ɲ�|<�;�#ES~r�a+w��D�-��v�Ų���;�6dc9�px�QL�#U���{W�bWg�UP�����Rq�>�m��'CZ��R�i����nfO?��!b�җ��&��X��E��ش�sL^fB3�%]����SF���M�b��zoțR�B�1'�)J�}�J?ͳs��ďl�����Bf`����2Ĳ#vT=�7��qޔ����R��tx5���5J�9e���[��Q�@�r�X������35(���ͥeN���/�{#��ڇ����/�u3z#�O!�^ˇ�#_�H�X'2~���=@ �fߧ����.��U��5o���-Q��d��Nث��SA��(�?���܌��~��9��!�C�
.В�7hs���v�	{�<dV���NE��+м�q��]�w�y̅�[MB@=�F�X���^����L�^���+9%d�Ǒ5Zv~�X�p ����+G�BN�JjR~r�C�d�L*���:()4}� �b�葀�{�!wD��j2�������#���@v��}'����(T�����$V)�`���i�KWv��	�� ��R5?//H���m����'���`K�˵ނZi���4����f0�X���}�u0�>.�}���&x�Ԯ4=	w8��&
^��Y.hl`7sr�}4iW���=�ңD�����
2*߯}ɸ�lV��;G(F������4���y��羔1��q���۳�Jx���T���f_�]��⊑��1W��s�޸��x���%
�m(s�A�5�
�x=Mxy�~R��B꤫�baQ��$r"�$�!{F��y��ub��qN^�ϯ/� ��Q����Sk���y%	���1Ȩ��轿U���=���F!�\�܄�w��]Y"��P��u��e%�ia�+	�<`��h���Q-��.u�i6�Ѿ�G��>	nA�����:��k=�g)F��!���֞'r1A���HV�46λ��M�n���iz��}�p�-;eO�P'
�e^�,�jwA���U	�1���Hw�A`*D�Xt�J�L:���O4���7��X�w9�xsOv�̌����)C @E>ȇ��$u#ʘb�8a`�׽֧F^���Ѱ�7�	�5ɯe�"ٞ�j�����2��c��~���Ȁn��]n��Jm�4m_�'��l�r�;��k�SI\����3?�_����|s�Ҿjʴ��Ou��T}a��J-��I��mKA���Q�Fϯ�c���j^�5�d 8�c���%!6��(���M!y��<ˮw*X���4j�wg�=�6�������j	q��s�3�8�Q�/jqb�Ơ
E������\=� �^�I���%Z�gT�� c���:�E�޿[�O�]s=K��w�'�!"��Q��(l5]L��_����3��e �lU�Y�Ee��d"�V"��	/H)a�N����T��N���<e�i`����������ۉ�O73͹4�k����ֺ �0�Z�'=u�w�Ұ���֩����.,"�: ���[�mzu^R�f�;Zx�#�c+��#3]-
q�Z�",b�ғo��L�0P+@ɰ�qxP!>����2�l�4��.�t>͕���ؾd#����A�o��X��F���F��z�m�}�ɺ����$H�����ּ�b������\A��P|D�D�p��dv�Q��h����Ӆ���^���p�sB�a꒝|�=����ߞ_�ԇ$dN����bߥS'|�m��%��j(���O���u2*��v���.Xi���kNJA�YȈ�$��"+I�t��� ��,��JV{�:��V���C�!���.~�7:���Z��2��7��� I��ٷ��� ����VY�%�-ai4n�x�J$�4������4R�qW�"�I�%Dt��4[��L���$d�m(5m@��P�=~���}Q��h�b�?��V�g>,�L-���[���	=�Q�(��X� m/6�>Py-j�$��9�d�HwI�[�%�q�e-����e��]]�Ir�b�T�=��)z������]@V���H��ҕ�g�q�g|�:K����yr�N�¾z�]A��QQs�K�(���h�`8h�S,�XQ$!@6�O�x��� v���if2|�;iL#�S������9�a*J{Y��M�i(3��� qV��麧�Y�^d���p�`����iB5ݴ�9w�k6�&��e��y��Ъ�{x�6r����t:܂<�:#�>Qy����tI��h�Rߴ}s�3dv5P���Qw�#~��CB7�/⿕˅��U'��-n���gV��m0��sΆQ6���]�D�9g�!Lm}$�lV�;�g�V�4�l<��J��z�y �R�??S�d6�g{����,DƫuS�A�li�3�E�Q�s�2�Aը*������G��_͓�Y�����n{B�6zcP����ONwH�vL�M�����|
8?�qzZ�Qݶ��2����J���,=3�t�Y �zhIvV�<_1hx+��!��|�1@H� �rw��A&~�bHA�d��*������g�rD�O��]w�������B��o�=;or�ufز��%�R{^$���*�S+��j�/�~Z(z6�#�3p�Ƌ���*<y:�!)����뵺m*��]�\�/f����R
����;�O�("��s��������YSd:�Z�
T�1߯L�L���aꅥV�ΐ��V�V�D'�S?���gN}��,�vLsRQ�h��i�t���*�Hz��=���MIU���x���}>W��li��k�K���ã`a�3C���b��3�-$�e���[��2�,>���)�Ƚ�����x��SF˸ �`�&�`I�71��*3##��,D/p�bo�b�3x![�ɿEô��s�J3ܘ<n�yW;��u��;_"i)0��1bf�8�O���3	5j!1r7e��]8��z�U�0;�'�� ْ)?^%��ʂ���b�vO�vҾ�2��1fy�&�Pn��R��:�,W=31C�El��]�,Y'�sSl�^�`\���rBӻ^h�7�t�Fv5�7�[9W4�\@I��پ�霦b����@�pbͧDBRs�������3QLo�����N���Qd��OWD�A�V̅�N�v�e��Q��Ҍ��@D�Y��"DW9j��� `��<^Y���8��r?���a�Ix��PS2L�JkS�b*�@v̫��߫Mq�j1oD3������1+@"��b�xQҾ��W��(�d���g�f�������k�Rg�*\�x���e*
r�pp���xI��n�O鍕����a\QQT��I6��%��7U�}���~��ؑri��n��.�bPh�P�Q��*������'x�\�6�p`�G�>Fhz��K�]_�|[1y��^��R}�tO���$�w�R����ì��tU�D�o`����9�<nùOܬ՞G�%�틸z~-'!EQX�犝x�Fc�dy��[ڦG���Nˋ�Tz$}�"�`��ֶ{܈�n$1��jl�X�7��a�^]_'�1�M��-MxO���!������M��<��8ߨ����!�4�W?mw��pH�+が_�f<�c�	]�U�ŗ j�~X��UJ9r�jy����;(�9�x~|���˝���h8��ؽ�n?P��-�w�������n�����p.e/��1���r���������t&�&5T�J�sː1Mî�#����.���L��6��|/�'?;�b�$�Z�ϲ���1��0�8���ҏ����<D�æ��q�69���d?��g����%_=c1u,f�T��Q��wC�p����L���f�5�������e��͇����P�jᾗ�����Zpƾ~S _]B�Ι���<���j�������?񨶧MjP��V�4�j%o�����T�z��}*��E�����5=��T;x���nw˗�&����Ln[H}t�*;m�?cr�f�����!::%�<�s�ΣCo�þѡ�R5dAp�E�	�9P	-b;��i��9"h�u'qr����!R6��-�B����Q�$׈�E=��soZ�r�WՕ~}�u�f+����ɁykAd(���c��?_[m��;P�Ų���P���k���Y(#m�-Y*�e/mu�KN%d���a\?'�).�����Oe�̟������%�iKEɵ��V'C;f���Y����qݭF�A��/M���%� ��+��i���;BҜ��+��P��H�^�J	��[�l����#sAK�/�}n�^b6�2Ï"�2���S���2q���8����GX���#��.v>����i3o���YJ����䇜�p�A_u�'�9qa��;*[^?q���5���~�py�:fZ}��}&"KF׳H�u�9 �v�RC)�6�M�f�?x�t�����-ƅ��6Y"D�D��۹Y���b��nQ�����(���5����%r}�r��R�͕�J�g����5���o���m"|Q:(�5���9Adr��g�1;�2��k[�����n+�k���_hE�SB�B����X���xrW)ͭg��?��N�6~�Pj�B&T�*��f'=(}��ңˣ���2�H�z/O8�� q������9���+��F|���T�l�=��K��: HA],D�O�D˝9�p9y}�x��w��+��=)c�D+�����p�#���k\֊=z>�[1��cG�x��V��"���`o��k=�1�ɽ7U���Pݠ.2s�%u[�	G�q��V�'�XV�������8��apJ�,�g��-�p+:h�ch��f�;�����J4bM�V��zOL����	ʍfS��Bev��A�� 9μ�77%��k�T	(����C6;M�!���#������㤈[�ҳT�l�T�F;�P09l�k?���N�W���T��=W���������#+�ks1
���y@���0�y����iTm����=L}�NX�(
�Oa����jo�ɻ���s#B����rdcհ�����;��մ��Hh��EMU�3 ?M%]/���[^e������R���l8�j��W��MU�v�ir�� ����xa������g�px��Gm�  c:T�h��:	��c�Q��Xc�T.�����k�rb����PM\�S�!#���Y!m��#�=�T�V�1�C4�6���r���b! �)y�j.��R(���0?X���']Nd�#�0��"1���\뼗E?a(b���Vߴ	����q��D��)�f�?.��2K�t�EL���Qg���1�ߣ>0�#],H��v�!��T�g^��p�=��UC�ev��)։�x�60�өWb���l�/�N��v�_*�pNj;��H3w@pa�r����0l���w_�B����_�l�s*q7E��W��/w�tI���h����_��3�B���4p�#�{��u����?l7��?d�_����g%y�c~���$#����u]x��4��� w��������e�Yr�6Ȩ\�'X��v2�
4�L�/�%N,��Y�����a���(S=%(q;�h�ؚ�	��lA>�bP䗆���,��'
�V���]�4Y���TX�G�@|bwr�JW���7�w�f�3߸�W4o�p0��]�E�]c�\�i��g�Y���	�Yы�T����:����/7�( �x���R��OX��ņ:Ŏg���� K= ?̛���&:�]�3�W'w!��qv0��n$�G�c�Aǆ�_���u��ph{���M��i؍�i?e&	2��p�4�u6twX���a��z�M)B�ɖ��O'
G�}>���Q_$�1C�V^�ij�eC6OSh�C��y�l��xPG!��$2�E�1F��G�U��Yl�~j�`QɁ~5,9XiM;vL��d��,�gk
L��-5���oX:E&䗹���v퓴�]>��(#�Cz��+��|y$E�b@�G�
;���T��<�fB�E�S�?(��mF]q�C��ILX�k5;��qj4L�*�3WǓ��HJ�y��g�/$:�r���%��ئ$��3�v�Q�v�a�3��>0�exx7��b���y�����S�,V�ߖ�67B���CR���딜П;�A@�\ �L�U�V=�0K��k�ĽP��r\�;w�p�:5]7�c9�=�	�Bt�5�7��πI�*�$<��q�f�:ߌN�?}H��~�p0p�-�� =m\�7���j��O�o�`B����?H�F�$����H�swj����K�j�7
~@�f�{�k�^M�p�E�V�P*�%�\����� M�t�[���6ϴ8�5n���<Wu�7@uV�(,�����DMLz��C!��6��S�h����ѽ	�5�8�����`�h��}O��Y�}���L�IJ�X����V�q?AJ�[K�tz���M�Wt�{�}g���@��Է���r �V���QU�Ze
~��z���u(�����"���˫���䝺� �!>�Y1���kZ���A!������h�4�D����Ɔ��-����/^Qm��͕���/A#YO�}^�wa�Q��N��Z��PD�*;K�f<����\f���هs� �5�ic�@����wR��uJ��6Q���y�6K�'�<I��y՞�΅��co;�ָ@l��_h��ө 3_�M���1�l?
�^8(e,���9�>5`���[������6�7���GH�s(8�Oi+z\ȏ:-LyRT�[�&G8���P�ѓOB^����[FXf���2j�{���YCf��'LorG�Q�	^$�w�}�1ew}�La�.S�n��(�����mO7�.&@Xr��A�c��������2��)E3u�F���"���G~O.��"�ni���G�Ֆ�veE�>�5#�*�SΨZ�8G�ƿM}�ү �q�I"W��sD����,��A_�T{Kq`�/�i�8�NF5���`��+iEP�t(x����
%��@��c	J���E�1"I���cv��ί����`��^!�VG��g��ݼ��F����'�1 ���f�š*��Ǥ{*�8�TW��I|������H3�'Rȇ�"�0��\37�?u��%�0�fgO~��媲R��Z�K��t\MV˓��>�;���YM{�]�����t�Ґa�f��J<µ��+Kd�y�BԀ�A��`Qz#5y�5D��r�
T!��nB�v �Ki�m`
�o8�]Z]i�UK�/:ʜի�鸣oSeQ�N�o�;��j�"�ƀ������#�ת�(V���:"Lq��J)�Ov�l�ge�lq@6��T��*I+�]IH��N���V���Z���빶(T�>�$��M�_q:Y�Q%���i��]D�ؐ�@��1�+�� ��MܑW�	b�4��sm}��<����V���b5�WPJ������lR؃w_����'�,,dH�"�g]W�˽�E�T���u!�D�dx�nk11Ȃr���R}y��i���`�N��"�4�
7c��W
ÿ�m��)�9
�lP@����)nQc����T�hp`c�H��m#�h�z��7]��.�jVێ$�x��h�/���o	qNu������{쓽|���+/$�O��A�a4T�P��}�i�v�@*G��O�l4~��ٔסW�5L�uE��H���ެKu�D�D�������¡��}��>+/���>�jb���r��l
:%�.jG��	�Ld��5g�݂W��W�e�ϪR�R��$T��,Bf�ASM6��,ĳF�92�ˮ>���5pƿ�ʉ�#E_1����(��dn����w>ܪڐ��LrXP1�x�f��C���@jL��c*�=��!B�w�z�è)��;�ǧ�鲮i�)??��ky���j�;j��t��JP��g�m�2�,��Zfp&��{��p,�sG�^�������Ivsj+&'�P����q��L}/�V[�_�כ�;@Z�:>�m=�s�/��
|�zЀf�w�0�u'�Wߵ�t 0rd�1��?=L���a%s	ع;U�"�bc1�W�zW�IQ�FN�Bfz��x�*+�_�?ϟ����;�ۊ�a�KV �c+��.�]5!�l?��=s��n��R�`-'��N�|HyQZQ���� �EJ��Ô�u$���n!z�F��6�<�1Y)�q[�`�Me	��1n2i��u�{\���ks^�t�k���Iρ ys��A�aZ���X�V��i�o���jU��������(�k��(��GB*W�e)���'�cV�`FJCWl"��8�����+�'������G��w��4r���<63qZ���x� >+�I�-�dA	�4�)�ҚH_����C`���L9(�Sf�s���:o��������mw�p�{�dW��ݟ�/��>�ګ|r�e��|V��� �I�*L���Z%��RQ
D�dY�JLg�]{�{��Qt>0������f���<=9�/� ���a�|��pp)���V��6-�`�}�47�e1~�D�M47Ȝ�hO�Ź5�6��rl���q�����(t�wp�;k�P �̶���e~�C��OWm��@�2V�y����ٯ�c��ξDä�'z���n�	�Ϻ�*��4w:��l����gj�� Է��b\���� Z���q �2jۺ������,%�|�v��j��;������xGm�לg�|�|���2�k��B��Y�{��6�-�2�S��4�(GL�yY�5Qj� Qs��Fo9	�Tf^@�*�����v,}ҀRk��z�w��l 8�;�~���o�dbT��
ڣ���{aL
�/�H�E�G�Lε0�)���ҭ��{9^�X3�*�[T��nH7lCc?=!D�/o⑪k�k
�]>O�˸|��Ah# jJ\�uI�<^[����?x��g�z�?˞JyfF�#��O��N����$(�Щ��B�~pqe�A�HxT},��N>~ݥ�yí`��FJ���WTw�Ӱ��;���Y�(�~���ߋSǛ�,=W�{p���"Dڊ?�UD�.!,����y�����!#���U���3ꠉp�s��-�����0�s�`i���k�炝$*4u��׍�#룿PϪh ��h�F�x�C��i�|��[K��	���|�8x��b(�ֱ5-ڛ��!�aC|f�>�{* o��`�Ÿ}����o�����z��c��^�m�$OdS�"a�хEwD2��?��w�ه�
��B�dQ���F��,Ͼ���fxk����_����c6T��7<CeǎK8�P�t'���K'h+_�@�.?�C�m��
I����m�E��%�}�<��bj�d:ƂE��Py
2��ul��>�S=g�B���Ea�>��*�6a0�ԃ�)#��œ௝J6 ��F��k��'��Y֪s��������k�-X��'*�R��U��%z�ڽOmk	ͤ1�Q�]�XH�Z}��F�dp���<�.�:O���҅�������Pu�/�,��s)r���Ҝ==>��Ѡ����#�I��HK�\}�!3�Y�dT���n��1�G1�T~kD'q�|���,9X�r�.+[9�ZǛ̚�\�zg'��Gq�䧑Yo)_�m�	C#g�����)����K9����v��Rm��#��J(�'5v�!2����\�/��rL�?��������������t�D���I����]Z�1bZ�T�2�sʬ�¹��-�C]$��1E�rW��hi�!yd�5V��0Z#�]j�K�R�I '(6c4�5�a'W���i�Bz��qX�ɈSS���^��V4�\�u%#�N?9Z|Pٮ�ĥ'�մD��)fs�!��?eە���׹z1N&�;�3����e��g��z�7+�&,0B��A%���ƫ2;�oI��Uq,���P	����4U��nj��>�5;�6iצ<�R"�=g"Q��
D8O�cw���'��J�si�!M��#�� �*��{�
m��E����T���q��<���zd�;.�=�x��EǊ*+�n<%�L��4���}(u1�چS�g�f���_7����Q�zN��o�1��g����x^��)j�!s�2��^TGE�
<�"k``�m{�꺢}�ќ,���-�\X|����RA�r��7@�~���_ޏ��5�Jt8���V)�#0|!�v�-0���G�1\�m�������ä���xT
�ř� ۘ��)��/c��sƲ5�Pr���t��S�d�� ����&yg3��g���������+cmtC�����K{O�1uz����; �-Hh���Xw�0�Q`�(P�e&
�e�٘�-��7TS�]'c���'02���A��Y�όTc~n�p�`R�K�7��L���Iv�:x�:|�H1����GS3��j��M���^�px�H��-|!*/�&�[�%^�4ʕ�nUV�á�R�3�Ds|c���\/��}��b�bt�P?r՘8G�17�Ֆ3����>��_I4i�%D-X321�k�y���5�l<A�9�ޘ%�ze]�Q)��~�IGmHn_0�O�L�,������a�D'Y�+R[�:� ����J��Ŕ߅^�F�&�~�D�Ϧ��A�F��S�{�QB�������a�E�*�RK��%E%S�k�E����ŹN?#����g]����x�#4򇿟)��R�",U����6�GϹ�
G��#n��dr@����sݙ'��|�u5�om�{��)Hf`rE��i�����u���!,�N�P��F �?�
�Y��}�.� �c(>�b��&������z%��eN��- -7�ʇ�
$�
-�c+])@1zG��i\[r��#�e���t(1�����Z�ƀ<��U_�=dz���ɒH�@4�l���@��ӳ9?Y��I�쪱��[�TG���*;-n�Æ���0�B���l@�; y�.��`�ȑ�w�An��kv�Rİ�Qqn1�·�����+c��������Ƀ�c�!�p�@�����ͺ'?3�o2Z��6.��G��v1k�%������/̱Y[#��x� ���
����D�#��cԚ8�(��3���seuC�6�̐m�E�����J����T��o�$09-�Z��U ��8����bl��:�X���̡WPS�}�LDLc�n�ґ�k<Vפ8�dVˈE_>�BT���4p�a��\�����w�қ-O����43M�85�u}��&NDK@s	�@k@`�M�Q�L<E'1�OߴJ��X����I�Sc��g�)AK��LL-�8q�z�.� ������鉶Gk��R�qb�
Вl��c^J{_Pm*8�R��9��.�ؚAUq{�p-�մ�$�T�$�0��%�w���-}<��g���OBk���(���Cw@�`z
OϖA���w���)�Y�+��&���j]���n�{e�]�sk��0�h�HKԡ���l7��x�������,��QnZG���;��K/��@����硨���L)A�S�".-���� ��9��RU"��<{���M�O&��h�tfO��؍�3�Cv�� h��R��y�mg3�8��QL����8���m�AE��M��;��c+�Xh�O:��o!|u��ԟ�wg�s�z�C3t���\DFV�j���p�*��sD�}>�3��ʹȪ�m^Ț2�0t����T��e]�6L0��3�����f�L":�C����7�'��]�6��^br���B��z�`_�cۊs�E�յ��JK�X6\�Q���s�	�n�?��߂� �b
={{�?�M�By��?�;��GX�<�0=y���r���!�ǌ�=�����w´ �L�4E2��4�������IӨ�,FkDwl�������BUe-b�I������qw �+�{,���r�MG5#�S t��o�,jW�MxAР�����h���.��[�?�8�y����UM�����P��nV��P���$�tYC��K�*��~�ӷUBXl���L�"��0�gn� �M��V#��F�!J�̅ߢc���F����E� L�'��0�(Mc��"F7��=��di����+s�H��$l��+�S���?��
����D�V��\ȇ�FؚP݉�9�R�@w�WW�
���;�6�6�+7srO�yr�S�������*�gD��������������U�`^��܅��A=���Y���9�S1gD�Z�5�m>?5�)S���!y�X�Wj�uݣa����K�eT����;����Mw�C�/m$NajCtlj�d0�Ŗ��%�h��h �c!Y��2{nt��`g�]q���|�=[i��Zer,Q��J`�{d�.)��V��:��>���@%����Pֹ 5	��0�[htb�ި���G&as_�h�U���z����N�3E3�Ͳg�8�����S��
~D�3�i,����l<���s
����$F�d1�1�ز�����|��-��+�V�R�����D4�7v9�[<��p���e��Q�US�C�QS0�~����˸0�eG�
[z�N�n?f����(ş�3�@�Ҕ�k�nHz#d3g�&O�V�u���0l͏���P���0F��gb&�����!@�2��6B+G���R�&��RZ�(x7JJ�������7���~%G�'̾�Le\�e�������[�He&(��ngC|}��ے��oG�򥴄d��V��j���t�����>�o�^3�%��9^��3��3+Cr�ٛ��j��ۅ[�Tf��.�m���̥�k�?�<
��,�'�6��5�Nd�*m�+XW�Y��ߢ�`�C�����>�>��kl�?��R�4ƥ���aa�eE��Wj�_g����w@�^Ѕe�tl9�ۋ�9�����}�e�H�a�kz��?����W��8��a��ʚ2�[�sp.���n�e��k�:B6�0�;-S�8&�H:ު���Λ�P;೨���`J�g��x�'� Qm�Y�^��65B��i
@�{j�:d�+������v�f6��Mλ�ųQ�b��c��z��2P,euQ���&��������Z�$O�r������9�g��d��aS���=�M�q���
W^N��>J��o%�� R�"�$%뜧���g�?u�
����c�8G��N$h7�^��5>�B�P,"�q��y��~��H{,1���d�_Ln��y
�%&G��{�8���$.��"6�|Im*��lY���>�`�'�3�^�d�W�;j�j �b�K$��P(��>Ҝ�SM��/e
�=�����@/�e_ib�&'<���֣�� �|��ʘN��TySe��T���	3j����!��L��p��!�P��m8�4,�198BΪ="�oɊx�����kUj�_'����m��sP���/��gE'u7����6f�Ce�#�@߆0���X��4P�UWR�#dP0�ҋ}�9/xH~?�`/1�i%�=P��^�����-rd�a dl��1�C����y	+��b{�`(o����O��S���8����$71���dKh�m 2S"~S�6(��uuCq�q��.$�N�qh�˴M�ZD)��OlZ�;�a�K�5������lO��?��G�	J�x �׺�v�I,���x1�h�~���ڌ=Z��rC�)_!m3�]�^�_�푹�G�K�؍j͙m��"�
��`v�RƑ�S�ؑE�������:s�KD���|�b'}��Z���N���m��x��zF]�Q44=*3®�b:zOE`V(��6��~
�"�p��:��|\vj�*�t��Xh0Q� dy�=Iӑ��u�K�
s1o ��S�@�{W'>'c�F��p2�(�\����z�m�(��»[�Ց�9x�#&?W�r���#v *ֵ�o.�J���lbP�:a�Pt�Y��3��#�Dp�n���,[9W����\��*�vT��҉?H���3�|��Zz�Yx��i�[c��i�Urt=PZ��u.��|��"ėկ����c
�N�A��EzqJ��[���n�Y��'Ys�x�J���9����֥5�~��G�K�w7d���/���W�����L�uL�zK�KH��ҝ/]nR�;U����÷a�[�pE
�<k߄�@G
n���^��3�2aCg�b���a��5 �ÆMe�ݱ̷*�U���T�!��(΂���6�Ē,Lc��!�:Q�KN
�M�
�RU�M�,�[���-��P�j��(n���tf�����~2�P��4�3Ԣܲ�ʼell<-�b���+�O"��4�;
�(�����N�Ґi�9:��7>�F�tU+L�4��Τ��|0��LoO� G��Fg�Fr!g��W0ZǤ5�m�^�|���s�nHԥ8Ax�p���cEq�;��C�P�N�s���Ll���GF�[���YA�F����<�|S��}�7���X��4h%w�d��X�R�cq�̾&d�J%N�]�q�z�6xN�s�����8۶V�oj~�|����~Z냺LZ4\��-U�,��@7]7��v#�u{҆�qSB*/ܝ($�4Z F�B�C�"��e��ٗ�7����W��|��#(/��j������UH?bK����������>���J
�i���,�o<KA$��e����=S,Μ�=2B�֦�����z!+�n] 7�X���д��1�QML��9���ݗ?N��6��/S�#�o��UBO�җ��r���� ����P��b@bi��S�_�n;�.���P�p�b\+ޠ���c�i�|��)~8S��U�8�|�դ5�gt�ǋ�������>�P���9��A@-Q�k(BxW-UE�T���3�TD�+k�y|�� �[�f\����jy��Z���8lj~�_L���������NG~C�f� D�e-�Z�C�7���<c�pb����\���z��K���,H�_��ӕ];(��͚��Wn��P�@},��M�	�p�I�[Z}�D�n2����O�3����TڪT��0��_ݧSx*�Wk
�JE`o�S�8?�!_�+� ޽�C>s{+���ۖ<j��}�C����tt��V��A���)m�����63B���V��ސ�/<Rc�6\8�K��_|U�C��]Q0���/��kW�{��Y��*?.,��L7 ��+Õ$&��ۜM���H��36+�&*���kԃ~"E�6�)4KQN�� �W��0�LB��8H��
@�q|8D���Ar�j
�}�;���b�ƹ&�(�B�W�|_�X�:�ny��A��v�-�	W�%�iX2��� ��!�?����B^�13	
�.�L0���IH��q��-���FN���g1�:H푯��3V�t�wuy����]���m���n$����e?
�X�D۳ Ɯ���_��+$��8Ǭa��H\�L����iAo���>���Z�4$��DQ\����@&���e,��u��v�I�H�D0;��������x�Hٜ߶�H14q�����(?�[U
����x�w�(����+�M�m, �M�,�HfЧ(��刼���R w4ah5�J~��@����\���o�H Edʽ�bw���~9T���!��������b�=$6���r:mL�PǠ�~$�_���4n~�h�tw�����)AcU���E7�`{,}C��2zA�>Ԩo�
�����#ik2��4A(΄�w�X�X�C�Ď�顂���Uv����X+v^�HiQdo�ydY~���J:�Ď�z7�9�����C�����/_�Ŋ$X�m-��H`�#��@=F��e��D�=ɝq��nC��[<��~�̄ ���^�-`�<��� q�Tw������R�FdyA���������p,��U$D��2�݅Ie^�&=l�{M���S	ۃvl�	qL�_����K�� �������p�� ��۬W�D���{RL��a�&pqg�ڊ�I��h��[m�{��K�������0��]91�pU���P6)�Ƙ-��R�l)_���2�g�Jv��Z��.m~f�i
1V"�����,��w�����x)�=ڮ�?��C��M�z�	
��E,8��C������37 W8'm+���k~��F��5�As�Lz�@�ុe�|�+��s�s�3K��p|��
���l������p���:2Ԃ]�;�t$4��-�1� QB��(�\%�q��Xt��:�tZ�Qއ��'
�ΓO�W�G�~�����OF�P��~��aE55���ڌ G��:��E[�lL��3��n҈���U�4",hW��r{�>
���䛠��b0n,�h}9���5�P�����!�[Z��hO��-~��%[,"��L�	Z�ľz�n;:�a �GK��c�j1����v��U�%��y�l��q�
b"���<�{���K���[K����D|ϝ7\�U7���1Bs)ß�N�E~��dM�=a�yOUo�\2[�N�/�������E����Z\Qa�����ڊBK\M.J����R���fM���c����b��H�p5����9O����m���c�5��wv[�'��_⛆�F
�pU��&x�&u�#�����L�Ѷ��}�a��˱�5_��X���P���_��{`"�'ekȭV�&oG�J��m<P�5^l{�EqPn�U��>1;Nˑ���#z�[�F����+B�?�l]��s'�ߌ��� �T�ה�����}B��YS�c�M�E�B��x�X���I��X�VG=ŜO]�p����T������o]j˒8��.��0��l�+o�Ut�>��&��X�6�:���
�ѶH9:]�C�:��~H<Ϋ�͊�d��B>^�����ō�C%:�&�]�>�;װ��5��ș
�����c�S�X�ݒ�0�TEC�(o��s���;��n��!�cu�/hW�TI3 g��dE�������w��$%�O�`Ȉ�����"�mH���d5A�U���n�C�F2���D>�	�EV7E�_�'�ɿ��%C�8j�ϰ��Z��p��`y)-��8$\���܇���!wCBo�O�����^d'd*Q��LWد�#���c4Dz}�p7s���"=�4��#I�U��p�,6�N�D��c�'�<��9/�;`���}����]�œ؁�?�H|��L�O�/��k~�6Ԥ�5���%d���:�4P�o�_Tb���������D�<��&E�G[ߔ�$��'V�.*����K�m{%�]SP�/)��X�xīu�Aް��M&0�PBF��,[q#wW��U�M��,�htOE-'���3� ��(��_�l
_3^��2�o~5yޅ#|!S���[JYPsy�`�q�T������dVn��@���i�a�W�g*C��F����������q�nN��؏/�w�aq��H$�3VF�f�"{��:^�eA`�n���Q�ҥ��anJ2�k�VW3۵���蟙���+:8Y����K*�� U����5�hfAsB���d�ҩ#����#�*�ƛ�fػ�O:��8X�m�~�
˪M��)+�zYP��{�?fNԈdae�̑��[I��z�	�ߢ")��~C0[gf���S���2٦��G�h���h������#�E�;֊�\���
�?�e�9��At�{,���K�GkL�Q~�p��ԭ�7ff���f/����K�Ȁ��K��hS���B�(ly ��Ɣ"�JÝ��~S��|d�_V��7��n�].��3g(�<�A�ѹ�Xs���_��*<
�-�g��������w^��2r�B�F5Elf?�\��>��u9&�aU�-���}��˭�`�-���kg=f�V�;L����wK�]F�h����킪�����^��J�;��H�/0� R����!b��'�B6X��>����و킅 ��Al�z��^�y���������ɓ%۟��| K���������K�Q��3��$�>�%����,ě�����<4��}�t�3X�P1gō�S�:ē��{4�*�rg~�K��]��	ƅ��1u(�ô"���Wُd{��x��w����|�o0��`��娨�a�)�4F�S�qZM���,���r�������_�xIUÀ����E�=�~y�M��K�@�5w��S����(uAuzU�6ՆX�Zy����vF��r���軰��ܠa��ҙc@0�?���>�q�KJ���6b�����%�`t�(���� ��g���r����M���	��T��t��u�W��7d�x�É���Ҧr�Bq� fR�];Fk"!t�������a��f�v2c�#�Lb[G������7Hȇ+����b�~��F*R����:�B�4��>=�}�^jY���7`�Fy�ra1\+��{�G��h�u\�s��?�_��B��t�H��
��V�"�Y�&y���$��c�e�h������77r�i��	ƍ�oS�D�-����&ǲ��E�0��S�U��V)�)O���Ư���(5�.F�v2�	 ���[�0\27�Ϊ:PP$� �iJǑ�R�QB�	{v�]���_�BGk[k�9����9�ؑVv�h}�0����� Zer�X#�_��	f��2��E��c��"��Og��Ḡ�k���5%�s������(ګ��.V�d}���<*��X�`��C5Se7k���on��f����龋�gQc�h|��~�{?A�9���X����h����g���#S�ͮ2�3���.��5�*f�d+�B��Yn�q-��p�����I�WS�~��K �׷~$N̂�`9$��{6��c����nr��.V���
�\(	���n ��[���jc��T�j�
E�#�z��$�`��\vFgO�Y��P}�#�r�D������E7��:��ӳ �#�J�C��]�ߵ~��U�~�-�����T�I伾z't3�S�3XA�K�6�`KB���z`��85a�4}	+��L�bRi\oK�\RX�u���5�U+6�W���E�j�8�fAD�y�@���G�,��[ �U0��7�� 2�*���#�bQ`7NzY��qU���3>���=��`وa�چո
B�n1k�Z��À�LL�2B�5�����i���q��@DW�,��PE�>�?��Vu]q"d9�>�ٔ�*��ɇe$��&�L��9i��i��q�@}w 8���М?��ɞ�>��)S��A��8�b�"	�S)2�f�d�&mǼ��5��	@�j�/{�$�_U?��h7\�2��\����s�)XK%�a��1�D1�#�D��q'��
j*�\�`?ȟ�b�OĿ�����l���X`m��X\��F<#F wD�N�]},Qc�AU�6m�v��f+�'�9���W��	B3�L7�E���m���xS�'���hl}�{.���v`+��N��?�m�Y���?V2FH/1Q��6�
9��?�}[U"46>	a*�D��&LƓ�B�b��Fq�nRp޾�H^maM.tbE؄\^�VE���z�P�@�C�T>���g���l�^NXw��b�57�I�`9-V֐F�X�A�I�F�J����f�i��xM[�~�_\J���d����H3	�N��<�Ƹ�@DB���N�e��SB��������r}r�yFVy�\J��i2qPl��ߔ��M���&uK�G+A�5:�֒�x0�� p�����G���}�~��'�G��nq��z�"�Y�\�Fn����+���>�_�1�1���zD�_��!��n��c����:���x�������Ԩ�݊��,q�|�^��	�^�C��o��P�׍SԌ� �^0���bA�kKJUE*2�y�5�d��\Q�f���E;t��AШ���:��"�T������#w[�BN�d}�y�g�z~�2���x�B=c\����o�(Z#a������5�n�����ķ��S���BR�˕DM*|"q1~ǚ������@X����S��!Y��9i�R�+D\�:V ~�ʒ`2�.#���7	*8hq��z�S�(���N���v��NV?�^�9��������r	1�V�+�-�Ry�g$eLhe��Y@D0U3P����TQ�S�P9Ǯ�e��,����Ȱ�����N�j�6>��N����ɍ��Ն"�>r?S�L�-�i
"���\� jW�}9K}7q显C�U�E�R�P���ўY��o�&��C]��抜R�W�s�0��u-O������j���N\�5 �����Ǿ:�&���C��,��%aj�E�vZ�RI��EZ�6;B{�,S�fQ�h�3� ���;����s��[	m
հJ�Ѭ���
v �+Kw�s�O7`H8ֱ�a/�#R�= ��M��.�I��B���J�Y���0yS���g����4m���._���0�J���屳�*��aH�k�v#,-��i�T�Ś�?;^�Њ�o�۰_�+D��B�"�f%t�>���}pY��*�g[�-�0��#j3����u9c�\=�l8N�@�]�˃�[oZ�+�2do}5k̪��/@�����y����c|�]kK����P ��{%Zi�_=X|��L�:�h�jh��?6jpi,� !�n�]�I��#Z�����柤��,��P��+��Z����PS�ͻ�֬5{Sm����P�����b�p���Чa�`V�tՍŜ/0ns����Q]�c\c���`�����g,~tg��j�礥��qZ��\�1SoT��g y*l��A�"��6H��78�8`G�I�A�"�l)%��L�Ftvr��_Ը�M~�}�(���u<����`���]���9�����9�~�k8\mΉ�����Շ���Я��'��}���@E���6��cx��I3J_��rq;M��T�+�Q�n�Ԭz�П�Y�P��:żC�T-Mg����h���a㉃5�fS�̜�o~�6��5w������YܿN��g�m��,(�߮r��&CB����`���d���Q,#¡��k����m��'�t0d�Gw��u~�Zy��<��?�rp����-�Yj�!�� ��e&0r�`ѻׇ��w�%�h��+��?_�%�L[��@��=Y�c���Dq��)����c���؞`^Oj����d�`|�$6[w��G���r�
�����T�/@���n�$*R�ROȚ��`�������݃��&:X�iˡ�Bq	C�dF��� ��U���eפ��s�d��Z�y(\:� <��7ΌW�ԫ5����>�x����9�@9��=5�D������� w6���T�?�W,7��1�g#����������Z��3�Ja��DQ��b�؁���44�^9��O��]���X=۟��`T^e�4�}�`�����������܆��fƜ2
����W/�;�OR��B��.�P�����m�nY�A�jX �N"͍`xs�V�fP�I�3���E�C���(�D�p�������꥘V#�����\��ׅO<g���z5?&B��*ѣo�D�v3E7��<��=��?�к [���F���C>��*9��ƶ=��V���$5(C�Ï��`}]#z�*�n�)�	_�H�p���#-���'��r��Z�٤*zh8-�-�l�Y�x���1�i7Xŗ����0!�xFCF��Ym���ƹ�L�]�+f���2!c��?����P��h
���l�����w�Z~�7��:)`��2�������\��U�؜[={ʲ��>��sT+K�� ��ߜ� �@�J).aW��zX��_f8�o:+�ѥ�qXlwG^yӺ�v#�Q���Hx�￨{���p@���S�3ƽ�r�P6�@9�a8�~	���ܷr�x�Z�j&CD���z�n~D�Da���b�$��z瞇�����B��U(t��P�F�[p'oކ��K�ؾ/���Bc���򒨻�]*y��'K�֊PFIy��oz rP�*C6�<�t�L;���Ox)�V�uV}/u��>�I��9T~�[��Cg�R�6����so��-��\��]��b豐M�g� �`�{�@N��%؃cL2\/4�6\����?�i@?��cY�HE �<=@}���9�
D�j|����3�B[q�Ň�4����i���u��@�͗�Ӥ�`��qP�/5ۍ{�p�CD��i�RE
$/���(.��A����q�N���_�t�Xh��QN��M�b�Y�+ ����Ee�FᏧM�V�R�J;��n�H�}E�3G6cHRWz�6�D!�^O���\^y>�p�������ژ�`��2@6:��׍H"�㐨(���q"��Rb"�is�V��+�����%0�����\rZ��>����R��c]l$���*h���ȯ�|7�=D�0:_������HE�F|ȋ�r�E��0!L.E?Y������
�f�6�I���S��l�AU�zUSCh���(<�
�\�O ๩�)�H(u�g��:�XVM�R�2ҽ��c$�ޭvH�*�NG��ضr�P}nP��*}�;#��y%@$��b�1g�'�o1���|�<��|��l'yz��T~8l�]�X�⍊ns	��{�)_'��#�rv�-Ҍ�V�>�����vpf1�af�ԊFoB��s�KDWض�-l�#����VE��jh�>�w���drG���Z���:>�Lȯ$�3|�,5v7��wA�$�����Qi�1�g�Ӗ�g��N��Z���R%C3@�}4x�L�]#qB��n\���2���p����]�'�%PA�}B�͡�6?P-��D_P�r�	8�fȞ�۾%:Er�T>���??��21`���h|\�;�6���Ţ�OjF`��=q�_�Ч��H#��&$E���K�ds��#��<�4���%c�n���*�k3� �����B*ϭ�d]�.�1u��x&��2fSЩ�e~?ZiĐaM�����Y�.|��[8%b�04�{O|�W��Q�{G��i�uj����9�U.�����hi��<|/R���f1	�����2Cp/Զ�"r�K�ZNp�W��?a�=�
��[�]4�tN����GY*�#W����,o��L�T�oR2U�w�[�?Z�"|jV)������)�ke�{�����!s��ٹ(�����fx�V)2Ne곮�d�v �81�.��� ��nGé��lZk�9���;�����\����h��=�9�ʳ
Z����C#`e%@�W�ɛ��YI7l����%`���"w>�L�3h�ՋQ�.8�̹;s��K�b��%��cQ!WY���6[hBb��! �فqRJ�q]?�|t��n������d�7ގ����.�a��G$����0��T���`�/X	�Q�Ts^&��y����������%i.����f�yJ�˭���Ib�z��H5c�;�D�����ˎ �qsś�wa�Os�y]wt�O��H�h�x�߰�O�����+l����:�%�@��X����@�Zu��y�'���\�eTJ�64r����Xf���wu(�t)+7b�4�p
4���Y�5@4Bh��6�ȷ�S�I������M禖]@�fsr{�)�b�#&1�p�;���~pYY�&٤�Z��Y�~���+?��(+^7W���������_�`����$F[3Ry�DW=o���P��dTt=J"{�'��х��oz'Ot֧P��Ϣp����{��᙮b�>剀-��u�u\��+~ȍo�Ғ�.�k]����7��#/��0��y���B�o�{>FD9$/�ެ�p��3o%��*v�q�,cҙ1�� �Ɋw<���Zj��m�q�v�����&�3�XY"e"�;��3�ٻ���iM��>���e�x���Bf� 1��3�C�,��rԼ���:Fɽyh8ק���Q�pE"3Qr����@��?���{M�3�3�J�v��P��婧W�yu�Qy[k�+#!B����"Z|K/��w���nͭh��$�<pԾ�AN��5/��\��k���g�U��..��ܧA�i(�ו-���t"ʌ
��\�έO�6�Ys�J������
�yw�w�%y�����駶�Lsmy����x����nS>�]up��>�W��+��0�D�%A��M*E���iޞr ��� �p����H6/�40'��s7���7i��ŀL\�����ѹ��_\����>��-��� �,EL�
ES�4�D��j�4�;i�xe�b�u���U����[2K�9�����?�������4��4c�q_�LF�r�'pa�Ll�\kL-̣�b���%g��l�=�K0|�S�O�="���Zߣ)�%��c��خ���`9���W���~��Ӊ�#�������X����4u1S�-�`Nd[t!���6F������oڤrO�6+���E�v��7�1�Q�=O�Jm����c`�ᣱ. w��>�9΍��U�*rН��4�ֱ�����Ju5Չ�7���l�b�@��\�(9#�����ѷ��3�[ڍm�jۯ�o���*UO�m+]}���q��x]E��7�̱yjN_"&!x���Y����z���OX�/ʊ(m�D�y�"�?x����z&�D���@fg^��Ov5>��
��k�Un�����:�I&pW���!��l�l\�L��q�r4i�0���_FV�(��!�Q'N�2)t��d�z�1�	w䚙Mm��
��`�D��D�/O�k�x��)6�N0�M7�	�&���Sy�fn^���[�ӯ�a}�E(�v!��iZrq�^�Gn��u����T*�>�����y�xs�b�,P��rZrz��tBn��+?H�W���z2��vU�C8��F��>}�[�t�r�Sh)�l���������Y6����DY}L�V=׀��D��bɑ���B�/�}���r�7P�`�g�?!(O�e�2}�>�P��Pe��.3,/��5���"�t����|MWͶmୗ��uIĤ޻Q��2��}~�Ù��rE;�*p��=�`(�k:9��vL�r�4WE��Ix+0u�4�E$>���m9l������w7rs�lfu�l8�)֊w	 ���I����P���k�$�?�iY"c��{\�&N�Ӱ������k����0�u����Z��n�0��6 ^:�}"�, Q�F�`�z<7��3�F}+V7����@��6��=BoU)��˫i�-��WQ�[)0�6�1Y;M�*<��B��3!���!���4M��2Gpؖ|�����_�&.ԉ���ln�=�_M�F�	6�<��}�J�I-ZI�#U^ ڭ&N	^�<���6�\ ��Ȅ7s5�A\����}y�T�D�i�}���w�rX��W/8���ᛞ^QBJV���C~���d�]NȬ��t3��|Â�%�����NL��lv���l�m7��U�n��'T	zE�l���gm	B�3�܂h2vj�Y�,�B�����N�ى�F=����0��A�}K�p���Ĥ�����el<���'mJ���$������k����b��ay�la¸�r�0HU����/�=���\{<��;";ј��Ѭa?~,M�U�7)�����0��ŭ�tV��+�c�c,25���yz{/���${�Y\bɌ��`�;������쏍��>��*�tޥ4��h		����� �v%PE�)�&��*<��F���=)���@���,WQ��fV�	��I�&lzqrR6_�4n#�#j���Ev��?��՞�ќa�2�:�ϸW�Ml�17/k!|�֓��\2+�����#�x4������O�2	�V@�?q^�Q�9��ߕ:�r�]��aV�����+h��]����q�'r�禖>ŇY�~��l�ⲝ�9^��Ϋ�~4���e���YS��)��x�{�)^��������uNy7�a]g�k�M�my��G������,�*q3	��=��ҏ�L�^R��傋�B��=-���d�!k��]����L�>dYT�iu�����
������r���i����̲ܷP	��z*#��Ïߐ�l����ʷ�Ż
�n6��f���g/ zDA�i�X9��}T3��)��!iU� '��]���Yi8�.U�/\:�ݸj���n�c�/[6?(�|��s-��\���75�TV�H^^A�B��ÔvxO%�����E���l��\�q7�d�ODSՄY�]^8���e�[��u����P"dZ�,^r\��j�
�Y�=p�K���Ax���j���qH��s�r}xJ3!3:��Na#��M)c����p���Zf��I��2�2uqo����$2d��=��b���B�3�z�	lFw1	�ָF�À�&���U����Hb��A��BCTr������u9I5�ߑ)w9�2�zǻL�*��y� �#s���b�{m�㇊v&p>��G�����e����YW��q[p��:|�5\隳q�ªy͈�X=NΈM�Ư��wr�)1�C��s/`p�:['B2�v*�0�hDe]9���1�>�Ї�mu�]�r�� leC��ƿ��M!�ki��Ue|4�A��n��=�éz�O"�ܥ���A�r>^vq.1��#�jw��>�v�r�6
w+����(0'zw��c��B�(�k)%RԔ�~7u�Æ���"�14F����?/��e��>K�xC����l��1o2�j�.�D��iT%�U��F��͌�㿑K�u>�����G~���Ȣ�i�5\��џmI$_=��]WP\�/ǐJ��'�G�P`�ڼ��B��������U�&�]+:��
|�$zG��5��h�CE����I@��6��D��	@&�����͘f}5XC?%6�\.p�ٹ�#7fW�`tQG�l�k��|�ga�� WӋ&*�BX�(��AK0�2C�TXT	�[�n��-��V%e%��)�/P1��?+":�"�	>�[*!��mY�f�r�Ǡ7e-��S�bGO0oy�~!�rpA�􁐐T5�6Z��P6iY��[w������N���r��#���7� ?�l��c��[�Nzx�ռ�92h���g���\�����1nH�ôS}�'���}Q���eL,^_,v 	�#P�-��	9��M�q�y��o�pL��멓;��%kTp�4��!r��l�vf����