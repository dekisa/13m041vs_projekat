// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
gf4ZzBmHcxk5hAbT9goOJyDYZmJFYOFeiDm3iqKztRAQs8zZXJmb7ag6Qxxz8I7MX351OooZC3FF
Q4ogd+wHY3/jRJuB+lpKfEeGgF3xEA1dYMvBAUcK3o1NPsrW6vKSLo9nrJ+XY7ui3sn63vWW31le
9vQqCz1L+b7DnWLxvusXlNlXBx01L/jtfs2F9+bN8s7YnYb/rBsBC5UKEoaKzcIiIgL/cjqkBu19
wrXwz5nrZw8fRO+rZMUw3W955uGw5tFux7tX0x2Q/x8aKWyRu5TENBJwlRPFDIEUKLOE5ENfX2wp
02OxomUB9hByi3xd5LmzmR5Yum3ZixJQhEIEEA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11856)
dlwG7QtrL2/7G6wH0PbGv59beqNbGKQnIRTakTuskVkGTe3EcWs+RTXkXbfYwqsh7rBwKabyTX6n
P8Wh7SamAxchoSyDCm8/hDFt7FnpeG953BblIVqR9C6/liBp37me/mzorPzrjs5efzJVVQQ/GMse
Y50JuDipPdIpdQjo+YOW3UvhrSt7v1hZJ9Wms6FABlvZ9nGNsVFf4ApgSLK3t64yxjjJ0qxIG3/O
1MsYCnodU55oYAFfk/ajQwDF6j10dOc4DFzoetAeICgAaIxIkbd+bNYR2lowWx03uGWlERxq6Xaq
QlroRp02ROvEAHKRk3S37YLjFpWvYQRDNC8N8mQ/JFjFTn1r4Nr/PKtRu5ZRKBsb9dy/oTY/QFB3
p8jrA7Hhik7+IAL1BrJKwEKADnxduvH9ipvvUvV2TG5ZnyH9uXXKp5+4TfXbspL7uRe76M6I9tv1
JkKnTXaO4uQZS/Dagwkf1U+O+wQFYgL5N8eaNw9Ri6kt+XU7L8gSohWHFDaXeRzASJHSXUCrGeU5
I2ayRVC+CBX7MU8NwTsKsdZ2yduyA0HupDg7SBeEj5y6jhzqJYz5TiAMtSsDI7sEKjC47MHaQz2o
dO27Z1wcxLlrZWkqPWW+u99oeTcaQEbgBKBunLDDeSPEwAlnLetOe+P9+plHYACryBAI+dSwnLgw
PzKZHaKHxQyDOYkkJsuhJYVZtNiT6vlerLRSRbkgYJxhzaOHjJUjIcxZ2rHC82gti48Z1Kkixp0F
ZxxswtBBO+duKCZUtqkW4OfNUMyW3rNkAziHpIEi51QOeLEcmjZgp9Thg6+ho95luKxzCvNbvHAG
7hlcgDm1XhJWExVmPxexWcN4EG0KOSUzFKN/MqRzMUXhq8gzNoyX5nHeRp6eW7zRVzK+s73Prlc6
aYGrHrUiJowSaxKUg2qr9qNgNtWquSCNGJGSgOIxKwSS6HvHql4A9ZIiHvCeh+CphDG6LJN0KdjJ
Nrb5Baw3gNA7QrxQk12+pZbcAiUTBRKmS19SIfLY2NwpAlXBiopJxPXpoko3U+ISOO1umXOhfB2g
akuQMmW004E28kPYGUQLRrKp1rpIuXcjqVIyWisR9TRFNV/B6bnNr9EDY9gjbl+wdtjpyEgC+RTH
cvhnjWXz05qZ4dFTZxd7MoUoMMXyrbLcCtnZR1Lb7pWlPCbsK2MgWrGM/WQ9vVhMuLojJiiPA3Xd
g9MhJ8Inc1lRHyHXA622xSbcGZkYwlvbZy3oPTHU3ZA0639cdsVofe2RyYlZhAJJeoMvXKT3ptP3
8DZhTimRVS1OAIaLzSWWHkH9Zn8SLUQxTE+PUleSHSRnVrkb8upigdkCSELB9y/GtsPloMeyokk1
Vk9qfInZVngSNDInSL/S0g11Mtqev+KLieN+C0UPffzWpPAfsum3zzKwZUgMBEOc5Uw9RgM4Np7R
eMcd/Lyws35IwM/QZ/37KsklJqR7f2yvV7FgkJ9XS6xzclG+xyjhAvOcKRd2KDMFRoyfZk2wWlSH
a78ZvG42+lCcy9IsRm4rlW4C5u4nwd/ROV1T26sZURUr2Qhenk0HIjfFZdXJBex8RkJEMMpjTWu5
uiNvE4VwlkgHFg2ZuX9nxvM9D203Xv7HggHLIaHesxjLsA1wLaGLMilXRho1DSy33RfWJtKzwbPX
D650+3hmbUpNy2/VXi7iZ/O59P8x9cYoJKOTOoNSviQwGWz0oUNlBumb92OCLt7IXCcIdWdkR8WP
FNMmkBOM6MyCA5XvX5d/onOFUhKnAhjD3yIeWFDeRld0Q0sSTNvzbIv/zfxqEBb7GyU+Ip8IOgQt
jkcZTdj9GgL2bnP7+5pfieRN1TJlBIPhqstUtkcsh2IReeThGJRNIMK09bdbAKi/u72E1rgSJibx
Q3+Za0Y+gCwQ9EmZF0WKdgd4I6LICGEP5etL+e2mO1NYkIAkmm3xlE9GHCxfAS8sWJCqHMG7cJQh
W84ItuUvsa5Te98McwlW+EtY+FSXGR7Ntl5a4peOPBlqGJLA0EW9OKLHRXovKHPj+2P45UQ1VFRb
b9G44aI+yTEQMffbde3nCOKoMrkPjFy/LyOyWuI6Vv+gEvF1Ai3rANRGTFpl6tsvWwpXWIKT4J/+
piVd14vm/3p+3NfwoO7rT2ul7NX0aHJcc82p7YBUulrzcnC/yxcxx0edhdBI96fIX3Eh2omtULTa
MnSP9PY0NipYDlqB1D17jIyjvn/erpMcHr3O1Ftz2ivfVvO2T9N7qOaP9ZdYyKeNPUGa8sDm/D84
QGC18calnT4zOZViQs0W6r+psVn6JaT6tw/E6bnXmT+jfWuPLARwnfbblhVANVQNbVisxjzJguA1
nfnylhbPrQ+V8aiAiNUMrp0VgP09mmWxfRkTa/2g396S9/jM8pJEKa9S/6iMDHtvYb+p5gZaMYdW
z45+KETOBXRwsO+Dzo7XAG1RLAI6OYM2HhuUVv+6hT9fEn6d9/80Azyhq6yv2h4SDRpJQVWrqa1Z
+19ps6zkSmT7vwv2sHHnZpNyNqM7EW8dguJtgxW5knnwBUFsnBl7I7NxUKlVjHg1BQi/S0q2bSs9
utN6QWVsAFcu/hBYDXPpc/2RH366JMAH3puMEGtMJM11+BYM8S2xm3Bd/T02Q1dPJHrylqZDQ7OT
mU6eIv7DLDnIFzxcqozfg2Z9r3w7FiNr4IkImcUHfrAdFvz542HqKrBOHlA079mYS1vWBO7OAf/B
Ck0Zyws6g5NQ2T61wLa12rwaeW0zuoM1Sbc6w5vl3/tJaLxIrLXBsk7/JMEyC2mzXjgIcDCg1uMF
lGWUbz25vcldEIa24rqiFXkK1nLFlU3ET/LgXOn001TaF0gOqTU2EfeElGbmXWoR3GPb/EcFLsha
wfwfYAYpeDLKrsyVR14lbr6zdmw+9bf3tanEtT0W7uwJ+VhUdBEvUJgRaUNvco9wbcOYAH1Fmrfs
hHZnXliPpZGHSOfS+ubWNXK7EGyDMfPa8PakXGcwgPis2K9agutzJHRO5nTTeXedvO70Lzi5QWmo
xVO0Yi+hW14XjWT2U6G2gGSvHvsl6Y8YeassdMqCHZN4/zvJTPQcmfkM5L5iHzLn9/tN2QDgkRzc
zbaj3N66g95Y/DYkfs4F2rqDo1RdZwDMLxObcmgkpwfxDmjeASllqSpR6BMFBQf21oSjETzIuux6
T8SZZwUfbi2X4bXHcQPqDthcAKLsbG6MHduJMduYywxKxpBm11SB7syZimNJxQv57+fMSxoJqla2
BTDEXsM5b8ctFkxYHS0d6BzMGkET7Gxz3t9M76bcT8Nv4/R2GIWhYFSYXLH0mca66yWt+kXsiMwH
EiOcqNnZpcmfLGFn8kCWJRZ0Lfw89w56zz8cs8HL5rMn6NRWglKOeQiaZg8EUytKfUXwVaA7Toe1
5N/LoXs/6t9YquAi0daLZ6YU7AHT9tbGAEDTJkOoS9tf8v3ltbh9AJHvJqJTHeMOE0GXthsjFsKN
In1bMDVTGLncTl7l/tTGlpbnfF5e2qhNSyPYmozKA4Db824fkh6tNgIRu3if/+glPegnH78gdLNY
SKojsHLHDX4JWYkB/pYyrHiF3u64rb19f6E9zKX97BgYjPbQZi90lRvUqLgLR6WeTwgvNLRzcJhP
Pjlj3a0IZj6hzSdikPBemOvvmzPX95CvoymdsxXRT8uReoPiKPWof7S4trZVPsPbrabJuii+jNhv
/ud6QSJ1xERA1j9qub6EjZWtQlBERF+xpMVvr+MT6UeIWSWqd39dgSovs7YWQe5PyDEEM7SlSzxI
L0ca38MN7rcIXMFUrdV+3ySGL6aowv4MgWLDGVIxN0DcUvmpa26qmF/kBiy6oMIzeHkpdcwXdTgV
1LOo4dOjUmgxn+8UFVrkTOd6KRfCinegbD3qcRm0eRjAafA9ADe7NF1kDY0DfsiXnnyBQhjdCQtR
op5QAPqzYd+87SBXiCD6F71JJJr7YuKiD8dRqdlpQERqTrraw6QNgjD2H4sTpgShDuviy2tv5rHm
1fUMsfVaYpJXd2LYN4n5MWLV4EoVBnqq1Ko9FmtyFv2jd+fxyh2moWfFlqGqonmXocTAcfaRhT0k
0o7++PlAVyvrM5bLOOqSphndrXZ1oES9wguDlQM7btKhzRoZ/jXu/L/F8YKsJIAw7TKvLB1y0tuC
CRG4TTnr0Hs2kpGz9vVKasJ+oMIQwzg8KmYbwEEgcaxCZ0lQobtciYppMsmDz/q6mRY8PS9A7JkY
QPZG7+HEGHJYUMC4q/Vg62kFymIrINIacqp/9Q3XkrbKRTf5sOx5StXK5n/zW7dtWfwS6ds+7i0r
iVDlIi1CMiYHhacmNvtqnc874/2nw775pRyToAmaDnRfkFooSW4/y4HxAdqBJnEWYWfkn9lvZyQV
YRtzkCKjO9zSttF827OkI9PwQMTRZb7+wY7zPajhI8+vsgfHRo6vFbcB5UKXLuLn6plWzuu23S76
ySZD3HFOoEW1qt8R8b0aKCgVp76D08/FocVw58+pedCjbyl8qrh2BE9RM0KHOii8Ft90HT3j7/tg
EJeOrHdq1YwI/BQlx/JwTPLFaMjrLUtvmHWB1XVQD7LKJF2Q1r7SLFW315sf119Ts88VwqyE2HJC
l3ukAAa7gowMloQtFEFsQjk/sH2vrFno35XBAP/0d1+wxjTrWpxIXKK4uCnaPWHlkLq/vN6pKgRL
sZ0E4SrG6lms0N0C91ZArcD68kPrHcVkaQ+w6reUqnRY4zClG7F6v5Q/9vXhYKlFVrb3emjaoQl1
aRSLPZnemnAih9Wqvo9Cob9b81D91cA+VKCznLR9OgSPEPy0Ip2gv9D0gL/kRbjIeY5U+jSdqWq5
5SrMWfirO5QPuRPwOX3fG12G2SrvKAYAKqhLWI+pE6vMEMBK0ki7FK4Hf8R8KqeIy1DrBIfxAPk8
DZmfK54VEx7W/lgka7Q0SKV9O+7QFqlMDG0n/qAlqBPneLW+Eg21kJDYiQWbIYUbxulDqSqPScNs
F8/9upos4PRr15iLDQBzk1dD9P6PN76vym1legeuoVB7z7mP0dwAXhoodoHj6sskARElxXVsj1VC
gcN3XlinkGOe2KnohU6bg2CvjkC1ZMgZKRPWlI2Xl7mbfGYWxXIVBbV17PsTw0ZFehxw1zdy7Q+0
4lwt5mtNLlaQjvpynsIlOTrNNe5/+U3VMM8QU8WHqL2k+IjZNC3d/7D/kSv0S79YF5mM94qqpbH0
JiCaZnIVMnmRYdQVPUSN4HTCf5lt8En5TYJ7znmZEwFa3HJ9H4I6GUklpDOM0wguOym8KuaDJdQX
r/7xAdO0EufFLxzHdf6I4+TKCMKykS5Q03kCvQIvCk4MkzM0K6btTUC0SlZC8UHurwZsECLLyEbQ
kuc6x7B0Aq5nFSTDUSWb6jLUX/gStYGv3uHnP1PUEuy0Dax2y+4uYZmdneXg0MZMLZqLLSkJCP5R
ZWl9SS4HB2M/KZ8Ep4RCSPZRs6hV75uOuFXRabZabhRCPOXqVC6veXNjLuIr2bicVQES6MIC+5YI
ztiUqk6Xj7hl4dACvI+SQ8+wQv9K2PkWHtPfOQhgo78aMbGzkquC07stg4E3NOiW5crcIy87w4/s
bt1COqYVOCwkmAMu4N4F+WP57Zb/r0yEHrd1H+mxj547IpX9CM7OcjcE5pvga6fpz1RD7fAjOdfb
WlAV0kF4qPWSRrGF2HgUt85vprFIpihdAbGreks0sOIP44vCtWRMTc9M8OfMHIzFmEhyAx0mHHdW
ag3K+bjo2+9GkumCF+o9dHrh8J4Mf+aaVvu93QLJLUT4rwUGUtGt3zTMgVHv6ceeTRVonZZX0jE8
cRtqSZY//8O2nZPUL8p6CHrsuTXow9s2e/2I5DBRr6UqltJ7eSr9jGQae5rgefP/EN346nlyEc39
6ZEjYjok6HGqcS3YNVPypOZa8YYIETAowvqfNCdF4+fPvconO+nBdhLS2wjz1Isq9dfN2oY2In9N
2qbNldXUraEFP7T4h5g9ukn0+rrCUPqhXXRFUzGdTXecdEN0L11tq97BlYDAytHTgyenWEONUc8K
8egUECr4/QoydSmOi+X7jP9gEDZ6uPsoMr2eS0CG1Qcx9bY6nQjd09JfWNB1xq5hSbnZj8F1cVp3
E7ebsdD1uRyRmFNgM3OWCskSKS+GrrQ51q11zJNGRqsWGaeGVAeA1L34B6WFEzvgZUKLOcfQcsx4
lTT1Rep/RcDNlBD+zi9uPCG3paNqR2Tlg2FqZY3BKFB+cP5a99NoGthcf7E6Yc/beYBZ/4H3pSjv
NuDfr0LL8tTAJfJ3jQ63XSj2wU/ysUr58mfmzHAN2dMpzczUIOxpZZjQFuKLSzMVBIav2vggdYla
WhqS77iLI25MTqncUQmdoTA2T6iZUzzZJJuWOkpsvhkeJFGZ10U87bwKk6tdShU1JKEoZAuGuCiy
D4cLtTY30EqacTE3vG2RUP+2pPNQTyUs7jlmp5uG3p4KZb+9wyuR8OA3vbhc+dh68HjoHEu25BwN
L7EU8IZePoJyzKjNKNheZ5ekGCo6yLua1SRQqOdPHFFNhbueM8mD2SSj55HfJ9LyzFQV0TH8JjmB
vm4SR+y2GWM+3Q3tDiPBYTBPCDQhQSM5stxhF7HhuJpyjaZhmChMtUMJZCT1rmSopHOZMDHa8g8n
8RTknpyR+RgjwgvTt1eRW8HCON9406WEu0BrojFCxDOT6FgzrFkhEKALPpRiaAca3lLIzI7C5tzR
tN0bvo58NSjtS1CpFh2/vytYsZ7swYoeR7mH3fLI2v4Q5Wpr/G7a32aYOuy5OQdDee+WnEZyFxPR
VwLT357VS8ItEumJ1N22LkJfUqyVs+pfs47hf/WglD7TYeMONZpYWclfN3WohLiZ5T9eXWzAhrGR
cMLZPXR5kFHRFd7JSMsVrRPExy7W3D7LYkajZHGDHBCKtZaiPweMlNU9AmmUf4+dkp5REe1Nru0J
Pg+t4DOhEVmL4m5ayXQxjlckPbaepodUzy1pDhuHVSKMQVuaGppIpUrUAdx6XKMa7iCQicpTA+XK
Igakfv3aMqk722aKQjNN8QeuQ3eQbehSe+oX61/ngB76XyoqcK81/w4ea3jEzZ+0Q8E/dWUhPqZ1
+bocPV+KrZgGzUYekeQUnm0xJh5n7Co5Zf7XccKtuQHCU6LDPMuW27tFlXOgKtdOeP4lbtg3Uzr4
dkF3O9usyW2nxa0mZlMASR7Rb0oCtg8vTnvUxgLjUYNgH1kF2Hx2jI54SN43FsSaksexn4xhjS+X
4iV4ubc0LpeeKnXY6gp+hgIyXTmtJrrrCj13IjAW0DM7OGG91hkXfdDXTjG05z5Qbu7dfPuw6FiI
ZuQZ7NqFiUmHhPkN3iFhrh7dW7twOUGhqF9wbfK1MLiJNaJBTtmI2HUGi4vOJs/Jl9woNe1zk3He
IcXNNHy+cmvT8bzab4M+O9Tu1gUCTXr4SsDWVg3zm4UktiqYT+TXid3tLc3NTsu6he7eaLcTFD+n
47CmDl+cu1RPxc+td29cRmyxwUJUIfqswutrT2YSbWdzT/Z4j7SDJZUHOELUZQWKO+CwktslhKLR
5yUR2+1AgexZRANBlDWVTGmQlMc8Y9iU/Uug0l6UzsuNIIu6CzjGR14eK80MbhhFomNGCF/1WlUL
Bbiv4kPiDdAsLqvv3EPiRaxaxxxYa/ZE71424AARORjXm/dgfn/fy0Gz6fKLZ43gmNcpFxYwSPV0
O9U1FncFiUUrCVg7JQREXODGbFQ2SJmog8rx6CrxK1jO3zYU6KXrrIUD5uNtZuj6X0ZvU+MW3RX5
XDrQ2uESmwaTx6aCuiDn9LxBITrIVSENjvN+MO/HCkMMRyGe6HZrYhMBebFyKa/kf7xEC1RXy/5i
GzJAbEV2Lpftw9VTs695jHhwNcXvuOY1IRCUYrJBF5J9j8SxhoOIp9YtphyX4DgPjgVtN7er23vt
pO8uOnzzg21UUIznUf6aCKZ4atPQ+uv2tgdYTROtzyQKrdVxmyPKlbt2aup+FL34JXeERaFKbPZt
QHlS+P8xlMcGi9FjrlytLf23VBwcSNfpgvchsDt9HXBSEskvEhq9KQMLATqFRtP8311yyuNn6ZCz
qmf2LvOxcbxSG4QPNWYPvZZfvUPXryYdXn3bEBEzVInZ9qtzxkeumnId1s12fHAlLSYAXWfSEERu
EMA+LqgeyKjd84hzA+QfBHdnHhhSYqT5AMGSeWa1No3AoA6u7sdPPq/1dhM/xBTmUx5/dnVdiEMZ
+cLW/kb3m/ZDZeYt0sqSWHoDfQ182P0Xs1V29brYg/mqPR0O+XoZHGqBOu1UdrczHpwziB5YGlt7
DexEINTB2OU/C2RygIYQw75xjZdA3GcoF788SPEkAwYjk7HK1TGoCBbxiDRaaBel9R8z6PVDp9Ra
BKiCKG+gnN8D12iU0R5O3/cvDCAU4gJ2IW4MhsTSTY/Fu9MOQHT0GoCW7sQNfqcg7ewld6OIxPZN
5JNnYdutjYdSAqihxC2atvZ6XKM2P8OD5d6ElJM2oeXLo3GK+ATuDpIgjmVAcjnBsWura6f/M7DI
1jxp5GzqgSIl6d1cdevb5e/9nd8hejM27KK0AbdDnFGeV2a3GblhQt6m2ofekFLfIZZ2cQRn0s2/
Kli5Ir/FXfOxploNjK+8TIAFVTB3S7rf5PzvXqq3+8vpiLvVzLKP/6o/01RldXxaxI6okqjZo0MB
odlfq3Qf7dj4BKvD+5oVgcVW5UGIDB/EBwJF15QfqAsvcnwssLZsXLILI+TyZEvjR1/zyBBelP7l
OKgDvNao1wnWwCny8A9Z8lVXHqB/QSsBfXLKcIOMmiMCBwHfQMzxsm56IQ/I6g5L1uJrh6DxIDYf
QhXw7uzrKbt1mNgunTmxZH+DPSZKXoa3BVJEBL5VmI6TIG7/cONlprd9Vw4ps45O97jtJ1hz6IK+
3wqabfLMkGaaYIsbG1oiuavFhrLqILrl1IVKVWV1K7JdakyahF5aIQNQKNRZeMaK3jbIekXaxpRI
ugqSBay2OGCUb/8i0+NGikAtEeVFvkesARQBG8FWfwEJUZjv8wi8jt3PFYiv9cJNYl0JlfBfcXTs
E6mPNKWJI1AU5GNYbmzZ2v8GnzaI77XDGeaXqIYdq5n6wzN3WW3AfEVX9bL+GH6nqfh3jqkL0WjD
VF0MbrYorhTBuQ+zbdCshbHgpLkksNnSqY1xAY2xICd5lEsnV6Nz0I2WMbTulZLpbVWfepgM5qw8
sv2EQZvyHhbeyYt9Blh7WdkhvzY98x4tT4Y1i9o/BZzmtGofU+Ni1ErPYt+h/2RTyxaL6n0y23tj
k+8EgvqmQBRFUhKV60ex+EXIf7ZuFa9gExfdoFZVRqhng68rBiT8XKSLQE2Y5sO9fODct5PYpefs
oY0fSauQdIyTwJQCKMV9M0WStuAODy8fcAZiapVT+0oaqJCmMCDy5T9xqPN/pb0pAXMwWze2ATTZ
sQhO2RuJKuhIh1skZgFOv+qzhL5rGtrUZOM+WR+AaDuG2/FGYvvO65CQjDiYjB+H1hw+0zcYBb38
RRxoq7suyOG3ymEoyG/fZbtYHuz8FAacxoUGX3nVOT84QBys1Zb4B5ctjd4FWh8eT3hQaCJzGglH
NmUbruLcgTGd/bCqn2SeZTyglhqkXUi3uPT0E5RaosQ2odgODW00FEgSTnsQw8gNSabosc8WVv1J
0zU00Ft3ZCerjKfbdEWhEUh35NOuA7C4wxDzPJXpQ4GzfBMOiV09VZE6ZFMyKSa0QBRxmE1dSnEO
PR92JUgE85a5FASXRmUfOvyZ/Qk+LtKJhky1qNOPpbp0Xyfp/FSnzsTX9q+mZYgFfGKt8kTWqTpZ
bSoW2EZYtp9gFmrebtMoX6K95N4M5GmwWP0fpynKsXrcjN3BA38BzHtVTk7LskmPlm8Rk5ytAqyZ
Tr0Nq2dmeXpy+uA0MngUmd8rTD6vcMbMIxDdmdKi7kc2qFagGIKCXi2ZvvvXk0VMTIkKQNq6Z6bS
RQYZ4UacRf37vSh7yfK12bwGtToVHsCgvbPR65+/Snjt53OO+duursYmNXU2Yr1fPFEtasCEFP7I
bixrtOXtC3SaiOlJj+qqO0M6LtO7AZL6opkOTzLfqUa+H/en3whcrCHdwfpOD/7eIZ7dKK7WISnj
/vNCRL5LbpwoXG75n+XZu+FP9y69FR+PrbzRjqik/dvPrn6JJDKKwvCRivq56CxgM81jBbg+WJ3h
pOl4Nf1hXNR+aDGal2yMRky4mmtkIdMHbl5IJABcQJs1i6mg0bO8/8sbQLrxxuVwfdVXnEVRJYK3
QLuMu/f179LKsP7TnMFb04qkPigSpGaRvpWLy4SKQH3N9ZCBwVN6FGNmdiHEMIos1k9uL+BgR52T
0Nw8oWVTXiEjma7evMqYKf2bwWdz28YETUmPbnFwm+Z+XGBxsceMdAz4SBuFN4bO1/yA9jxk7yAQ
LRPitmDO++GPMUq6qpyNdEAcoVMsgCv3kmBOCF1lxqJfRJ+AN6rTcWxw6F3yudcP38lK54caIupY
wzvTFodHAkSVMEA1MSQlmbwCt37p1Pxc3wUmGF/lQrYn6r3v7Qv8XA0EkSb+8iP4hEmOlvMLYKJR
/HY5SGpO3Y4IfelC016GUf9hipmgCYpfPXqdEoLYZycEjIH8iBLCppyMBr7yFLEay0fFE63A/bnx
GjfiKN4W1HqjhBQJtueoZlMmV7NH0UhfIqxraokhYXtPT9rPSIKnxxOF2VS/aS7bJtSGY9Aqub/I
toLz3kaXEPZYYmSDc393G6UBOgRKA2YDWjGw5pHkc2wRqNG8iak9c+2g73ED2DgZNxeXyiar/7or
218ZKKRxXFvOTJHJ3oGfZ7ybAiX/YTkunHVDxhqB5tIB/L0OsiCiVtx6tz88KledLuNZk9+Q9sGV
/wAF9YSsmAtcctSXfVuIHDcxyo+6PTRQsA4UApIObXhAYCvGyMbWagM0p40CWgbJaWvVTa0pdc4N
6IPXJtHVmXg6yOLfwjRtaBR8/t2c5UNoxkHtfDU65YTJfDDPZtKtsIcc1OYy5QIPQDXfltwvUm1s
F4QMkpHfJHvZGaYgkiQ3sYTVDFy+FDt3SqXjhXquT7MWhieoJqbo0zRskNzfGgwSZwcKZcwsWx6C
tn4VgihmS9f5mGBfIUK64BDg/8kt2VRsBWfKn2uxvCzF7J3zOVo/KEqIXLuyR3/T295uuRws+0xH
1b7CRbQo7ojLiaT5+moJTgzrDxZZ3WP9GC6QLUSj0ia0VyUSDc7pVo4B7Q3u723XZ3UbaGHPhLZe
yjELMHJmqlc6EOeMa0PW8pBN60df4EicXYLKjMuyDjiuKo4WZ6IMraAOEiRmbNMdt7QYuwjS82pM
tHo91u+CwvlyH/3ffjoCigBEJm5ad31aFfN1Dpf5FyeUDqINv0cYjeykBeeCIBDQViWhgR6scTSV
ihfxYkJJ0h0nJhaByto1jyH0u5IUbp3/LUwSje4Ie6VUSTgksEmDcguxHyYWSQgft7m/XgoCOkGF
/SI3RmC06w9CCmRfiOEcOyNNfZoO+OmAedmHvPKie8PehnHtzS7C74z/stGSPqpWERx0jPbjxo7R
ycbSJ2G1fjZxMUJo6r+biSWv7Gon2EDchFZdS3hG1AZ/baPEweCRND5uirvUcSC5MmelLZS1TDFM
O4UWQmtZxXC3BOZ8Kt87lb9Gdcktu1ZpNwYycVw9hauzRyrfbg5RlbLkRmclMvMh1YqikNne4KAn
12KmMknNUf78AzTR9z6TJhQO2ov08ROvSi87SXHMASIQpyXvniPAi93naqOHFipBmjRJF6O2+IeG
LeoJkV9qUg/3qKR/Ru2QPj0fVeJGZKfDBW9kV7gy7dqYkgIq0j2mk0c6mCaqwrTeN436AVFIcT7v
u3dZib3YfVPCx3XTkpC/EjVqhDkVhps2C2Afvk381kxXk7kCimffTHrxtqYQTThBxWZwXrX59Nuu
1DIt9a5fE03xzjML+GCUosE9k9pRhqpRJjEHAzN4YmZtlaH9eCO7du9sZflEAJqNvt1VPDaU3hMT
Uk+GaeRFDvl7NTXSrQOlUODFu3Ynv0uaooSuNkaUUmjnaGZTWUCCIxhCfqOIiiQY7BlhXPOwRspY
GKHcBzm+FQgHU/1DprE+voomOzntncyjv746XErXiK5xA4qQeojl9RJ1yoQnh5C8boMDDEeB0+JR
+1Elmh3CCqVoIqNGuGB8qgd1kZJRwV41Oai8dnGUy9zchpjyM8xtkVfpcN7kjzjDVPDUuilLVYM2
QL3rDk7qo2daI7Oa7dhHnmRToaP1vQKAKu6C839h8Hj9vygyALKROYvZRQws7WYK+HXXQQwMhsCA
wDEk5IyMkfk8nj2y/fJpbB53a9bSwODUih2MJJWMiZWM19w8UoKeX5OuGlBLXkfJQjq9CHIPnUaP
8/s2WPxpMHMaQ5W14tYRZSalri6TjHHu1cpWZ9r1uxXge0BfbvlURGQyTf1m74CHnuSbYPyPsSGq
AVkhItesZg3lNoeBG0vDrcjMlkiKbbQZjyca69mSuDp+EucZFl2exkfo5MiuykdlINa5C+0njJy+
GhBsAjHT7RCi9+pjhu2wKBYaqWmg9A71SsoZy5lS+07S6MSpdF+fw1ALEPtgN2tMHab0nheLhRnT
ngKvexi0wn7S14qSdCsQ2OMg24WfJ4f9hYh485WmkNyav42/b8BKhi1u9IgTbRAwPhFkgDKk3N8V
CcCZGYRI+92aD3D6/9TMFY038fmSmowqlEeNl5CEuHrfl/gIMIbat04C2y1rW8UfCZybrOG3ddIl
T+L/Sw+ciAxFCXd7oruV/6MveqPiI7c0agpiYUdzIfIH86muxmb5pV6WjpzRPTYV4AyC3ax8o/YX
rYuhyyU6ea0bjFPrsUDcLVmtqxsLwyqWC2n8Q8MiibKH1w8AqZcgkrBFmr5aohkyLWnSnAz+06yx
SDvdlcie6DtPxZPffzcanIvzIWsiL5AVU6bkjIZfA66ZxMEubEfrxJaOcKqegQru9W8dWdO7XcCr
mtuZMZmqLrPjCbnQV13lY1uKfmClqE7DQmYCq5WkTyfBIlt40JqFWhyCiRmwrJM31drmIRstQu4q
QhZdAsagT5kCcIwFsfkHP25/ebqvKYslNBV3cxyRwvohlvZ9aI0+NwnHZUqwk/lCogwts9CEp47B
jmyYQ/eCBbbTg3DG4/jdFTMfdy7HELQMA1gIsk4msjWfHIUqNWx3O4yFDD8B6r0qscfGCpsGrzCx
iyL8OTbO6LUDBYGVBt5LHF2UsrTQaPT4khC9D8oIHSKGyi55gxFEdk9MEk9S4ni6tS+kI8Ik3sBi
DVwVis+NW4DnnuJURnoueKSjnNdWtvLNLcQTyPV+RpNilxRTaoYqgy6AIhQJKk+D67BeaykUGqPT
MvrlvRg1k6uaiqwkKxRIzPsCGHjfbnnF9gKbyZJWcawmYUS1FInKd0qZQfanW1OUP7YNxu01btdl
sOPMhJor+97NrTHpJO+ymznYiUJzrhnH/twWtQFLBGW43lsCvST/5PTMM2u6tRwvz1giVCIoNSxa
0XVNpIQtz5hZOCzo5jqmGFA5ktya6j9WwIB2Ls6R8by3UptxDYHj/GhL49h+6KXVmn9rRoj8dVb7
ZxfnWEo6xQq0HZ7Lzq7ddktP4mEruxqJQ9KPMfBVsiy0xQS/HArHECm9O5pwLndWvew8z0X/SZHl
rxK35FN4P94xgmIj/KRtTum0X/g4U8DSycyAJUybraUg/FaZLj0fNblcFPWpdLWRogI/FUdbqIuZ
MSNJciC0E+X6PUggOCaeDYkUgyCM7GW6Lxn0pyEyPjXbncx7xL3M25clkiQwsS8VZ8T/7hREMgnv
UK5Yyt3oB+I8/zLrceSOlgOZPJiUio1WhDQG4i6LOR2H55FyoyEY+BKTHcoCo/FQTk0n9NQ8846x
j25zrBXOnoVY7DDAp7oSzcr6ld6RYYfdJLZRSU/w7Gfuz7c0oPGRbYBDPHIjGupuQWAi1XDsmMyK
GjtH18VXdUGaT05EuqaarPnJl7bSi9s7mfRoanoYmcWdhCEyeh5zggzZ4/zOpENLnCXrSb4wfPvG
u3kc0+1qUP3VP+0WUTcymuzfm/4V8+PG6UJ3wrrKHuCh0GhDcRllMpK0h3a5yYEuYW7VuU0xAIT6
1XIMJdoAIsIc6JJUqUvQZD7btd9tdv8Z3xHwF14VShXTLBXHspGVltN+msU6oo4PUuyv0D+Fe+55
ZN71CzrBeV5eVBTYk7PAOtzq9iDYp9yatO0Dh7i+EVkZvd//odRrWRnrCYh4fcvYAmLn9GFTX+vR
qVFpJfbo/xvJ9Atq3EpGZRMrz8zJCvUs70yxuLYHxami1h+7rX+XNTTUI6N5FyZckkykDx+xUcU5
Ox7LEcQ45rJBYf0BojeM+vfVYKfj5jlRDyKWg3mqcj2ApTA4nWmCp+VAE+wzu3SbKksXc+uYU+ck
YIbSoqiqKaO4oSu7GFXUu/LA0JffgGnkzRlmxDw4QIrYtGWtEZ0FOAfZ7IGtlHMp6DHBantWMaQy
keSk8cfsQ05eIlaDuw1KC5nIsQtX2JTq02qH6hZbBwJMouvQu1HHX96r3OwrK01iaO4C7Lra2ykO
kv6ugWukB8iy4qJTrYuLHY/UiNBR0evdefp2rKp7UWP4VXf8/HPQaJ47bRE8gLRgPsArN1S8te0C
g27uxPdTbuRm913OsdZDrbxts1NALRPZBaTo+babAw0wZ+GI4qK822vEYB7No1yBYj6gqfBTlM3P
+W4Zge3DrM+Oow0zrm8oSxXDvpFF/emW2KNXvYWNrF72TuecTwotJNCmI3uushtekcc9r4YKn1om
zQS/cfIClWCRJ1f+WT4FDcEgHGX+3Ilys1M69BNfWhXjiOeNeOkACCIEgZR80UDmFgJTEY9/mkar
0MzVaoJLfvKSS5codjOzemarbZThlnEW16c+R98C0aI4qM2JJ5uJ1VMXiZ4Gg30UKAYB/J0O2TbS
7k2OdXD/ukOmjjbvsEO8CdFanAYJX0J98YY9naSf5PfYD8lFxsb9OPhjrOviOYDv7lDM16OOOSga
hrIEPdr3je0HcQmJq4iinkv4m/gOtBOw3yEbhmEvhqeRuCyZyLV+bIHX5gKyXk4Tv8FX6lELrUwj
kUY3f3O+7TIta8uobTHL2Z/wu/pGh3yZ5JR8gWJ9+dqBFNvwrNbp7YK3MkScksewScfxVLx+3jBD
FL7dumLt5ilmXq2BU2m8wnOlgLeOgzfM+hzzyt2Lp6RtRSnYuzyrUKZKeLyc9omnGaZRg/tHY1N8
nTME/UmSzPhf76eRB3tFre8eeSlMID3GLbVMj4/lDyiGTcOiI8f33TCFAICsqZvLLuuM8wHXu887
0cndJ0l35Bv9syx2j/mKKfHlQlAcxWaOIPXqBMWzlydJNu/U/ukjZPusAmIIEjfh5+dyWfElz1RQ
RABp0WMgM1EIBp8gcKJouM2q4ulSn9R1EoyxObe5FqvLqdjPx+AN80XrugpB7z2EAT4eu0X334VB
50gwKDU2jseQ90QGzXE8RZEKAozaJ2iZ/irKa9CEY1FTbDJYi+eUVURDrUkkjeDj3N9EKCxeyFmA
FM55N6WngMmnONPpi/339Du+3ONV5+5cFs94rxYHTWD3hF6KulqMfaTSMCOe68msjcfPKE/KdEIG
47x9wx93WdFlznl0bqe2DNOopwsQP48FUoxX6Dc+azNT9SsfRX1L9ReoEqUZVgbByQJ0r1Cfeeu+
`pragma protect end_protected
