// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
v3y/EjIQvlS+XmjapEfriuOJ+DviL8yQFYvW1LiS2VjwsdwEnM7BWw50bQCC7Go1jEDqSefOizcV
T9ZgxvcaXos8SpM1ryECJyzKZ2rp99OsT7s664Sw80ft7HOXjeSL/7AH+RkK4eUav1QsrOHACyzq
r8oLKBDxo5c3tNvSvb5jtIFXRc5QNuJ1n7uKs6UrQemxHTxwdUnPEw7nAtVysDng603J+5x4k/M2
cYmWVnEsdEH+8hxawymoAnvA/e9ZUsJnprh3E6TG+xVh6Lz9jnyC3pe5Ydb6I3t32JZ3ribvca7S
NetH3iFmrjr1FHLazZXaMKEIw0dfPxMkb98xtw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 25824)
pKo0C8crJ+ZQKsyctvvKQXoR3L48H/fTR3FDNqWe29oEoWSs2KfmFgMIw/ckIbyov7rAkBmb/C+o
B3Fh7S24zXqDK1H0UkkQM9XTRyyFSKkX1FuHiS1vM17P6tA4p8k29+k9L0yqNjttlhDTWvmaHPfM
PQWzLniUkmaFkV3XsvOYKwnneH3RU0MJQDU1XWA4gT9vWAR/HPvUkOCyjFsvYMEy7o08uUZ78q9z
tqAbYJKXDKkdhdVE9iabvbWyiI2V9XJPY4W6E3kh1Sv8q3xSd/P7hFJZ3L1EQpXeDLsfMNzluGhd
wunzEwLpm76AgrFa6FQK72th/gpOqeEvRBsHSU8nurADoBNfFD1/bVpYUebwM63fcC9ln2DXwpuQ
Fyx+BkYCt1C/R0C6i/r6figsxb3+6HoNd17+WF1NisuQuUVUf8QWp1L+d5Nh247gIVjQVmQ5Euzp
RYUFwA6CAMPeKxrVWyJjs93Pr/XlieJ0B06sfd2M5MkBuwTeSaRO6XvZNqfzFzdPXtvZhUymI+TR
PcyIqvLGpnc2LYyA6fh9lInvdI6Ss7FtjJru+Zug/5V22vOpwg8N/gKMxVuC82cvqaoKbFU7uhDt
tDchFbo9MAE4kAxL0jU5nWwc66DEPocyRpwYeYopu8FejYFtacEVCXW4jOdgv8d0Oc3zpSxL852a
ZCNR9IH+pwonEZIovYlNNuGaHwbdr50dvzGp0QyOuzFtJQRhhCEkcPW6fOevQMmV/nECbKMTtUAD
XcpG5ld557FKMk9EY+mNPpcW3mdQtxRo8w8EEbzR94CPwhAtNUtWPcrCxVwRO+JgY1pvHMAr3nd0
eSHuvaB4RTVvPYLGsVcPugtBEc3ocLIN1eG3K/bGxJSRkiI4d+xHGtFfKvMwg0fxJRepdLb7v9Lz
ctYIn2zHojlQKm5Sv61A9o3O9uVHtuidCuDTOOzy3IaD35fSHo1iz4ffyytpSixbQEH/CHJAlaOo
ABlCFTc/LhZGA/qoBdB5Rv+jybox0/zbxObZMRwVM79zCdZW2UjhO7xZsC+MzGYTSCqUy7EpG6yw
YnkoadWoT1Mp6od193sdc9Q9zZVo/BHAWbfuZUeps4RmIxE7ccQFuZeKnE7Ec8KTJzCMzl6xuvlr
lDDBtGkRFqLd/+SnhQ0tYv9FbBWLKpd0VUiHaxEQsS6NJxnx+w4uJergImEzo6zi/IGiiOAMhxwd
cMnpdd6wG/RfW9Bv65UltSyPvdZtpqOHUJCR5Ttm83MNKBPtSLR9wKiXpHUK0SNK7DqalBRJ3erm
usA82UooXx0Rxbj9GvH2agmU7Xos9/T9FYQ/nNNOGy7WRvIcNY37V73WAD9SZQKYh+7LPFmWszjr
iiL53etCZLKPuRidHIytf5Kv+W3Ii4idrJBFupwwzNHEhmVIdp9brHlN1gBHuYZrfGUfXLrCk888
nwQNOzXnghurFdFZqVrY8lZymRK3CLn483aPzec+nc+VGUImmfn9ADNAl7VxLJ+W73KAZVZSrT7p
9UxIv43o/Ci98Pnhml4QC7E7f4GofE0TAInwhBJketKfPJyI4gK/xwV4jkLaVoz2VbXlThzahuh8
dMNyrLVscHDKG5wUIRSrnxbuR4xiGUTYmD4mHKy4G+sS/4o9eATvbg9Wd5yid4l05Po8/SH6Urek
dbcom3HJUhzEsmNZT/hgEPklUBQ9rXt+Xz7R7xjJxFS8I7/WPZgKnJ0/CtGPEMl5WM8y+h8Twxsw
6zvurGrQZW3Unx8x1DG546fKEfPr4BV43A5tGkTmYtoqhD6LD5fpiCaO6X4rAiezprDPHe7jQfnu
mGpcXqAiijTfYexBBCmJfPNVbKzId3T8UpBzErwOut0mPAJTbcvBmQNqC2KCL6NsV5loszEdnQNx
JIy3iPpLFzPcRRhQcYp1wPKfF2Z1bZi5G+lZ6SAEd4tSxfciG7Rdy3OtkElkOa97rigZAh8eO9uJ
fDpxJEDr9gAEGW4qwi6HyoNcNvE2EAdCHRIARV5MLbhYYew8hmqd7QKL18CVZb0TTY6qA5pMZTYA
2ZeDqjFzjKYAFQg3UGlaisUV7q91hFwyR7BbqBF3Lx8p4FrB7+pL4M7QcDTxAeSFnf0MwLuF1yfJ
DSj4B1KmGEHHva9r6ubThGuVh0YO1ZcwqeO+Hmjvhyy29sNffIrU5qyjPCw76TeBs9v7TRuQjQaI
wjlcqvBrKqI3wxYhV06eeFnt8isosvi1kwB3Z/hInDkQLHO3KOK+fb7BlGNCq79nrhET0DUdoYOO
ctDloHrAzONta/fgox8HjZrGGBJor/TUfyS6QgN9iFOOpHADC4+vOuZGRJKJtrAuDTfTajXcZGIK
Y2Qqz9RZhxcDIOENVa3ro+szAqnUbzcZ3/VddtouoiOjJUpyK7QNLw7ZFEvWq6bSIPAdSgaOfVQY
bJMLQh6ozYyBWe+Zb6eIpU9JKx/uPzSOSaTnisrPtG4jrbiO/ke29eh6ss2wT1u5ggGNiz/sJ3ak
AS81RiSx+/VFN9tfdeDtXmKV1asL5DBu9Tovepc+xkPTd4IowdxfC/AQRXQOZyq3Wj21QaICkSI0
4go7HwUBPa30IzYYpoSy4DoNQLr2DOpm0nYaDFQt+nZejtIi7IP2lARDfGp5oJwM/IZ6UNeQ0lu3
YzckR2rcGUdIctvPqnwEfnGXWG2m3hIefi2ldBdTZN3e6OEIbBhIZzdrGofFwnWYBwfmKYjXkony
qCRu5vhKhK8Pe5qCO3G/5IFjqu2olu6binbdc/62vYgG9yIxQjKgqe34lere0IyHcX4VlboTscLk
ToGR20cRSgIxTsNZMSMdp82RmYgXxHAHqPEbGF9vGya5mOilzj3dFJG3eeNF2jA8eMrNu9s8uNcb
7kmzHCwi+pDNOQGOQuRaro57fX3GxZhdo2wqPEAExCH+N8qJnRcEC90KKjvCw/hL90bQRkb8wmtQ
j4OUbX7d/heFCC+xIvfpWVRn85h2NCTntJ1QNI74sSNwwJ6SmetpmWI4+Q08oB9OrhuShE9Jawux
I0ZG+4WZIAsKZZlUxfAJ5X08mLIeCNVtxrZuhpCAUIAR+xsJ689ELcd3+T91zqC+FjveaujaDYIc
Fk/aUg+IawYU42VrxapsHEA+9+z3vpbF76G/YmWJ2QIvRM1qpXQBkfCHZHET4Huua8lhw7OoTHrU
ngmSa2bqnVxKd7Rrc378VPziEDBAR0sx7slNAtaTPhV5KkgdjwYKVT05Hj6BoYv2JT3Nw1rF9X8t
fBiiM44OBiiQOMrPKsgZM7NUvIRIKxw9xkdfzw63K8MMt0aKFHDPn0ifWorSmA4IFCrGAxh2GAPu
dk585GOrVmvKQ1D+yADwTZcKmHoxYtH9sroTeJMrnyOP9AOASWb8G2Z9miqCWwshrdRjfsar4486
aK6/7m6jIVfdwL8maQMfeUKGPrHCEBlNwU8kxl/JQSNw4Y/SeaNvP6KeBU5rcifdXoCzf68oo03F
Jlg6Cuko/jo6ZkuDa5nrbmU8KD4vryDu8TPHEpHOk1zCKQTqnXTuwzF3LrthjFKu7PHSEhveMqD6
0/BcJkjD+2LrufJ3C6LlG7YbJq5kQcZ31wWP4GLY0FN+crVHW8ivzWKkohln/zjchg/+1PIAWLVN
MEdCE2naK6tl/d5rInfOAzCT9cdWbcaspOaqaMnhzNQwVSp8yx5G9gHwckOWadXwrix9ugCSALpD
UyB3n+okciEfIl8DaNuF90TsHn2+rOcQYR5MR5KBQoIKIPdB9OwMnwPFJTiSt97eFm5q+kRqEoK/
LEvoXuL5KMnCiLPcpsDhE1ObuML2/C63rnI1y31gFzOP2mOUVHBnhI8RzwC7CnnWFguf9He6OpHS
dSn217CDz4GhHykpDMDL+khEkFngS5PelmHU9V13NgQkvPL7NMh2AnOCICvibNSL5YmYMLbATVYK
pPfTyEEmFajkOuSvYo63iQJkiGScmKk/GVkNiRDw1dUgvUvd5yQy2Warecgq1Zawb6RS7PmbTywQ
bKNzuAfdWwY7xPGTEbo9GcB5ECaTcbTZBQpyTDpqBR3hCjlXRkVeWHOJg9c9X4BuWaGSTNCmMIE7
uNwC4xPlgBrgbbM9DgGMXsmEvOAMsLEIAEJe7OIEcWMm7tK6DHvX/Umx4exA3ShaaJcyeYLXi9ym
Bk73UPnvOZ2mORkuh4geDIkM50kpJVwOGaESgs2T2UINzOEbkjU9cNV+ldy44Fy/1TeW9YW1V5FF
D97ObjPEvlNyJQGRELXYVvbfB2reDs7fFHh9tYekGt00zHeK3reRFRGJkShwQsduNRDBdPq1PVId
ikzoFGioMViiospfjAvrdZPc5UyE3OmuKjiapzC/9ZoV2w8l5/Mnnj1pTWuFhGQw87UZ1CJza6vS
Ii6BZLswLPXt3NTqJCR32JURBu3d51XIPE7RoKVKNCDzM44dVVhKa8+eL8AQQed/q3KHqFAUn0Iy
uubt9SUj8GwCeaiYU0cr56d/O2Wy3nipLEM2ju1e6+o5gS7gHGhw8qNJKaRw4aRyVozCNmCeyHgw
V6aTojcC7u601nLT0ajjWkUuj14X0lgDMbs1FLeGb9YgmuGjUh5fcqgcu7hJIv29i1d9RW+2N+Fv
B/JTqNi3mVUTY5bWI9Njjlf2UE+3sFn8GF270AV4WudgHbZkFewttb9cj+XACWqG8Vws1yUukxiC
tQttpFZ98P3oBoM/HlQlw7kMGvlU29zAPcD2zG+b83uKw4v7odNl4iIcoEv+4FJXRWN1GbvLKTBZ
zbDYlEli8szBgmOCOW4RIyWNtJRyR/1ZVZp5T2SqEXwnS7B5gcDtH2z5jDHa0mjrhPnb2zYWtz34
y1Q/6pG6CmZj43BxINMeEP1EyIq9CVdw4Ej5LRr0LRKg1KcEITnez860dRPFv+siSFT8oQmYZkxs
AG7PyNzPQ28IvQN475mUQ71ojACNQWfj/l1HPqu46dtc8KM/Xzf+77NW8nxilNewP1qF2arq8XkA
IP+8dD7NsM2Y6nUMUeHZCxhguiRtD4bHUqizMmReq3udO8V4SiYx9y+2fX/4xfCeRAa/3qmyc+nS
vplRg7AigfP7RKdraJ0g0ytWMTclYjL8j+XIHQtZyye86BWhfGfPGXmZD+DEPjgD8XIlu3mc7dCC
x62QUEh3xCZgju1fNqVO9tKYzF/BtuZPJCVbseY82bm2L7HhjE3USIMVgVt8jwQhJCR1nvp1LDaV
o9jRrFWx2FXpsdEJCFtM6a00oq7QKFkb91svyp0USVYj6Z7Tx5OWPW+2iVbja0G/m1vxjbXvZNnO
tC8oz61dNBM3s14f5n84JmDEfnL3/B3/sN48uZzxVO0Es06dADKr2S/CRP+M5mk9ea8yoDA4NjXP
dHRUgg+MZLZzQ7wckCT/9jhVd46Cyai0VjnwHM7mcmW2t+0g/Oh3iTnFwvwDSQ8vOVh9qtqgphnE
dWVsg28SF7c2CBnw4MqWvIkQkNpTNA88HMQCr+wvDziqwNx3kQzLENxAamri5LPAA/jXg9UoFHW+
t+pXGF9OBQoVvliLnoo3hiC+AxyVhWJWeGBsoDSk6GTReyy/28EnxYlFiZqB780YWHPvQvg7o17R
p9OzFf88I30no1lJsGjoDlwv8kjGa2FtuuiNU/4c83TC06/zhbWfFoo5QKGVgKbK3k6d4epMEnHf
rQrrtOP59IMFxfKHn7kyaZt/ttBthjinS0SuLHD3v+1MhXeahm1W1vbcAHRF6xLqQki4ObtDM/CU
834hU+gmjNvA8Pmu+/5dEqPYyTfdZ7ZHH56x6tqLbOUr6ZQYZk8IvkgNqTZFv6SMNfjFpD7ziiXg
tYGlH18dJFpPow15+4scA5Wnvyt4S6szp1rRde2hl9X3boWbpIYBCwi2OxAjc1Tw4uC4vCOtlHG2
z0ewsijQ4s+Ajfvs1EhEBjp+RHlGR/Oyak75SePfv6zx/PU/EGgmJtalotv5xm+Q6v/4B+wY2sa2
jOPpSescQlAp/dRnaHPAsr9VxVWBWo1QOcT1GkkG/w7RyYKF41SfBzr3/QdWcDGTWNwpBA1HLfk/
VLz5ivDTMYwywQXAVLA/947SVxEGhf5uzPvdK4xcI0XsjQHNk+JpdWsqZBug5Ndsgrv264poXPUI
4L/+FQjY9GEawibY1ZTN3AauIY0i1BeD+mnZuuWTo/i6q+tDXwKY2JIMzxXHITsSAzAYddBjxua3
Dsof0/vNGrE8+OVRQvwwRTTx7o9wFrQLAYJQ0CBywfpHv0AeH/ewVzIzbIA7eUe3+iOMYlri0V3A
bfEu5MCqyG9gpWgztMnAwp5Q+Av9bGj93X90bDBUhWISwqNRbjKdl3TGdECD4FUIF/+O0YaPwvs1
xX6J/pIVWFPphOi2jS8gP7Vw7Fn1bacj8WL652JX4+dS2LB4TtnrsmQONnx5sldmsxOo6R3IgWxu
HoCp65v8Pi5O2gUz8eXN5raC7CTAUZgWpwrfUmIMFAAHNumbdbBQhoOY8ZjWrHetEMq5NlxLmjc2
irvDhqWe+9dRxvtK4gGvi3/7EkSVNapTaZaEypRBi/qAEhEhmPWuROFZAGQeqUXEmCttNyMslbNF
bzzLdiubbyZDGxb+o2xRLzV2LhbBDIb1nYA9mymhcQtdQc5iMtR3MbY00MaLHvFXQZjFnwC3x+NF
Cv9auSuwzpqHTgnF+E261eodpg1+E6bhGb2Rv25M8gVrMTPq1mKtV5/OD4rF5RVn9EB33XDm6wOt
i3fcwpQmkYL2TzStKxlb0RHmjlIOpUYBntuUFSnD1H2Ez6gfeTY8RPDK/zpQM9Enyjd1PnoKs+du
U0jB2nYOkuDW9nJioMHLDz5HcQzc/+GhJRaXWRNGX0DUIZvTR5VT5Wg6S4WrNEFCw1rZICKXZgSo
kLV+y4yqFu4ajVDw7JLeTf7JE3AjyVvs0Wn/bpTtX2Ago2hpR9CsRXfEnMUcfz79Z5SimNEH2Jmy
VjRyDmMgiJDFtHqHbYXfFIG5PDCmkALb296mAYJfOrObmTDYTFnQFYMUcbF2cbBLsLrprGpxAcHh
JqxnIoivFhuW1KkxiCJUF2p/s+KzncH2IazZ2KsrufK3u5NvAbN89AXeYo3m3U14UfGRgQ9v7M3N
0p4uvH410V35b6LX3BNokyXtsdJ68LxJo+gaAdvm9uLlqMrjwF4F0ZyeaoNI2zb1z9oz8nVhSBVn
emQGLOAvXk5SLjlbuSYSd4bnoPu7caOWU1MiwnwLdvGCB7gtBdCodWO+YPM/Io6iDNjL2Onpivvs
ujYOYKnQDjFQK4G/9H3hSDpkodwRgqBK+WfzEjxml6GzN+X7dWngItgiqQ8KkepD0krKFScNc+m9
6mgWGyYjKuE3sqc8kFAuPbsNIjfNArBXbxYTaFiCUWkhddTi1sXdllLO7xT35wu5me09lYAmWwd5
mBWCOQptddamwLFM2PNj4r890rKxK1rKW6eFv9fMLeHqgOiMoU9tZ1jA/nyOwgl49ojUKqe50siw
hSkfG0k87nKxntSFGp+8uIEvhzcEGx7vYZwJZJsdWpFZEq9uibcu8JCxlip1l14snN4CQECqLfpO
cWMfYrkh/x0WJG177AQrKga05MIdgKNbP9H6xHRI5p0nIvwoTWNA9F2TT5quuCAzZdDDTVytntbS
qinLRlLUsr2EPf6gaoZdVKmgInmLFN7+0KwsM/awXTyQTmcCDXNQOzY7zGr/c+VYknNaK5/2EvY0
ASWMP1Jyz3Zkm+z06Dk8cg/ZTQvhW76C2w3NoH3DXLYH/0XH3KaZtNRRilXzxAz8wwRWRdmE0BoV
oXVl8Xe9rhFFjQi7UZaFmY1RX9MHMKGVboVZAh+9z37q8cNkkQvqEoTLEkeoiNYmewVjl3r33HQa
FyMCWV+36KHyjj/DLkOmWGYivf8LMxLi3hcoQ6uf9KJttHYMdYFT8mdHOTEELFuKF6YuxF4T704D
vbl7zf56ASLJxlcAOVIZckfx6GMjpEf1lMEdllEjzw/u2DEE1cPXi1GMgCYHvc/M5w0KxwhuPyfv
XTBtVB9K2gpyn8fNTGXZgM7iHc44vwbf6jr4zc4F84Tx1KolvXFtK9ionjXDPtcdXoslds8+Qs96
8F0ObHXtDYFbz6qUzl+++oEZrWY7scnopTb2Z/h1JRhvChBKG3zMy+YllD0OYydXA0n1WUCUvC3y
1gZCMioJko1QJ/rN2icbe7fUbx+zeNHaw8ECmO08RaGVIxxVmPy2WjLxFjzBlOjZ+0MGaDr+Q+mi
G4cQ63+otOF3OskZnbowMW62OPZN5uqSACNueKFB5RUwx6trf9ZHIhebZwcwD4iPVvg9hus37Rqm
pcU2x/MlTUNAcvGw+k7NWEIOp2mX9RJOtoEvMLH9tPucV0NyYAZQzBkP7A9z/qli9WMebIjEvO/A
NEYto+MyW4eyLu6xfjxREMMv8xHBIv9Xi5kFc9p4vAlEwBV0EBPooJm3Bisz9so7UahEPamoGPav
M8ik+NOxMRsaUdc26W66fArczH/nJAeWyAXZqrZXdx46pf664Twjdj1R9KULQJg5JTGyl0cOVuyt
Zq5RMmHh7+rPuCYE5JZSsS1fN0M86Af6VgLBwl5Pve+sUm2dTKSzLO3emBuSADAzybqOQUmiH7DV
CAMPmuNvWmfi6/jYRKk35etBCzz5irfaDZuSwImk9xGScsWDlEXZSaYulYd4jXok02TZIpVgWVUC
J+ff1I8HK74c6LdcdEnC7X+cZv8RGj/BExKDBQSUhZzwOAovXNGpzIQxBjAJk3VHyFECsrFSsc6r
ucDMqeYUVQ+6LBswz7cO0mGmr0xPWetEcoFEdb5oTYe63ivJnkMvEg/lx+WWr82WvN4sxDF5tTpu
R/ijVnO6pVYswOGqOP0Fhom43pBm5ji4e901v3CNEEaBcYiF74+N6FMiDHX1p4sh2o9Uo5mUbqzk
vvnRonY6IwOHlR6ESeGqaH1JFAt/GEgvspJtAwghNyQl0uWkrB37Cee4ZOpSu4t/4gUFhXEhhF25
q3nwI/L1fmJbnh2fr5VlrvbCranX9WC/CKNtolkg4oJTcrj3z9XEVc3gQ212bB4lHM0K3vjJTIK6
PA7xppgmeIbVziToWv4wy9ZLu40mLfj6KPnsUF6CnFoNuAH1I4b+erzscHG/uKSLxNIWYNwzwEW9
bBN1Lc9sOOKauwKZRgs/e5tTy/nEI0UOvqFVj1gRswzaTYSL/PD9M1fNvi2/Z0I25QOvI11AFrY9
1yE/Eg56JTzPgHHYDVl1FlT/qQIu1a8uE8XQ7jBDiO2Hr2Lokmam8hDox8Yb8WAkMS7h7Fgfw6v3
U4ccaO4pnOW9zAMnUlBDwqMEujYfolp5PJEvwKNPsa+uQvt7JS8RbjcJVJPlqn46QB2FXlzO3d9C
YHuVyWRWO8cg2RIFwtY438xCUUkreVguBbJmkGsO5c5uI68+6XMMwcky5lwXET5pVG0lf1jha48N
bKng0V7ms/WrRvxh/CzThWWovVlD90PwJyzhzTHdve+aAVAL+53pGjC9yN6Aa5cjVLpA7Hrhb0qB
cMEnKQMsdLbNmPsUqYJ8MSVM9KasLFSUQ9MQfL3/bEzQ7SSeV5B7HkwfZYbM0LTCicZdweM8sJD2
Yl+n+uiQhYjpKfCq8s9Qcq7M6VpL6PBZlJ8iaCnJwvtymeeeBE9WZPNHb4Do8obbeS7uOjL4TPxm
kP1g/48lDbRjI7ss2jyFjZImcDJOn25vjqi/kgSL19eiusGlTp3o5y9ZS3ZzK+4JKAi11GtqwQEE
uE1VRe0ajln8M41KixkWY64sdAxpVcdhW3L5aiuCGNbfExSfbbB0eUBex7VaP8gGMA8QhteIuIJK
qlhrKM4PUqyXmnVJenm48oMu0WiMBiLunEhsRKag3NqCAqYNP2DdEGvaadVypbG361dHyn4SCy1p
fs0pO9Qxel5eQT+gLsqfEI+2iwmJYRG1BKA2vB1e+8ilY2wm7e28tXLWMl4fxuVREpiq8Cp11i0y
Q32aFaF9/Im8I54CeGtObHvSXBjmCt10rnsssgLF4nMvEJjelF3aygoUK5Lmgnbj+DLRKEcwHzLO
h71DQjw1Bc6ycbWm4Mzg8M3/vhLGGCyZFlMpKNIO5ab06l+1J7lK1AU0xo8umQwfvaoSWaiKuPRd
Yc3iXKuAU0/o7/FISNFm3NhVVvVBJD9e9aMhsYqBZFNOmih7KWT+nsOWmhuR1Xpzoln7cls78sOW
v39j/1zqqLqltVjHB0VNFRszJCBrmV9vuf5up0iwI3OPihMWaI5CXv1vGWXbqJKXlwFVle5F/1N/
k2vIE+BBGKmRQYoy6k9cw2yNNKt03q2jqpi2Ot+moTuqOBwg2YgGHSfArXvCxorvDA/SQI+Qx0Qo
CQTMfTNGkZBCXAzR/a5z+WGIpEBw0uIGgcz9Dzfs7ki3OrZC7gAss3xF4aAZi6t2D711Dv8yjMcx
Q5iEeiFL2NFJ6dFKP5VX3t+big48FgkViSUicJTDbczd8OXY1txtMVJwVFCrtrqwytjtGjeRevem
n7ukTzlQVJfOA6Jy7FIoVukvV+Wh3Bv5uJBiXCsR9bPKaZxJEgCTOhyDvaYNeyQ65MhznofBGkVe
J9Qal0f7J7yEc2rdsWx9e7m+2KUnLKX5mq9PFB/8qTNtjGwjzOMCKvm2QvvmsoW2jLA56vMy1UIZ
2WQ+nMxUP11gET8eib7EAOQlwttqlO3Rs8fUy79naCse26W167UnZKVKdBHQg+eECTgEZJZNxRvx
A5VedOPK7Yv2ITe3u8eBH/UCBSKMvPmBJCjvdGdzfz87zSWm2IX14RaGHUT5DoEyl2bxHDQg4HIE
hjZspW/rE4Ba3k43qaL7+BwkdzRzTd/htOds2mBOkinoymGNZHyZNdQnrpkzkBV93xjOWdz+tuXb
y6A4CkfyAwaMWpD45YxEy7ug6geKTSq9e3LnunTVJUzakeZWBro7ZIUgEQVUY1OJ2D7MOKSyGvRD
HHgtl3u+AF5osHmygtjJZXSLRKwRm3v/Gr8ZVhBcJjJQeVG07bKXvuPiEoqLb6fB/Y1qmagw2ljm
XpbdtIrxdzly6GfPuzMs17LG4ManhdON9te/MdlfSbC6dcn0shWTs8y8HhktOq/eD6LUasli3JXJ
PyIAfASIQ+bptTYTiWdSUnZNZ96NTsv6ISAs3K69Pqxxcflgofr3fHDKEcjQ/D3kIRlBRLxliulL
g0bAAjBkKCIrcQ94s6VX8FBu0BJHeamzpZSQN0MG8e0NwKMHfvxFGyLuSf3H1bGCADaUeSFOPomM
f0nseNj/1UXrPNr+iwHFrq03wdUwulixlXrVw1ioGJXPsvh75icmTjQ1UweDHpMnFr7r0/VZevis
g04nIgratVEhY9NBFsK3g+18K47Xh8CpJ04vt0TbKCYU0M26Flk50DQsahaNW+B7FVghudSlf+PB
paw4oQPXg4DbHGUnLJyv4E+8DzDy+enNvWX+MtgKux190Pi6mBwAyl/gRgCvGsse4eYg7EJSe5XP
EfRlzORTFKqwVwL5I0+IP8Aza8sMCRmhefQ+PtbsRyHJR9YzMMOhRXpnwlAD3+LWyecgkz4Hd0W3
O25jO9+XBdmtMilUcrJbV4MtyXi606kG6dS4AhrjCCvKCwtMW+OfOoG2aKnvOIzmqqQArPUtWFpc
Uv5BGF5PGibAXyG/p56tIs2qAOZA03nq2MYNzwyWJbyRsZXNuCOsObGHbN+3+aFEVBMwE7EXVfjV
7MiKEGdI5msmj73raP4Yym0RDsmzqtikElRK+nGDyon3sOZDRi7C4/aV7ApjABfmqCvNTBicr/Ni
aLoSkoyxxIDTrx1DZ5jATJ/rKJ/OejfBBAIF46Br7zaMMw11o+2Z5qsRMG3GrGrgyJGU9U9VcCvt
2lsihs2q2GLTYLvd82/HTvORas/pL8zPbfsWEJAMLB4CamKr4YiUq3GvdV2NdcytSV484pT5v1o2
KDeifvQ7vv+evRCRprJDL2hdhdlwtSViP/kfLEkiSDqAwnLO7Vm7Y2Cn4QJUs8CLcy3mPPnGr+GE
Bk/BqdNZ9Ij+vaR3/PsZ+8Uk99Q9Yl801vBlfFQ+DBycZk+ngpvIIEqNfQr7ub+GIswNooJqSydF
6BO1QYrgzl7tSCLI2vPXu5/t8IncDWsC83rHR7+lstIGFGylEbBOZAuZZVbVr/fMeO5N8QRjaEb9
Qe6lBt6xTk9dc7IBLIyP2zsEPgVKqlWfUt3XftoGrf+yQPSTXTUThcivFp3ZcTrBudjk17qOLy76
N0IZv3wEkpBsfi/i1SdETCo3rM0OSs5RmtlmYbdGUqKUCWKWZKzz53gcjEvT4YGTHhxfmJ110QnL
bsniZDM/h4h88ZVpU3BVX0xB+V2CTtqCeQFl4i6TrrOSDMik8N9xkKpMUXC2mSXmiN5fnMtjoVH2
X2PJ2QEk1u03jm3csH+DYYD3sSa1cy66cJcz05EaUq61X4I1HL8xKPAauTNRq1SEFtnuTNgCez8R
/p2nReUmIzgFJGS7M81vuKcZ/6yVjuRKdvfFC0nZeEFWVU/PA6U6liJ6H9cdQpOygejfySO019kX
88YEo5TrshaO1VxWJhSKhIjqWSmBTj6xuGuY/PzyQUMPlRvIesDOixt0m5N5pyBueEou0Q9AjkGb
eXScjmnBXtKGkU4O7kshve7vdaeSC4mOMWUaFZzu6ig0TtoCJ74P2h/5uMGumbldbSH01BEPaDkO
JUIivPSlXg8wBHp3MDgsP0u4h6sj1NtijreW1v6EY41xLGy4wsei9IrtEowfgITkCpi5zqwk4VrQ
E+Pm4XyYOE92tLhLzogniPPHrScHmies0KGnfX4iZc0Xz55P7hNB8Zx3mZpRZg4mxpuwAfn/tHvV
eYt4ce7m6EWVq7V93CX5gN8VShPvCLqCnvqb23ty7SuxejDNkxPE+tHQswIYnph1+7TZVC/4F3Rn
zKOIYVhNqS0eyLTjWVdw76QiMI/8I/fVKojXwquLI0gDpTkU+iQRMveXj2V+aTDO8bcIzFep3vdm
X1AzWO8r6PGoJVxj07MSqr382JU3HrUou4BECaUatwCUHkI8lkm4p1AUklermK91SR042IqtZZpn
kjidMv1oj2H/F7W4TW3cai0NrlqCFqQZc0fVth5KjGylB9S0g/ovcl4/098c+6t7G9HGjq26TvdI
cEmMnhn2lOrsRxLn3mK86KjIKA/g1AnXnLuWDqGrZ4EjftK9ltoyP6HkZ5bMVIblbGrY8CXcD/xC
GZ11dy0/hbMneZpdrfyA5diAc+ZkvgTxI4891ZRRtxeh+HSpqckncUBkOXjoVxzMnhpyJCVg88St
YpAUy5zcFJ/M+pwtb0F94kAq5+7KzRYCuTsMnwOSWTZqw1Hfpuky84KrerTBMqC1kUjnfvI5ycQx
us71fiUjSRrrjW76tKEoos/LReq1aB9veBjUPayvaVstIF+CND5A5A1dcWLGeJpKJUstMFSuF5u9
Y2CApeeSGoanjrQb3Gb7Dce0BTGRiTek/oqLOvJT+VAgP5ZGns4z2Rt3a6DFjPt4Mh2madHB4R46
x0Z76ggW/8Q9kaziu668hmbcYtv7NIs6cRXz5JpFxhNDrzsXPrKLMfHPtIcdWgm/+ZdiRu3jSfzA
1tFDo1zspTSNuToP3GTrrprWWCG4k2IXQKuDcYQ3JFbO8acxVRBMXIoUvtOGqBQcjq+SAypwm7RF
Hw98+bGRDVFX3HMUBxqpggiKI573PNDdxDv8f9L3fB2DsOlb7vyJU2Qs3ufrKJ4pjzQIsHAHTYwZ
EllaOlPvjaaSAOhx+5Y9VHzAcsriTI+XCKDFCUViTnoayUj/p+VoDToh+mac5jWyTYV+NHMkpd1b
Thvc67Vr4RM4zoXRejTmMtSgBclIjO04MA2IMjdStorPrnM8WLAtXysMKx+X0OH5qNGkea6yHNnG
AXCYFY1j7ihP4Ua1uydSHhEfqS0yGZPDmqkBYjjeG2TfalE3zDK/NZhlpenxhHKIywiCKV12ZHJR
dcUMjPE2JW6+lVhvYU+xdmDZCxNVimjm4VWyHaaf4XAOvNDXTdtEGLRM0QxysBfYvp4yRV6ydzMh
48SUbhb5NDw2upbrB0OEHXbaiBMuh22+PIBdjOpcE7LFfEtZFaOGd1VL0XREPElg7zi1LSfhI3GN
VKvRRLCdsoHk7C3jMH1PYQFnwvKm2oj10KcmzAwC2KOpB6KeHXWol6Yjanw0+mn+ARVEaX8jgM73
tcOnw4jLeNwmzWBFOca4zMdNrVxK+MY3f4g1kYFmtb46l4g/r682Mla99pOyQZCF+X6QcyhHOMJk
u81YYmhuWwP4Vx1voA6F1YVZbupOBNK51kt0BkgFcksGmxchMPSOtKIjqpoxPmIG/yP4jLzgYwrZ
SPlIz99KYwYHtIKNvBaPilDXm1T5zqDq2amsAQ0xER+RMbxE4AcBKTSdZ0HYjAOsxd9rQN2SOylX
FIElmSit6AFvnJgkuosdOndAV+OxnLIh06MLEbKW7sDP5kSrelhDRm30afCx/fBYk5C+hPUbh/Hs
oLxVKj23P1CaX4zBltpUzv6XOQpaqJ3zsqLMb3Zlzm6GDl7yAOyQTAyH7SaKnxWaoLPvYWWPkKOt
eOubSIOMwm2tE0y2i8ZtHPxVNlrfAshLErePepE7BOMdDzVkL7OpX79f0vx24wvR7q/f1I/6QQDv
4qaJPSUAV3NsQ9fiLBmnJo3Jx/gV0pHA3kvkp/CotVXhSCr2jD2VtHFvTlatpSY7rc+l4GT5Aod7
Ekg/T1uLXxztKlj7c7OWTPBJ4YP13Fw788ONe3raNFYEUmNQrDcaiEghwAUPgew2+34qfhu//T6G
9//n3OYefjCB8Jx219h0MUYAn1VFph18OvozY9I01AMRhtSpTSHHx3DWhtRWo18A+iZkbxdMsAgj
cbmYoxDpzwTgmenaaXVKDJjy1YQHug7nzxMvvT1UwljDCju1c+Y7yAMZmdkw7lp9THzuzoZHZhg7
/r/YtvPcVM4SON/r9fMeOUZWq5DV8Zone+EDD4g+4kRaLhjCzRkmo/nY0WOHsSxBMhR7UGUZRcFF
VWq5PL54+JqmkqznWbE8R8axJpjz+ycQfO428OF9A6+FTZ9QKplAtbtoR2Rho1JpOeKlgXNxHdJ8
c2q8yy1fwRfX+FGqKyMVn5dLNWu3+zKakn/rYaXXboPdcUBdktyh3DN5WkYa7B0/1EeH41tg/csy
mKSFiFBu9B18cfxB8ewQHLk+gKw+jAHjIzSEWRAKH9QsJoKuGcaM2RbvIKiMoj2G5zjL0CWzsVv9
9SEvrg+KxFL3eW3i+LJ9ZVrWgPujVzaG3ubXCLVNyhA0Dkg0eepnnS+5n/ZfLdFQkn2lAwnXiQTN
49Qyyk6RJRM+BcuXYwY8Ygm1WPPqrSpB06Kwc3+0PrScjNfvxHCqUP9r0JTpIVFvcL8tXP+Ro4kp
slyonmvgcbjiCagMdwVRb4BPPZ07hY1wIXir+yXI0G9J3UXW4AeNIjD99NXxLdNOunVPgcyY2K5t
eEWBUZhngRzT2iuKhDG9QX5qx0NILKmE4evcK2Co29Br73pmefPY4X061hewJN1IC4fwwRlhDpvQ
mVXA4ZVT0wlPqYLb7T69N/yELWLuw3GDrg/nCmorhw/CkRCSnf05ic3c/U886EVm/y8GPBLOTtGC
Pt1SbUxjFNCGY2U8iWLc8VsraYPK4/kKYC2IH3f0r5N3SGu0j/dc4wmjwatU9GijLM0YlksrW51t
bKLzMK0xNcQh+fMST75ROTdKEFmpWast+Av0iBXhJrXZqdwyrPbehJz98puIRb5eoa0DXMjLilDU
syjb7IvxZ1AYrLdz9ezEB1KBqpf25+602q0iXBvOsq25LyIgdY55bC7TzO2a6TUkWdTPPq0UxQVB
sLl92U11Fa/LLqpnFirgt/cvSNhcv74lshMncYEDbEjqadTHBR4kfqP7B9DwVXQGuZLUgFxF5Yeb
I0Dfv4aRh9oPGzgpf1LuK5MsBdCO0kYB4YOjsJm21fwME0dimewRlcLe5uYpMZj7OyvC0L6hO8L6
go+E1TX16ovhdDDZm6pCyXGPFuXtDzpPEyRPcl2HY3D8PTCF1U8wnLb+Cn8kjeQeVo/oY2WWhPqG
BJxhFz3hCDftambUqOkPT40RKrm8B17rKhiNzIf2PUZFRBx5hmApFmBAQViubgWyvX02hmsWZZCt
fWpsQRlRRKe9jKpLMIIWbA1OpAGXrOSUzN8LelkIItLFpBthE6PGkLZF5wBwVeUxERqjJOEL+9tA
ximNxZSn8pdYjVaKjxcgFUfUipoWhrwuGsMCnnaHla2mYclZXcVvmyxXS6/wuSbB/sN+9iuuoJ+z
pdhlpfUEsI6RDoeNXi7I8sdLdZnfJOFVEy736KDUNZ5xfW7HlJLCsN22kFCTIaQwCbpz10Dz7cgC
Cuu/KPMZYS3YJoOOlD8UF0e2tsWDAxaDoEDE7oyoInq6B4C2hXfFPPlDpx+yaILYfNUIR03dyVRs
YA0z4974kcZMI/EHTBZ8Iw/YL/KXt2DYu2KA7pGySxXigqDfwwDPu41cPTaurUtJ1yLR1zxBqM5Z
JctSVdge8UtPanzHEi3GylYG2beZiyqoR2OT6o2dukbBZZ7Y09uJwTucrMEdtdtRay6K3E7GWKpt
YVQUZmuCh6uCKolXc8e+z0KZB+jxlOTBWjdCVcOECp8VwkpmmBU80WAQeVZfTnN9Ip+ux/7EQu+Z
3kAlhecC0GQNNgtRQnaSAz0tgOixXPw//zLJ4dnx2SgGDIfwmW9kIH+fhaoAmJEujEYMLoHCT+VP
e9GnF1O3TcvDRd8lNio6bldpfueIlplhBDGfCEA5hR4ESwL1JoKh6wOUD1L127u459h3PCH/fbEi
CrRjU2dOxwcuqyDw4EdFar+HRcDCgDS+PrgCoCPPrudxw8CpleYamoKjBwS5yZ98DrW5/l9WGjog
FRtEZx7iEp/ltVUDnQmZD/kgeq9mdLXtm8gFi7ePmCs1zwrxwxgiK55G3Q912Su6PBynOA8xjRxs
iB9sZ2m18ul5vJp6Z505RPAJqwkIk0CfepDI3K0Kbv3grpGe6DQ1OFObjffK24jAG9PgkdOxftJm
Efu2V7UlD5w7PIno1fv1Y7ONXHqzjwBlLnaTajFwVyo/H2sYMxx84CjpgPaB2RULnmoXWMXIc5mF
7KpUs0hUeT89uR8arguQ4V5K4XJ5wOVH8zfYg94HUlMOtKxpJOiIJavj3kdWRmDE/Ov3aagzERvf
SuzhFkgCAOnaDOZM2pWGHNRbSL2HZ/nk2hyLfoyMJRtjQz8feRjUWFhaAulxV4NACCcYzNUkBFkt
ZdZufAzsbKbnUnBh0Pjlk1cAX3A9P6FJuGG0BsV0WCuZN/lzIrIbPJxrlDY+GjVRSVKLXh/X3GXo
OY6Vnw8VSoIA+N+rX7oAXjjUtb3Tt/dUqyuhAIFUyoNTYYUMwgfqYhFV1sgDbsqZBO35jUWxxO6p
fUNnAiYGRa8zEV2b+ahOen2fgNMmZXJAcDb9G5pU9b46gee806luo+bKcb84Y+SC6C455YzY1klA
PTu/9FozJWzzNCiOEAqrVHw5J4Ely4dJX5eWkozwTgQLH0FqTD1KdcZ2nFUTaPVGSGy5qCTSTHWf
PwvPM0z+aX71qq3hdWTsMGFyIfefbFN3pJdhXnOTS59S6Z+5lUPBO0ihJxSyW8R6MIuQIRQonbaD
c7+gNaNthPDZG2n5nYD/1RoLz9lnwp0np249zgfRGHj2X6GDWefL4xihiYzKqx2rZ2zgFTcjtyXu
KSL9dcMQabxfkGqNFLLAv3IzeuMyK51I3fnV/f0KFctCT/xa5nxrjX0mii+U8/xWyF1iSuAp+N6x
knx6NzgNHChARPAGGQ9ovWaFtDckYJXAb/PC3CnW6k5J4Xpp0WgyCW38CZ/JF+Fwtm5jhYe5RwYY
TtDOC7XmHdRM8/4WCdehYOm2m66IeXcjrRmG2r0uvepdw+3pWm1fV0+YbzfaHlmj/fvd5uBrOuU5
QFFTEaVTrDMzlh6NujK8o+xdZ8hFxhwPEL3OgmKtYglQoeH4bZ6Rc7vVWBP7lo0RXktWp/8+brM8
JP89XguGQ5tzd4cPu6p8JDQ4B+7T1OKo84tQBT13GHkHy9M/7WPcG59d3MrE8TT+SWehMU8tLidn
wInev+lrykSTW0rW7Y0UfAbPTmei96CjOJ0KThlpw+43L3OQIA9zVg+CT4lF7bwaVHmOQfsSVSNb
1KMEfhYlvE12gq9Dv7IpXEnfDij6mrAV+TlW38cKv1RbVEgzITWJaS61RyvoY275tjlCeqDioyeh
jJIxXF4BjA0BhXJ8ekolrOsI1QmICcxEJcJP5WjogObKSquimyON+6WXu/t2Ht9Ujeh5EShVIdfq
Dj0wrWu+rD/9JC3Xgang3pBdEatlEen0SdlZlHq9b+vVRUrxPShBJNy7j+pNXvUEsvGW/XrfnfDC
+996XIHfXQiSjV3vuNEXSw4qb33Pg0stlq5/HbQu7IBzRqoYNaXbQx+9zp7EnClm/XjVOWkUSY+c
ZpmAUd8H4NZHME5HHKU+pjQlxZNtKgBJrdN/k9oiF+uL5CP6RvQ9ppNJSMGZOVqsJbJgpWDZtC2h
eMirjBmq9d/ypsBIsrszNyr8F5uPXrK8AY3hzbjbTxFHyeOzhQixPj8g413cbQdIueXNRB84yR4W
VBinnA/XU+ZUOQgrp/qFh1ZSMEalnYfT+0Lwc5wbFT1Z6CLBo4Wajl+/tz0wCClWFmsx6XhvSYB4
I/LzNBXgizkcTxjHei2wUPDElhawwddmjyXOU3SWE7ColB7rat9MmgXljB06QO7O0qN9y2NycNfH
z/OxGmVeF0lDhaM4yw+ShpdX1xnaSNYP2KyPWcOeybTvkf1+t2j1kVu8FLu837ZwZPppY5IDWPQD
GViyTnO1D16rt9rHVNFSn1CM9CCW6vZYjCDzpGKf6hHLHhII/fwGOnMxG3dYeenwdih1bkX+9i+I
COpGii14Yf/XIBRl3DzGvnnAoWIVzHlgSB+cXiulFEYHcA6g2BiV0JXHCit52ZPala3EkarIAxV4
KhkCjz/4hcdU/Vx5SsaLi8MWJLkqm+EQ0DQwX7aJJO3d5w6AEMEmpIV9VoxdIM17tyeHmoqt0HFj
iV2b3NO0hRRkv7qRkZJq4woGWN1Swu65/9O+aw5Tyzi8GC+TnDasoJzjA0Ni/gLbjKQImJ9ourDQ
at7m68ZVPqEHbiPAXRi0Lzib1+fCXlri1rED1GiJGtA/kVvaf4tfxnWMgjy+8gJaYKp4iuqcSVM1
KBlii+844SoVEf8ulEJ7R7boCt0BmLQ7eKJi39sBOejcgrDFqzT016l2yyFHtmRkfjPO6zskK1uk
5H3MYrsMtcspgokXtCEHKxSrDCBuKj5655J7NHfw1TJf9LL5vm3rCAPSm7ib4K0z+VprHPrrTCAK
ylpoxvqTUaX5RU4wYDmjJk+as5kdSzC37qRNOFFib7Y7sA8UfO3uhqsX+8xnKb2h5Jc/zz8KA5Xo
BnahNJGe9R7HEbfQKsQEYm1YfLBo7cyxMVfl/LSUEaqZFk0tODk7Z7ylfQvRayDxuvxJi6AJkgjc
U1hlahwMH7XM72ouGnyisHXJc+HalWfqojwKT3uAMXH6L33chTGOp6I7FD49pYKgXPaZ4r+/bJFm
71s8dwyOqU0C7rXG5j8KUNzWBZtpNBJujFf3FzSrWG+uHzMQjxhzMMwYcN7OYdN60stZiduq2UQs
U1wnCKqG27GEveFT+t+x7HKQtgn15gg6vte1KxW+e2tQ0LPFl6My3ErJ0kuA87Tc4whFrNDkAAg/
+l1dSWpglK4PgcaQRRKx0Ie7gDM7ILzoLSRZxTO3BpFS0HQluwFQ0/a5nwEphnai9LbI+ZXpm2K6
WCtHuHzJltKTg1Vh/u7ZTdFvc2b2peUfsbqRQ6PPryGq/HKoDE2UV9Ymgt9H57BYR3C4K2Fp5COX
OV4IIBV+S5hfqLo0qWu9YYbnEahZCeHHTaD6kPFNToeRhLfvzmIGIX6jLxtGZjYvzhEbEYjMA4AC
K+7CNFFsnZhqkgGk3G/D/ApsRGiGHFOOs3L6WOW9pjGOsw1jRTmdQDa32zMKbQ/p04Mf24sKectB
ZtEayGCpSfpyUlmRMr93yZIFvIg+vl+0wUtOD6qtos3mARr/oR2l1P8FK2W0GxdNWSVQlNSSWfov
QiAzzJGSH/smr1BRApKONw6jBylQGaBim2RdzlMhmfImDDgZ9uFbp/jRqeMcno7Use0uHNj4vpra
mrq5gUTsi1YH1r6kxAcIxRRyMS3IaBcAfSc41mJ6xugy+3Z58XjBUqji97LvvlDTx27vm0wwTJf5
qOeJHu+nctyQDPEYmo4/0lZzk2L8TY759dmSDrInwkVwawFjmotzQ7bcVwmcMNHMM9vEiz2zydlo
vYG1VVzoJYxTjvFiLREhGycNxKVCwBadIW1NRQcjYytcQvcguQuVoXqgnG9toAMYoABPEKrx0F5j
fhg76igeudc38XLPra1gzjDWY2fZIlaAymxbTfPiIrV6B3IhvJGYijcIy9CCYMa1D6RjLtCFX9mw
57YQAHGW7ZpAy1A6ENbrlUY0Z3s2dwKvUnRF0avuItrKsUcRPgCSbwe5KEjzS4xOSOTf3rn0kduu
qOBtBnxH8gQ/CYETKJ8oONLtOKpi5ZARA7cBBeOOT5D6sMUPCeYrsRWzuIbLIJ1V0offq9UgbOSD
IlnzhBJvGZsHjatSlakesQHdjRM4qN7/U0cF1vth2ulN7HNMP9hISgXvVSNrVRxG+800cYwhdrlO
1sUC9eLhplWQKq+gh9hIhD8zgfdAJyRUK4wh4Gb0KhpU7Dibcf1QzXfOPtGlsuV8Mk+26porUyNO
ATfLW1a4Qm7m3DPxDk9QOqe23RWIW9AcYKhFYnstQwhikrNXCNYeTYN7C/G4+3dWVaH4fQhxGcgP
PQeK/AAlj0xOGlxHu+ZkqCX3IeAsr5f4Yk+yiIHOMfxmAIQQFmow3i8pHA3Gk5FZq5+yRZ0RuBlT
BlqqJfc3d+E1YgEz+8qBJB1tkKr/JsEBpp0XbyReiXxNR8Mig3jeQCCugSEs7l7B65v8//ztmHhG
zzL6lXzzafiDSxinkSq2lVe91N2/6aU8kKZ/DneSh4E8AS9juXimW0NdquF7YsAX0NoOrIDYFClQ
1WDfNcv9y4t1GP/QWU2F9OCvSbhYV7fPpGn5cLw1k7cT13QM7ZpK1j/v4ljDvzO8YuAJBc5wccVC
eV/fb5Zm7XDcS6dpVxg7ce/Y4v8FTfcQB7f/XqViUUfMqL4Ix68NauzjDxF1WffWwq6lO5KgSJAH
P/nXzBpb+v1wsg6nQtvkesxJUv+2D7Bp3/yZoZxY3p6katad1qavAoQPcAu8HOgmkCcxIwQeDzl5
isbncugKnIGoqwLajWOA1xiZTON2+ZF46kchNuo+f5Yg0OX9jmD9m4m7n26jE4X8i80nWif0pKFE
ZuHxCpqh0cddsVkWKB0O5slzm+pjKrEuAoBfdPyDc2EhZIR1eteStw+TxsYNDrP/gs0Xo7qDdXXI
LGh8yuezM655VCU1Icb20P6rE55yhrDziV3gBr9f0dlSPUhcMXRACPK5gNYOUJMBegsgfC1oiIEC
M/3U6rb14vBatS+Nf3pBmNDTIZ3gkOIXS9c+VbCHNJTbbto36XnWFYoq1Q7BUSDumr1A9OaC/5P6
BRJu/jq2zYs1WAKH5zTgNcZGCSzA3Ubcjo+B3iAC29vFQFw70Yot3Pn9hJdNitPjMyM3qUKRNwhN
1QQthky4RC3XaPbfhfEnXbuVK5PA5/SXw94rdv2/RvxuG9weGgomldAzGmP6HN4KeN1AmJh1NItL
HoLmzeIcn1yXVhRwCdnUpc+6EoO4RPYk3XijFFkHdOyZu2uv9OC8Jbd8X4TY5s8zoT0QlQQVfK0a
TbNY4XRqk/DcQPMGqoqmtw//T2Dx/CL/TL6APZS1+HSnKA7ExQYRySOqpcFhP9IQboKy6t5xcndg
g0o0jcS/CrLRQOElS0KbO5SO52QaYqJV1xyNpZocsG2ocxYCTSzpub/wpMYVg941czp1EedpEQmJ
GTPit/ctjDfWT/v1ILueKGNxs/mU3hbAOFDnN2EKcaedFCRXPl/EZU4UvLsfXMChqFSCuij5gSt3
FqrHRIeMzKqu/GaAwfjUm6yAQS2XynUzQrBJ8aomidmfuCDm0Gf/L2NxwZoiAfC+l2/z1sWAlXov
VwYX5c14b0Porh8Uf/gHIena/GHN9vRqpuewRniegwDdMbJiSKRp6SXip6Y003C/4wpVEFNjAmw9
31jtsoYCWhfZqx3e1TIk8+AsyaEJqI6i+3S11OTxJRRXMoUKtT92ZOYlXRsbuc9D5Thp66MGxLWx
KFYnmgCzt3BsHdQQMSk1Q1cDcrF6jOpqYjvde8wDXC2wWBua/xS4zwVicX3mLapfNk343t8BKdZk
E8btDo3XLcnm/82ZmcyN1HcdfBAImA1C9rxZtstCjv31NoAWo5sxmVuanadk+IodABqVOm8qgLPg
Fx3r/Y/DXhYYsG5ERpClk/OAJBQbwuGmYwlEZzi+CewdpELAw6UfWOW5u1EITSGRGuLHj8wuwV9z
EA22Al9yc93nzkCeB58vry0wrUauRzzi75+HiTidOb1GAyW0IFJNVgicWHVYAsQEgbOjrp/D7BS1
R040jU++FqKXBHoGGYspcaTp0Cdiq31H0u1mbu7dVr5iBQS6+sfw6Soy3/8lWBMrZOrdvFFEBYQK
K8qOj57bh+UfWG27CBWu25iQnbmM4vHX+k02cNCbJhe/G0Fgm8tQGa+rRpVWgHgEyEbNeeTOxh0e
zXFRDRlzapyPY74xHeF/PQRnPoTijnRLQj1b4B8dwv5E2GXEk93VoGONsCkSK2hdlzF6MsWSm5MQ
deXOPRaddWtPrKEKBV/PkU3YGuhwu9GMZ46Aa0N/LFjGNYlSbH1texoXRqxeCsrtEaSnf5TvKxfN
AWcUQGbsLM+lwqFBROzidL3H/F9RL6+/G3w+FisL0BTpreelaIigkvlFgqQifFIdImxzqk2JROqZ
AXCtxFBqQrzDqegF44DNDbLGjG6fFl44YvL+PcgbuPvfSsUd9O+FXDgmXsr9AT6NI487kWVaklhi
SjBdg6SIYjt9gi441IOwoWupQLn0T0oeXyk5eY39Y5BNCdt9+Pv2tuQx1JsERiRT0NETKFN8UzvK
iUbPYNyg7MM2/ZcAVKbMbzdoXN6Lw28Eu6Dyj41rViKKq/pi1tlFYhxUPcMm4qHDEmNDh9MorBCK
nvIVceau/Q8mMnERWz8BZgMOOPj1TyR3b2c5mkARZGOB5QJaz0R4opGBdpmzB8fG39Hm7zKlMtCH
1pFN5soKJchF1LKEOQsgONjQnR8Am6jBLmWl2/6VvVRlytvia6phh2rA9x/T/gSVZFJK8ICpvmOk
X2ODGd/jvZbeAfWarCVUh679PG+lX1jbZz0WTnq0F75/D33c9iHHISTMARrN1FqV22LHK8KX4a9z
uDUxPfd2Ain3WcedkBtl/ulsZgmJO0zzE/2x2zusH+RtO2to55rPi1i/lpgyoxD9iF9LhcrhxtT2
WChytgQzLeWqTwwvwe7Xpvy2ZTm29BxjmJ5Tb6fRQLJoOiJfwwTSuwbSyqsrKUvQS6uQdZnmrpui
ZHDGY+9uKFV60fcCIV297SvjgBzr/LbQOCWAX/AuCUHgNJmm/jyYDb7zpnuDCgxAvoIbTdeZ5nvy
Bk1Tn7RWs0hfnbJDzMyVjeY1ZdmWL7ZQEopiM9LdmMPZC8pEBPLJMUwNERjv4iNhvAVOmfgeSdkR
d61NPFEPKViBTe4k0IK7TfEMmC1R+4eReZeIL/pnbD1lfw+TelDfXOxDNAt4Mw9qs3t22N3yqYUj
jtcJpRhcRxbs8VNavPPJq3x0BIQimKgItwXWVAWUWgazlTIYhrW0IJFTZmIABDCpfFDn+AU9Y18A
K7OUgurKRVUBJ7mZlaQPnGlAz4W6Lo+/JcZioUSh2LTbuip+0zCeFWaU7yHLZrP64gqgJYBzMY5r
YLaxmNRPZkAN6WaYDDkcpjIH4yBPgAJA12InbSsXeT9gxWhqfNBmTg1HSB3k3G8rdstbDK7duptf
wNXxARbZYH565fA0uV9wWhoNNfpazpd/Dqp/Y5surOGGX6Bih9T0hNTNOP2TfOLWKqZnlCkUpSGs
59HkIi6mOX5i1w+n7Tlct6G2MNvsuYiIsNMFHA89mKncBrU1dC13kfUWc82o+l6l5GbGvspQGFEY
e8RtUXiBExMV+cFe06a7iXnThAkh1vJNtj8NO0nXjU42uRo4kxs20tSPHj/Tg/ks1pro3zD1mZiR
a1V7418Y4VuCZfNu/HrIIiGnTcYk+4/LiNaJVr4Yk7xzyWwmO4LIbWIQ2dMAuBzc4tzwgSobuWtr
sXoFG4sTmdhnxlHzyyhY+AFldzbmg3ykefL30Yk0Ly1FlOCweOaPvc1wJ/D2T3nqG+IWId6Ch0xq
lAkz2h5e78Lp84JwLnDbAuz748bLBWayU5q6OCRa6rKN7Ss5CrsPgWkRxCRjdNU++J9V6K/rfwSe
ly+3DQhtLiqKQqdeBnAIqX2/y0aMMhjVn8j9xJOMGz/2o9RTrWOcdTUgqytv+mkykkwPeAqRY4UW
ydqPNYL7YsH2wNpS3H+fo2jXFWiZtbmX94et8UKERwSpIlhUgPYVtdQJ4sTFtNboOiIgkcJOAMPF
yn1iKuXcm+mQFZPVRGcBscdtPgFUMI3mPviw8Ec3kofaf8cfTAGdVvVV3eONFYOGxIKFjJvzPrb7
BPvdTqhnIT1kpCZzJdRZ0s2n6z2URApFqiwxAKFz5I//PL27cp9nXAV6sh/KoTInL1qgw86CMv/0
WpLV7/3pQZtb7aLgfHt1VsyLGJ0zVDl9d7g2S60UjDbW25Wc4TMSVhqSUVtJqyYBCDVwXiPH2M4r
bC9td7b5gboMiTEREBkf74tnoExQde/1oc5WsG78FPNSSkCTVPe2vf+EWYu7D1bW0wXdJDmGgnVO
rgeAOnMEhCKCfvFAUWgAUywAX+6YMf4+J2/3nW1TLULi3/ikxeWefMF9C4TOoi8Cz7xG3FPbhJkE
GPLMVSBBkG8x4KU/BBRa+rqEY2bD5WLvBFIqt/NXEi5h7u5ksJD8G/+8xMMe6c4Mtn10s9QOMUg0
0+HUsjteuiMggeOXNGVxU4oWylWHFIpSwt/pHkovKDmofnba+rMjiV54E3rer/tBRi2FfERy/VG/
S02xXIDnxhWyRXg1My4W/sHfiTTRAt8XnihuSsFeO3Cle/GvDZMlM1+vEH6IAUecXmC73nQ/pqQp
YD+bA7HF4HLRAfTncAMrpCvHFmISv9B4rbSFOq64je8v9FXHqrj0/XG4v6WihTuRQDfZ4DP9NQ8M
BUKQYBBOry4PypYMq9pvtjpTM3Qg3HJkinfF5knJ2Dv69B3sw5SGxMYqtmQb8gc7GnCEDIorH+qb
JkrA+dDcZeFWnXltTLn9cpiRu7/ThDHapMgDVm9FhpLQzLK5U97/PQo5v2lB+30p6q4PNjuNG4ob
yzWal311DQzLzIYJEV0FRMcabd7kJW403bJiW2G8j17erdUEAv2XCpwDvl7B2nsF6/AQr5P+6xet
tSUTruRECyBxHghEFyb7brxLYkBGRvt9cSYUcMp6DtrRfbTFCpc8t9a1vjappxOAMo3IPwtdaNLN
+gvBYvphQ+Rsas2BSlizmfj+H62tVmRCCiEIKaMCRmrjKsh3HO44LhFiOCCvKBhUlTR9H9DvZzHK
mnHCPzVUOpdR44FY5OscEf1Vs76fuQXt+a7JeJR7uNGu8RKyZMXBPPQQ1Vt38vUS9af9L4t4w78M
jKw94Xt8h8RjU6XPvQcBswCU6EASZ/YnRUV5yx6VFIrh+TBQHy6Vj4gcmEvEl8aJ2toosiv5D1vL
jTlngoucGwqSR3Y1sTOqGfhkwndJNWxZ32m+45QQP+Q1DsxhCISpqfiBvHDptgP3KNErY7eWhKsc
Wzc6lmStFSVV8Zc351ov/DgHnGITjFc7UXgTQf21aRYdEBtBl+Z70SfLlNA+klOLm9vJW/CnkzJs
sA7xEYa5ZKTCigejCfdpYz7V9GCQTRezZGjClqej/8WtCXqfbWmVGvZAtrsOpLtuCyl6lDB+xoaA
Gkvp12ZEoCAb+vfKKPpkQn8hr4SdN6RQW1U0r0h2nf0PWYVdF9CF4aINAQUj6Wee0XVmkm2MbYik
bMY1DoDnBmEnl4dIwaUjS1wa4QsFVI5km2aouvH+ptdVs10GUVEdkxX31gPSjaQW3DZSV2NpD331
FAR/Vx00096jsq6Kpbc6E/o+T0sWax0THCd2l4eruw9rPYssz0wglNDT+uW+2UzLWDIA3Zke+CgE
NW26MikE05tuhcD29Jvv8+WBfZfbewL3JLJSx5Z1AzOxDO3MZrhmx2sFbTh4HniUgbZGk+/m+GT0
SfQgyyZYsQ85t+RBezK8qFUtgtBTjvVV+8DuH6GE7tvaJu26R1tbHQ2wvIgkgnUvdsL3fYQfL2Q9
lu3233l6yHQLiH74+OaLgD7eot/cCJobMTBD40O8fwtYIxY4IeDFhFIVYokLaFevEgvzoqeBvxdc
YyS6fEUzgwPjHgtT12Je+BVoou22R4MLYhcB8Qqo5MWsdBAilBGgxJ0MNRsoJvn32tXlqUOAHos6
y13YmhAei60or79voUjW8LvuoLXxgQRn6kgvfBEbajbRZHeqrsJt7IOs2rasSGT5Jzd6q7LhhcgN
pdchhTuXq69ZLpJVXTRtaw/liziMSbmZqgMLVI6YhqHfl5xtG0t6hiXVr0Aev0q16H3tYPUHTAbe
2Issqw7GNOCJ5RH748Plof0bmc9lU9pLsHC+OSBgUgTIZuZakrZ4dDWekGZNE/VZ+XdK+RtxUUMv
XcvFmitxZVAZoDbHJplvJWmenpqfu9apvm8cJd68JmUp5JO+iNQu+hJmi7vZnuqvr8MUsFowr7fh
fyEL6H8mDaFYTG4dy43l8+DX1R2/fJNd06DRACF9g8mt8n9qJskn+U6QypDAzK1vWvwckMPmwGPh
o2qUS5l9ZNYbftIWkFIvtNPWdvIecAUikIh3DL1aVN5XiOEdc68D7ypECC1/h6D+VZpG6wN1PnqB
vJOygoGtISUnvwA2nxPBKheQLKCLxKbzCYxxQC1NcgRv0bK1yTOdsHpektqYZq/8YR5mIFzyUDB6
k+XcXpIuJb1fohQVzFUyeQhJnIKoEzm1dNomX3yv3niBR8hqGDzG7O4wL9ktAK4Z2ZCwExQeci40
uB9ZSX8wnLixALAxl78a/4tyAwr5eY4BIzuPL5pUxYPyZyp/K/eND27iSfb9E91IkYH5osMHmRIk
XRpCOj/TwMUS+e/98ziPTiunc8ec7LhV7neSYcMqOfbahMfvY7hW70MR7e3aahQt6hKkgtPjhV5Z
aw0rydIq0sm+/E+o63DEHZybKRFPjPtoMKRC4SjY7kGfNgpH+6xfWk1Hm/8XpQSf0anwlP1AIMaH
FL6QA4LyCJELc1O/k+YpP0jImiiFDw+1z/IyVn5JvYZNOcuIKO4vSQ48IJgwdFELHu3/kCpk6tfQ
Sq+chMSp5pEkZbb3D5+cL37mzXvUt0QthbM2ylguy9w0b4cI56i/x2lvwK+JTAwqfckNuP8fGzWf
5kuxe4Yjld6GOXkU1ZMpio4kS7It60dDQVACSGDcCRGvLZNHgECTX0FhptXE0BzEOqw90dfsgD3g
SgW6P1WftarDZ9OPflfCneW2hFa+WqLborf4jcEDSTEfHPwuxXpNRliJZpZj4+8EAt1/3IIL4LwM
1mynvFGV1gzio00bm4/4OyBO/liMuh+pfVw/dFj9OWgDlKhVLGOCsKI0wYuf+lZohi7yUnLwaf+g
lILTfg6qb3f9MTvo2Hu9OkVFQYK1LczWS+QnYLckbF1D8O0qz+tF/FZaiykdGR7yPZGwmBtH34AT
NiKaU9I/SXXExXFDJs9kj5jhNTjGKJyPnSwq/ZjonVKWfW3PZzCoKCR5D6CpASlgQauN3r2zBPJ+
/geoi9XSFF0rHMZFahjYSoV6Gdqs5DWUZ28OQQ3GB1NQpRxbwNa4s4i5v167TpOB30eO/n0blOGG
lZ0ilPnw/65R2pHoiq51ABhp+dU1JdOV3o0iQXj70ufBsjfF5CnTK38oO7AtExmxjwjdYzAxgbnA
IHHIUale90BVZYipZYmKaqSzYhB7Uan3sqNSF5tQKR/81HA8xifyzQ7XLJhwVmtp76rLTkpRx9Ub
u+qbKwrEUpE9Ejxo7FAaP+tuii/Xet6IylmnIIMKoBZMpcWMj2ZLSLyKVS/Q97cchL1DIQFe58pS
GiATcd/GxTXyZravs35UHuPq69majrlvkMA+oTdg43sEHRGPoLTYcOXj7vaUAvjG8faNAUQ6yvny
W1uRhmNvYLwR2dI2J6/aP3kaH2AB0+BZcZTdKczDZkWIVGnTnRPInZEWayhVsHlF+E71u9y9ncYc
Z+mn5Zg86xS64hDHsHD99edBGGOljmfKeS/vwp2hTckpC96Hk3oqYBsLT9sqP0SocQ/BPkDUDBx4
jlSpzt9cgqlPRTrvm8AGnocy2T0Ss8vBMDYT9iRuQkFNrvSW4/2/4ImYLo5AQWEIRDTc+jxqCwzQ
KmXFM2iahMbMVRuaAkFOv91DKX58FhZLKnXtENaMvOl6PbXT1r1+tou2u43A47SCayI5xpdqUcGY
RH4ssmz8U8gaXXbXRFna3UVvQVIXMdOKlJ+BGq1R+PFUCcOKLODVC366GO9kpMIay9tt62ghFKyd
ZdEaT3YYvjjWhkm/G8QcMDrPoD9M1dkhud3vNfWwCWML84oj1jFgmljoj+IJb50SO/verSRc843+
5jl2eZmmqbejde6G3nqSaiNxt3GCPQ8q4leGHAFY0IQdkRYLP8MQoOPKj4bthfn3FZl7S+butxDH
SWb2+AeBKc55fdcUhh9j9/n+ObtabxMtGxrzhlgnF9IOD5r6Hodl7Xm9K5j6IHWCFalEIIZdkvmB
k6HP0Jeq1qszK3vKy6xtqYm49LPsE6x/QsvP4r4AvXrA7zXFCowCqlgUBHI9fYOxYxItQFRY7lX4
j8ggPDTNWprFs4YPx5p+9LI5xVXrVb/wxFkeW8LbdhrG8SfbBg7lZPxtZG2GbprZvUAPi3MIAh2g
Nv+4AdeWshqafVd7FBm76JRRSTGeajH6OgkJlqiJQBOZWrr/vsBjPzANDyYd/1QaLnrXXMgCXdGH
g55cloHQxRpHyQsvNyNXEiWkIO9uyWVeVzshqv6dR9xMRUhYm6TiJ7xcKN+hZTbADDRYBlwQTYHb
YzfIfeExuFSkpkqFEV4C0hBhp5E8b6/cSx/jvkcQo7SdiIHvcPCXmvvfEns0Ir2PH8O/dFDSvcu4
0iyQCx0s+wHXe3iyqWy/M4p5whSdtxLlO+dyk72CCzFzs0Gd6tx4l7BF9K+XbDetaOBd4koUedDF
/VR1T6J1ARK8f3JuuKI7FfYMjr2PVlJDmCP1kJTMoz0qn+EHAzz5ldCYeVJJQ/o30qfp1w2+MDVI
Vjp20WYAp6oMCKRIYPb2iCcxK516rb0MBvPndvNiSquazckHi0JBzDJgFhykklvAfmjzRu3tiGSY
rRt/Fs8tVEth7h4cKeUp1iA31wNlWwpgOe8fHstm6zJq3jig8uEwI2SYdO1yuFLADL2g9VBn/GyU
fdoHeAW6Ggt5Rq7alE+VGCK/VF/5EAyWTOgJW08P4jX4JwCkcOkxRRaqUXDRo5obZWKC9RwjP17O
TE7UZmbGJsj2TxYMc14wnNu9bW92mpdZXSpg3WXpukb5apXsDBex2gDPc4+Hf3MRxxrNBdw+K0U9
CnPNJL6TiBYsFEnrxj4edIHpGt4Pn++9QIPcU/JFJqsqYDXayvtRDnsqIcksATNAVpvlIrPmH+og
Kok2+/fH0BJXf105inRNhgxubdaJQVTw0AmIHulXUivUqIgnJs9QdIlmakismViPlgmW4HTeHcC7
8MdqD7RcXqbLZhXeGWa7Y7vo6pPuSrNvQ8+ATA5du5nktJav9iDDktCJ9gLbJqssRu2weFrgFRAu
l1f5Kq+/ZEaq1tu7h/G9QWpaG0g0wvNJCeHVWCLIwgGTL0w6DMUjoQMoUjuqNcYLWjSNE0uT3KX6
RfCOdwv5ytoQuZ/EZ9Xglu9C+naycDwo3E+FuayrHwsyrIu21jIOjrvjocuilFji70/7UpjgzONB
NikHNa6nnGfRW/yP6xzEbrlMHXs9K7t0vqGlGDDAwazPIdnkk18RcQYNnf+RFxeioBVtiNpIEJVP
8Ju9bQ7/T65bpKdi2hqfM/8iW+Lg8doSizhbWQ3DWXvkKEGxcSAd2bU4iWnu52fsBWRjiAyLHtX6
HylE7fiImGruazsJdE8T8hzisK7s8WreKUMc7k44eulPe8UYfnzf0QhzKFvPhBqmch33IAKC9lo4
3cnLRm9fGt02mkraLDrBZsYu1423FO7lW6T2MaNOI1dQoUA4bTTq3Z9HkcYP6Rb4bGhF+IkwvaUQ
mfcgvHtOGVs84qDQWgQZTwM3LvexedV4VKVoLHtSyA8j/z+TA0zxPqMNd2pO+gl9Vo3bYrFdpc7j
CSxPCJYdlD3qHsUEi3J6sfy40+aFCOQqb/hJpOvgGNEWbBOwSBVrnwMAg4D5yQQiNmmwHu8rTgpX
t4eC6iMJ9kAkn0R8j16zyVv0J3Y/TwwTWg6zY8ApAg5prREdXhYcjI6RyREgM3SvBElMzWTbWJGj
KvczU9I2YcXPVDGBdAOX7S1B0sAcBzFNiZ45vQiZ6uH03rpROL+xXAKNmdF0DEvfQWSfDs3H6Laz
4PloPuxiCc0f9MhzYPilr5niu0BjSOELeolBINHjSnvrqGiv6orjmzGwnDJbRtiYos6AtkvmXQMA
FRvBbfI5NPJ4B4eP4H96FTzfRSn5oOf0aU5ukh6pRVhEARSq8ezzbFHMJB4Aae48GFqLM2K+c1vu
59knD0kA85n7bmRayKqMZ8+9lI/XFRwf3wchn/9slS8cMiIo12g752DmUq55ywYciDU1tgWEb2mk
bZiP20xEBeBvaZg3JRSLJKCY4itKchhzRUiewT+Omf9enhlQyLyXFg6iztj10j1YVFDFgWWsohZ7
/9TwusVsrIkRI7ifc/RBNza34mlUap1d3FpUvJ0LYiSxmFxaWUoujHBj8CjazD1/xIstMf11G8OW
L0eMOPSzHeiDKXHcJIyDWmcbV63q8ImBHyNt0XgSTpNQAZy/DsWPJeCDKixJliHkjQ3mYg3knyPK
UwiybQvDAP5bRb+Sb4WgBESlGwSma3pSAqqxa3bPVq6tKSvmiI66J/nglpNrImvjCnHtaGzJpS8Y
Ng560B6pJpb9ujjJVY+jSKfYRJseRvjw9YI9csUjl5jm97tAB50Tf/Q8pmNMdp0Mut5KEbYMMN3O
Kb+OAqkd+nfZEK4314dhJOH1ZM9zyuXZfk3oIl59tp/trLHjX8HIEtP98w1GNNuQ0rDdFFHs6Msv
sshU0V3jlZkfxvugpVYSXPlFylWwT0nK1GIKtfErXVV/jYoTrH5+lQPMql+Zl8pG1uWVFvUx3Yf0
B9A4ezo7cNf8sLcGtBaHzmXY4LHRu4uiDTBJSu7eHsxj0XQFHAaRTj61Rom6p+0JSpVgr3DjDT3m
FwdNwcCeTVLM+b8JqJWlx643mAJapaDjjk7gyckW/hzsezzNrIZIvjZzF3oePZfp16Y6rIQS1+Nu
6bgDTlj7YVbvAL/OH8p1F/Dc63O9BuJraapefY83MGW+Pb04x4zQO6Yl3aL95WZycksXKJWq9+5v
cn1Nm/svIAxHvPoOS8WPjPLSrk6KeU2JXgntbkL3xhOAaKNNCgaXl7h65p/bEPMyhy5kp9/Wo12x
QYMj25yGJ9dK6yAzrySh87LzdSj5fGsKcd/QkYJ9J/a/gJW9cuhb3SGP+8tHqVMqkctEAT8oi7VY
Xvy32fztj2YA4hU9OG1rq1dXrp+twBQkYUJ+Dn2F4SLc91OXVZ3HWqJQ6SFhywoPhfaroanCYjyL
SfnkoY1l9ljxtIOFdW51SCwOnWMhsPJW7V0hZUZLMRacmbTY1XiAycNoV+plAwv5RMMrXJQQsGGq
sL8VAdiTvVz25Uc/JPF7X/O2JMCEKf5bMhy8cfOAFXDsu9ybmvXTs7S5YnNEZVjJTiwH96eWLxFn
OfYKa52z/LjEcbfWoc64R1168SGp1f6XbcdYeY27sDOawcHydzzkBhB78sYhk09H1W1qkGfMIL2E
smHTBg/t5NJit8YTp+qGiCSvmsEoKckOcFmWDc6UcMxDlSXaELGMp870VVD0T2E27xftsp+VTMbD
U9lSAuAjs1oBoJJd5KxJQFkhEaHnYPiqvJ7086t9qgX9kKu8FfE4POnqxufw+5Rei8wk+wZkUfER
4AN47ERxC/ZO+2ECc6v3PhxlVYy1UwhusVQFwxx/gp6pUzcppb2vMu6HR4Dzqx2BZygigkXn9iY8
PoUDK4gGaLuHrKQJFxBsFbKd+ymAMwWohhrIPfRYmYtHhNl87msy2AmdPKjIZpjb41ZmjFvBrVcw
/Ah/+lqEx/uNJk9rHYaaDujE7DglzK9iZDf3JvRQPK36EqEs2+F/WK3g85SZxtcVCF9BnUD2vhZE
wIUqtAjScydMfaHqQ59EzqZsaKl8GstQfjjqa67hlEg/XkXLNJzDcgM/bIUHV65eogRynrZPjrBq
B7YumGfUuIAT8rdvDDaSqSOSnDuBtLiTxzIojasF90/9d2ahSdFzBW4EI9U+9bFCyhWJIA3V20Dn
1khg51EWGxFsDcZKChGnmlTKeeDdE9rJVOfj16OgIMFvZvM25yYwcu5sIjcKl2q8xRSgQiMrtJZf
WBlE85PpY1BgBT1V0xe/wsl6X8kYd5FWqfhc/a2/e8Y0t8upbIHqd6iBJX2w2qQSq2dPiuDz7PqF
AMJd9AQbn1GMbbApFrlqt1zsD7CZyOWJlCpsgQIrk44jOO6iRnNA4oi8/Kr+oz7dRJIf9enF3Wbw
n/zoMDvDE8cYl6JxRmW7HMNXUu8DBTBHQ+rJwMrEB+nbKfQgAyOwLFpQ//38ybE7Rks/VP3R3Uoe
lGMCLya5RbA4AQju8rkd9NNSF1Gb0IdJNwiYKLLwwkPtdag51gsCe/SElADGZNNru53PWe2tXZ0O
ODs0ORBhXJalCFZZDkX5xiCyUzPpqoQZuHp6eRgM3Wb2K/Hc+sluhq3bjrQTVvQc8+En+oAh/sui
3PS6UDaHNO5dsDFqkwPH5XzsyUEp0Azr1iE4vbxLyWBDwyJK4UlzwTZzmBYIUZKc1mvqjRyrTzGr
Y0wlxf1tDPNsCKCAqKI8uBoi7bSdiA4WEuKOr3zOsAxRhcqI3oGFyZbvbq6JfiCuxrwQNkjXAb+W
tuNcCuGW6ZZ6WMSO/JPO1L4WH/V4O3XfzwrgwMJTWv0Saj6L+6WuouZBrwS6ke7stEJ/07wMWCXA
sEktslRHgR/PXfK5u4qwKGB1is8bwvH6ODy0je03gMSSul1drKL7oH8a7ICcdUT3h2/0rsy+Myon
cqEgVfJqU6U4qYmlNTGk3+6sIxMGJuilfA8bLwZdKGO5vqv+UH4N9ScbryhwdIbbZPrYnCr7MwWi
9KlZHvssXdM3nYwJuACgwtPlGyqEC8KA4pNJ8Qmb8Gyo+9LL1A2z9zsyu/pXiZokQ/MCLRjrsN16
qLefqzQA4dFCNvjZtOrHiGVLeFeqvrTvh5EcrJchqzyjv9OVhUTptnivoXPuWkBtcEcjA6hagIaJ
XvTA8tYnfxCF8g6qOeQ1FlDomHe+ZohzxIOjM7tWmN7J5PmalSLV2y59SiDkkEsfScwcy9Oepuxk
jZT7FTD3MSvsduDzFV7T6RCszpupbEoNNiFy+vXbS2+x0M+g5vBHZFsXI434Dhhov1eZRxt8EJra
+lZHQTw9QHdOVV0qdCe+oFe2P1HLgYHHAdx4PgpJMJJjmAvvXs++yEOCzYZf3pRiIfo2f4mVJ4W2
DJ1RGCA4s1hg0iKteVjMicEypAYddbivYHT7J99R5uBSjEzxSPvjbl3r07oZoBDro+u58Q416S2b
zznh7EcyoEZU/3XObP1ra/FdXn0tw/x92dSF3w6lmnfQ5BxhP82XU0u1d6Tn6gqIB6BNN5y+zySI
YyYLrpdABJcGqxT6ev3DovyB7MSXyQ0TfzjV9oqNRGg81zbOILKqc2LgD8MxolLXvY2iOa3TcQZA
gXi8
`pragma protect end_protected
