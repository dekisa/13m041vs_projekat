// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
VRvhOi2ekKmUNc8RXhSCJbjxue2k/tSboBwd9ll/HCTYQjO18y8vr93LNOb+TDRVFY+ZXT3g5XJE
Sj/dlHho7x3B6fhHRJZNgfNeIhD1McvxEXGn0O1cM2qO3xWkaktmfO2klp6ZcK6SPu88Mofk03QN
8LxHsCOHFDJRHyoLPlyiySH+idmusWy83S5W/Lhyiy1VrDH7Y9j5IA2XViuBKrg9MqJg1VAnn6n4
50g+ABmJbPS+HhZ2IHjXxqGlnGDQJLLKL9cO6ThEzMOHYrg89tQZeTtSoof1hZylKW3ZM2SmtNhn
PqUOmaShQbgYuXh7Alzr2YBpuf/N/+J3wSCMhQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24816)
PJV/Mv5lYeFeQqSLLdxKkbYJejm09zNKWLQQPn8xGYyCoItJaQsKcqt7YHHSt4+sVWZ0bs4vbA27
1QNKTReVDf3Yv/+TdraMpUSBI1ygOo4V37cwJfQOYx4YrHJwcfQ/3QOmTKzvKF+LyFEDEdJ3s2Fj
GX3Jz2QkYOQIAxJsC851ebN8kHIA/YLQACir6ZnXC6Sk4kXD+tY2+r3/6griov1CrCq3wIYjxocI
obnGTeIXwJMRzqJYAY+swoXoVpjLmN1piBM+46S7iGxN6gI09/zdMBPeiwWAa7teE3v/Sws/TWAg
MNXxbzgujMXsdQNJLd/q4WZLH+L1KsQLBavqAZ9B54D1TC2jDC9JWjmL3aXgYwxxPFb8g9bqJZk1
NM6Q9ASRt5vUTqLKZQMo5pHWPcZZ6MBOwNz385wR/j4ZmptIgpxtKkdiCDirUkSUToXZxKE0pv/b
oxPpPTfGADUit2u21KF+o8E7KPWMK7APrRXdG5CfsNkJo5FwOcbOVqvtXfWmiSeJU+aDB5ZMYrEm
tnCAP2Lba9Ek71yKVRu4BQwDcAT0Ipmr1UdOOsBCuvV2+LqgBNOVcnD+PQ0x0ZQRggds5oxIbubD
z7zazMpJRsm2m5XU5mtsufIZQDRCHdowR6VYP30K0tnP3SdpjlOfRLPu5aKHxZ6ZCtl9wMQ1RvO7
Ynr2CnWzEpv3aP4TH3ck8WRh82goguCaVzX90zzNVnpAQvf5nmXDaMyEeNjloeV3ueDkPIXstlbz
+iV8rr7Xc2B58lIUqmFowU1/5lg7+iNI6z+ONmSRn7hcHE8DGregSxhFIZYqyFC0PrCmUyKqPVoe
bZ899veJmxj/ar9cJ+ScARe1v2Gq6jr00O03KP4iad+cgKfIFjYJ7AUUslUoptggFP+6Zif57A96
nfdp/VgsS+lLPQyHN5scSUBolLaGHr1rdn/fgCHneynQQVlpT56seZaQLrGgGLbiMFwviO1OpVjD
essA1ESAfK0VufLlAy5vp/c6bHtdzQklHCULQbznnQppTC0WoGQNidNAze0QuAZjVW6yaXHqWKOD
64awlcJ8SIhC9Knodu0CNhTqmoCqnvv/y0ka6/4K7oAofCPq2dcrnJpaHkzp7h7XRG+TG12KybPR
oKkLu3WNUbaojzRB3yoBQFIaeIu4q7ybqxzVy5LrNF1bdDXJteyR9WoMmJyfXmfBp2Kl0fUNgGzT
lFw93dsPdnGvDsfTRgQTv1VdYpRWNNABuPcNxkOSNjYnFAbdJ4DMsypEMj8tOiBWZcAYRtchw3u6
HO6duvBr5n8vHcSihGQlOdmPJri0ddcSg+ZLMn3UPvgbiJwkWrL/JfHDsK5zpmiFRbgo+sC94G/M
66NuJLHjh3EXGi1uFtH8GeQ4OKRVmOVw6kJF5EHKIRp0c0tY8Qw4Fypv+IU/5DjO+L6sZetL9ImZ
iwNdLYJ4hhbTgw1MgKDGuGhBPOZSyAjK9NvJdb+b5XbAtR7udeimJ62gFVpsSk3Hq6BgeiBHZ2NO
bVQEryAZryKZVw3DeCEFsJ1rF9OJQQuBHtn5B2Nc/EHIT+OEDLfVcen9whlzVF946J03KlqhfNTz
xEzfIzzJPDoiIf0vRHDSSOBkmvnUqF/KCej3VD/4FZ3gafB7O1PkoLZ5yWXW+J0nfgfrdskzVQgr
FwWSOv1QiAKJ34Y1GE2TXByxko4kU6Dw8McAPe1WitQiFabNHYCoQCqKbwywhWTwHuEezoL59Q1R
5LT9HBTVwSuyaMClBn2pAVUsOL3SJFVpsHGv/SBvLVRukJIvJDpVrFiWFpxxAUTmtQ3q59m6AOKT
uZl1jBzwojp1yKOl9lwjEm3tHbJvwbHFzQha2IPFn5uyZq5IBIwunlRyvQdQ+gbXPedlGuBNwcvr
yAHnIr5D4NNd0dXUVW5NUI8j9uPVpLh4eW5d3thkjnv7+24sy8Y83P220F7Gw4of189t1LYPzpoy
6T4N22lOHZ3YgFbuq7wh3l/hcL99evwGKY27ummgwKBdnY70+SckaWpt9kmWhlaRlpWxDEY5S86q
eM5N97hSxL0SiR0ghB1wqaZybMXSjmk70+URQAouXQduGcWUS4xV8IK6cQ5BT/A1YJ/PvA72Azjm
kS7JMquFtEb/U+Tog0ayrZ8KotKMWZOkk4vsLO6iZx93+1RZTbTzDAdAgyqviPe5HTmR3NnGgoWe
67YaSkQRo53xNE1HorgsQWssvpWvZy4vfWmSteIYt/SgzTvImgd5AQF7JYjWKgeDKHD8/UUUHlYH
IMA/9u7+HC4ygOvqYvueJN56y21bc0Z+FQydm1i7q44nRlO2TKOkE42EPWn7GI6cG3J9JaKSW84l
kxbA7HX2CwFuihVYwDgVdd0p4Bm4mpMltJqX5lS4BiIOK6Jx6UqpK4Z1H+QxDz8JJyv3y+93gdE9
sANKa9y7CXIRDnDpRtFU173GvzZ/43eeNEOzvIA7nvRY/YsLiFR7WH66rYx88P8mGjBxx1MZ3zrZ
WuJHIyuk+k0yH027sMWsf30lHKTEpuq9RR/dng2wPG7cpKUbDfXaRBG9mbktgQFCYSxEuehnCAkF
Cmow2D3leiSyfGDOJ8uA8OgY/bPEBfAJxQo4g7WsFh2Ztkv7q9qYSOCGTAoAO5Sb083lQCHXDzd2
W6f9zJuKA1dRlL2AgVkp463Q+6Iq+v8Y8gRa3mNZsWSMSuwaDLNXlQ/E5Pnw9gGUxBgZ6aDb4S+N
2BzF9lQIkEMsAoOEkx7dEoTWp6mSNpXqTGDEuo9Qg45EGnA6ZWoaV9Tgi1Xzt0C4ObUUesXY33C2
njVHiM58Ynv5y/ILMapQ2DO6ite/XzLm4X6Ypvdwvbgrcj6NN1lwRkivnGmgO+XN01Tv5tIVP+Yl
vpjQk8FgM5i+kGfDmLRHFfMEUoHTQKJJXt4YzW4ghspIbAYblHP4gZKEy6u0q6/z6MfZuaSb5FUN
mx5jpdEly4TZ/UALoPRgQLDOJbROIK4p1mr20C2vGGMwvCU7j+C0f8hwAN5TFGgVFWYFw66N5NwQ
uJqySdrn/tVpVLk02qJoU0Nc6XEO06T0OHELtEBd0MNdP8YLSnlLPhWSLUmnwYuHar9gj0yTnqJv
6oozWE0ugmgvyAf0pK2dAGWf5CWoUhMOIeMwBV3252JtSkiqsvpQP3Fgu4cWjnkeuOb2zAxmuxLo
DmuIxOcAodDFoeDfkbHP05x+g78cog414yHP6yjzN6tdn+zx/8jbil44DZk6MOoW6Sr19RXJ+D81
YYNp6G3t2Wz4LIWGDoxUo9hAdN4VkoP8UoVGhwDTtHPWWtB997fRD8pI1QagPAY+FNF+PwkV6HiH
LBzxJef2TVZZHwkfWJJyBhsU45B76Azypr5b1l4tNSFeevgRmIVMZg2GyASx/lCuorZitOlB+jDv
ZUDd/ErZYO+PXhup9EvqPla+xCWrfPcjeNVJjP+PVU6uyJKXUTZHH6LB33oXsPbfMnfQubqwrgzE
2IFu1TBlzp8Tnu2eST5MDjJhV9GEiM30ExGsoicTiFtue6lTSD/r30xlzHPeqIH79OPvsn82SQ/l
GX6e/U7cxFN+qGZAUb2ozm0zsZbBxYy1N/MJ+aoaBrxc2ANHlCj/de1P6bNQpw2mjBIZlwjMojtM
x9Y9xiiuj2wykPl9nrm26m5YP+lblIO6nM9G6rKFGjSLzTHZLSpTI5i91sb+Vr18ymwoA7dg2xvj
7CraUmUxifLsXCrlSrgS5IYSkz8Cv84ny6CbXdxnSWqlJ5pH1oT4SMRnF4zZY3fpIq46qnt+bVMY
Rx5/oU1kJfWtneAAZa6SVWKNGOjoZtr5/Liu5BHiZnRH/uWNiWRte7yh8jhJlR8Wiw4FmJN5ndnl
F8qbXFLCKCu+srsFTBFPf3oHIMDrtKZOb+Q8X6ArFAKiCJ47dsS0w3lOE43g/uZAZWfqw0Phzq52
c+ezzHct9YSNimYd1w1TAKWrkhipw6dwGHub9gvajep59NrTbzmitymr0gYlbTgJ8OdrN7A5MdqD
xONfQVfv9hu4RWgOTyPKc7VWI0VNjc8lUY9VfEKzamoaqEbl0KkKEUoYWP2Ry9ks0P2yvtm0ETxd
6fCgs2lA46OWtoFiemXhvzwrcOU7SfLhc8xXR6Gy3loGYamgqGzngVI7Qg5onegilwWasXpK8nL8
Ox6RqhKFg3KDFZupt6ZgqANOL4mrrhcY6yR7G5XvrPFl4VpAfcFHbt4/l/nBBxcJwDtm8Pbr2BtX
zaRYa3idocyMHNVdYXXYzcr1mXkhuzYvij2hstw0+7iDSZuTpx7fMrDOYkz3yPoa4EWd05BV4kos
TFIHaTNjv+8WM4Thttf/JhhaBxZzT92MtlvTcehInG9ilAx37FthJb/O7xUDdB61GysIL1xuNoxW
oAU36S1wymvQQ4UMJbZXqKbPg/M5aSIzEOQ6l98ZnuitgrBV2Ad3N5QuapoJC0Ju+EnJ0EZKb+a9
1aEQNglVdx6DoSALlM4e0cTMT+tq9ActaybesjXIQ5i8kAunpafTLYrtX9ekRwqdA9s90YJXE7y6
1EAlsZFDjTFcPeSAR2v6pK8DkiXHsmoYGXd14arIrV1Q5osQ2u3w3ebVZmbBdXSvTr+bycSZsK96
JLM3iSzGNC6xYliMCWRBVymXnu/N71rwA6enKnksCyjE2QNSGF/0Z3liQbDawTu3+UBKmU9LLlOb
94wkJGstVJFI6CS6n2Mb40w2dPwHDCqQGncR14AHP4QqbPWDD9j4toiAHnEnf7FCk1EmYjTnobfm
go27Riz7JKXSB2uFU9oRDr2a+NKOd5YzyTD4mLYOiq3aToBmIq1MSjr6J5JwmYfPqb/3OfoABGi2
jMilwa8E7cs0dR0TP1dvq58Qg3BIZ0Teru33iYDiQDL7UGGCAwUt0oGeGdt6u9DmAo1NNqTvoi22
A0xJeOXAO3EYcOIS7Cx0zqNcEYEZmhYFO5qLByJwtOVWbEKHu7GQgceLEh7IwjioowzuYp9f2Q0O
uqxwSB6O1XhaLbm8RNCdsRmUWU8YAGqAGFbgqp0zUzjovLVrJrPNluTtsxI5f/0MiTb+P/FoA8sk
eaSzRgpEySSQ9ROoF0Z6ktIVEK3Kz6+wgoVHEEBMNjv0kSSpQw8YXuu0ZNoEYMwIHYaLnoWhiE2k
zsGm5o1Z1E1g5SM/WhHUOJmWVnzrZhqFXajQLoaA+P+yvkz+qXaWqU8o6Gtcq96aL39aSDUVq5FT
e4wDIsOcX9wwqLM6HqT/26boJ3ilOT2SiPYc/UTbYCJWtzuTy+hNYHBWKPybSzWRGfpBc0QGOPMO
ef66KgjS8T3ujTLZ8eBqBmZaYVa29Q9ddX5y8Xj4eztcQWlcJj1CEGuZ4j65MF2OlsDhV5MdDsyE
J/zvXbybXdw0kq87nUrlDwHS27WdVucDdp8KLOkYm1gsc56lSGykqY3Acw9GMPuNFUCPEnMtK8sW
VZX3nYbbXoDjMy1tbH04C2er3QdZAYj3mOzfppZEEqN18YxBjmxriTnCHdfubbpjs3ho+svbvnYZ
6khM6ze/cQi0ULdlJ/INHhmkCC1CoHmNOL6d5QbpecJeT8/wORbW/kS+Miefbs8HJ+NlFneDSwVg
cLUCwYnlCLJZthakdygs/u0yCZ2QEBhB1RO3lWGmEOb8GFWr6ITQ2tQRIzVUjRLJgNvDoW48hVjk
do3oBcr1mwJ7N26WSASgsVsK8L6Iva6FdX/hw4f8MqZvy3m4AYjkBaWkOnt13x1u4fGGqjKP+Aqo
i9fShScw70NSoWtYGK0F7fWqxD4N5b4dtWVBjQEugD7sjD4bN09M25HCLvr/T8C5pl1Rl0r7yEPG
AvMvig7h0jePcWixUqAZEQrzYUiCrqFr9xtNQmuDtaAb2CZWy2GF41zucsQoKMsWJ3J4Dpko4rfL
/sIW9/kdt81OcGuowScIIEqioaW9Tmno2S26u6uMjz4I/SN4Y0sAMfie2BD67HrDsKSyvSgVgKsh
LAy733LIBO958Dh9k3y6EyMgtjb+8hE2C0KVA19sjxBt6GJhwLcLn8yvKaKGlHVdoHifqwRgnXi1
EyUOsw85IeZV3iQFSK1f81eeslqLuCAPQW+X+Bl4eALvH1+gaGuT2iC6ELb7+MPgPnNfPVSbaXW3
fU3TmxcRNl1LxbrIU/atAdCceeKGMy+PfCkkl88sDfwNYWznloQPDeLdGJCfuM+2vyEegJN3lltC
MCP6ignz7MeNTwlwbcZTIp824jAfYxup3Ukq1T+Y0aSeGXZ0qGHe6CwJOyZnDccs0Lo+DJrr/7AC
PkIt8FbPk1Eo0rDw2gf/3i7xntlmp3rtOpXZYUO69FB95aU4/gkfuvKS1CeDmBMeRN1c8SLwMmV+
a8LXrh3H2NZIwRmpzI0OcIWODm5G4OgbqmpPee/EkJiAL4hNq+t08/CVzCS00boI/Vnm/dBU0lfY
vI9HxewEJScTFbFTP2C2FdMMv0V5otWlc/orOQRHhYkWUsFWEfuiyVKZBquHM1HviRCaoDB9U2Xc
mgdYh9cgvT+BnuvB5dBDf5Hjic9URuUui1tHYCPAl8ZCIYOLuduR1Sh5lHbNYN+Y3TyL0sO7spoq
Y5+12S1izAFUposgPGKkoVAkt3taXlHhFA3esDHxz1XwXbZ8fvQa3UHu55hrMApXxl7TVNUyzIUI
BFnoJ2p5KDMxNepRbeeRJiZMj0Niz0Yh0a9NK9DQlDEg0i6sjr6zxO4+LMN1fUil6DmlJC0m2muI
x/CbcbMhUVptUkytGd22r5gYrLcpFvApBimEFQ44wYBq+qSmLBoggRAEHVAq3oJ+ObY5JPo5ywrD
7bbdX97KZyu7bRgR1eYj1qedllr5m+RK9SEtiDrOSGkULKTPA598Zyey000gtrHlfwCHtNNJucsk
5K3ciXf6ay0rhF84dqJLdmtysoAak8eCk3KplbBXZXhkU5n/fd5+J43uMbVXpxtADiQ9c5tZso73
U0nzoyY4TNPxc9JIQ4RqaVfogKjGoAdAb4o2YHkwGPiGRCT3M0p63yb2E5DNdxLzY9a2am1B4Bl5
nULMuu7dKsvuFMQnO2NaGyTn1QNvEnvTWzowt3KcGfR+qdAO88f7Euf0iAlDGwAg4+86sSQDhq/v
Jm/UQdPBb3UIgLTS4xNCruc8FyWxBXxKkdfv629udliPQMQoEivubce4NhNHVGyQZhqOZ2tw5iCR
SapQKhPMPhy8THg30AQlkqwvCOKzgj+LewgJkrRVRlq64QS16tDLb8DWsQYFEbBhC1b+w5AyI6oa
d9DuJXZR5FYCz1IMc1CNrmpeNCCy2Cf52CCj+Ny/nHE5tZEKT0uCp109FBW2LP32Dv52W4NdhilC
8Tq1sU3q/D+Xfrn5h/jJZEnr4Hj6+ug+7/WDLfxt3Q2Y7xtSqQd2BhyyJA8o7ng2WwVs1aQPtTZj
dOvzsFtBQCkYWs+yqGorr3Taft+c0WF8z2Hu5C42KrsMJlZ4+MwiOCMUY1L+ByrmuSzqIqJikXxU
dL1f14JUzzqY4Bx6h5kFJQWUBQl4P03mS8fZh44dGAB4M20EqmEdMD7ghkpUyKpurk9eAIv5SaaR
YLKVSG33+oT4o5FLfGz025vqxmdveJMT+JlXLzgCPtRvF3SmXtc/pQVudvf81a2WEEJkymkSOkih
3TgtMLwqghMtqv4vrOyJavfGJm2n6GAzHf7F5XoQT61JxrhowqBGrV1B+WjvZS/2haC+/x3suODV
gAzPNBfcFB0wLt3JagAB5tbNURrP7hv4YQULX/mox/08/3PjHB5A4e6D0Zqcfb/OMyXwoAnUfRJc
FvVzimshBQXCrFrn8Tb7zsrYx+uHhdSllHdGCWglpWNYaeVJhO8vh3wJAMYDfaeB8JsyuGWEXimA
77k3YQAPUDZZ/g7/TLd8OAqigXQEZcMtvUDNA2KYqha8hT11tQpHaa3oHaALD1JxqLoESw8RAzRS
IVpY0YQbWdfAi2je3vk1qVeDwBQQxxDFeN8H+fV+ZZaWeZf9+7ZS7FBWFzi8RACu7begNdyv6AhX
tIp+07ijvl1jqyExwpV69Ss2oCAzsKV0UhcNUuhonIuHakljOpeXx8bSPYcS8Qs3YYBv9esQuz3t
WzNueDZuYwjSkjcOF5CN54M5rI/wrSlUajgk5KVWv2Oxzy4larGJCCSj4OOnolDrMhhT5ja+iKaI
9c9ohvk9ScKmLOc6LYEEHSHtYt/3+FxNVZDdQouT/TfyPte39hF9FywfWEicc6UL981wkJP409/+
hpyXzvKZYD2t5Js1bT958JB/8xBsj4MGcaforTFUxOfXsEHsoe78805UnOVKDtB6NYR3VholaD1q
rTJ4rhk9OJ2NEaQ2ZfA0d8iw2AtTDIFEk51IllVxo4NycsoiCtM3Yox0PvMbz42TTuVADs7q/P02
/hRi11Qi5UiYnsiiL967gQzLVQCe/F3RsVmye3jqi428zVROfPxcbUsQje/ZBcDKkQN5FODt3Yml
gfnZJAFu9j7mb5YqOUvwbg5fXCoQsX5pLnZXouPYlFrTscsjZt3Swt4qWTrN2ZPKhQcLHmIh7Axz
qgpRaUzbeiNNTAJp7/Hs183zYGe2Gf8HLG5ZzfUE5bJCsbFpqvhdcQL8/LKcU4fAGe3JdB7Jn+Oo
pXVZ6SMUE4Q5LnGvwo+7AyroFvFzSoWAZfXos4zk4U5N2V4z5FgAcoqjolJNz6J3kZiu1GvH0QVc
Ftsff5hc5fFDXi5t5F6guv3zLm8HwrEWRBgovk89CIkO3KmMiJ8HU77iqf6LAhXNxz2BveKITEqR
8k/hSslGB5PwSR2ZpdLRvm0AE1+QTfCBmo8HQ5tQU84dHQRZELtzFDbUlrxo75tdgl1bqCWIJP3k
mltmwgA5BOsz3s6rP9cJ0Wgrrz7UOXb0akk25+yQe1KDXBvoiZiUsE3qUJYB7GIB5fnFNSmphtlc
y+kDZ2WEf4ofRHLx8jgBK8RlyjuCuWlHn6vy3Dr4cD7NCmI/dhBfWO/LPE4Yu4rU5e+62Kchx5AQ
cymTOUuoqt2QXF8ZhcH7HDgDo25/Kq7gvU3BnaYqPThBEeW+ZHqVbbrerX/mb0NNl9LvvxNk1sJg
393PFd/NhQbskHNUAB4TFIReaFOEkqc8ivXAhTyZqBIeFzEZnynNiByMIm8Q+Xf3UCldNrzCR1p6
HowMOK7l9EBDODVWQR1ITfmcGBsEMXuMDCnYam1AZvFCbzmwRVu4LCrOZoKG+ERQft8rbRcuJmjv
nZe1s5r8WrH6hxjpMC2I9eEele2E9BVL6IApH3oltRhhzJda7Kxg+rlNF2Sa19cH5kWaxXNfOSeI
6nfTNQMIkNrquuD3MOwMCwIOGo97o8u+9LDCHmLdyL8VvZVRw2Mwc57bXGIZXhmpCIIF4hPpb5fu
c9DnVxb1DtjN4EsETmSvCZvti8DISy9d2MyoMm39wuaMx0/o/chgkyQr4wiHIUiU/G71RgJYST9e
BKBwoPqvvBZ6CkVumrEe7BEQVVqe7GnQ6vjZkZnG6ObTc8h2pThY3LYhFg/QDUKKHvnot+If+m2Y
l5wDdmRxThYxN4ayxSaNe1KZhg12JC/qj3PSPkEeNEcJnYVNtU9WzWNRTKZTKA9C1zgbnfpqgYRp
6ySn0zRN53m0EwxPxKD4DrVRZjf3z9FiQgyqaN/a1ttQTQb+LWRxAAcYnCAXtCrCdEorKY9iAPYj
pj5aX0U7bu3ABRBXcb5cfkAngeSYPg7GtFetMwECruPtso7EXD2HVpU6G5EEAZePWnHgd/03rNv3
iK+YuVQT8dL32xX5hdqnz92gMUZq7zHLspw7YkPM/3Ao8aFA8teITlLnMGWdPrARpgyLHYvfbtLa
qAK2FI0vfurdv+nJ3lwTSDMxLWPsXnufszc3vxVZcmbEh8bsVlEwKHMHlIOiUrLijmopdxoZJ0+P
7+KRbe52TOju+bX2cB/70jZft3EDiuePZ7ph/W1azu162ij1tFT3e6toSi6eYf00SF8futTBbwct
lB9dXDs/yFmK1z2CWqE/SM/Es+LgfqC/DzOJDcFW7tcxW0zb/hIuTWnujoBmxiR3CWRbXYjHtgRc
GwgpTEHmg6MfghEgnfNr+rwSz/4g3dEheLUmw3LT9OIAfYbQsEaNS/oM51ol6bJ/DnpaN6YtLGgW
7UkCC09xDlPIkalXeo5rGsM45hhbh0BNr0alqGjJCXBiMenDXjriE+SImirTcKw/SxG/AiBx+3Pp
BGO0+fyP7sGurZHXzCSiOIeJXwtTkZ0sNzWbtyFWWIXhq+4H11pDy/moIsD0fH5nlFq9oVqXBxLR
9UoQUs4pTqdebbGHGsgl778vRXuHG+0P398ykMrGl0x3AAESJ3idGC6VtUFDfmoOGLEW9LEjDZdv
0z72B2j/uHsEPqGxy3OyVdXqmbGJYuKVwL5w9WEHX0TTWWxuqrw3K7u7JJzTNsNnsU8R4L2OVytA
ycAAWjmxJODTYbGx7/G9+QIKZVdJPf1HLENIhEaMOe+FYO+YunZZZVPokwAVBmPpsm81p5eETq3s
jbdTM3E5rEZzTjcbc9IWxcDJiUZJOnelTouf4TmjJ/Er40gvUp8APGRyk40yFQ0rAn+lEBAAkgiT
S1Ali8XEhzOKApsbmfVyddag/jfCQLR4sHqcA+ixcJNHYBaJdhGncsPIrTCtmJU+uzzpOB8jqxmx
LND9pNOqpNeHz0rq580PP3RFa/mDnQ2T6iEcqjLHAHpC4F2qpDifxnVjZm2tX2zqJDW25nZoBDEw
k4A/YUmUg1sY+V8q7WfHmbbDmunqRrBrP3DnKg+5xb4/8jrZyvHELu4blJYAJuZq5y0+hwyAnXCg
pYoHiZAi7mG7vPLDjChl7XdmHxFPzKTkkhjDiM68U8vH47jDGIqhcpBms5E9aKdAAzl0SJjiK/Jb
sCj949sdJhAa7huLN1SYOWxJOdjkrdg9uF5rbOV85aPlc+0KIbMZz9NoWW4oaMRbNRcoHicgO/Jt
X3tCg/ciksrHwozRMNKIklolr2Z7Jz80hl1+dYQbUKDQMgVoRofDaCxTB1U0TTd0Fc+I2lCds+Xt
83LAaOZTGrPbqkeDrnevXJmn9txJotCt4J7XthU2sMBvBWLjXOLneAYq81CVs0yaeUCoX/gPORfK
mAiEG8AQWVwuTHzSmZBT7xM4footzcGaCRQrnrCX4zYE3ZxqH5DGJUrDhWx/eUh4YeaAEmBEdMRB
iGyBy3+st9rYi53K8Nbq3L/2f8UoGWrhklpChWGHuR40S0DMypKS6gOoNZNqqYcgolM+QI4YRmTW
BBizXZiuFA5B+8PJfuT8baUFokon16M30uWwG7z+O8GAM/EE7TEXFYesJFWX5PgVlYJzWA2yXCjb
2y49BoGBt0YmoBBwbpWiGhvV6QHcZIvp4dqkhSNf/TzvtSyQe+soaIYbwCDQZ86QiHm67bmI1e5/
4PurGbvOyhiljwF3jPAn6QKCbLZlmcxrF9vxYoG33LlAp42VJ7IKCvejL2SYbxy/PzFUUwFmOCXc
V2lCS4fQpM028+ZmOpnYNIn6b8JhJqFrtCfWGupOC+UFAPxwy5rXc6UXuiweuC43hUy9HVxqFLgJ
zVfHCHuRW2YGRTNg9n1+E1QT2rpxrVQaXUaofx9IM48QdeHPk8WHq1yKlm0iSfaCUPx5q8TJguwf
ScrX4qbw8MDd3Ckd/cZFQwFRXwzsw2zhre6cbMrU/Wy/dcFDrc3yq/jmSn2rzvRMCkfs7wiDuXTr
1wvN13JQqhf77Zewh1GHDdJdVrvAbKP8wAxXMmTtkFNbPVzOL0u4046t7Xd0SceZUmiNWPsm8oRz
gnHyrqs/inbOocyRXYw+wZPQo13FIqwvZMCQaIw4Oa8ygXHgJ9WtbRqHwObzjz9j8Z1waONt7M4k
IH0NGA+tddumN4OYe2rCSLv1Y3A2Q9dGVmugT6Jc6WEycqWVTIl4S94iC3ZQBqxwON8yDragxV5V
Ofr3WJTOnyVH5wV7/Eq6AU2JockMr/gB3w11wJ2WxjI2+v4UTyP3Fr5csOHAlNE6RMnZbEJaZEbC
aokgqvibHy4mwX2Imns6qaZ1s5oBWb/6XFtv5+bZEaSlZXz5AVipM6X2z1wl920r8dv8I5ewvJtD
BSU0K/2b4m5l0k6mfrSqyuOS7iVpcQ00UFjBa9histG599Wtm6pC3qpvnnf8N/jA/tJA43Suztrk
Xd+WNONrAhdWIRZ+d14jWLbBsMZ7mDPinTMMgKSxzsxkZvBkEfZ8FBl0P+ZC+BcyIdqVzjHEnS1Q
5whMqQn6KpY9agDKaOppw6+e5wxy4TzvWQKDiwhZ1sTf53ZS4EXyGV7XuOyOTjbOL9fkAtNcqBkT
4sgOJxNzFVmZWRaqicKZj5IaAF2A5VVQIOFSnFtWLUt/jQGQfbP/17I8UXPWHSUR6JxeOMGYSGS1
DDFvqZlwQi+/r2u5PY58DPAQNWNcBTpKtY40wiYWMMq8QAcLY5vfrWfIrFxezoKSQQL+xWGZdUlS
EbYWbV6koNfcGK7WEPqrsF4wc7wAGiI04Kwb0d8IIGNAdWMrJRnVONTQZbbNP1NSnIjOZdUQiUEx
sPyM7naN7djmTKLOdx4Kgv+IdUwtYKzLeWddcgRnd8wAnDcEVVmU3PZJJW49FrIuU/vr7MtVzYTD
ssX7432ehebMfbHbT7CzLOjnk5BGzPgDfRGWz9pKOnsLdBJzpzzXJdj4LYwY74MNw7s9pxSpMOQY
raoY3whBZfswzlxCBBn0AB5rS+a78CHFjILafgGDlq0Z4tcKmnZ6SBCMSYqcGjjETFHxfhLU3FU5
rKMvNoh58AmjSh2bMgRXj73BbL32hPETDSrMFM6H1lsYpN/cYtlNcIaiETt2sNw5aLF+ayyBZ5Pc
/BZygUbnH6+sB6+bxVcboCeSfefutMsZQdM3kCNgoyWPTH4BDdK0LbJnrp2vJ2onLyLtDfJbC3e/
U69gvudqCowBCEzfmlLY3bwG5go2tYIS916wdR3JVIFx+ddBRIKOKk9Wf1Kp8SgP8fl69uhmtu2b
2lEg3tG0i7HWSFxDYUZgftFd/hYixt3g5xpVBsl9leFMHVtO2FNqimI5enocISI7O8/KMk1kk8xu
TYs9UYAi4NDp7Q6nd2zemXmzti4hpchEab3nj6n4CbFVy4r+/aKv/7Qt/5TSUzjNm3B4Nx8UlhtH
D14OA4xcvtZ6f8F1jrgawuFs3/sNlIrLozB3YdkCjl0j3o8B/QmTTNe2L9Y4BecNKxLzWDE89tRI
seT3VMKQZH87YiPe5B7eAsNN7QwrCP+nvmsGV+ff5zBnpuDCy0jb8zJIW33k2cJpYNpqf+0FViz2
51CYKonoRrRuxT6DrZsD5n/c73JqFTuGKApFqN6M5XluNkMld7jeA5zXPxER2D4yYg95srgsqrbF
S0V3CYeduEDZo4nuYzoHVMOH12OP7SE05JxqT/3K8IqTaaReMrKjrZsRRgPbFAnrwCsmMw5YkJV/
Up1Fpmh+Y+WdYIVorItFrIsQsoFQmx+pSp62QijD7kIxhzQxbD/aOujAvr8RbNniXn9GLSrz022X
tUCcZ9qdORicw5YZ6yJdXRGOyGuXhwxf+FT/OoAyOq4cc6GBw/f/xW72Nf/cbpPMXYkr1QPas7+X
71LEk1qiQ1gCBQJR5TOi1d91CL4STXGQeccOANW0m9kDrVzdLOG70j+cHLP9nPeDVkGunplMZsjb
4vKrWZHDYmXeBiB9LqtknkhB3VkZXRRZdZRiGQwdPAGYU8NEnR77VMPZS/7h2lAvs3SC3JPDVL5l
jjAAQ3l62gJAUzsJbKV3JKLzdgfbdAAFHnxDmrWkrm8z2fIa7rHVUJUFIF/Q+u3i6iW1n1D7a6E2
QdmkA7QZet+xKYR6KRE1cPrgSuCyd4SrbmxcEi9y8m4WJZRZXyy9ICymo71N4fhqBJM4F0hMyaTA
cNhBBTP9mbvlKjo9gB+szrSj2GLeVAgcM1ZRbm5Zpdel8WH+hqQUVcqNnNQywlsEACyLa0Dihj22
fGkj718buSGOryIVBimnb9CDeZ6Cml4OzfNkomsMTb8ACFnDHS/LF4EzTIVeu9LFkTkH50p1OZPD
jYcF1UOmeyZxjv0rLtmAEM2UMiSH5CwnSjTnClYA59x0S1OtJDKkT7aHgyyCySgnwXkp31RgTzGg
mQzOVFvGAsld+6KZnd08tehlaJsJ3QpCKqDH0xaqDYL/6MsDVXVyBuzySjlQOBuJaQkT/ne+V6qe
TCOB7cevZUvEAmzM6ygQPStavzt0g9ZApTqk1aUAZ/1bvqfBBOHhgyS9jEwyv25byxZV5xnoZyyO
TCT+8Hm87wUn6X4O4H4eP6sk0MZYjE7TN8STagUdqVG+lCxEPhb/fxS10SqEsFPwZj+8qgyuQY3U
8tDEQGbgL8JwlRxsH9jtQFACr+NJNS+cjd+qXKaZ39s13U3RdnAPj2O/xjKwfskvpMVSdMwqhCLI
ybQ0STagTNKVzEhIZiQS2mIsgcBLRANOPD2ZGca9I00snyIeb8xM577XSkhhMPLp6+xpaO2+0grb
mLtu0W7Lg2nbP/3PYIsQJUNMPwB2+N45z0j/ERMQvyB0euu8aV0ovjxyT+fWt4IXKI9a6gLz6SSH
MR/aNOmiSGNrppQAqK1Ui77gX4Nc7KOxKX0fAT2quFYmHdakXXYDoB9aR3d2gKhMUpysyrDyeQZD
EKwq3XHwaCIBdm9ARoG5YSiOljcQk5k0CGf5Bgj0wWZo0/vzbWBKRFLyrmpx9jq8+oK4vxmMRUom
PJ3UicpTVVpHuzXY00baUGvrGud6X/ceVAsctZpCNXEIJ9zAB5oeRRWnB5HTpaN2WJ6WkVKJ+7ej
uDhcyINaJR82FT8ZB3UU+KmBmfEoBjRAyI3FVD8CrrIC7vhgIM5KM9ZJJMrPrLtXmvS+ltkwhCz+
z4XILmcrkbUmuNtjCgiRXy93mTAbHTtjc/4Tobn2PRgWEV+BhO7Ndh+qV4Pscx7isvflOCF0QlhY
oaaNOOeb/WFwckTkKHdSAPL8xEYxemyVfT5or8w7oDSvHOcDH9Bs7pDRj3MFCJJ7n6zQSF/kL9GP
+uHfY+DWiRoeVxR0lZAH19A9WFdR5EtkEn/tsIAGjBw0C++O6vC//j0ImjKW0C6viQgFBkc5/cDz
T2yTOM2mGj7r0Kwa2/dgO6YgMggI+RUK3Ef8mb9SQKANqgiHw6zW7xHmH4WkQ1gnJakAbwAmawRw
HV2HjRmyYWePjae0fVkRANeyEzzsx0+5YD+8zreySbrNHWmkMkOIqYNbrQBBFtGnKUI3+chon/rf
tB6LbSS3od2x+hKYVl9gXPYLhKCENJKeIYYBu3evoQAnnUOGVFQq7hA+xbix4rccEooCXyML0Fg4
z9ztT/M/3N3c1pb7o7flxvbYDG5vY1Qsyc91t3DxsvdXZLA+F03F0A4mzQh3z7qyrOrFFbO0Ozq0
eB63p9iO0CrggbOoCHY/6Dg9L3y+CVeP0P+0AJLAmSI75dLKfi6wmZKzr19lLLx2F9PUUAqh6dNf
laMcsBVM4AhgAink48zvA4og6RD+pOByvf15ss2kgbW/IvEPh602BXmc341pJ13r5rMq/VdwbPr9
2NGOqjJEPf4lu8Ej+OojtfvUAxwJ8V5Lx5UvcrTjmSgvk92cMZPgdhebNgYXr4YN9x1fahhZ5ws+
0ORMTJD2+F/ocHqW2+Ae34TvgYascvF/cj+SGxO+jVQvIf72ut6D+qEReMe+nmUDdLFK5Tz9XjCF
LeDX31mneeqZeFQptR0+BYFshP1nvnqhA/DhDbSHAVyYN7LVFbzFMZSudGKWkcHwwqgV+KUjSFkv
swpp8D2FES8kdbGN/7Rl9ronNEuzYok4+6GbOCEYa4iXpqc3UgmWTDzcMOR3mX8PKDoBttMJUhAN
P4QqwwurPVxpd/NJNaKbUdfryPm8Ojfscy3t2Lchg3igsq2UryIzq8pCX5lUd0SHeqbjIsaHKLQo
yWnL2GfAXOZoaF119rDSiW1FG5qGsKomi5Q7X+RyYUsShPCd9kstzeSKuJynV5/4qORmn5oTD3zm
Tyr/VBKo5XpGsMLv6x4FV5yEU1VzxsY1X1LcZxF1zQTVrt8mVilwKmjE7PCENvQGDxbDqJHpD/iE
nSa5FfjMBS0/HQ6VXCQ+TtPnf6/6K7Wsv4ABUVmfAJS6VvCDY7yy2JTQo/8n5qA5P6LUZObwcu24
ydiJqTw9AuBaNC4gA7Y1l+8Fpr7xhCMNYyMIXyKZjNwZvZ3qb24vEL8kPjcZDDvKj/HFTa9sXP8r
XVHxnzFGO4cTMsz1RCv4JOdXayVS1vlS2gpmnz7LYqF6rF6JuET6W/Q9DAIe36p+VgJYAUKCtYTM
2tTP6otBV5TEj9Ouu33Nj06ErG+M0JP25XRBl2gUY7C7Im5axZQXAEAnTAkx9z6TZCgA9vDjWxHt
Xjx8+iP30IWKVHUtoXFvpdkqAMIgBrc4UsMWBXGz9m/f+u+cgthk6OL/oOz6Zth4usq6Zbgw7wyd
9xmbXgnzrRhVteuLxWj/9JauXE8AUQkmPo5JrGl6tlMuwDzptKH/VmQ9bYHWMc7EWDYmLUkGPH8h
cZUULPK+hTRDJFUVmB+InrVzgf/XpHnykZiQGujsj03g3Py7TR5ESSRGfat99TFOX5y+sdJBtFqY
pnaOjEfYBPA1e5WEA+2g+TpNalYnoDWWlrtH2VmWJQxrZ7++0DXJ2gPDBNLn9d71K744/ca3rXre
o/aUp7sJUqp6JgWdyFhZBo0lZ1sa4b5nocsK7eLandQCorR3T3/yUrhExxvkwPavEj1MP3KuZU8z
h7ME+In9L0UwTJZwp+HM/evvAcQLZ/RJs85xQJfac3456zA212lSeSbjfATXOBl+p91RoFCsfNfd
joqMPU1CLvxDPTBJUFoc7KyqzQNl/s9WcpdxDfLxgR/Fqr0ByvSjswP0aY+MxRiE+bYJmaPC5PYn
wEFCnkGIwN3yPu1eTOt4fojpV/CpqdrbNIZHnBzn5U7ycEBQqYsI4OzeKChVMYsJX0T9eNlPOd7R
M6cOPPeoxaCW2e6/dZ/giMYHRrTWKI0ZBm15jm4WuhjlV1uRmWToH1uOtBMU3hhCMeX3xqhtbuNM
NRRQxSmPrQsDdvokibcwk1TxBlwY6edaFyAq0KxgKLk8gU1wX4CzjLzWdvBX0ESThVKjH8mEyen0
MtkGfxN9nEPfiqX4WGhZc1DEIabVrq+FXEoKS6KdDK6Oka6lM9/huc3I2OJxWf5hhuQsxiR5ydHD
+s+8gS326pzG+51jyY+AMJTlEa3zztdUxuBea47cxGbr/cWHjxrTy4glZ7wQ6HcOQQI3c6ZJINkR
TOowaHsLTVtcSX0jH229vIwSXns7xhVr51SP9Y2CsEueK74yyvz9xmiFvKw03JtEbdCyJzNxZ7xW
kNP1PEZHolkymbuUjFWuAlJBIwFP800u1NSZYDp79fe3srI19uA3en7Cs9AMW8t9B4137wLtSHlz
8YsMBSVEf0VPJl3LWF6h1h4OXgPTotfkBT4A+t5lISvEW+aXwTuCexqVyx8OuGZoU1EcD+MtV1UX
L51NtOfdhHi3vjWmDtqAI7kk0Ut3faZ3oKXptYpdWiV9XhXzdBS0oIWXDtoSxz1wNS28Ua8MEsyi
AXoNCbXX+CdyNKQ5leAQ4Xt5DgSM9vIa8sKQam8X7Q53pgvluHPAFGZTB8VFf5tzqWvDZL2ZKiy8
MEQjKwctW9hDOXTeksgQ+gAPxNB+wOpoTb0ICwvZwZopofMA4nkX258lzG9D42ps59PhO+5egqas
tecfrpz4+XTpKzIWhBJ5veJlX2SMuzjrqMEfjzE0qCRyp5p5Lmx1MPZNxEosOicGkO50zmff4m2b
EPikGG8lxT4St2AT+h7LD/g3E0Rfb9ypfagWA1Lh2kxpjJ6tsnnA4fWUGR35x9m/+9wWg4WGgsLm
WmkG2xPLoL1eC4LxO0iPf5nEwc9wZ4sT7oQQQyy0xlyUMJ4uJb9IfPyTJh7HNruvP5nVXvJ6ChdO
sWJbIZCB2jDIXZVpCDPKz5BKHugwjosUmzL8yS7Ti7RrANNixgTaHnCd9X0nX61TS4K3oWXDydv8
dmf97eyslNeJkGC8IOZzqYYTpmmBRem8Xbswp3ZcAeVUCePg2XfzM/0K6GIqiAZ+LpthL8jO+omz
+cPedlQs92OrcyTxW9M4gSAgq6vxN7t7FRZO5rjpPpYkYTJATJUSysGhfGeHqEWljPLobuSBpX+F
vivk2dIjKJhquYd9SuBJfn7kwaA4sk0I3B99q+OkhrCYWxueW0xRuoUkilZtWd4aG2G22gInXyUA
dTln9+U7gpSheKTgZmnttszL4qxQ6ov2zflDs8svTug4wsFDgZVgt5v4Zqet1/i4geH9BgH5R8qG
2mFPd94EAcqjSqupFKAXm87YWyD2v7uldKI4O9mIkJvaKWHb1TfTti6z0TORV5KAlfpzx1pDOtku
QBZe7X/FzDfc6l5GFFICrlYGZCm8G5vRYltqRb2wF7bL6XvomfCmV83cAfwsgwAislOR3uc9V49V
jmc4LfrZStCYxaeGdHZiv432L1AgxLpf/HnLyqxrFos8OTsg8Wm6f56+zRwwL9qx58Mjv6sN38ZF
Grzhcd5g8xUFaMFgJhasjxnnh5bCAXfTCCSxzfE5vq5/vB2iAOdNhZuv4MgkVWTFXFKGH0RSj7bS
IV68UTCDIHtgJeFOAnv9uq7YgNtXfJqRePUy+hzb5VdJ0EXkxxQ6c2ZqmenxhYFewuesiB1UqFoz
gfjt9i6ZiG0nR6ioF5GOZ3b3SpO/EpNf2F0gMaLK8j41bvQKDBsg+tskpbulFdmN26lMMbUPLAai
CQ+1wun88VSNaOPL7uIAAeH6W/i/EkDvKxzIsJeBIN1+RSYSDRSNkd52C5TwSvy1f9Sc4RrD7rDM
kd3YSl2BS1yR0SS6sQiStHog8XSHPNJdKpaBu6j3aVkD2ZgNC+RA9sGXUv+0HPJKxUSqdS0qe80p
H1pb2NoGZ6hOpHmo00x/6qcZVhqkjvvEQGhwzQASRMZ+XVqzsbNclAFB+5W+55HC+uvRX39HYTVT
g5zrJE0ytoMUwkeUflyOtEdDvXUczNsXJyXDUAB4URT+C/qdS2nNX2tx0fDVmWdMij4DH2QqpxJ3
qynCOjHUinlcNbzRIaIjP8eaYs7KuOZAS7JqCjLMV/Sr2F6SW2WjbrPKF1t6mgyOSgaMdzIJqf3c
IoRREGHSXSkqrguDIpENj3qC+Nmo6TZ9FMy6JjbKSx1/OxK3qHUqQRR+xN+6neZQ45JxwOLMfWhm
oxxGglLJ5nWpITNmfVOwu1s/1jqAK0QRtO+CRrrLTP7S2qaXjkikSAxWfZLdC5iPWDr/SdtPaAcd
AawzqKNqGYnuY5yR4+5HEESmrMu91Mqe4ui22SjA+c/2Q9rX9qcFVlwVusigRxeq1dnwekzw8nh5
ar5tB6wOKayHgCB06WifPVitn5r9Sr374fbQfLZuwOMODqEYTPwD/mMNhUHmVDis1/2UXToLb/pS
puy18/ElDafrRXNGkuoKfkEifWgSYqeu54aTmuHHEhKZbCl0OItCmwmeS27gULGlOx943i8w9YEo
YQFTXnFIvjYzTT6tIgkGmrLsWXSvEdob74BBHf2nn06450cSdMYkRQQr2RLU6lg2Ni3w84Gw8pv9
VXjf4br/FuqD9b+/l7cbkSHHc/vi8CgHughw5Hny5qOXk2NMtvCg+gRJ2cNIep/6E8qcrAbQ0BGx
S/7N6fu+FPY6N7uAAo6x3fLt+fiVUzxLLQtqaRsAgslQ7WF4WpEgN8vswilfNYZb7SwgURaA2Vhh
jN9HEFhoJEBYDjSys5hzUa/pE1ixs1bgNUV9YKLvfm8Uqln+uKwb9rLyw7FItXTA6qVJ4XXvXKUK
nkjudxeQvxjE/NgYTbnKmcUcctrfqMka/X0vs6iABYxx+nd2t2G/hlyjsWABfQPQcjKFUUMXRlh/
vmBPUtkkPyztoAz7SrAQqUJcEOY7MUvAWCd9C91WnVfAQPWLHrOLPvrYnpH6fPDMdVLybE+VN2kC
LsspH2AfVlu/owPxFCqVc0LuIzwCPCz0vF6ZpQY4+V+f/NvqLZb/X2tsq5HT7I5otdLY9YXpK6AW
CbkIGM8IrXKwPRA8IMGRywOtyZPd8fw6V6KeKs7/hnSqoM9eQQrHY4cxNKt0PbYVa7BviqAh4RNM
h85Yz9ebAm48yBst1SIe11WdjWJLGjXYLhkB1Dhu445XVm+PHl+XcCmqOuwqU6d8jbmmaWC/bRsf
ZJo4FFhuMKT7KrVjslqBLIRLMpZNio4D5yW4Z5hhvss02KPfBraASdg0Wq4XEo85twqrQZtHGkQX
P9RLX+cI1BbXaXXx8E1NJdnL7FLvblXxhldoqVoGD3yU/cC0dWqgA3j55kQOBfKZDpvNjejbYz6R
ZEEew72SpOB995WSQ2TbDk8gBj7WNnKPU9lNMQEELdPM97uI9J3XvFZVZTFfWm2hPvS0pVsTyj9/
0Hw9sLMIbaLTSj8K2k2FpGlNc4FBeo3CJelL1vAL+WrZI322o8sY1HF+qRb1vROZb8G3dLdex/yy
RxJY5lncRM7qYpM9JWlYDulY9dUwfQV4hLyRwH/zRq8grQ7Mu0aGPrGpr+fYb/RO7Q/+tIgBbzQo
DhWPNKLi7vG3abrNRtsIuJ4QVFFANlKV+6Bvj8E03TmB/ZeLf4Ix0rCpicDWPbPTCP0Zb8Bw4GEy
5KoOFAhtYtnrWlMc1NpXCpXLQ3/GXe8HMONXLAP/icBxuGvdD+xlzpMs9aAqGa6vmVXq3/k7y0+7
9IqVY03PsNmcVDXCmdVLHR0F0ah1VeaCo2DbRqCNgba26J/uJu2y7jpASUXDiWA+lesX9Lucikjm
E5TNSf6yv/Otn6BS7W4iYFjDJJ9lQK6m94TTlgpmA+kIvsB06zN694UtS+cQkAIFiRs214aDr9ZL
FfCBRLENbCEn6CDj8ZHLluSWrkbdyUyNUTaOzie6nNwIdveHXCN4iDm4G0uq9zgsIkkdSwdXAysT
sK18sSIEUutmV9oZQic0pRgqIa217KNEdeosFNMBhvDWPlDlNOFrODPoD75lCui6tknNQTQVAUib
MaQsv2HrvQiUiDCynCK+BJzQnKqh40GjOE6y0tTJLQpNpDpbcQrp3bI8aTHT4gpM69laKAG49jkg
sk/vO60nBYqPGM8KeHMg9UPDxFk1V85+56yayhxMFbY7WV4yD153eYNXIA94eMvfX1aIYOJEuy7D
uTPSnzG/dLja/Sq6bhQxfcR9vTsfpUyKRLOXGr5+4lqMI0dKYqs9g+x7Dd54UThH8gTYdSduY5vJ
filPfYin/5JK8ePiMWKw92BOM/CzMHdxBSCST0IRhv9EYGB0sk2JjWSzok/ZKSCs3ViClUiQN59r
wD3HZjui+DPqg9MEDeKFMYh9Klc+hAt+utfT2kvKeynoY5FaY9yoTJmDzaCFwpfimm0FATYmVSZf
2bF7TA4/uZf3vCGa/6MdX5JGDKbeOP2TEfuiS4wjR07XZYH/z5jUwbtcCegH+KjSHUZP+QyztybP
DEfvaQgX4yXAceeV/rJy60O8axI0bQisYYUqbuHLCPosQ159NMVQF5L5LIBDwsr/MYy/N22nyZkK
Qnzqq6M8SXbOoSWErCmr9d4piqNktzEA0LbmNj0hm8M2Yua+qtx3e10xCTiGgV2yVAoI5VE+dJaT
KICN+JSvle4ZYANyPBMd9xBwhBHlYTuXDLGw/Q3wIoGgtBaCK8Nag5l8xoYu4lY6ljjJuTiv1hDc
wtoV1PDG/i/TeIBGfpRmcMpvwmuW+iOyAAMMvkmQHbgoELaosmnyM7ssyo1nrvGf2rhNIMzGUiYD
/5XJLVyGVRLof+U100eES+Vu6jzkod2sRirjxSuRuCHFZn8jkgvLKJ/t2bY6HE71JI7uqoId9Lz1
4KlCl9btSBjuWQ5n+XzdEb0FMjlg++8Q62Oh68q8XGMMLz42WFbPQfMrAxcc8YnDe3p7EWAAUgQ2
ra7OJ76FlLwis0i988rza1scimRN7gsGvef0xR2zQLi3V/2OL3QkaH+xTBgaib3K9skF6U9UzsiY
RuSSJkmWfLeE63jUpEleCr4lTZ/KwKnZbaIdOuNibpUdnf8D+TWoWrOQMpK4wXFDRQovHpx4MxxM
dEePUi541AYkM9kSTUb6jamEDa/ZufVcSTUOYaZOJY1kIXz2gLoZ9NarQsCwizMl6HSqhhRnREgn
5AmOIuZxXRz8YTIkO9rSg/dJrOHiXZJE2xyllulS8Lc6TBGYB07sdPNLO0P5riP51RYTfbj1HAt/
tw5KsdQk+Wbm0lotUsQ0D6MJzOvWHgfTJzIy0GsSUrq2v+cdRPMcP96YInxDQtFMh4gLPXnB8RYU
xt46e6kwRlG/DTcW+F/SAcS2eOeRuKRWZR2WTL9wUbsjXgAvD2fSAm9gZHrXuXSBDwnaoh9Ehpd9
uOcQea2xgZH77Rc7LVrf3RX63yWwn9yyK2uZHSGzmliHsQPRs/Xta01rY0wpm4NlqGygq3n3ghgH
68xqz8o/YB78UGsrPianvbcWoL3enEwojbKcXfb7oBn4uEcmlY9ZCIC7SI2sRTYJ363abXlUTGr0
vlqrJS0C+zcOTXKaGIo4T9O/Exe+Ok9ePp6/eRYYgbiQXz/sSEp13q6Vzwu9sKk6Ss7TUQlSieLc
SXT9T9JM3+6C7/7a3HAic44lMazZywfF00xe2YJdvDc7b0Dmz2F9EOTIHV0Xmb07Phq1Q8A17AI8
3egEkMfnchGorP8Ql24IcHoYnySxgIloglP8aDIy2+iadMUcznQ1FbcPEr5JawmXj+wJoAWxdpB+
QxzCU41EQ2EpSnbkhHYyBZSVdYxETIYGRTl8GVrSW0nTRmwy7PSoiq5FmIwi0jRzdQwgEkEtDGz1
0svw1UuVsYNqAHmPpOAmonQB1WpMJt4ZJGfQhrftGdvSlp4b4UB1kCkhnEIgVXNb+/4NlkL0OFwu
IUM4vrpzEy05gmavnmbxrkoDVx064Snv/OJL3S7pG2hEkdE2ax/rygrx2fI7uekrdY5dsPrRd36l
sbrqjxeQxMs8e3h1rrAfRlL0MSMPoOvNUn4V3gDSL4gZvq4jPj0FUkKDFjZrnLvU2lI4RvAmmzYW
mVgFPN6EdjjFzYbFgJjuQ5oreX0rT/DoSaqpkX5HxMUqzR9zQ+NGMGcQoQlNSwnDOE5E0xpB0+LR
oeimQS9Wm7eUj3ibtO6zWT+kFhLP9wYiLFyPCgp4pNLWtv4Oc45zFKTJ3GXvQEsLv5cAuIzTH4qS
/kTvcFQIcD7KSj3/panqn0euN6PXWFLJk1p+xnw4HTxh7bylW89s44ACRPzij1oTclMhc0jSdzgc
JFC1QeFWFw82/VQWjR7G7q/QgcwJkA5z9kHPXKhdJ0nrCXg12tozvB7+J1MvPm1/9/rk2SqaJ2Gs
+/AM4eCNxPVSNaWIXFWFy/qTi87yU5GZ+HyQjCTlCfnrmKAptkDiMPVLc5orQhFuMACQA80GCzJj
1EC/BT7mY1Qvu8/Y47Eyhg8g35ub0XNH+aBxWTzmxjouhKNxANJqgdaTkLs3gNTDEg0AdUQuhYOH
SPTE2DvBVBMHA0TseZDca52yo/u6ZGencXhYC0CX/NYsw54A0hb4L218wVl4z/y8Tts8xdlMSGPW
9qhFiB3KMjBsY0izNd2S1AcZfNamFujpEdiaaZWxbv/PEqY+YE1uSNxIjB+4xAM0bgae8y4CN2mR
32bJMTQ44qFnMHm22LR47evrJUd44MGR0Bd2Ykp4aIdjJOXOD/JD72EZe+QvIs3flOR12jbtc3eS
cEp61JaA2BQTuKZ0OFI5G6KZ3E4XEFn37dF7QrYw/MzcnOSv/koRC9kpfIZpqSWBQ68aZ9EwfUee
5wHbpWicZsqqgAtreD2XE9goiY8QC80kqLQXsFqlO+rUbDpeMhMco5Pb+eziipQz39uRqTKXRANh
a7DGsbuClKwZf2w3yE00/xw67tjvm0P9oSP2uH9e6/GNYgxjnWqoRpL/n399FPnlAvJGRQmdqGyq
2Z8pwFkU42H8Zc5xlKOc2LhnuLez8NhwQFrL7b9JWPKjPExga1uwIUjjM3erGSl59r8lLQIo5xgg
F9pucaBcCjm7JXGwI6H8KQltZVtJvZVeeCtY5aWyeZu9bDkwJ/NYzcvU/9uujLZf41+4TkfP2WFL
uW3gGpEBTls5dLFMzXolHcShmA0nJzjdFuCXoJRLxGbo3BZ7irSPGHWapsxFoCvlkv/XDeDL3VF8
T2ZjPlv8JSHusaCSDpxdd4svCZF2+cl84j7L9yCdX5hwnWM9DvlZtS0uLLUhAruvvH/ZMcK4GkOv
Ywmz99xrHn9f5H+qRz4Ty62wYu4ynsLmvS2y/49TjWYX2MJKAR0JmM2omAcC4kGaNhd+iTnfHuyw
tFWgO+l0RPnijUxLBbjy2B2L5iFmBlpRTHqxDsprVzjLYlaUyApC9QSj5hdBDomwMWhs4vERD0b9
jfVUc8VmQlBrng+Tif4yWhNfx4NToZAjIg+Mt1OufU3yLJtnYCPBjLX1Nq5z4Su+7v/aVdd4N+jD
gwBs7Or+24iAJktxvEhTd13PlMIrFPP4Oiu3/vMfot2cIUC18Xu75AwcgjAe/o0MIWJKuGuiU1Ue
VWeIf8JfoUluq/XuCXPlwbrZjwDTxf+nxHvEk1kQVHzASmZsY/F7iw8fP7qMXlttnjguuVZIH7nm
dUinSjzSKRlSGAP+GS7QxtHXGXlzmRi8ZdnTKgWjXPppxbfd/2i9Y5hWzV/e+2vrsm7HI4h+ufEF
S0RaL86sDNYJwyBNYH5wjGfjlvwtExuyQD3cAMAhFc8INSwa5URen6rq/X66cJV/ClaeyxC9EIrP
8jDV0rh1bfh68eguDbj1bXSgjwNmyQp1+lMXcD1L7mJ5HRe2WV5qCBoJBDCQknaQEUtTa6TsUDrJ
HqFeQOmEBcllC5xDsquswPBD8Oj9kxcmKs26E1owsmSrbDxK2Tuvnn2cSRKq009xiOP3sAGTMEKs
peEwGgvxcjrPC0hThKkEHf3LHG6rcPgUbwgMlpgI7Lk1vapHao9bvUsRRXvX5kdW/6zz4ruvXSrr
zIevEjxLkja5bvAwcGw12m3aYlzVIp/DbzAaBKFl6pAz7BiJ2mpCk7Ed/MNnb0v5r8YizQI8xzEh
9XfM/zRBSAVdtgD4tOJqStSL/1jDOeizXeW6V1jhFNAQmocC6mlTJkbUrAF+uMc2tNkAJu2Q1Qn6
n4CdSYWoXRltCqijvsODt+LPY72tfquS/ljj9/e8eUJvlcG8S80S2HzEkWa8vpCTUrseiRMx1sTD
2VyDeNDoErZVMdjtC7tz1ler+MMUbHqAXIvvBaasGbeEn/s62EMCh9Pzn/YZiN6URr5op6L6jwPs
FBdBYdj8n9cqBavxk0ucWIjGpp81Uy9AunHJctNiemtMRbcTyngz4HCnKpaqKLjLmi03C4HxnY2n
NbiZtpnIJw5rWmf96O6dTYUMRytGh09Pur8eh6V48Y4ICdVrFlj4Xl5xDXgj9T+VGrxaN7YG7O3x
YtBpyYNQTw0NyV5x2fQpas1ELG4fUiCVJh++DX0S07SL0XSf7llfHuxZQdyzpgIKFwXWn2qQHZk8
tqyJ02m3JwKNMf4EdY0hiy/1dYYPu0pNokKa2Utl2Vjn65KxAvb1qXQUkbJOvQItlb76KN/UlPGQ
MrOoKZbSlZjtGTAaUF2tZIaX16spK5DtbfSguQlAU5OYiPXUOLronG0KLy4/OsA9xYIxKVDOLObi
u8BaQbWXMXZmxzxufNvZx7HPI0MAWRNeX+OQrHaQsi2mtrcqK7yv5yp2ipzIiU9XIz7UjUFRvg48
K7oZEGeepxB6tkkkYADnBo11UqXZ69OcgYrQISZypYB907Jt8v4t+vvf/hVjyExMomAMD6gAFchc
3kwWrqwttJRscYTGEpxJB/UNOu8HKN6/LfdrR2Rz17RRn0ioeAPTA7avgln7DBMG/VDDcRkx8rhf
5nbnICRwH8VqCQ9dMIf5HEJwa+Gt+NqQh++fEvUhNLm+6B+M9WFvMrViWleDrp/DyMn/VkelokBQ
cOLs5TQOrVjeTM7sMelc/c5W7ZdIKR71xbfhMlWX6cPtPV9MaXNW0/Zm4drN7IqurJvM04IlqhAJ
AJDQHohJUNqjuqod6ijE/PpprH86Y/lUtj6KZcNryy85AKgCGPhQu1Md6MRIBAZxXL1qqXZZI5Xa
RDZ+DOWb6ZXlFE2CovDoJiAjFAR6toF9bVLM7sBNEdg+ZARRSTNT2FbjAIAt+qaHPn0geY4gd31G
PCv1bBzDprBIP1AGXucJCEfat3rJLEQbT9Ngo1SXqaBv1Bx+KspZyFNCTbiNZdQCTiOgJZf2qJSK
hnaXAATZ8uy8U5tBSJsBkpAYQsLM7w7vj89TQiDSZrUbVIjQ6jAWrUWp3UwPgSN4qfe+/xpACvmm
gZ3sG8SQ7nL09I+P4VY5sWhMHrnaRWq6AZqvsVfdVvbbaN2uLxJ2OHpzmLbwiEK73mFeRZySZmU9
GRp0TdSANQjbdJJkKWP4tHuKPQEELJhcBYeVhbDELzAy6mMNXfA6DoMHtXBWf1SZcCJtcuzy4vpk
FKTt5qfW1Wj8LRxBSvaIps59m5SSQvCVt6Q/pEx4JoiCjFQIjRHCNykL0/nD1cVrJZNKNoyCoZCl
q7a35Eq5+eOtTBLWX+VfI5oRExJgDFjuSxHHfdkC3RhcCssBH4RnIPInwgsDNlSUhlZqQX0+5Ylj
d8+NFxKirgBrhgF0nT/Bj7LTl82XYbKCIMHtt7po+0IlySIrvpw8hnJug36Np4D/goS5Ve2LHswB
2VtHj+HtZ/R1qGbqwjRcJZiPAln/NoQ80NqeXLHRM1jfXvw12VIfTKEJMnLi9temYVkR1bE6HRhM
ewf5ZRSjctHbbiwM8D4jTS57ah6lIJahZaPsUwsiOmGasqe7iaN9yVpAnDKMHf1vfVXmZzgx0DcH
Ue1/30Otbr2pOdTm72E8nkKpBG4cTZ9pEHe1qQlGWtq6ohkEdUGvcDwrGvw6D4gVTe4uP2cr0YR9
r3HN9CgRcpqPYuHluz7kqTxBsRysnFpZ3bY+Qgg6oDVyrR8FkpPEgCIRJiQSRLn8uSsTTmYQpGDE
phbqrCtdfkNlPbaMPkMKaxCIKFoDMHtpzQHHOGNIr8G6XZEOzBR084pvePywAT9LChW2xq91qgtG
SeE+1pnehtzaqz7/SByz45y6Iod2sjIuHPeXbRz9L5P/dVYJOjOtZ34LwQnbM71t7JrOv6Kp0O/i
FVfX7ws18dTOC9eACQjxdDAk6nYiZeJYND8Y35zEaQ/qG+BNFuHLmCCto0pBKxWg/1NGXv559EyY
FwV/z+tFPCSJhkUar5i6TOussTJIOikR+sl4xen7Jfj1ZWgEFRymy7cYdMFwzRZZLbYa7PVH9JQv
IJ/8VYQB95wsxYhBiPVGOVydo/dlIZ0mLfBB2a0jTbE+r/GKT0kW1fysZo18FfvmBDrwP6zbd/7g
ZT6Di6d+HuACoAL/eQ9DWjtlN+cKWVbgaWSN3p5a3hUpvjxRGklpI8JxZjbOYzThYnL7C8znp5I8
1aITu0ZBCTex7WVeml+GkptIirNFaXIjI5I0ABq7Ffg6QbNqEznLcdCZcNmad2+pZqcxEdlWCAO9
YP5S63kXbqBsY9cj/CufOQtpCp1PD3lP9+Y0KuhyQQAbpz9KvZ2xDJfMmI+bgJqKTg/OamVJGVOL
iU7I+3JF6MqvuEtBWG4bgk/pUtSl09r4heFVlpK9qJtvaMHUXOQa7/dkHFuIdNpUqOqf0EDrRSZT
eINP0Qij/DvQV7y5ks0DQoIE6XQvdKa9ZaXtA3X5RkR+dCDAeVlttjQnLt6/9KSi+rJLcRMG7EH2
8ZZj/9I+L5pE9hSQTygIXe8XKJIUpcma9Ql9UKboLeYEnmJmwfLlWbMNeN13gFBWfClkrzlq+jPG
yL3WWwVKPUWcc8m2f6uiywl91oo78VSTobsmfmt0QTNd7vL7iGVAYwWW1PT5oxVHxk2P365mSYQQ
ySF6lVBiKiwArEExk90PNNxFhxHaoMomJh+dU2UWO14HetnXcKvurBNyoRGwcVQSmNjcSD+PA0bt
KrZjaBps/jUfUAeszrNOiCs9JAOWq+iN7O0Vdp4sCa0U8qt7u+cllGAyheKH3RH8Ku0tv/OO7uQK
XXiArSrhjDp64zY99vtFwHTIQB5KBx/oRmftiAVkfT8GDR2wNtxweX66eZQV4iQsoIGhV8yLzvt7
GEeuVwl204PPRbqgIPlBfdEL4CdbybM095Z64FTLFKLkaOPeui2SLKtH2xXvMP8zC1KhFtug7GWq
4sibwRWtb+bSr4ndNBtAb04eqRmKMVkq+PZHeuCn3c0eZuzjhMlN66KV11Hms7TOy/8YNpUlU/Vv
ofKzA8y3q9uUba4A55kFh7qSw2TZec1C0w/khf0utcDEgFoMCqdtdXAQ0z4/KoCNk+Ig6TWEX2QQ
ZCjQ//Utjv9GaNOI2mYZsTg8Xqeh0vOINXPj8pQYh0Q3igw+qwNszHQl2x64mSxQQOL/1T8Ms6fe
PegI77hTvIL5ZF6qWFxI3WWutVF5mrobpZViDnfylFiqWr1TlcGIHenikZHd6qmpnAgB87PBkrTF
640Zs+n69fv7/ILJTNLACXJS2JvRqlB1pYMNzjqyZAZzgOhR2DQ40k62UPopnIYEkZ1KHjSbUTP1
TrLwIgXMRv09efSKbfyvSIufxILRkymfx1MZ0tUxbaGU29s06qaxflkSVGg3F0FJOsrEY+DQb9Z5
1pwC5sLsSb044wAwXCK0iDqgj+LCH9LU6vM1QrqBYR7N69dwyZTkIGA9nO8fQGgGMMo/5F5s1Zo3
jNtTNC/OkrNI8at7bOKwDO2fFKFHZzyw7O3e2SqaswVS6e8VaJozq3eJ9+TMVEkGEFWXhiOmwwze
c0/U8BpSRr6F8hQjIFox14/u7muQBh+NDkKREuv+R3sqhbx6kon+JIDVsTBt+CVtmDiY4UvzF3f2
2uIDKXJb383VWOtfEH6e2L6CluL2BpyZzwaymmzAZXlYy4ABQGzT8PaqPQGwz5H3q/v/zBEaTki1
CuD8GqdGSyOpPmjqi1QWskNiEYiV6GfQq82vwvTiFcaD6g0dozVfbRBkIo1inJns4O/7su58La9U
xSyiYFjM18Psmndn5UFytNxvaOBk+i+iQtN4JDgvAY1grPKeYDNJAyxMx3khXraE750e62iFBhWe
e529iNoli7XQkkQEH5j6VJw4OQ8YYMQ7lkXU2XkWYiWe3Uf6Qmq1V0jBp05Pf+WwnAmBP4zSJEo8
ukEUKK4hVFANEmgnNxDWDS9+JK+EzbwzyuZL+K/4JBRrmvSWw+SuImWd+jjzLEqjAxNUrePAw1Sc
1+nlvFH5CJl94v3kjg9+evE/PLgIHFRhMl7xFDXlWoynzpZwRWwXD87vaoyOTqs+aofZxb5boA3h
XEUTpHrgdj5A+SxY2TzsLS+Cc2RyptVVVXRnROX2f70CdITGP6HTi7W/LmIe/PhLb43WrMzI6D/n
RtdD0/bIeGNVmJ1RBg/ZErLyXshVJv9cR7z7+70oP779YBWK1Uq21qYOYtknrqOuxy2W78ai6/GK
eTMaTxHpXWiFIMJbW1bA/KJNlsRyYMNOe2mpgHHrOSbMnS6dQjtzuc0meipf/dzUwsXc04M3u8zW
xTT0Zm4FWpEMQVgyq5x8/+q9BoMKI4cr9U4vPigej/oPK76nvp+kNasdJvd80lo3zwpNJuWAcLZ7
uBuWTJqAWBgjVzyp7thacsnCTPKUaQt6c83gAGt3TsG1v9EDsG1IlHrkKuNBuyvBW7R9l1Z3LZ4s
lmwQWZxBxU4nF9LvfvlNCoMrVy4+kD6gVt7uyeazrSX4qLxmtcUIntn5kiEyrhwTccigss/WpZcp
E/m9ieqQYY6mPF0orVin86D7+mv9K1wsT5SWa6um8BmaeJnMugqwnzKweCBdJ9dxgDnWrxN8K8f6
lG3EDpsA6wEHNyLlybDKFkfjuuHepCSrN1vufBagFjrAKAjNu5o1CRfdHyGJ+4cM/tc3TugGZwiH
2lSYpCw30nPtP7lxlYIvgp/ryYCZD9lxVHZ6vKiiCcGBocmSyPMpIalwG19QMUbav5fY5+beLydK
p7Ws3QYnqA119G0iePjp0tN9ONztq2KeU73frgQqV7f7y1/1Wxz7Ry1EjsUth9rq0t7C1Yt9Er2Q
97uVdDyMIcN0oMeExW/BN6lUjH8FRuje37AxY82LsxQKAYPCmfEZRh8QiyZCTO2lbis8LP3GDlPJ
Rgx14HXuRpeYMpX0Y/82WxGwJ3lxw45XZeL8+ufasTtyAyQZnTRPx26QnP4jGsfMcJHiPzGRsds9
nxZHwl10SW8ft1vtR4bJIQZcSo8awcaE/JMGWvzFKsmiLhN7mke5fqgiFa4ETJ4nSViZNBoLeI6v
mIyCKe5LAsupsyzGrL9MyJCAEV1GfhLD3NLdXyNfaZ7HD0ri7vIvcwe4VNcfYQHZifXSlPSDQws/
lSW73YXzbKBktGx3hsPpJXm+bjYAjh1hvhd2NDqQ2KLT/oA4nv7an3tEWDn4FaGwV3VRYJJ0suUU
Jj7+iX2rfVmUnFUxiJJLyOl3FCFD8amdai/3eVjsnhfviGlgMA9iSJcpOkhWzdr8HWiYcAOW3bTF
y1VKCzwSvmSqrh1bM0TzSjfAOJpkTX82v2Nbc0HnlH92Vfl+KsfH5N0AORaoxxgB7vaDM3VYHHRb
yF2sWwyOC3NE0z0IglZOeMpSzhevz4r5LkSDv1IsODNqi5hMiMiR+c95oIZw7V/n7W7VhVYkjSmP
KB1CtmmL+UkTNVtgqj4v7CLE0xzS2WN5Z8/XZJtgxeTjEKauMOvsVQ77i+BgjW+8USMiq1lV2voV
BkuHhD40/E+MekJy98/8ReAJlw4vB2F/M9fZNosrTsig5/3L2DxLZAfGUQdiBpcfzlescbVAPUMH
sjO5aoKmU3fjHCWuILDhNfOq+ox1BymyVvHpaeWKImxQ4bZWnKNPzLtrNFMirJQYJlhn5qVBTiAn
nAcSvZZU7X1DDVrsaVmhhLpelrZBz091HZD6Rmh4yhbEBQcKfK0Uj6H6C6Feb14mlJGcNxxL5i6Q
8qmmVp3MC+aj4xQPz8+cAJxVjv92nPDt/Wo8xpeF/NjfTtcTgj1i4a5expuze7Ui0MyIj5mdGivQ
yPMFBV9NB2o1sTOhW7N758UR6PwLmG1DsS58Fs9lg/2Rx3siDs9D/GgCYi82RMq6ZEVnsTqd6K4N
2j32LJV2+6JoIRLRMTMovFMRyr3cm4o6QqY663Wv1uiMpYCriKgQO50f+oTvv9rVJvtQ8whOqxua
c666r88edEmP9Fwx11dqCtSfa2TciKXN3btenV5pv6HZUDa+AglCWZmiigiDsFhAxxEUSg4/CD6D
SJTlHdtsrosktnuk87+WhA/HmHmdJ73ikGk02kdMD6mOh7DpEBCf4RU7TT04OidpEF48lovY1Aff
qkMiSezcVVouG6Wo4uxQHVlkjwQnjTOqnNciDLhfyhO/etPFeN/9Xm6wR8ZX+QSzz+6n0/NAaHeh
Q+AudsZPHkNyB43acTM2So8Y7k3pyrUGrOBpZvHGXcuuC2620mMdymgGbghGf5jFV4IyUZ8sLBoI
qj0ssHE3meW/SBHehJfuAk4qPdMtAO7Cds+yTV4Pl5T6Qaza/qu/xZoJ17rTs01EZ/ubAYCZfxyM
4xOs9Vu1O5cuGh7Y6iUKmHiyA+j014JXPwzu11qOpJLlf5/Uw69rbwLwzXJ44rN7h+ujs+3nR9hQ
E/tBdZcMGBopeS1AAKCAnA5vgTW8nRik2CvasM0l+U2mZdRlDiePA61gNBZDzKkPjYj9rp214/1D
i+h3sfPOd6yn5PwodM1RcFRjzUgiqPHpK3IlRMsKCGgEX0hLugFTlfiChN26zKTSclVXs/7pvv10
nuBVY0Wyjtq8gviifmcA2glnH31DCKyeLfqfZeiPFqOhFh/e7b2ClQ2mHsC8d0RB+vcwPI0EP4Yo
rEEAYmj+BrBgvdw1RTpghqYLa4wc2Ug/aJJteEUzcONGvhB/Lj9t0lR9/WAvWixOZmdVmrX5NjFl
19/wfaWJoPddU5m1q0Jp+IPeannKIm2L4wW3/kBtKLWuxrn2eMNaFXj//lmAJzINfBi9Jjnj94H1
oL/5x1e0tBTHWmwwGm5hByCJ0n1IHHFpoUVfMSoe55I1KPmRWXlK+l/tOZcMYo9JM2a1yLGOjhWX
8rY/qtXMi+xuL3j8O8uWBiPPcVzLRUtn0vaNkOgbbmAEGCiLVP9IhweWEL0TbT98WLZSshCkt9Y6
J9E52MdDyOln2Cd/juDkGi/haZkKj6Q4TJbTRj46twz6Xzmf31NCaiipizMrKMlUaw1v6eRyFFwt
Uyzq8uEJGxtH4Rjh1zorEHJaQze++jyryDysWVKl/NLaXNPJB4BGoehFOBNqQw1HT3Et3FEpD+D5
6Ggxb/3Fb2fegyUAYQa9LSuUtQPLt0VsRYOKC8aIF/6YqxVTMEXwOAcqydwBXzkYinO1x5YzyiFM
nRTPGEFDbl1MuZv4S9rMqv7fBHE/sbrcmB5bzwht7xKa5z3osloTEzoKi05N0qOiD60KIewE11iY
t0kQOnMN+TNdTollYAKmoWS29cj/lotM9R0OzAVsxwv/T06L8l2PGt50484yilPbrEwrcqO/myrb
wiHKz1h09vdf90SFxW7jENMsPjisYZpQUF7Hptdl5j13cJ5lnswVrRrzz56uHkuAa3g99bFcprJf
J3D6km7aAcDwAO+7TcGW3PT7ZFmjCJmGKqVtn5Vt8YgGYreWeKgR8cVx7H1UmeNcQT5saeNAfOFW
+6+2rGkelU0enOHD0D5NXDgOD1h5
`pragma protect end_protected
