// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
iUiSi7HW/ZezEhcW1aYp1SC9CDLIWJmStpnp4106y8mxKlDS/B85lbO8KEtGPz+9HH0ZWSJrJ1Ah
ekaacT6l7qu6VNKUFzqV2PR3/X+srupDfSRZRjl7WIXdcQ+X1RxKVGuFw9oBKVkFAvftuHljcziB
eI+P+IDFP+7AdzDqytteYCORezo94R5jZRLeh4y1e6XNDea4GZJS0qgZl3c/98nPy2LV6WsKIxUs
bU2I9+ztZrm5BRY4gnBrJsEOeEP0azHrXIm7Qq14DcaYyE1K7mc8lpCShO0rvUwXytHYrKaxWI53
cTFp9Y/RyLwTKuA76zu0Y420DI6J0vIOfTytJw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14912)
UtniuKwpdinPxFYym/8LdAqLzFeA23A+xltGJD+/M3eTrfoPe+349UrhJHIgM4treRZZQN6R3Y+p
8v0LxeAR3CKxAhCOzK+H9ZYvvqzKKShJKv1yOKwxng8awNbHK9YtpTzb2D3upCmNuCWqCPnkjKOZ
E+f9yRIMcNT9uDrF+4cGgJ8hj5KhnW6f3Bg3aHASf1bdjr/u+UXOHDxiOI3lswqN6o9lfYdpC0JL
wU4ufrZQqWc344MdPRuiJ3wbkBp3CtfjbKUfBRXY4DNrbM4S9pthNEpgDEIeOy0CZCOjzz+xSY83
/dcc0Ib+CCAh/FmQNaMOuiRk6dcxO2BJuq+Xz88YMk8Gj8gLk1tDP4PKhD5stYYeBP/fYsqjSO+I
erd/jiW7vh6Gagl/hgjiI6pQ/j38d4aKyxGgD2Ja5OVUsZmzQDiAAWHOV4oLD08Kw5pUS06ZXs9t
IdyZwNfYVUP7MlU6RxvQTQSbfUkuAs0GkgC7+AsprnwMFWJ4OWXtlvK/eALzPLxBKPrci+H52Bb4
ay2rMrSL6bDpyxLoUYRvBcYjenretiX3XwS3gvV3sJEVbLC08K10NZ6bz7n5X0qDfg/c8JH/Qi2n
2pIsOKkhrOvKb6jXN6T0Vvq+W9BIxIVBrQtIr/ZoBfPeBiPhaYqwb76QDXZH0kBjkDNfy37NCOQ5
jsUD5siS+eWT59c4d1+wZHiAu97fzSRSrG0vffIXWnPEk59e6xF5FGgKafMqylkQ0xcVDxsIkeyA
Mnw2g74ImGxc53c7kM5dBadE6lTrBjbksD5OVxYjgqKQX9APTA59tZ+4SFTyeYOeIKyD/2tT2mFa
zQbiGKg5y/dQeTlMESVlG8LGdzWrAhh7oWoRKnx0Dt02RfYWcwEHSvIoTxd1aZdoHLYf6Lw7oFdL
gc9C9gUP6mInnHPoRy4r33k4kJnYi5FKWCSVMRU8Q1XIe6/0C4TQtWbD5QS/jxzVu8TKBYp3pHzg
V4mNbdOSZu8JRiffrGmh0gq6cTU+VjZ/xbB4cNFmoGcTuZAqsuHE11w4YiMk5WaQt3xh+UFxUUWG
5X0/6VBrOUWnGLYNknZiSPDCkbUUUkxvGrhjauEkrpezwERRgMvX6Gf+INdutEDXoJ6ou/ZLMAtL
l2/DVFiyAFMlqbawSKViLghU0WydTtHn5wPjPIi79WLheBahAfswkyqu8VrmI52eSMGWRQeve8pQ
OsSPV2G2vRve2RkXyMwNfhAfA61x+QimuXXt/s/XYBzot27TTaGKmq17KO4kVod5+EzrjKTlNgBY
SQ3G+xRpnHpVPbloYKCVkv69gWNU4zrbmWU9O7QjlKxbVXTe6bEUTCTzgk3nqFzq3exPsZY+5LsE
ff2nKzmWHGcXGhKldUaOMPrYwsTbajbv7jYHBSCgnskX0T2NMrizdePG1hS7kf4LYKYSrIfIpMUz
QaX2QyRYZVC9cFgpn3brDCunY2r1niq32AWa2dYs5oWxWRVSsriULjUwtfr2vYKwtBKV3Kzt9YKt
tOWhOB8xZ26qGNhiWnvIgXfd9ANa383r0Q47BRQpPfUU1vxBZ8L/O2A2Y8KpepGK/gh7tWOBXOul
oZ/rVWItVjXVs/GREBO/lP7pC3qjVXP1vy8bNqkEf6u3V8kMa1lzE0J0LgftSHvqJbUo9vgyCTn1
TxieSFMfu4bJ11IhjUVrEEC7s0TdhR9V4iaMecd8RCtDTs4ovk7lG6v2zFeyRYqGdzapoF35O0uX
jRISzG0LXWXtfh+gK0edslti6aoSBMsO1zWpp+aD78gzMuSYKtOHd4IR1AdaS/OxZ0O3K6TWGwyG
k786L28Hzse+szek+eppLDvAR6Bp7t3TQ0WUlqqw+UCCjPyM3ne03z8G/wnflJVGYrUrmOt91J90
SMOwGp0dnGR4v0DhUCTHRiVHVC1QaSM/H5lxG4aqoNki27aUaiFWgQGkSgf6UpbgkEMw6PdJi5Ea
asV3Afy/uwi9BiEiUOW6xCkXtFsYIsZ/MIafy/j+zo9LwqBHRRqyrNsHwSLVsu0thE93IhPBZDzf
8SIGzgtN79PO9SodPbfNN/YEG16krI3tbkFCYVxeZFMLL+whNRabDcbT5lK9DWwGEtNL9LpBgHup
KWHyAAeZ0WCWDKFhe8mTXfmrhum2S+1JZlEjQou8nXUc7G1VPOYp3qBm70Pc0+NuFNUD1Vmz1Frr
0aE8d2OH48ib6X6OVgr/dDJOJaTeuKymlGTeUUBIVrtqVwqQmg/QApIlc8aPVhTia5rsgZ+olHxv
+p30FSFUmL1VNDGh+2QbbcR7YjBwA9dAwfSrsG4hD2V6gk4kxngwNeZlOJgcpn8Xz4TURbT10VBr
vWVq9S5TOFcF/zagBjrcJGReJfM8Jzzu/3huKGkrJA3eutngc136e1Ckb4/e+GfXqwTjIGFXxCcs
0SJ6YlrFBTSVh0PpavQFULPZV9D/fDYeQNxkyKHj9X3yhpcAvUZ9lg9wUsBXB6UKfii/KJ0sEzTi
8XrfMMufRaJWxOtUj2/OU+tru6NACymxoHtGBuDn+qUPbFQJkfvg3co5DxDJV0kver4HmONcQua5
tTifxqhxh++gdYFJ+O+RH6KWv+X32GDR30ldpDXm+/UzUAR+yK76fKq6f119Ee729vIvlD4SpQGt
n/c9hCZAGN/U1Zht8WeqnUXDI1ghl6GkJwIlVbXrwjT5Mls8emgeYtbxqOVUShmzhh6LNK7VG3LA
cN8ig6LXGHHDzmS19SWE4f+Gmrq9je2HAWHqs7SQMDH1hZkz0w5VrpK81BIfD9otW9Me6H+hfqs4
86mHbEShjKYjEcr+vJYax6Cbs8HYmcDCiu/hyKZ4qmJvtbD0PrH0v87S371cnnve8UIyRFFeMezE
D/nCRzkiOHF2x9QM8RarEvrdjeD6jl1ys/KJYjaw9F0HGLnAu64LpCD1tX2YkJRQ2Ha6C7aKe9iY
bc389zZ6e3iqmXwKpHkzQNNdiR1cCXpvPkTkWozKpU4Mny33ifE2oQXj7S9YZ1uP3g0Kc4+Mo3Pt
o3ncqomAqCTkF1hXYQKO1nye2hO+wp6RUU1FqnQ1zJMx7Xc/X/WddBnDZmlLHgmTkfb8V+lbcuZz
hwJZ65jJSJcnF14cx7+FqUstlwfvwcjaf9ovAJOpHqS3YHOu/Tlhwg24mWCnyYFbYalRC30cUecs
gMCc+L4Dwn0ZKadu6qxLPCDyAvN7y+3hI2F/UHtsCwKWxJVQE7raUuVlm3+flgX0mDXWAsqS7KYV
gUUNce4FvaBNcR4n9xFK9RoDmhwC0bmy4yt2macqi51xXwiK4SMR9uhDxpcLQHK5Rk+1GCLn2fb1
yM8fTiw1DPTQ0n3hRydX4pgGVTvu6dUTrYctfOlhRT1SFhubw6kJitwBy33YLFuxuksqZiflxu2u
j3O1NW/4URd6gFi6JWWZBknq7lVeiWkUPdauZRo56mLeCEiAO1eAijK2Vdox7zh/aa9m/tFDdlt9
+f2duKy09F34oEzU66hB9UIWnGvUNNBJ+d44Dttya0u+bqL4da0llcrqsfzZUnDEdFOaG3wbtnjG
2I0zMtG6KZuf5qszUvKSfUIOa09ucRDEXJxoHTTM2SwKZHTWd8GEgiF+hC3WpRXvMggdFvxvjfRS
Sc+hca6m+sLpeOtdAFrJ+fm3piX4HygXSr6hIkDgzMxpZbbTwjgm9b7ZTVpJfj6XF5Iq0zDnDXxR
sp7/Eq+IYfbg65OuOBV8Wjbr++2R0G5nkURzbp6Dqo3GK91QJWXcNnAoCZ4es20Nq4ZNvQmjqNsv
EmHoVG8kV1p9syWJkhcsE0yBOjNypKcX/zwMMRuV/NwEmr9EANksJpG3Tw+0ERYADq4+1xwRjEqM
NMsjWui0CiwfobxSPTQgq9ekz8uc04V1YLkdhKLerVkXtUxGsovouQIGPu69l8LpCceMQQAOiJKG
sPl0Ma7ix2ArAOtGIZaYAhLeyoijWnmR/YyYHYnBbekvSSvEi1/9pVJXbx4ZoGmQOl4RjOez4uUS
stzo7zDRNPpIykJw1C35cv+Wd0q/QQYI59KJ4K7hLLz11ysiDCvu4R9lHackIZU+LSxS9sjtRlwl
PLB7SNA3ZwbvlU1YVDEQHbthyKIwA9YLLL+fctrv+Rm4dDlj9fZ5E8Ou53XVAQ/T/LMAmRAWXK+r
g2w+d3+zYveklAtK3QZIoCp23gaChHgpzvniskatCmT5xsyn28NprR/wPPGwuRR6fRYjfbjGqBnc
bTViaal0J39WQwVpk4v5Xr4Amrcm4vWwmizCY8sipdFToroXHKYPmkMlNnTHXCJS4ryPAmMLj1Lm
KqK/Wnr7uj8W/P0QONly466Brw9VKGPlRK+237xkfnU/ePrxiWBfXKhn+RABBi9jC+56RpdC95J8
WWzzAtAcaXfOaibt5aLlwOkRCk0TXNpwdceb7Z1tHT2ocB1HO4Ifmq7SpbSf3K0YovNnYql7iHEG
sjLyRR4Ho/sD1sI2HVdupAexVsdVLdQ57fdX+r2ghhKpzLADneNa6KVmHkoNbpkG9GX2UmRxf0ln
/EzF/3qyPghSS5X8gM8+Gk3de/cqTxnNSS44H9b6TFrTPKpy57Gsg2apdZBsimIbZaS84B7oyIEA
XwZKX18ZEgeDrk9Okmkma7NO7kmj17O3FYL/8nQqWOapsN+dohlfr8g4xnrajXycavnqc/hpGyXn
QhXLBsTlIff6XjBG0/0wNSSv54Cihpylm1FxD+9V9n42LCXOI8kwhvtgdj8dvWEngrEVA3WX2+fn
g3By9CIsV4D6oxAXFtnJZfGsfYzcZoWtXf8m23pfXK3LPJhe+qCsIR/gThtiSEFKi07Hs3YMwcrj
yruMnvFMPFcWNOhOHW527tx3I1hFHAdcCWPgS0CWIJm9fp9KDUpTEQvWjwWu6v/LUZhlcX6gREoq
RIGlMS9ks34I8X/71En4fiUAFV/lq474guNN16xl00dr/WOtyTh3FCZBHe/O8gFUD5iceeaOFK9u
E8lXQROr1OyfbgBCan7OUid32umJ8pf34NHGiWJiRbcvWXHAQojPkCpU/cBtWUmIlGoaN/6/P/dN
dmQq//YSLT/gBtbefWmDwEk8ORIU0FxQMLFZt1mG9uJEprTWsyp62fYxXW3cOhcUupodacygwa+9
utexDqR1Du9pi1a0X/tMvUcLUDwYgefvDu7DizfN1B4pLA0v5Ljv0K83NzDgBN4PX4e6kvvXtDUO
xGzB2xI2H3rbq6nyl7BPvl22czBfbH2m8yUyIuqaAggAs/ZhUceZ68D+grScPOJQfHSQ0heB9PhL
api6imVbpSESCiNHNoPtTnoGcqF9l96aFF46P6q8VQ2oP3aoQQm+Nova5nHO0SDUpDu7AspOf/3d
TzvfmruQJhjhqbqEzIJv/1p8CSD4yVZJ+r1gHcZvLRqs3/PXbSCBvTRHuuIIs4YbZEJI4lq92iJZ
61F0g1jOU/LUQam3shH5asGeVNR8WpPGVBtcUn4AbZArLvQu5bvseX1Cs+xVE9ulcAXfcWBKFmAz
CeQwsE39RV3WsoOEUzhdK2SJrAuKL3xTk54qA+1BLvWHh1I1Bnn1+cH4FWNL54UFpv+pRyGRZd5s
uMqBJCym+WsFjqb34xJm8iHhnaGGc8VY6yEhkD2dbigW69P+yaD4fx2SYLYWZr29pA9j7fYxp2RU
d3+GmogQIPoVWRqegsbZocBT6755QeJ9EgmsO3HmpRgcqXMy2yyfqmXIVk3uf8VAqwTOs2kexUL1
MFS7nCfcS6j0PWP+iRQdSZ6Y2S/JPu8vog+vofXiZf4L/G4k9EgJBbfkgnpRuiDIhmDK/CH8BFLh
OurRruhZqeui9u8HM0sju+o0GXioj2442SZygZOLrqtNEpPWn5jCWGmxzgbNuBQDRokzUm8p9h/w
pb9Zzyi2lkKBQqCDSzZoBrs/aL8ggIfY5K/uS92EvOZ7j3Fy3hqHTcTWsMYlsUdhoRHe2kamW5D/
7yr1oIoXHqsFChKhJSv4tz5FBNBACMsdcQJgcKPk7zQgtV7lZyIPetQbouBsew9QkkUpTDZ0d7hH
KN4fwkWUaBY/oJgZkvEdUf/7SnqExly5OAmbubnyaHF7WuVcWB4fNX0xEqHQ72xY8AhxY0Lgvtx5
ZEaqszaLzcanW9/NRYoRXHD86N9pAzs7JOZghYmjYCCop+vcw7v9ijHbSBZcjAjPRlo48Nlf6pVG
FG7ntX3cx45ixBDfYQsbIaOFayBihBQr+ZKcCoJPOA182em5doB1Y1dYqBq+ecQBzCWV1FUfC2YW
SHIeqb1q6+89j9xdqsbpnNTS1Df7zu5gyFpJof0MywGjJwE5CX2LEC+35e+lVHR09QNcLcFf6UKH
kwiWMihiGC5PlDYSZj7suEIp2CH6YSgy3povtvJ2gJlv0Dn7CYA/8CTMd3nGnWjWiiQCi6skFhhP
HluCEljffPJ8kQSJNAuVLaL2wajChRF0zJwCn6vVYzpnnhbpTEbudPq2lq05PJDum1GhuXxDmR4l
OuTRCuS9BBbLdSxwEU66icFvebRCeS3pNgHQcbFrv7XQOAanBT+2Kv0w9kVq/LM0SGAqoeb2e7lf
8OKTR28g7SK2Vk9Vzo4/zOHr6LeNyMGU6vQtfDlDC/0PHSlf1Lr7WG3m7dLqzYOhyFEKwTSHQ/ve
XRvbB78Blz+E1HtaBIRuo7Lng/tiGCGEuhHhUHU52fWbG+JdilqjCHi8yi67YqpI0OmzQ+N86TgY
0OHCo0MJ4GBJKjG/X4NBLpEk4etEkQ2guZTU3bGvhIs2zjzN4VlTH/A2TfzBXq4J9IzIBrWVfmwk
WRu0ldx17k+maRtQEGupRSa8Pwy67jSfjytRzLhA6b6lEAj7uooWcI86k0vJb1KZVmViN2Dmvvq2
7ncVxkH4hog1OqWO+FTjgEH9YKJEec11nRNMpZPXFliup+qqk428sCtQmjnV9g4/lJ4AuUJe/mlN
/k33eYubDIAE3vZNT2FeGRToYzgeTwsjw6hJK2dasrhMqbEie4JkN07eAOPnES2Jy8LQt/mVhpxu
gUm8tBNTi5/QhygWs9siiwbJPHbHeC3SNHtLUzXvbGeUDzDvG6ssoynmbQoC0p7uoRJfor1qerET
b/B97Laz0Tu8yqirkIk1f/MZKlv38PWFsARtmm/P6Gy4/d9Npx6Sjs6u58xrsh25uwJDHY34s9Yl
w7uAE7XuQEagE2ZZOyquqn3nQgNMbqqq+reM0afh/Uw8pvUy+geUFoHHvoA0gesTt8CvH72a86Jz
KWb1tgNFvCfEuGtIztzT9MdVKxA/XRiMxOGK+GBaz4mylV6QPJjZD0gKSeBtuW1Py6qYwYpM69B7
3f75nLjHWPeNc7WnV6RzAGFu1Re7eF69QE686W8zlBdP70jMfGZOTMP0md/ok08ohrDT0//4IZ1h
lVswQmyEpONLfsxWkMDC5SnBi3DIx6593cExFrRvzpB5oSWYwdbeq8kTkm+rVb4o/KFpemuHqSYS
xi79K/JxS6gCPW0nTNXVgrqQD7E7eogDO2oGOevVXqS9yRn+e0FCxxd8jYfHY6zONYYj9DzrALm0
F9ul9Fl17o2LeGDD4kikZxEu/yvREto7IevJcEhE6tulUtz5jbQrK7GdelbJLEVLhMzacpq8RvVF
lbzEmXN7t2vxAWRj1A87Gs2BSa8tyCwg47p5Mbj9lFF99ayE8v9792wwY/V8exGDW7SNmTvsiSZE
3o0ujz0j36/urJ0i3oWQxkF3oT2W+rKxp6gFBKaBv9veOaeEgqgcK1OgXtquk2j3oDHQzuVopLnw
yzdoRMr1QI3wGIDgjkxhkGjI7CdxPh/t/ut4O082VKI3PxJLgM+uBscvusq4v6n95ldrIIIrVrEU
rgXkjzfKqq2yqi/eD44dNUMJwrAhLNC2RmvWkreKtPJsCvzgcMyR/qiYJPQHuj4NEOj8P6/m8yNc
H9qcNOtYJ/gdR/ZJRoAace+NLVZTI02C8cKrWEAGc5JvR7YFnUCXJDNNF5L1JO6O6cLk7xBjZ5d7
1w9G4ev9hXfP/9yuN7R8UT/iZJkZVStwFgTVSY64FRdizzLELjVlyq+XVmGjqqz8X1IOYKGx42sI
Kcp10L/DEr11yVxJcnv50eYQewGg+BbMgF5t5c19GeSQ4mmNC5OX4hzYQvcOWVfbBBI+UWeD/HQU
a0k5n/LmnacRoHK+66XilC2K4BsGvUIwHlnF0pf0JS59JhyzM1Kln9WGpMrbfAc65cijpyKeBi41
vOC0Z9RlFoBSQw0hpcR0y4PBwZG9MnoyE9yZFyVIkm6tJ8USfNmkkALOKtRihYORggrSUcqD3bog
wXEgKHkEgOXFd1VvkbUi2H0y7/c3SIGIU7mRy/EUGG7LcYS3oTJX6UYDL201P2dphFeIlcnhkttt
854z7+tsBR1hnMkinCo3b4NR+v4XbkmZDy6WKr46dlrRigKPYC16ApeXxvfz+rnSbCGkCvd6azRf
773zJO7Cd1wCIdd+AeqjATIschUy2bubFHybZ9UXWE++jRcQZ/ZOkT4FcrWbkuPqfavPgP8TTpnu
+3Ge2OZ8wgVmVEOPXncKOmXUPfVg2MSCqhmJPtK44yQVN8GWOjn622ocyzCGcK9C3FPqhhG+SasV
IT3QKa2oxgczZ/kp03UPxbWUWjI8sz4p60TfCT343O4bqgordQF/OtZVCo+EMscvXGNpnZXP+L4k
JyWswBdWsE6jVJg6Bh0Afh3sQHTUKcxUcU9rhwAe0LWGgp9uPaDL39SQC/F1y56USsLt0leQtvGS
uZubF6fEYZukIi0ZAL2zTibMxa3SY3JlhXhPLhdY6V3m+A9nNY47e+PDoMgHs3jfHK9kvmGArrOy
xZLqh61cojVEcWqTe2/6267oR/CjlNkCVWikX1f6P7yx8ww7njODu/tx1hYgYxT9K7RZ6UFydCZw
3P5HT2M+cbyvg2NA0qc9NLROQYz/LY0Z9ihvnIfkncA9kEeUurNdMdj0WI/Fqw2XiMQ7OAX0YyRL
7FVZlqkL8ceNfijuNaEKHIrKZwGo6S/VH5iNtBB4dex7wOjtW9yjZ/t+qr3y3k6xBkkaCWwDMP2X
cO8jsclRG9IcMrgvpM2jXG0dGVUCpJzn3TIDZ18ySIjfInpRJCFF7BckNIGRuJ09GRhW0V1Fnt1Y
fFt6BEW4cNBJf8+wyVlMa30pFC4vGUqGtzDo3SbQee6x37gNwg9qNiEEqqDArecsTna7aEhwhWkA
FdBUUAmjfDhkmntL1Ns/0FyjR64+hIPJXjLzkRn78Kp8DSd4JmQhbKFFd0n24ReeFn/JIXQukn2y
Yn6gMhIuADDl1TX0McJLAovGR7LWGed9joZwV6NtlIEGUXk1bSWSzwJVCstbUDIqHz+soZrpu2A3
tZwJWvcg1atsZwDLWRwgUULWaE2/JL1GqCQG6JkzKfyCLF89Di231dCAl7G+pJwShFYdX7TSESyt
QiKNh4yzkavxhfKvdiiO/C8ucONKkFYKta0/0OB02SSaOeQjv1d1AYLZcL/vTEvQ1fMT3CJXvHbM
8KgfneoNcwlU5HVWc7hripMJ3P7s+Tcl6mEE1tK8cMZ3ZnzhlG/oJ9CFK7ZLflpNN5TareBK8A0y
ERHDcxSGf5pLksXsqn+WbZFErQSJbyi1Gu/LtvWPWFqBgjH4Bcv3e8qzWxM2/t9/PAkbigg2JLq0
nbgrvZcwmIAeVWqNiL84IzfjaqJOYCu7W+IffXVjf0vi3xHutqQr4Zfd+YOUoDzPFL7xrdNwBV7F
3GXW0Ag+mSlZGO5h2itIURAsGSCWx7/YWub+QEHXWPW9Hxl8s+XSN8UwUcHEtuyE9HNfqigPQdxA
adcH44hMceOn33oEhm5/4UpdIoPRO46i5omL6xcjlHLFve8/og/LeESq55/Ob9Ho0xFgKh5718LK
wqqD89+Enf+lfplDXd7PfTnNh4/qaFVqC+gmR8AULriTTtwqQuIy8Ytjl+2PGEZyKZWdjRu69pQv
WX7DSPCWyS3Eknq4qjadHYQ6xDI/eR1x5e60YoKLKqk8a+itQrdJzDIpCPiUS9uBK7OPzR+lqll6
xfSZi/M/L48/rKxZDS4TiYDuVcAVHwnYuB3YB4xe7Kf7hzP5K8CIpra7Tn8ZhE60SDD7A6tJfwke
eU0Y1ZX/Qo0mHrZxaPP7P7RKn3O35MHSgExK6Lr/o0ws7BfJm8UNe4S3Kjwz+m1/sHVIhLfVs85x
7HLspNZzx/fmQ0jlkkGu4zkhWwl7+Pz9/JydPeAtfzeN9xN1xczMBTEp4aFY2TO9UxUw76x5WRbN
FTXOGg7OFgFQPNdSIZA2usO5txH4Ka8j6xqU7ghefJ2b7V0p17L9FJ1IZaPpXqN4OXMwmGV6y7Pz
RtzZIiwkiCiUrebHN+XXQ8Tk7dBXEdxVjzvw8fAKg0PgzTd1n5tR5gdJ3rUhVrlkDS1f7ApfzGi0
U03Ge6fG2rld2uZZE4QjAjm8q7Yw+2MopVfKiZZgLrg0F0ygc+l4qSC1CXt/b71SzKwalVubtk4P
VnUp6xncGksE8lZMrXt8hVmX0RxcwfSljYiyoDCjxmxNHOcHhDdL2rjksakgS5Lt96UX5DvSHEMa
/vuQl2MJLRg3n5UZHaUw8gQ1E/MyfxfyisgRQGiJphoet0/4ZPNTJ66o8FDSszZmAMy04vKP2/1G
Nn72SbpUqrTRNB0hPcrRQ4YwFhFCjH8kIIV8ob1kmifd/SLMK5eyvRqqQa/DyPdmMWZSN2+KleO6
zIdV7bXtngt2Owmxf2pbAH/rQMFLS5PfcMCubl1BZvYKCVnyp2EtH1cJPP33YMsxfhVACNO0/vd/
CLXrK1oAnGqtMPe4pQzPYpPbYnOwVnxDZ3Yk2ZdEDRRiUaOyINdjVEPUt4/2m6O6XtoHIX4Vo/dw
uhbYo38sMRqaXzrY2WZliLsAIxLWvaqLvm+PR9uQxJaKLTL5tdM7Jyjm0Q8SLtUlVWcdFdl499bn
rS120zh0jZrRIv62dP00LvQ51RuKhD8qXMh/FEbpCIrtj3XvpfHf1AtX3/yT0JMbVpo0eOs5WlEk
yXtEt2NoV9hcyiD+GlGslEqj6BcrtpU3eqii0FuDD4bFPH8vAZpiNeJOLsofu6Ub9w+YfFj1b27O
NTNXU45nIVwnpNQVk6VMbseLRlfnCvzrnz7oRsD8LptxjdytFM0fflND4NSRXSj5r8aoU4cJs6sC
aFhVyuZ7ZRlP2Hhz5ZaUoiBG4BGelaIbnw01g9ihvI85dPsh9b4pcyEMdlTfcCMOWXZMdjBtR13o
un1+7Pcs0I3DNeJU7kK7Bat/rBXNchz+B1tdpG1VF8jDHhQM0nQ4dfv5wBDt6sqrImw+GNEOkCBK
Hoc3x3KBvRAkz6M2cdDfvwmOuJyBLBlsOiqYjtSnTrQwnIBZPbi3uQTwP7FSz8zho/+ua2wSZqdV
w31d4lbWYZm9Ppd8o2ozTZ1O/VO3q/9lQu9/f6azsjYCeEWp0wu34sWgp7+mGsje5FK03kQe5ShE
Wwjot3YnAoaODeTt/6Sc16sExGNp8fHxmjNUNnaaMdiNm4fG5ihsgEDts5UdkY6SHA9NyXciIENI
bLdFblTCzIyS5Q9OQlQG5ydNxzCL/vbYbHPBp0HG8ivijXOj8mS0qK7fsplaE1acL9ahVcsKtSyW
4iOBFTiT0uISRwJDzg8kDQ6P0XSFgeW9tJ1K035/U21P1xAOtBvO/sydEkbJIiNgfgcmV3+aO1rE
6hbyS4XTKQ/6Woe7Rqfg4Yk9W6lJCPqowI5aECCQvLlWrUdlS0Zjv3PmqGdFF4f64Z2s3VJQ6nnF
LlhPY+xPYvHyNUmBqzMPH0pmnlmClguBBFKXP2/6e9vjeZLtINNwRiOAkOV3OPlucbnspdk0vcrW
pN297GLaJmHoy9aCnU5TLzMkP3U6xuv0TPwCXL7qicqbo4mJ2EkM5KXVD/Yd+QVXEEECKbiucu4c
Ox1Z5n5RHyArWywjOQExpqdGGOhTIT3gw2PZzAne9/BSEBK4zIh0IIK+Cit+K+D90zsQWmfhWVOJ
3FF2ZHUNN2U6CPi6kOY9uIDdZSNZMfrgVgB+I4P5WJ1mfbS/1aoRYw2gsFFol1xzEH1zzw+tOfmW
K8TGTjFxyeTzcOg7lWf5nJysfF3C+iB73w3Wqnfe9VWJCLXXzTgosK2+CQk0/VmmVUGSM9zgQRCB
NIWNaKUnfnWuvDO2X/ldYCQbcTd/GAGDs3UhGNojUG+uvIO6zXEZKbWlhzBbsmdbjx2+HKNgF+do
2jy5J0wRXAEwJLywrxVbZ7XC15brZIA8qwY3pfrkXiyLA7QvrL8zEW/pLt4eHX2HQ2hL0ZkpB/Ot
TgK6JTdjzFDtdSRLbt8gqhEJZQEe+Tglt+bikPITjIp48/Po1Cbz87Yzkq+00dDLsetgq9Vgw7HB
d8MnYf4+e75SoRZ9iihzOqUdSVA5r8PSC1pMRQNwmmctvR5ElFPQeH3AoMzEdnC7wpeeqz8gn+hf
xEil+gz5YpJeVsq8Y8hk7PeaFetHzAdoJjmCyzXY4t+3Q+I8/4yhzOrp5Le+0tQkvDMq0tFQ6nxP
LODCHWMO5NqQCqNQngaCSNCmq4+7bvpeWQqtZUlw6NOCGXLmeiDlFx11usS+2/LqchTwnAja0K9e
wSlpeiif4UFvPwWrSJ4Xtjk/G/CTzc/ryhlsRuPIUVfgY8nCS0RnR8Tz15mCnNOM8nHaBnoZs+tx
oe3bO1tjid5w5bg1NbhW/B9nkVO6kMqKOhLneOHT+Tdf3H/31TzswvnVC8MjjKqbSlo+nBui7+Gy
S4X3Dr5ZXlR8REz/43Se8f0crbYXMxstQROZFYtlL9T9AomD/b0FjZuz/o1Q98sgdrbMVtEgMjNE
aDwTtLDjSPVPbYBrt+uTzeUnEslgEltR96AxDjUxZTzIVRF+mLzE2cyVBvXz6/tiQt62rB+wfFrD
UxfRdtGm1VwghUQ7AwV+w3woVVDDpLLQODasD2MjgK+B4/yEdiu9FioXkMtaClBAK5NlMN+3AcyX
d/hGtWP79szpJDvY3nIGeto1KPjgztJRztupLDsFfH2DbQOUasTQMQy2VoUaIyMWMuTpTg6wtN7x
SigX9QtdoFkiin+niJdvwf+reuXW/szrnX10+FYoRMbgUzIuynOcUgNpjOHO6DMAfF+Us5y0NOQr
JG0ZzwA40zTHEyyiBMyEbMSDDkCmJHZ+Fii/uFCI2H+2x2LGxbqTFHqApi/zUTV0lEt/1ulLsNJV
9BGIDl8UThpxDK+aYUWJ3rbTAxVO73PwlDPvcdWOiy7UQU+UsWtSSF0yJRHcN6jwp8DnUEIvz3F2
U2RdBPTl9GfYuGGLGg7xs+PDMIphDuWwtgX+zr+2VqtqJCGu8dDZWRHmSOS5TInIVxWE2eB/qdA3
hT6X+rVwkNoLyq4/gPvlwfTDuk19X530idlBbcZK7RZ+TzS8P7C6nb+sf7miBkiKgocaw1ncglQ5
s3GBbdrHZnJPuM77sF8CCny+N2e2BgkxILUmeVkIllFfCIS7SRk+FhT9UYp8zvOM2bQelD4iAVOA
1BXLSmLTJAbSAJ1uhzOb4Iurz+tyH5gMz1tyBT4A0oBVVawSczZerjNgZPzvqLbXZHvmitP8l+Bl
f+RH4/qq/YKrlsJOdYST1nvJY63/AU4Km3mg1hxWLMRZGjYzg/YZBPBXe/54aiCe1FoAPaP4Fss4
KpnA3Jsxnydqt4lRBwYjAZbLJm48ayUQmlCCA0gXhbx1LKkL8nHtlJcnJI//Em/8ZGnee0HTcsdu
kb4w77nlRd65mAgTzl4Sr1H3VDdNtnBo0ABrR9laPfd7Cs3fDPTxMXUk/QmKPDrXU6brulOwtKre
//8gUf+hEWlKpj7aZMyEWhwISbgG8ddUcgPKdrd8QpMncV2OSQMTdWPxvtcQyno+jGs8E+LmrWjQ
W1/0vV0aTkozRGyWzQDJ2+cMUNIQKULK01X2mHnoPNYqdWHjZVxm9+aBfYiErUY8rTSoLsn+7nMW
qZp7h2q5a4UgfDMP7li9acIYdeyTCphJKZsBrVTxOUa/atKAWx2oZH42/6SfhSq8iH3LvdjXRQ+A
x1eHfhyZqrvPjiinorpdmQaa3EAZ8ijbJHi1rzG3xmX787PPPtVXSO1yOLblcWXpT0iQ3O/BG5x/
8r8bRTgpuc+ijWDi/Z1xFFsarjFqEuja5OXWGvWO2a1FKV2b9WQcsqzlY79aSeqwJ8DEeVMwMQgv
L/v6dcFF/s7aMnSn0mTzbCotbcUCEYuzec/NdIsFSXTwzllpXMJl795J7D/Wg1/HN662dKC14ccf
DoatvvUqSPhi5CEAlZgle6+qbwdtRyXlV4t7wl7kJLgXz5RvAWTV2URVxl/oD6d5Q+Oj57wM3jNi
eR7WAdjNuRWMZCoIdSlq01wUPCjYaTf+20FDo1GWD1THus80ynhJZOUvLPUP7jtpyYIlf+Na8cHb
8Cw2+piv7dtpvJIwWpnynC3Ze2ZqT5KrS4GWaitb4moFeYOUmHa3Q7PIQbiBXlw6z7etdIvnoWTR
V3bau/3FJGWkNhoQFU47QmE3Ar6EmhF9o6dUztgBBmlkWTiy55jbRkdfhx6pnMEnvXTDs35uyqBZ
N4GDkUz5bW8nJd5oKlus18Zk3Z+vj/8D4PxPd71biVfmVpImRT1MuttDUcYbFdXVaefsYT6d2aJF
zu6HDtrmU8TDu6VznXE/MrTnvm4nh56dEMtLzWQt3Lp/isZwCF2x85+026BwMNwmgqG5VPwa2STf
rogXFK9skvBGtOXA8Cfp4GWcFEvqW6vNpzXBO1xXzjqVquAdE7XW8W4zFYr6RSe4lzoBB0E9Pwi0
30AkGTt7BbTzvY2aJDecf7S5Tn/4mo1AY1Xaam6zdy7xHWpNYkfDs297uxippEXRaAemHzWHfBuw
DvddHvU/W6d3cbpWp6M2rhXzaYRWTwzudF1SoyPdL1heUEx5fY6YAkpFQG0zJPJVNp90Zf/KROU7
eOWhXKYYlwo++FCg13xTF3Ecfap9nfrC3M0hnltrGPfdmSFSymah9Db2Hrjng5fRDZn7aZpjRquq
hH3pxv4N+z7f/jBVlKBzvXTzH2RI7KmHxr7XUoYfTP4vFHOHUCns5U+iw5Xe6z2WgiiB4UA8KIzr
BhPJQ1cF2KSE9aytS84uvpw7NZbvAYRTbCewnd4dBLyEFaQT6U1q8sBoZxhvLYmR6/h1x4hn28kj
lfqOf4OvLwgQIJu37MaZ0wbvyPND1viOlVH8o4sLUq2SOGWBdLctiPVvh6uYX81wO1u0UafiHgIH
qs+3Z+dbZo6SqfixYINJPd/mOooRVZCSF9oIF30o3vjr8GZBD2ZONulME6Jlj5UEAE9UUh10qHh1
M7MMOOAMae9W5WIOJ1+uhrWvoebQFJ41S8Yn7jjy4zLKXEG34QigF/qcWmCn+FK6yFMda8zcpIL4
6mPphdUjKXCzzez3JAKPHoOHGKJBvbDXW5b/cJ8IXXgDUoG3zGRSJgmEriOxDj4c21vHaBhFBa7E
wMqRItiPJ60+XmndqcFgrwp8bKAudBGIKVnoIaXcl8HKgjDzTGScPvTpP3NPKnhGv8sgM+M9KNk9
HEvAwsKVLTZCEY4gchhEKgB0oHY2Z2MR0IDgro+pYfz85FgNQkKqVrnxTjMDXH5+2qMGWQoNbLFn
AwE+H9g+xxMMPqaQgRnZdGOOCSxL2DLQdcFHv4UaL6W5KtjrmDWQiRdCEFDNEuUKZDDtESbVRN08
LZqv0IXqw/0JEvcE+i/chbAwdTDKIuxoaSb1kHaMqMnDezBDtfLVLBbTCsQ7i7UArIySHZLZHYWZ
qxASRiHgp32NI1i+Omk7nRTYaHJFPgKmocHdcO92jiDWkIgALsshmgA+6dNDBbVr3iXoXMaCta/R
N8VzyuH5TGhbrDrgAXVAKeXRCWNl1H+FIfjngKj1BLlonmr0JVlp4o+j1mrhrK5D4HohlletGnc8
PS/1CyUvZIu/gDTYL+ACX+S1j8naO5OEnRTOSJ18+zmVlNiEXaV7UbWBbNS3LxabsSq4DFcfmlyO
sA/A8dRaYxcW1/+4gbQhdRkXASMhWFzMGg0QM3vKBKLtJubaPdWbAowHn9TtAVjbAKWleyzXtsDK
dS/C7Yxor9xG6FeUuGzi8duf/47xNMGjXjysYhAfAy1AGK61D5tKseHxOSd871JsSejgHveL57tU
RpAusbQC7GjDG2zfRCDJYkp7vr5vOnGT8c74AA2WdAdo0csaRTcSadRjnLbLO+JRUYB36f9HMyF7
2bxqAqOOMKXWlr8mSHTekCunlTs55f6M8z7tlWDM4zoFn8BeChvRaMDCD+o1KLJBz0Lao5EbGxY+
JVKVLNzhpmZeWUODqrJaK2PHfkKoAfRvJY2D7BXaHUt0xVwL2G106JppEbcoUdLZ1qm82U5tQd+7
0KHcdjEqj0wIaahCmXOvrxeHELHWE6qcqC3ysRoPKIgysCzwIG1dWp8xYC+wdlvCVo5z2/01O/UR
lkVWJs+6v0Ikosn23YlfZwRzJGySUSYMuKJ/EizwaI1eREEfzjJZs1vyQHGTvl2WZFzn+9xqua4F
HkI7X3IleEdBa2ejzh3P9zZ+GtGS6TWIl1jzx2jmZ6/FHkr/ZrPpwNDuu1rZRINcnqQcMrRJ0PDr
sgAe0MgNEMJeQtqxNaqwog6t4XV8u/F1Dsh8WURnBxGci1Zl5yuccYL2bRYjtkuwpAQnxg7GmvZY
TV/X/nlAbodNyWyI/NtPfgYq+rAfEUr6VM8KZTGjQtlJynbHETRLyNdsW1ga00X3HIIeJDXQxf2U
HAIaXblrJdn20G5CBxFNpjDVM6bjhhf+AkIXA4X3vtfM2fk+5c4lQVj5BITK7x14hkmhhQGYfuL5
/8OGGUBjqHG7lmsbkJLLTKe85LsIQKWjGZAUKoP8e9rtkiVW8Dfk15/aaG1HLgK9Rj+mbq6/iMCD
q1BLqcE+Tawelp0CFeNSqzl3qH8QgeJPTt3ngYouTI0mgREJxsIitMUmBV3q3aJTEUWPS7AHIWAv
NuXT7NBAaMmwU/BAa4ZmdqlmESgC3JSvBcKUmUYgi7FZA+lfXbsFd4IoqmKjYGCyufT79dg6UEb8
K39BWmcPojRxTJcceztaCpeI759nQcyVAvefvuy+oN0ROeKRtE2glRL+6plc+ILsFEHjJDMDpsKs
qj2LFMOJAg1g3ygNtRKbZwN838I9e/hSKuX5wf9eOMYmq7Z10eWjc69deg5jkNZAQGpmG7n5RqGB
+IHycWP6CxhsQMthU4qVBFkCedpn2d03so4qh2+h1WpfbsuB/VtRl9X/ckmH8KD6eD2JUfNoG5tQ
iSQ6FAJiwQFyGQDfHtF9RNBXkAxaGs9I1xESW+cetVTGFrQxMboMUUKUykXVENPARra7/9uFphJV
gzeAs7RB/6d1f3JFryKyyxR/o0AUQjMQhvUXVp+4OrFhOBT7VaF5gAz6gYD19aFLLuraXd9BVeJk
veBIM1RMlLQiEa1WdSSOIoGOHsMu1ZGrXCbZFOET3Pn8oX89qBaO5/fimZMd3sDNx4i/e2km4k0L
lxSMkDfmpCv9xH/i4Rk+7AmsfYZxp6irc/hTlaa15IIxFag8EELjtshoD8JySJ+JdPoukCNR285Z
Rd0eOPw6O6I395YDG31+ug4luEICXIwdPQ9lcllAtIdXU/b7GR8MQZFPdbQAhvXjaBhOeCcWSc4M
/2GD+kYQJIBLYPzteMISvVpqK6LTBfjNYkhLSn/nCwT09BLqxMqwtskP4EqCYyw2esu2C/cXKzH3
2FqyrrzamfKUe5NAF2Ltb8IGmHNGsNQaK8vurKxA38Xv07ZSCM8nWzn3Soy3+IY6IRYJFYKosKUD
hPnH1vhaAJF5uSqT70D/c2uhGvt3pcXu99qFsFSIK8gLs4h3zp5WkUVhjzBKxOcFTy33JtM24CJY
xGcsFuvp+yYz+jrptIe9r+S9AzX3V288o+/cv4Tkz1rqxY6XcwKmC/bc6bWC2j0EwBmvkkLPsmrz
5yw4RJTcqfO44WpaSHQGzos7RGXs3prp8+ZOxC6/0Hqw1lDNcAkDWWaY5vg84ZMGYkI5YHyW9+Ba
+Pnw39nMlkuOiJaNTLNQcaSuQeecDpMPH0n1c1QIZbGyVqEpSjVoOT5hdqbQksftH2lxSTutUL6X
IZWOp5ojwEy745cf/7IfbLuibx/uzxKKali4t4Y2WVFywneEqFolkDgueYOxq0syFjjFLP/W/YQI
ZhhvgyADlcfnfTxapDmj8I8gbQ5NgXhDzXPrMXH27mw3rDmYYJgzLvnrCHXua3NWBeFXqebR/LPz
jLDILwyuPjAJOAHUOvHmpTK8KuK82WUDSFnXMu7lBr7GYr4dfqJFt5rUr8qH7XfsqxPCVzUJc0S6
2VwO2FY+3oortguOiASKxYCJyACBkD90bz15bTJQYRlMFnx4SrWku3YXjsEujnLjE742o6ntTVMP
cnxSry8xanE4xOQx2AjPv9cDEGTfQCzDiKXamNpGLWmIc1bBpAaHtiTZzlHSYHmczW4O1kO9gvu5
1XxU/el+VD/+qglrVcAy/ItBcqvh7sOc6sqsZxYwxX07Nl1WmICsY/ddUQu7ICQUoZ2honY41nPk
qd5SBjbIFlVForb8Ihgm1acaEj6JabqGJt4Ra0ILopUxG9fzZ/+vY3B9ESV+JSOxVuUufQiLsWAt
kCdXw4wqS2iCYWODNT7I4vJrPMREjDpLfaN45xfKo2d/S2/CXtVFs8nRuGQpp8so+J09J1Pp8ybj
m7R39MCjo2jkxmtWfuuP4Qdtap5a+D+PrgeUHDRORO1a98HVLqQQNxgQFTcsviB6p4b25aZfqaWk
2Rld4NxtXj+hFAEDEwl4Qzpy+mMq+ITfUr2B5YcRCSVQaRKqtENCoJHfIkn5yCoTyPYviB4usMvd
O+HsX28OFOvP+zcdn+4djAzlG1UiKRJ6+fHdjgmzTnoURRrotPaq/uMwuwtBkTpK+M+uVvZly28n
1qxmigU4C6uarITo6N5UiRVYVlv0WhY+iAkBDptwuZ9KH693xQ8C6sCnupfcdofkgngqxDcfwcM3
MP4TevfLExRAEqWhghLA5bXIjia/7pA8d0JSp5me50wqnSi5JqXmhGZM/MxoOyQU+5LZTx1B1Qme
woXVdUmutjSkCKDes+YGmgvDXTY1XSBCEnbyfsDyX5LlrM4ph+iq9lkQyr0psuTYGaj5tuVCPfji
YUKq+c6Z7TbfBRLF7NG2vhRVZThbd4PCQDPs1B5wN3hRT1HoLbXUSigT3ywumvNE1ow7mC6P6mfW
EHBU4wAgydD3TVnt3M5gwfyHA4nZYEzSlIa3swUl4lBS3mY/fe9rPUxo5Ox1SfUq+rnaAeD8jw4b
SukE3WOa6H4d2DI3HrxLmfZGEpa4u57MAdWZqQOc1Ob0/yNvN7Tcb7El5WO78cTZHtksOK72zuUH
b1kVZB1xcSxGNA/SbSY3ZuWkeMKyqIMHV7Oh5y9oFNvAXzgBNz4N3F10S/TH4G40ZdylbluV6j//
WLLOS6APaRVi9Fu7sZPU8dcXUa7f1vzErlyBiKKtXNbK9M2rrrHSgY4a2Ay0m8LtDlUKr/5qZmsG
lv5TH0CNp/hfFwBJgxs5tkoWw7zWyfGIyyokceoZdIJosAerVS2UIj1B0vnCCVSMHoI2f4J2m2Tr
96ORXJV/oEPDhPGzrj+04k8R3a4BLM+9LpLriegKcE3D9OTBBKZ2htv4JXtYviu0ncLc2UhZqOE0
QoT0aChmSBkgw2UwbzfF3Og2P0wkc8hQVifYOYy3yu0NHg4=
`pragma protect end_protected
