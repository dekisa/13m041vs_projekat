// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
uBK39FkThwNcYWDTgaxM4JZHZ6h3pGN+i/IBtioqeB4SMgcBPLfODsl3GS+y4snUOza+okmhOO6t
J9URlpG+asW68HH1aLlp1nJ/EwGhL8waRUZjmX34i2fCZgl3Ak9YlE+626yrpHgnvHi/srkb32ek
igoK0iQ0oKpCSj+PewFEsIS1b4WpS8PoPOAR3BO4XcuixeHhicfRHa5G3ApobxDYpEcgbnVAx3sd
p2fporEuq4x9ir/Nahr5loHPpXgi/o4x3pRd2W0QTF3oKgW1JG3ciLK2wPCMui0Cq2EDq93VZHA2
gmDd7VmBY86tVw9k1kuukyl5PZDm0ogrokP4ug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 100624)
8w2KXHE7ndyRPrXP4GtdB0RBp0AAjOu7RvaQ+n4qZu2Ag1RTOFHDxk5Z4KOE429wrGKSeY9T9Urp
X0eNtIn8UvapPK4rguSVIbum4mMSQvV03CkikE01K8xssCK+tTW8nIIMBpm+jUxNiDZ9huWAdMwn
J+O8Msxc4wHO9EioekuiDrhEDt1z8Ox9sVDPqKfmQFlgj9adCE/P09p09Q1tuNid+Kcvf/d9TM3C
y8PsW6tqJXHq4cXYrHT3+ueuwauVQ1sLcD7W4ImeCumMvI+ZYLoMVKRsa4UybYKsMxh/T0DelqPu
nSKSNxoGZZdcI8XKFNqrh1Body2urhj4M4+KvL1XeXcnj2z0A+GFXTezTRdSKsTWxaMXpVTTcITo
NzHv3Jm7QXgZEuuJyI8hQqRPrn09U1h6IZXDOKihrmC2ozmd7x2FpW4C49NKwT+eFnUhsHxYhOLR
HXvmPOGljLeta4B6oHOKMu6V1Ye5Z3qKF1bF7rea9l4KXu787Yk33wfpiCor6XPl6ZwzUly/9T8L
tXzArlYhDWUBCbuIOS2g/+7yfsKiNtNBFcQAAQVzK1RbzVOpHsURbuOfvhfqwPlQ3nP010U+XZ7m
nfG0cVgTlkN5R+jWG7XnU/zc6OyNrS0W2EB6MWYXb/waZ1CQJJyxD3QD6rTIHVsn/sX4nrZs2HQR
DxTdOfgOP/KLBtfjcrEEJ06fjP1Te1ejlGckmmw+Q1OBqqFmhS0YxSG/Lqbr24lWRgWyhUUj0dM3
J5FLLKVXpBK3/x6M2a5v8vMLnGOnwrmbTIWLo3tNCAD4F/IJa+4p29evzeJaWRXsWz3aCzaZzAUa
+ICULU/djK0u+Omjx00BertjibMONSLtLg5Dfv4wr16Ms76lyIZrMLD/AEjtydd7DZ9DNBCgND+w
gi5lZgIpBl4DiE1FRekluV2L1hBmUwlHcsLZjJCzVeQI1szvpL9+xwn6+w445WYbuT96O5EP1KGJ
Jzzbygsrks1aQizIYx85IYGJXyBitH5ouuhzJipM6swIrVxVnQk3OuiCvDNzS4VK3/G/aeiv0bsw
Ypt0zcPErApKgNwcgzG3u1MV3yW9XFShm4VSNR4TXD+8KgS2RCX+9a5AGpMSRsqhWRCFuFbCU0Xr
gUbPkOsvlcFUT87e93wouKMV/oLBTFRoKcydHkjrssrz97P7IgEOHib6qmkFVdV9TOh85rdQ1KAP
AgPxXtFOX3SpPRSjEOUPdiAkjPXmNLWJ8+0Px7c2tDaeFbijQISEAFgqST0m95IvMRrpnyngL2Xo
UvRiQPFEHPRJpcVSA1hTAYM7uDxaIqwTAr0EmUPyCVv/r1LqPOlGvAr99U8qUzxNCxd+T9GmvMpD
F9gUQP2WoifT+dpEAsxuuonimpmIL+3ysslJnLEVCxvLqAzM69u9lu/AWA1/uUHK0wFcaAx8O0jP
8YVf70BzNsM9EaIvzppz79MAmB7/LGq4RRCBqylt0gCnYatyr9I8Hqm/Fr9/7gbB4k+t6MWZDReu
ckQX3gqX3OZRkpvXbQtanvVUoVdss/ef+1H2+rRIwCYtcDrZVkle9lDNMV+wrO9p2gpLwZSc+7h7
fNdRuhfU9b4qQUV15fY/WmSuXIkJlezxlL4tzBKvyJZ7w+cVP9BY/wzk+6sxqiGOO59C8rcbXdv2
qSAviLE430ihw9NinxTLH53yKUJM6dHulwmfRzv2xyP+xMlpU7XqKatXi1Jk4kbtFFEBgC9+icOu
5BxY8yGNQbai/3WfXkdw8ZjdqNyKrPVxXXopU6AK9VfXYIzLEUbLN2qkY6Oznb9f9fE4iRlOBFYa
5FDi3aLWvLIsjRxdnW4aFmGrXBypq7cERJkitmI5PiwmDQuKQnD34y9eSviuw9wqcCHbAAqPR4mD
kBDMFii8ErsWCiar9oIblxc9d9dzoujlkY12foCpcJx/BznC38iO81E4YpmNa6Zx31aggQo4SHWf
AFSNZ8YgssVaUkImE5Xs1jbmvlly0X4Hl9w1rsz5lhYQikHWwxrvKYMN6YxrKfmi8S+EQtTC1pcP
zAKbY1QQxOmgCNgWOkyXT5sICP5TdX9y+eniuiCHorc1tH9M9+XrsuOu33ZDOvcBqgllvc+IoeM+
D+OL8fc6eaMzYRrKkG1xytU1WbRxHKANapzR/iK4rt0DL/0QMaxJ9c0J/dnvtkaeSSHWbKVuXNdA
Cuachy0G14yoAP0iuLBYSetik+6UQoxQ8v/76DP73y81Mi6Sl0r5aHwLaYsHQh7uBW98GCDKJtHa
Z+kZKmfDfSjuSJUdgElZfhP8N5J2YypwoQpybTQdU23Whs6VRpIwhc+KcDvkRtGEIKNBfKNrhH2p
YvXfPiWJviezabym9Z/p6EqELGkKta7usqYMYcCOeZrslbZEKDvVVrnSziEo/ktu7agdm7Z/6qQJ
tNnX5T/Ry5cYuVGRTE7rygrGEVnoK55XXvv+oGAG4Oyt1aC/8pMtn1dvZYgY64w0FluVyZUGYcG7
H9Gc0ORUYrmNKe135iAs5En2eOKsNyVRfrWe/uasGCTVofSsPGxtr98PQTHLwtZ/8u3DckiTUy1u
/UHrFZ2JYvDyAtfmaMiVIBf0KJB7SdlqF29VU1Qew4gx77HZLX7FPIWoWckAFggyLhDPxM+Ekjzc
f+w75lT9g8UYINoFiJegbtxZfCNYzltLuSbi373X/tglUIxYbVZOkQ3OXFf+PkZaKAY3UVuzr8NJ
bcr1LQToP/O1Dk3K9jZLj4msCv+SyDCO9ckiV+vr67hFHt/hZTcrzilyMNE78PTLjUpSA96cWVeV
jtNMilJm91bqaezbIoLVQCbnUCwQMtyVLTJFfDEvN2Xc5Tf29oXIPA4JcwV55Mq8suDufLpftyun
LY53DO6TTeFSYOz5/6KR8lAEuoQW+Yo7rWhHo/2NDtzIp1fx6WnrdM7OcR+P3Fn0dKnTCkwDgPAm
Mh8T0eQZqlVfTKExc8XKVNn/ByGZaLU+TuJxhS9Q0L8pp1S0Bs4gieB9ACU0eoleIlgtL8fles5/
l/VKpg6f26sl5ygDf4b6Hh+fUNfEK+8FAUCqXror3ebHvK+TMlblfDtEreB+Vc+jR12lzacobF7T
M2T3COhuUZb2h95AWecyHQ42NkEpgEzZ52tBrM/lQi2Bqe1cinW0+df3ti/ebKK3tKBZjixdnt5y
suF7y/6OlJG9Jkjwc8CrZ1QbRpeQWI8YAsrk3GInXg4EyRwbpl+GFtMhM3CMtsXzCKcdqRIA51Ky
t0DiYH8MgvvBKCo5lelZM9CIx3SbaqwMMSTWw94R3BUE9f8KQ6/JlMNUTNOnNIVGh07wpbfsyk/D
Q3o/8OAC+oAHBi6TnDBMPjHiIM20sGb3lnnF1dtqKPpGKtnTlJcnROp4I05E9WT3Y19bWCrhCMdX
QA0YRNEFS82+4okPdlTON3t45Ba748GTTlR2FpIKL/KSLRChPEC/Vk26OXdUPTu82KnJgRSJKBq1
VbLAr5TMMsVs9b5s9szoJcdPdFtnIGNV4yi+W/QDUrYgZmb6hPipBFuXs2eSdEQmR8WG/cH4L3b8
ccD9tnmA5abuVIIyHTLqX/A1jiyUemxyfMGGcbdNtwKUNw73U6m8Dv2C/Z2mjz7GoN0NF6+XfKcD
E21ecoS5aWonqMw2eBhnEsy3jFYNcfqA92G4nLqeW8LyB41vlG/i7D+lIgXz+4gVjt2+SjhaG14Y
o7Dw3NZtnxqDH3oXlLOOCELrwuK4c7TkmpIB65rbok0atMacZQnr7zRDLW6yTuabqDZnAi++2imO
YQvIfa/aMs1XN9ARq+hBPSAQkgKZeBfNi9EU4rIS3tMntuQCDNj07XsMreOZX0zdqHdFeCT0PUbQ
mfvFPMFEZvCJRJwkuqQZ4Nk3B4dpQJS8j3zZlN3VE6vZ/5s5zDQDlCdYaYHK5vQdzObHRlWsFLQc
TfNoeE1QEnzGtexQDekOgVr82dYvSbim3QaHztC00a0Bl2b21BVn1l0Jz1MsBwcWYAdiqlFoLRME
gKulfeMSqPforep+vj/Zr9G2sEt4mv9K+jTJx1RKAa/Oah2P/CGYNuw38rpMWUlj+R+tyS8ZVR6S
iTP6IV8m6zqkgmcf31Z0ffLPJ4i99AqxKWBvHhSqfP4sbckUtfZLzI5V/Y+UUKP4A/uLA3JDXEoC
cFVGnRZBHfZr8GPnS2oEcKswcgGzL+P5cWEaGII0UJRvEhAvK5fOlCv8Rp/PkYjHtUEL4olM83bv
rrRzTCA3GhYubwTfazNoryEh+o7rm+DSE4IhnP+DeXV7AVd+yh58c6rqp+3SY3UF4F9qE0j1pnYv
g76c8LdAd8Of4ToDPTYr4q16V8N13hne++5s66atF39SwT07+DJNp4XJexUveHZ1Z7q2ly7bnaI8
CP0aJpyQRpFZ39v6+I/T1zfx8/KLyjZPFywQh4XiKw5rbNSmlJ43742N0dvZtflpPTij47Ef4LwS
ZNT4drzUBy5qFQcEYRSRJZYjtA1I2HR/G9uGtzTUSJhyhQtWvXebCLNJ+bdtQKN5mIkV2b0iKrJE
YaR9C2bY1/ssle75tMEQZTTN1RHj/toNm9To9aQSwaf8Xe8C+A5qCJUXDsAnz93msR3qB6KU7cIm
eomu/6eyqqY8mPzC6MK4L8TmrhRoBOef5x1LZ0q6l5VW08tX1MA1z8zkKw4Kzn7TRt+AucUfSxQm
hFGuY5PvC+wSqSOHuImP1WQu8v2YQ3J93clRrkxXfnQWSmLkF6M+3gj12j10Qfc2svXarZs13J1X
PRdl0btK/IAi6Yw1Ydoqt6rzKaCpyd8G+Y2Cl32XEhrz/a1PGWi7EeNGKoSWegIHdOkU11LOg7UL
eeN/pZd3j/Xpzq302FLdmt4MQ907g0hFx8BsrsquAT09H9+eu1VJAoOktEAcQpSF3jIVkUjyvrhf
r9/OpCAZ7hBNTJh5LBdSbJQUjDoOoFmnxyPN+BG13p6Q09mLqPSsPTKKkLsaPipcEnnBC4u4Pq00
4eGXI/j7zpYgoxJtl4CrbpJgY0oEdwDRDXL/WLW/24x1msNWKedpaphunzFYGjz5d0G06bbFzB/7
VyrmcJbTymisgdcMjDVo2P3o3cmxgTzUhNYZzPoXRdOiAckFQY6+CeSmwWIZXWdctBHASZoReuXH
Uj00nEIYNZEvxwUsMf31lZdo1VVajE6/NWzadc06D/KFqpXGfuK7hZ0QklWQavLUqn/dyVrjbvzW
v6mBMuUp92p20tod+2lkvMCMTu/e/SsCkGA2M45nJCQBWpbhpOPO6F4R4tueeD3swfuWV6PuL0ND
hFC2R30flbte6auA/TQWNljOjnlcKQM2MV/GEejyxe/tZhmjvh3+tn0RW8+iqj2zFLnryypjzVPv
NV2qd9kK2A69Lx94/DuvdEzt0VMz9CtZXCB9RZqBPCRrrFTHFgW1W5CNreVoMeJ++UKNTN8tBXfH
AZz1uZ1z9V95v9B3nhx9S6UVUKN7A9Vb66syD6H3Ocg0oPA7NVVL56mYolgV8jYt8lMHG4saYNDf
Ggv69WjGX5HUWH2nzEro5TudaenZkcpxTrA6BXi/C3p5WYaUSe0yJEHnh4gbzkuazfaaiLhhOrUJ
cmwJ4YzZAQYSt+UflNWx7EjeV2JeMn3bEqS+Vndx6uqpIiGKN5cIXPqMxUJx/x6kJpHEd2ZkLjxh
6BVMWd2QCHO/nuE9DdSWyPK1qbNWDeTCFZS9nyLrarowK9DVloi09tjzAlwYlkI2pttIg8x49fzr
Yxr1sPV2TjtDV5pNJUOPlSkUcdi5SXV9gngrsFWv1uKI0hot4X3gdNiANQdiU5mDfTtFdghZxG+O
YTlR9TEH1+ghlIHK3TpDs1h16vb5laKEzQBB4J73BsUPZsxsCqXtERCzSFJBt55rvfw2IYTFm5RS
aA+97iHYsZNcVvKEiJ/b1Qw33QRwUpzGJOTlvvcKy46ZSK70WluIe7wp3AFo0beuDXhfoVDxZO+M
BXGXEBaDRPIkvmYybUYX7oj36xvW5pA9lIT/cK0ndoyFVFrciSSfqd6RpR0UFcOda5Vsq5F7B8Cu
HJ7nS8D+npYP0WymqEG6SQ5cEwpxNL1bRgQgppMu+nm4Y855fAMvLgZKuFtsk045RNWdZL7d4svB
+NnP/CTqh1BlfTfuCZkiQZ/Bw2+8XD3laJPTcOVW4iX9GpNheD/YsUjQH4hcF3/YvLmWFf4cVa6Q
Cpo38SMwhbNh+7Hpq0fdxWn02ecf+bHuz49S2UZbT23ogBxHaGhZAUST4j4Bg8KnqRaIRm69gPGW
tFjYFz23vMzJeCJY3QH5Owal3j64M5Q7lgRfdeE6M93OgUnr0fIPOpS0yxP5iEgkeM0k6d5Wuhb9
MD10RP8AH6ax49Cg1hozu+lEWrt7ooHakMAq9hcbWNy7aszFWMDcPH/qd/nlB6JlOq3OVVvibUB+
auhvoHDk821Cp1SrZ8vmCo3G1sxpJsg3AJLepx3xNPOwDa1shoyQAEHbPP4eQB8dWDXMsokWHwf9
zMGekkK9MQNt/+yEjm7SL1z08Hl56hyaRBSuHuEA5Djm7NDLZqITGI4oUsi6E+rUF31STDRVDRkE
4V2xgbLvNDzDf/emJ0/6MCB0q80myMnFCNS/3HtpodeO3DPWFwo6BU6N7cQ76qhvHn+c5pe6cFy3
iZrVWzkU1Bau6Aegxdvpwe6dlmdtjr0cRW2GLHZYvuQ2KP53x8kQxUirIl8kbfc5zRIspUHENL3c
twRwPjlnnwc9+WYSzkG96u84l6E+6u5ryMz7uObjJIGwG864j8jkGz9kMf+uOfnz+lVSMSC80pzC
oaNOcbiekT169p9qH/ZfNyyoDtVXZqqvm+MpavT1hYtEg3oeyB6eDePQU8nkIUdG2qHO8e4h8nk9
udVSKxdE2Mg7FZRkqAwDMj4CnEzgGQ9j47izeEoqr9pz1K+A4bHrJ7KcQgua3TLDi8zCVkvCJp+8
JklQgqm0kZv06WPbi94XHE0nbGruC6On0h7vgDpWDcqK17+AWElrIiXD7u8LnLabLZRrLwp8gZVp
huy05Q6qvE5l7KQfBjKEFfE9SJNjtt2HTi5hHFuulbWXE2qxQyFTu5gDpsRftyTNrClWIul3AxwX
pOE01/2mYTD0KidqkPNbcjyvvLap3iOBMFPO7PprQE8kuFLPR1/0GFVBfTy3+Lc2XWKXvk00B5b3
MElPzNN882u3MhYG+69Rl7JExoXRLwYy1ItooCvdpBkPAb42/AKcDyYntUUIr+frvfJ0kS5+CiOK
l1zA5aR40e7eIfGcbQ/Wzg8JbR7s+KqqGbvsgy+X1VMjclgTTfa15pL7hdNM4YVEmDBqKwQp8zh+
xE3QR9kAcwmF9Skfa/F69mGRqBJE64v/HecGBd+N103D/BRCaXCIj11ZIBnVR7ctC86Q/0jk6zZi
j/GmIDKKzFurtJIQZMYILemga7z2GlfBmfSJ2oA4MPdL63Fv5nHs9tVRNL6V6yO51AgsV465S8CW
sgrEl9ZSuKUyNyzgnyUx8OnEPkc/UyLl9JgCw1a2gGU/kBxZ3XAJ5NVl02l3QHZi8juj1632L+2W
Gw30vOza553tqTa/zGBCqLCQIbNW9s0Bo7YYa6u9dggqMGOzN0PWDV37eJpSe+QFR+GjL9r8Jooz
JiJXQj1vIE1I2Cqmmx1yem8F6rIDpqFrMWnZ8iN+KRaHonA9xnn96lrdr58GMPCMvRSB8pI0j3jF
NXwCitUTieXMNsCeIRzPSipB27kg7Z70SOOQ5HLjnz4AB7EZsW3qBjGhk32ggTGeDPiN10AEUuL/
6o7Ms0YtR0FgJSBzqGaPtAI1azldSv20uFzx/sb6z9qQj00p4eccAFRzheyaDUVIQl1HVkSlcEaz
IK6pj9y6vEBuEjkvpf4agcK7x9cINZ1FnGVOdwlFdDJXFvcBm3fltGcHmcAEIWKdNuYLmNPANq4r
XgJpzsA7D4JimzX7CsfjNEVYtstvfRThc8uaLhFmSWDe4NfVv/Qjn0Dw133yVOyLgqbWeEb9TOS4
/RhzEdY1lqRH3PIsj4nrijJ/cLqyWiYVbRoT8b5j6RKrmSew7lWQ4wGCHFtiPLX6F1xJC5JIm9rq
mpPX47PlpdXcY9exGQu0urQ2fSvcpsyrwyENVnczFObW7b9XO+HLsdgiBoMHf5JXbJDKwUwBJdfk
2/PMuHjJuVT0pVoILWWcr8469p9XQLcHtjSwz1aNLP3z8uJ2hQE3tOxSMlBSYP4yvplALFd+BUM5
oZfiqPMdQdiY7Dq8W1L6oC6BHPXdUmi1q8q8fGNDW/qALOJPC8NhfIE2zZysLt2UAoe1lkbQUUDk
qPZUyTV7E0KiaSdNFNE53TzlYN2CpprL/TOyVIB188N7t9J0irUFjYP0Jl0Vo0OeqBVeaEeY7sLt
W2Fcqn2qSXRdcp/rsBYPTvqAVzd1FSEiMgnOuEBmLbYcKzxnRVVK8ifE+/d4ETEP7m+o1XSputpX
xdmCTGKVmqgEpokN9K0G3nRU7szl5XrckjM258lXaLw6H/fqHKfjEnL7ehICSLNhCfJ6U33wa0el
Xhn8MI7B7EyrRlUNX84RyEnfR3g8OjR6m2vm0+i26meek6gDOVEmshscZR7Hf21tjC95eAuDJBg0
bB5n3RiRjlD+B9wGTGv9SaEMUGgKnEh3Kd4qKdqZnuYfLMaJzxOoV61LynKmva/Lel0EQHSRoNpp
ACRTdqRD8vPQ48rQZq0Kjm3GYR2mBedTqwmVV1jUPgtf1xcUstvT1bNuC37nX1d352rhn1q62XkX
DT5Emy6l6wpEAK6jg1txA8NqITAWXu+o1JdmXbk01zZM1QoEwTd+llP0rzqfxHGjhdaXW0zFJifT
wgmgyQd04BNyzD1SGbOt+qaTqqNKUYZPVrQNcb9PkZ7hOdcGFkoC2OVzmVrn7nb6+pvtqOpkZZyM
QzpOm+MFZQsgsP2oqe9ztaA5YrUl8Wckp0ZTWgKDLV5PgoAy7oDv6UNmzHgnnloAeeaiusNeNHmv
6njldRQqrcvpdPl86Hb57ERqEPtZRigmGAAstVXrZlLFwppmxk7wVQtFRH0arN2VEqoPafICQzrR
VkGwbIZCtvhyixHOr0RbfqXsLW85798TM2iYvaExmjz2r522h44N6F/5cciK/1vcYFz04xqVI/XO
H/qL8yNMOe2ilzBwalnuN13shhHXsDUDf9E5BUdSmrXDQGwrIH2wbsDgM/xiKviMcXK0mAwmnaLn
Mx2+6j0pe/qfzJdz80Iw7K+eB8Y9OQVfanGR4UXnOIwPxFJUqQI0NPmyZLUJj8b6Z03VHzqqGdky
OYff/5nlZqLebLy2TEVI3IFRC4uNVQhtmcz8DiJh1CcTbaIA7EzUkYmmOxrGRnODGwUnkwiAZbzy
/IsQDACcnN6q824Ays87+VEwOGmVARDGatjM+ms5ZMJkexQvuXPYsC1yOmnHGa+Uw/mCaNCV09iV
y6Ty4NcqPuMSRdZKD+5gDiiexIUy2V0a00zmUIikgU6GQAwhLua0R0lN6Mir6DW2sBdR5HvFGktg
9SQhn44ctTfUpTYpEgpQAP1PNw48qEXFU7pry7ygfJzXaK7YNhgjqqTpa7SpuPGLXrMT97iGZZGB
5CrgTkFrkNIRP9IhUJIK1CHEQtRAxGAQAOVHreSDkU/NoaEDtSvFlqNfkpTX+6Ji01NNlQ9ILCcp
N1H7a8Rt4ngLgwE9SgEPwJefDevAeNT6CStHs/nOeIVSWQK3EoAhhr4pTNBTj1V7svRM+P9hIzDP
UVYctfjOABtuEg9CL8dzjVnW6UK4x78+i8UHaXOlc1upnbFcXPOLnnlbXp8UWmVCnDxc+SxTq2Z5
QsQqEM87q9o+ASqkVrgY6aTmh6eIlm1PLTMoDZeXnXnbkZYV0V6l8iwhnU5XBzCeg59QDgTisXzU
luyYNmn7W0eXmuUCZESZzpqhj3qEjf97wDIHuYZWfSOUAjpNqk9UrNBKHEBkdCjE4Wta6LlrFi3R
kDHR3krO433FeoJdjp9NmhVDX9PmjjVX8WPt8ID4Ossf7VeBZyAyt7BL1FIvN1TGAPtYUTRwolV/
5HB7x+0KWsuqnhzUk42gTDJIU1osEbiAzg48gbD+wUrd20+e1dtmEuP1NtTn8SgT9EIosTCJJgXE
V8Unu12qVvopfzinbneAu89qqncqE98uf7/zFqhDdRU1RYa/5mCgCiK3Z9rKa1zd2I+KnBJafjvH
2CkoqchMdFouQW+0RwNVS2u9KdAej83J3yzyPpmfUw/6b2iYJ397Zij787eahgmhTM6BV7JBA3sA
YURmHHv2AkfjxcJGfYSGTDgFuxchjsgWUn1PwmmxJN8P0GX0CwXhBzuwZ5G1Zn5ze/168kOSs74/
VBP0n236qtO9Bzu+V43JFoTvMtKB9jp8lNuPCAa1jfV65O13qGlU7K9rsL1EMWJoTTjKNACDPIJS
2im5k9tyyT0vPo5gmDZMTnbnG5oDc6vIzCFJv9lOx42Bi4s7Dad5yEwtSupSDLdYjrCzSB4D437i
veogVZJzFOI5t2po8SHRSYaa+5bG1/IQQoJ5wHMTSpBOTKiZCKP7XC8JCFzsNhHUZsy3HFT9GWof
s8QK8CG3GlC1LqWZWiaZdkIpw5qeCP2qzjflshTZwFaBmBNDQMBooFrre4WnxdWTzwyMoyK4PKDV
97zyfDrDotpz0KLiKpW3JCXUUVywdg+Z+ymBVazzo9mBJLJZ/QR0+5rtl/0smWHTwljRbom/Br3T
PBzRtc9ZiIc3UjNPG+cTk38+LOnUCOt4qFbqyhea4Z0AZwKT/Bh0zB5iwn/8FG9pHlCEsMabifzK
S38/rKHtlp8dVbOATAIMAggH9aZUqgtVg/6Vb8aq/abwqrQ2jrsY8dInepyHyKgL40vzpfrybvPj
sJbzdS6A2ZsscPZ74ilCzlU1crgY5p6KtrQyLEh0s++o2q9/RTt7czj2lMj2kp6Z8OR/PMtj6tsE
Kz5oGEcupowMcJy/Et8zaHmgUKgLi/K/UtNn6Nirfw8CGQy8RcMs4Z5WR/FPTLH4pUG1USV7sc83
oGgCh1TQgBGjtj6mS2QVJtaMwH1KMs+yCnVezG+unzGL4Q5Qy+3wJrxTB1tvy0/Xts0F+rcuNvLc
bQ9MYk3LDTqO4Fs9YHwr+VFi3hQvTJgQUqpKNr5EdKXEq6s5TSCn9w5KL6JnlVYnaS75ne/47GLw
JUd4YjZFhMji2FnGPCkX5PNfFW6Ab1FMHOV/Lq2o1AZ6nBZDhw0m988duoEocFUjaac6VStU202U
/Y3KlW4P/geD+DwviR13WSEeNS4CI59GiBpetcY9snI/PiCk9OyCgDJUfo7oFAXK/x4QMzKJvRe8
ktQU9CLHsVSqrqUDy9WPrOSleS3syiJZkbUAl3JX3xdlhpqb0gWSJSU/9L03kNeZIJf8Dix/rZCY
x9VirA81gJYnY/bYg1AL+k6xaJdqjiBdW9wrBIikDNaxXbGGWlj1G0x2e3OKsblWSlA5PRQS7vLW
x91qDe1VQ50IzrUg2a74Py/lDgPKLKswqUXDjlJ/VKSZIRvasWBGmOL5nFB+4C1Tr0V8jnNnHmF9
XW+C8PPN5guJoRbBN3/XoRZXcGaIsvk/N2hDdUyTIbkFRY8q5Y35nhpmA02GJ1RdCom9pntr/uYV
NMBhhXHt2CrROrkqkbFB43TtVxUN2L1me2SftdO9eXqOaFcvlVDrEUmojY8R4C8SfYnhYqfGZW4c
eqiajtGJi7PbXM6NNS0Zn3RrV+JnvOhHYuANAg+QnGF8k7xa+XESIuPTBCE6GKIP+fO5bPBfFCOj
fX4xg6WAxGUg2PZhktPYGftFWLZ46lzVMrzjGWhlJd0gCb4k2pFwg+tEctH3+hvuImBwTq6wuOVe
+XensTAu+zbu4zm1spRSRI3okH9DEuc/buzzJIy9F8t+0Xi4AC0DXWviqvm+fCQQiU3d+biyY2pf
IEjs1zYe4yagU7xAq4uvfw4O2lCrpllWPJye+slxaTacpa/msa8Js/MR+viyBvnAY7KkBVQAOfqY
7TxUSU1PJ3DFpLI7mlKgn3brMgjEof2jVbKv7AIKmt8rJKzu3deLFtWevD/psHyw/1bCOMvqwfpn
hr8y3J+KYMst46+SelOCIMqiQthUq44DKvWo1fCvf3SOCpu09j1kogmqOdAdGoFd5xEAf3s3D7ad
uhlrdV6YeQS0W1hiT3rKbMBQxgoYLWOnrlPSkeu7CCD80oLxcxowoZ+MyFL/OFOW4D1oYQ5FcAWJ
Zf4OokDBgnL0YO+L+0/Bo+aAK8chDV4ju8iBrBd1Ew/f3fFhFf4arqUyiumT93ZrqemzCR4M0yfv
3zGN5wQsJ+44wpCOsFHQEAO/wH0R43mH7BKOehee4nlicCF3tkrO2iPPPkxbRVIhZ0E/5Vo5vFSL
5kDWLCx57wpLguRT0nZDRrJ6sjYAZQeePFTfBOBW8neHeUrvKLOoaJ5nXAzizb64nlc5R2fy5qVd
uyZDsrwxKrlW5dNz+B6/pZ48aEEJQ6rg29Ph3E6pgcpPsdyv/jAL0lER8zXoAUdEVgvXNK284v6M
jtkxdoLFlMem89lU4g02ASCNGLgihGkDSnQ94HgVd0Iss4Jm+EatsiQZ4s+squIVGZa+Um0jv0EG
LsSG5ggmEtn00Flo15zdGfkv2r/swW+QTnlj9AZBYqzQBtnv9HehNZC4hZNyaRlgJ4BcaHN1zEqb
72r3Vn0+dPEJrd5pBiMnctgHbToyCK+C3YzWjQ16JwyDUGgjvl94P8DWg6agOkLMbHXzX7AXDw83
n6k92CKIfjTnyVnCnLJYAQI50rgb5Ryr7yjbYuA4W/ZnW7CEUKGyGnZzlGZzUM4XRizdd0m7moPY
+dAN2iRTIg+1sEumUUlIQieaxjgH6P8o+4QwCFeuSsSCR0EofQo7HxIwq1BnAGO/txSQ/qXe4CJa
pn3tAsgg2DTB9fQxvow6aJre+Lv5xaxwjCz2988M9uTOgKtfimO4CHECjkem1TRPqY28An2L1WyZ
O6K+Q9iLxlJ5WYT4z0jssFTIrJp/I3/LuJZGoM0lAYDCGURCIUMxB/zRuwEJB6XKj5FoLV4sS29K
2P3mywPa5H8ZXr/JMoux3cMYl0/Xq2EyUJSY70I7mFHIXifIa+cd3K5bwKC+RqJwdFkiT//Dznwh
z+7iH6pxk5j85NgPkcW4JG546mTDy0LMkCGVQaJGt57JWeUlogHK1WK2CswMEwt8yFT9zDyRdtU3
hH5+mPO38hE05smZRV9GL6o+cAZ6mZjr+73h7q/jUzovoSez6m0aV4c2IT+4wSnpH6h0T/AXTKur
QiJl6DTUa44t9q5WlwSdP6QdUsERhkKl+iJB/m+5cBF2sRpYr9PrUG1VmpTmTtQx3Bi7XyTJoVGr
heQDpYjlc9zrLYp7K1GJHK4lLomJ4iBUFquASqSMHupaIt4Jqg3Oi0uYyUFOs1oVrQu4NMP/RENU
U9zxG3ciE1I3G9kvuWg3RqVagdHre+f2fhWyv9MXQ4QfISLZgUBNNphFCTAwkGSGbN72mUu/I+zf
GMA0/iNeRHBO3J1jC41NxepEdOpT8D61UdGVrVLYlNAd2xO6WQdSa+KuvauRPa6pUsiOhlizrC4m
KwOFxNGlAOVjWpUiUXArQNxtbt4RFKbWtAl6V5exChHAIICzHK+Ta+N8mBFWGq4VebOXUfVXSXKE
MyaW5j2cGIKlI9kzzOgaVf3Myhd5N05FJV6O3PbgwoMSjUtHK/WuR2iGxFjiakGpDHtZn4I9IozW
XZK5bdfRhiX+MlbOJOW2UHHOj8+dT/nGaip6gC99wCC3Ug5PaoSNfpQ43iHVQrGNRBJaOkpLOxXH
BlS3yNwE1f/FfveBxKphdrra1ayULLp8Ar+mm5MpFZCFJv3HvYVJ5rv62wBmyFBIg2tSNoAXw2Op
M491hXLzL3hZjYhgjOOaIm+yDEnf0W4tWgFha9oj7xN2Wc+vAfbk6ai2+VRD18fkkNGj1AcDY1fR
OGQ3+i5zRx96ujbrEViCo4ktUq+JvLyj3qDO28mriAJEUpz3WCxhr1EpFnd5TicqQJ2zOhY3GYd8
n/BEViWt97FhFEBWqjxt8euWW+L89pn7rX+0Ne2uprVrnA4NslbU9sERZtuaYuQ6emhaEiwDMydH
WRXOfeT7VNzBP2JwZ+fBe9gau1nArOTyuuxxvB6Ri5ektBne0pheWil0tMz2m4LgZeiZ3vMcQQ3K
T2+CKVJ/vIOuyRo67TU8OAWF2mEqWAtYcnHKhbABzezC8NiiNFC3F+R1IgHQRYKE8yjhKMwHknAC
SWjy+nddLr1hNvJraonBd+4fC46vx7L2YOsySaIrwt0PYQ96sJvGs+SNWb9VtZX5wWoJsZb3ATWh
J+HdYIMSH+CKoTKLHCZWOHoLbjuOXmy00/AquzeE/Wuw00ZH0Soj6VxT89weFHPe8mYsgnJhajWR
pCJyjVyj6qXcDSNc/rx6pokwj2huz9325R/x/qBoTvLHbr8r4jt/IzKo5Zbp89bAbcTcSjRlRgXI
bXv7CsnnSDCTQcZd6w/b/yQC0ZJLh+ygNDt03c9NHaf9+BonKQ2kKBcnJVJ70rDPEYXjs9fR0N39
Kx1Trn8wUiu1NNM/ZqqptYGk1jzF2VPQZuBVpMIGt2dDCPzWjBqldr6pbsH0kcZx2lPxf/6CLfra
miPmUeOu3LVDudLK6MqJlAY+/BIJUG8zA1cSQ4Qtm1hmY2+/x2ioSP1OvTcDhQjoJTOPdXaA0/o6
bn9Q5hF5SDNwA+c+TNjGMYdVWKwKNYHtWljY+4adBBI6OfTcJh2BrVLy0BXe9g5Kg6dUT6gBVTQr
kLxF/gRvqjx2zGwTNkatbeiIJPFUALSK+5jTeQKdbZI9LXiUx3tu61hFnrQeBKNH+kMjlayHSVGl
p6P11rMHdHnegIC/8xKN76A450gTw6JQSE0hY3iHxrdAcWQmcW3WS0QyQig4/kGo4pa+e6bJ6DDE
z9j7KtrU/BBvvvnEHG/VkgHlDDhXpMPDiDvpMYUui2CaUpEDWihBSaC7XJMJjEb9pgzBzR+6befV
2WZNHNP4YGubuMUL7sqFGB8oHuZJx9EyuKK8cFmj6u3ofm3Z8jt5CsicVswSgseYtXIaZq8ePEQC
ZLb6h2lLMlobt1JvyNkgOpC/WUdVAsDtJTLK9+5EqBjeKKjzbbRDwAG4VgRnDo3jfJShPSELTmrZ
MxBhpNACq0u+2sw8j6KojPYJbxs1k7rCkEUUxHcg/q8V6FCw8nbEpylvQYyAi7JmG7io3iYv7zd6
y/AqE/1obdzOEcjGtdobWFi80YAgPb2KMqkXPltHfl/ilI3NpvozUFEepPs+DMFH3oQQuRcZmMiR
zBirSnwqFHZodrvNB7PZS14O9S4kzMUw0OFvePLHLOF+igEpRrO436dhPfNoLLa+xkv5LKRpWMZQ
v+P2rdxmo59JDlKyMoToy/1KRrYIaUfNRkR72gkanwtSkSWjyz6ScWeVS07YXvgXVhdXjM1vazCK
4QfyOXhihuf4EcYPv4w0Mp1NC9Q+qiQsFiiJ4crcUPS/tWLkkS0PvdOcu2Rpx1yepYk1Wg5lZnnE
cVAiIhmwhJbAear5trlhkqA8g6ZcnmcJdmMbYmv2BZ2upr5l+9tqOTxGylCPxzA8+X/G5syaMsJG
SewSypwnD/4Tm54sW7GTLrUI9rkN+RH1dba2CmfzYOuhvSik+pxIP8grcf3XUEL5y5IoDSR2EGcX
ex394PyTjRqHAv3GCvv4YLuvV0kKYf/Qz4OY4KSOAJ/4bbxr0jJDffI0BZiyxMYVH/078DduJ9mK
wqGgju4T7Y9jTRpnflhHxZCzIqz/Eev5p1QElfq2bsEgnw3danxwKCEhr/SHCxM0YXer7+in0cwP
dYAfdLQBE7eK8nNVGyF2r5O+2I24K9wLe5KryYboRDR77IlTO1smUEcVXt5lGgMxBABKGBfQSh2L
AmiG7RJ232g4nc1ErW915EOjaQLIGCYtMrx4IfO8RqbYg3pRl5/qu1Pccr94HRetejhe8KTeYwgy
ewfDnvWJXImkdVeNBUM3nf2/sD46ub3TNlbZ5q1W3nQpAYlWjwDlpAhhurnQ3DbAXGs22Jype9EW
d1V42DT1mfgWOvtrcm7/dToAIb6j484DmZnFJN2T7rIhO9duqAhOQ5WSqopPaBJwswwgS8RapVcM
XFA0x9DY3GOz9bENou1N4kzEaGv9/3z8aSOxLP2068DA8wBqqwmUwBHxlVJBmsD7lc8+hw9BYCR2
3qs4E1mJRUhtSszvDiVGvzbFmLgwDYH3k0ohT21xdmON/DsAuvDLsDg6NndnVH7RmXvbxAVJpW18
1WfZKeLoTdkSGksJPLLatDjOmQvUFfHu9MZlHKs2/KDKfpynws/6NpAvudMLZ/0/8Lmjw0+/BAYI
1FSQIfFLXMApG2WJQyJsfGSjGGT+kOcGjhUvv1P4q2jq+13reppiYFXjVw4qjJhH4iNP9inl37Cu
1mMSgwwxSfbDVJA84s+vyVUe/qxD4IvtXhGuOAp7suKw1GANPi+OupQa6Pv6eKtveOTygbwrdYl0
V5+GbfOcMGl+0I8lqSZ/X6ilEMiHvLcpGd0JkSU/UWdKSZCknCjIr28Cf9m5mUjNURz3q5OeRXEU
VZQv3aA+/L5NSVNCejE6KOtvb+BTUS4uYOxmlMPb0b1P6KJEGiMGW0qjBQoQKT20OPozN0/gNeZi
lj5eGOAkxWTd+QlOu15mBTFWu3TcnpX91OllEL9dguv792r7z6XlhRizJrRnQPUAl9PBM2LCwh0+
RQe4AAYypRdTN2YkoO40uY6FVUbmmR+hnwpAcLkNXADXUH2xipLxElrYiSbiQcGxsIdpePdBQVbs
UiOFPrZxyo6XxjZbM5MpMkNv+x9HYODObccweHVhLHK80cvYLDXCki5PRpPh4UOXpdf5BPsooea/
e2fnGcEPHP4B5+ca5Y/c6rXHEe3BuRHvwUWsoQZCUXrlhWe8yk1/W6/sSGKep+STSMdFij35leUg
y1thWE/Qo+xYF36suOwhkLUKNtWpgFerZLdEXTbs1D7+5fXLF1XKlp2AAweZMPsgQ1ryhsljOZKU
dZMZbQXiVjx1Jb8Qx6XrZeuU/BJ662o1XJ+LIqRdxqRfezR2kMV4kQ6395vRZUGAm1eVHZy5oE2I
YMRMmngM3hUA5RNZvwmGfF7iWdKzUJwHqoTRgjiGouPG0+jQuo9NAjyOdduTuBr8HkoQOBmVDSyc
eGUhiDZLzDgVwsV5PUAES5PWNTAKLIPUaAd9yZfec035nD+SwWXR1Ycpb/AViKsBSzCtq6HA15q5
55p0gJYh302dIhx9lfWUjcO8YF4IvA3ziACTdMb6KEoNxwDgAm0EfF6iHvoHysMpedsjxA/PgMdS
qhFdLc4CtDsTtve0/8a3b0QHYVz277lPfA4uYlCsVttowjGepKqYkjR60+HWW1Dyl45ugAARsug6
ak5B5erFfbJ8kFPaSa29bOmkOZMYzo3zCIJxljeaZw6od2j1VznMnGM+2DaIWQ9fVwtFfhgyM3RI
WgOZjC1bce3KLzNFSc5Sn+Brv1xE/dDRzxZBqFb6nS7U2zpx0klBjgwsowWbmyd25ofa4o9zw9vo
j00t37uJEU1xJagZgJnAOZoskZnn/Ci+TOtZc9gU1XguWLhQJ4AARYZVi28TC3G2tcQPmyqIVhQe
D0qNzVy3RV6UPUFbCMoQMGoQhsMAh2p4Sn1FUzG5sDTqCT8Zx3fI9jdSgpdbkmi6C0oRwumLswht
+zK2Lk3sv1qpFQsaHnUfDbDnq6YjwGCd0vybe3jUmuIfKROJYz94rbOTsae7LWveH22iUbfVpq9n
xI29H0vzdifE7oYGt1rmdd3TtNXH8fwH69+ZJEJwLZOz3hV4UxrO0UFP26/Fm4vcd2IZEqv9ubiC
Uj7t8flQr8WFBqy4U+HlmxlQNDztJ4hYdX9ByiSVswRp7Bb+abGzGfXRYUZtYvWas8FoM8DdnF85
rIiONALgJkHO7j14H0D1HzjYJ/wG6lL+mJEbW/yl4k3pFNGt1Y/2BuNkzPGVQNTB/bwuO7w/rwLh
DPbBJw5p5FaNwNvBDms72kgIVpNgpzyjkqmOQbZMh+9X8p3IlfjL6vWxUCk8rm16fEonXUrub0sl
MJ5kviIHjuCAXg7rN13HDvGJb7UzmkUMY7uBbNIEnl85/mCHdU/dl+sn9F3BqFs4xzZFY7i+YPoC
6l11eAG55Rdwq+3AcHp8pbCav12z6pqRVxW2Wd3rc6WJmh+nLd0O1JFCKTBl2LYbBRAe350EnqYP
PO6Nv2Ef5P/43TobBf5E9gvPgXpZqEvrYE+AzX555+rRO0D4Q8RGVnDDuZHOhH8DfN6k6vFR+UFZ
4xb/qiMjfhYTRrPyk1GjuavKyyc6Sgn7DkHyrrueu8FzUwJwX26h8xYfoJOTQivZbDYNM7dI0B1B
Hy01UFlwVhfnTp9WFXrum99fDJja6tALAFUTnpCEgFase2gYSMT2EWiHHIqzzTwFiDsOmKkstffX
36Yho6TRzQQnFg4N4FKvE6vf7QYATbfqhWvGawyLqeCbveXO+gdL6Ru3PhVqeo6VvL7BDYtWD3eL
0oeCLaJsRlrFM0CAgv7AJgAOOrgyptWs9r9ERGjjuWivHd8rsahO8B3eTRIW182PixHCgUWQB47p
rsl1GIqASsMJQDrU71Kc+TczFAeNJkdaRCCKK4NOWau0NNqmcZW+Qt3lE9m2mraUufV2rFvEdW7u
CIfS21akp15W+iAfY1N7UCx0wEkyLEBEqL5JSpEYS0mKNQcINzSC1tXhb7qPuwPG0ANL5cD3xmEG
vnQ3fLlBGSXIJeiQPklMyqYNZA/4XWkKtuXVy4cmowKxoOdIncd8szqE3ehMnwZSKKyTFHULwjwE
/DIidxaoIuUNlhxIe4gmdD6+Qs9MorLzjv1gpXjYL1n5ckQBrlVpuzf0NLwxBTGmk3ZZw3N534+e
SUyLHhabWycYMy7FsP2AWLZzTxZj1ktFF5L6CxZISrO8qqtmUU8wsJEU04DegwKHa+Tg1BPwTmOy
C4ahy+FkPbvYB/RQiyFK4gy9l95IGRTrLDqz/G/FrDEfOYDQpPCGKwiPg0emsUw4uxRcDQRQ1CkJ
27PrIndpOscrEsIJO/+yEDnVbTyCP2N3CWSqci/fD1xZjPz4VACotNPZ62KnXB4JPYssDqToLroz
IbdgavA76TRg/4BZKUERUqDB94DlgpdW2aACVfk1fEU0AE9/sp0QtylAI9MEpu3dk+vpbMUfY1M1
Wc7BGSDVpXPAkJJPCVv2vXp3Kpt2tLlGIJE0SFmLr508y0cdHIyOVUJZXyGzerOtQRRrP8e2BRwZ
1sfThcaGo+YtqwWkNIjClNHJoc62/1dP/1blkCBO1hYQaYypT2p7SrmKfKDxXlSvjbM2vTj3u3Ba
Ked5ys40T7J2Rzf2VuqlyUnvyK8Ux/E+kGyuYk3X+GKmYfYq1wcb4Exj8UIiIhg2tYA6FQ/d/Ma5
SqYZ7eBSZ2sAZWVkB29PXfbPgIby05tOjXauG+x+Mvhx4vNvNlsmtI5NfuB2VGZAjegCrwCPfq28
hmhIzAEeVzRdTPnnIK/B8po1B9dMufdXjwsx7Px0KXGddCBSdbXYU1Z53QnyuKqPj85bTOoVRZHp
gexv5xn1VcVvRhkN5ThVeiJhHkhfcVFznbzSHTCQgDdonzuujOQMYKG8IaCbFwv3sWs9PWTqQfwq
L/712Ok5VvS7uPTh6UGRSS1m02eVQb3SUwwLKZMoqeZwS4RciTJlpG/0//v7SWPC3ufowr6caEly
oxqmLJo535wci2DRizNVuaN+gKBNSv35ejYg4e/mdJD6/V6rlxj8EpPCbR2FfGkyaRqCmFDWySMB
7Y6GmyIA1Xvmjs8kd4TP5DAAZx/SHlyuhW0+DreudBOCcxtUgG1x8MI+Hm216+WbLmw7+zUpJVwZ
BT0K5ALMSGog20iCYAsQBtXxPx/6VefMReXq/FJNbLSICQqDet7fF6EiP+tumcxyxOkOd+t9UEj5
1UzfUD/6RLsaGV1DJCWQ5JG+X0Sb2+tGJ05Cq3HhTJZrxMUXxJ/BCnDTuYt0xRCDESJlmVAoTA6M
vw6UAeh4o4sk8zecjpKR8LS83YV7ZuWl9lHiPKB45z/g8XJ8ZmI1kZhAzK+EHvHAdFtAs1R1kNXu
Ak8YMZ3JziiXB+js9L91GMaNh9ZMD4Ij5fYd+10ows+ux38gGPzf2pS0hIZA8tf0ShnuOj/KvJGK
PYdmQO1iFsL9kAzh6Fty0dGu3d5i5tTrQliYN5rf05diWKzSZC5gosTvf7ZL+pZAj8B0zww66wq7
aGQHkNPHzs8mGMqWAujClSoZhgC8TDmNhlE805NF2PyY8jO5q6jWiMszyRfyZVEsbyz2fukEC+th
mNgooIwk58Rz7CgwWggrDaD+6K3i9BPhmZXJz4MDSvl/HsiZqItzH/a+czHsbMsMDHh2MaTHdeT9
NqKBbRNsvIwlDNKz1hHrRqUPssFoCZ1KgDMKqHJGdcV2P+F0CSLC5/enFWSUEar93ERmZrIedSbh
XZ2pbDSif9ja4b5y6LrYGbbUi+/YE8kgkhvl28d/S/bHhA4NBXcTJBMwRLRRa+lWuYkv53KqCfIL
fq+WNoEvG6sCygJMC2HV0wCyxBzuYN1uKv7HX5XF+vrJY2+n3ZNa9Rtt2bkdphzHAq918NZcOnVR
KFASKbMpLUp3aHI/A/AIkWkBw0MlQf7CmD7yInrdyvc9Mwop7A+LKvug+wiOaBMyB5QGJvQ/C9q8
HDGmV0p5CG7jMZ13tPXUc4ckVuks5n4eLIwSwPpL9AFMY9w45o+O6n2hYOZzanG5wpfpQoks2uy/
Ehrci8EJ+o+A9SDM31cAekvVfWHcRWLom0T4kKsVLqwtp0IHKaZ3TIEhjl0PN3SiMAlRBzbu8vcy
7OYeb11VAtNFemvRV15wpQeN5KdMYFkVEsDBbzXFu3fI8p0ERTNRkgor6TTdmsftOVGbgmJMtZCc
eHtz8KNUhpgEorExqB7axXak+x0lza8Yih6iuUBYX+nUmvf+l7mzjkVYlRTZHmWdQ6KXPrgN3P9u
BJrZKWqthNKuolPVfJcHgw7iK98Gduxt4n1O3xW2vgjtbOtalrKt3TWs35Bw+gL82SnXo/3yyspb
/5qOPyiJSqFyqyJTvtHbgwWDqfQnTz8WI9xdG8RPcY9ADEhWiAXdFQAmlDLGF+veOI9vQAtpk1xu
Iw9Pi5T6Ql/WXDUxBUAyGeCnVS/F8kgNlfM5qajIETqtm6evuVQzNOx9L0ROdyCSpXaESbRg+S8M
AzUxeRu4lnZ5J3myBykp2Yc0mZ54FTUnd/bc8LAfi3BxbLs0NDISuCTzr1P9xY54zoN3HsTmzZHk
VEkHq/0VKz8DUBIG3uRjZJWcShaTeFMy09+0aC/Ta7T1YCrNkIVr2x2dbbHM76BXFiomjJEPFOpa
5pnDxLJzbf4OhKncgQxX/DHegLp1k7n7U2IuZALi0bIzb+1I+X4pqD7r3QGO7Buy4QEIUfTaBFNN
sC9cHkD09qQAMGQxCQ5bxtLSJWuonRpQFTIzbUd/OTmB0TlMopZgoqi3EtJQRKVH36quU8cn2A38
geMFw9FXrMPZh3Dr6kNiSP0Tm1xdVc8jv0JryZkPXJEfiIkh2UspEuDEU5WLGHj0Hmz5SeGJDBX7
QdDlNsn+QFDMWdSXmg5v6B0QabqP0tFbjjQDHNbUMOhWRCW9xCNAIrNNdrE1F885g+gjJZb0Hxm5
7mvnItruIkKLEQK++OSRj2U0AGa/D3orQRg9KXVXsjQfcIZeA1ELAu3hvH8YuCFewJIZqgejQmts
BPH0TcJdOMHIM8DDSfjbbPCLKJNg5H6iJH53vm1U9HsWFDtqZnpLfIMNHBLzN0etPDgpLA1jbVXg
/FAUzArKytZMWHOCTDbjMPcznn75stKqP7DdVuR35UlJOKyiNfmKKu1+nRCfjuHY6R0gecjE4qDo
RJ8YEapdtmxSrBgkZKJ3OeEnwQy8D9rgKwE5OQXJNho2D6VIE6JjBcf3qXHqqyU0NlhvrLTKpejC
dKULOUMPijV9JTtbgqpAxwSRTH98FkWHv3egGeeSbX/fCKk1n/eyZ5OizKb64KdW4u2fQ1CncGUo
gaA2txgMFfgRgtFf87PzlnmHZR4WhQco05vfgfFCr1LjzBgo9CmdRpPM8vPTPH5HnbeWjGzFCf7w
oNmxFIXniQplcVc36zj3d7VpKj0dmljyqUxTIm0tJLOhQ4lp2btQtQFsw9nNItknbB6kHE6aFYJX
Nrl6pfBLMMi/iOYPXc4sdCTHtdMFJfZh880tiCmveyRMAnUb11+Le87x5G3rnIXQwWKDgh3xs8Ge
g2tjdWJVkkkfg4h0YSkx+6KSA5Ad06IZRzG28TNNz37alIMHJRigMH4k3CZILe+AxaPg9zsXC2BY
rxKDRtlWaYipz0x+Op8gCe482mCjFzmI53DZM1vPdYhwqSe9KnNSOZHKQDnIcCBaTDNmwUAfAY2r
5xO12EPdTsMMCln5zXdnFxUf4BE6rEb/P+KcoaTaSOGG4fiLi8GTMHqdvpORieuVpz3N54lSf50X
ASJXxbO6TlZlR0lW7NxDQHCVbl/2wQyL3pi1vBQ6hB8xUwREhoI1kzWWjirgkOpmVYf+9Qk4pGa9
t1b2Q6IlTb7mMZVVGunVCLHhwGCoH+9Op8P+Thg8ouT4WipqwljZNDW0vQYKsTUAmeOF2kT3rEp4
IPuAvIYv1JME80U2WqcP+rK74GZsHU5PWIlBlK9czG8ya4NdU0R8UkPF4O77/6uzLJAUT98DVJor
a8osXyKdvpJzWWWvcOiSbW4rWMnRw2ZJcuH860Ptd0r2EOW/s2xamY9E/G9EgyNXikEQ38+eJbso
5/PL/4CnxUJRnwK/kypjc9mFYj/gULOenWVhYRMEVP1cR0qruoEVGJLuuO1WFukxVHmw+WCcHAlC
D8PiByAQpuXFapPnYlUo5tc7FQZKSOEurmM1mOye5oewhtuHt2FirGR9syRuGE5groT7sq07Sd5s
xXCV9WcvfFzC/Zb5vuoigA1gvDHunxOe6awPtUkUsMwD3tiAZP2hWqGtwTgG/DQhUDgm2D7LdTB6
BdTDWlqFJVtbsUJ7eZbsuKpODcpVUfB+Qmd/yYuXHxPipk6mSXyGp2fxAspecEpH4MnyYhPKQsYW
xuDwKhn40BmS5GbCK21xWdSLaGoGto+RArQqTFy1lO51MrHFuL1T2NgREBaWn8msiaX2kK+t8BD1
6OqKrK3Qw+muyrgDx8u6NmiE3Z4pn7e6jCPmU8ErsEHlsSOqmFbyGPzsq2GKyW84PVphnNXrHwBO
ajsenqLlp+HabDFYayEu+xBCjF+lszr6crawI6uQmp/gtVGQv3wf2Oa4Ke5kwfq4ujjM0Nq+gAMH
wk6MinTiLVyP8LxPMMGn/1JXnErwM5BJYlMZScTAnENLPi+6LZPp1xB0Dx1b/gRO2lm1UvAYBgAO
/OnJ2uAlAkeTqR3dqPoaK9zHHueoD70pEXP+/jXf2wgtSjXUr5kYoKMETkNq0S6wn0IHnzutY2YU
sXu71CMjFPvg7IbqFiif3pMW/O1at8PWqdxZRzTNVjdEwn/04XVIn5HP2eUKXwY/TMPOU5tEE+P2
KxRfeWt6Rb/OqWcXtGr0NFsvJwwpATtyp1DQvVSkQOoqSGgOefzDuPnS87wrJW+VIGPnP6NInVUH
YMv4h/a/pJszNQlS2RQYO3JSe2sKS9VtR4OPWfrXjmIuTYqxgRI+MkK1DwcmnLWQ4ofg1SUFv6t4
ZJomNquQuLoDsGtvdh0G3+w8M1ZK5Y2KYZaX2jIX0DUupYZO2F4DnySZhmvke4BtR60IyTDHyq0s
Zzk82uUsbrdQuKLGm/IYGDEvbZrQBuYR4rhRlCktM2o503FGO/tnoDBTYMYjTS837BEgQvisNfyj
5xLBhkELHxyawng6JcIaDjinaz3Bar34GutMu5w2h1hlKXemUUQydaWkz37c3AP7rfM3mJRcqHA1
mtLyLCMyu/ZGW/ENGJQ6fb4L9u08BaotITQinHhQ48py78iYOvPnid//2pPmol3os/LFYVwse53m
u96F3jc7DoHd141r0UshE6AYke/iEtJXmN4Scxkizgds2aU1hfL9zCWFC66zjZeRkk5HYqR7jifr
ZqnAhaP9/x3Fi13EDSVue3GStYnwW9oMoE1PG8vd41dE0KWP3h5JK341liONszcHP0VuNzqKjz2o
7vXrxVej/Lg3DmzAVjw0HstguJIXSCkaAN+dkBnvgLiCfr6bjXoTD5SE4am/GYdaMM4B9UA9p53o
lxjgkTtz2ykYfzcINvC2sUJykoSV0a7QQWNjxPEKiWa+OrdJUH0ef1EKenyWthIh4XblEN5JYJgf
2uLjaGjuIfvxoSTSPR7FjXmBZQgRuuiD3T1Vjvyh7k9NTjsqUdIDuKkujI7RpnpOaxA82xTjPP6E
lBi3/LT5HY2HwkwEAIDlfy9E1q1ssjtRiEwUBhME6q0RLiuDPLMWFCy/7CW71t09eOFD/3qqj45m
qL0+dIxcryxovXproqe4m/vmrj+U9nYLEUR5wISEJghg5VBh+uT5hpqyYu7AcUum9jBXCLg04xEB
77qJ8KCiiDdlsZrncrnubRHHIHggtJW91dWSAm6gdM7xmav39DK+d+V17VQu/5eIHqI+VNTnbA/S
YzzBhiW5f7DE7FkvenWh3QjR+W2Pv6+R0p4bSAmfSpnComNZC7LHG1faeGH5Ab8LpB8HqHQQ1OmN
0Qye+eiQrKvmBSoVBz+rO6FBnWJooeQ5Kn8Y8h5AA1QtTbu1LLtQeDWxpL3CdWZ9vYDEqyG3ruFf
n8Ez+RcU8GWE14essGDHLBkyBKi+KewPx3NvNUhFz8k4us4tyz9Aig9rCJreLf0f8hngB+zKnQ8O
pML/bOUYLd+3ruOIY1QZUHstI2gt80yebvxFQDQ8WiUkh4JM7xpfRTapMr3MoPsYxvT8A58xFFYk
Y2p0YT1OQ3rd2N8gwqDkdzAxp5QDfJzEjZVbhfjT4Jx2L49WJA06gB9dn11/3spZb7CDlnwQ5h8E
lCmNPrVONlXa/YaYffQMcBto3Rq0NzYPqfTQl+ZBY7XoQddP+c5QXY+/b0b1nd0E9tLATEyKamLz
9px6guv/HvZG/Z2kywiD0577Oog1n72CWER4YNmBop5Ssn7y7K2nJSeeFh22mBqsms24+eELzHaB
YJbGqul1dOI2vKDOr3W11MVOoGI58wAj0d1ue4mVdI3VjqhbunJ7vNOxmrQA4XwmwcS52T5vSwV4
+KB7Cstn2lQNL9ZJarZD3iK1NxGzrBK5pDXB+zvsj204/WVy6wvEnssPZMm0vJPalio9i0wUpEKe
raCm8+vmAkhIft6ZvBoyaBsRawxyiWiuv3TNpkid0hF7jCUWT70PjGfVtil2fjGlDfoab49OKcwA
5W3HcdVOR9EY32y+0kI5HqRafaVDSx7MB4i09MJo8h/KNl6/iOAxZxk0HANmt23ihd2IxdL0csq6
pAnVqgBkCYNNMIcf8I+GWxlNPHXMPpGWWnDs5eG/nuKilkibS5AcZNzcWDCrPSLcazFVrdwMPNnm
Xufa/0FBPzRc7scP19cB2tu4GcLPqC55SSLT3UtU7GS/SuvG2psB2KsM539ImFPTNUEYzxja0lIi
OHp5LzO3DppcxO5eAN/F416YGiyQySoOiepnPu2UqB/Oj2cawbPl0qmFBzOFed/1328XTdKiojs1
xAX9ageIEDkZD44lIOmEOygPJFdFkrI9q3rac9Cm0DXE32jazWEnM0tx3BhPAVLCIRmHuC1tswKg
DPrDBnNKDUd0s/7SDoKaQkXgvDQKddNPbpVzBce9YxXl7r7AhG/NoaTOcZp9xMb2GxoWRuOy00vA
bcvq1akJtq8uYW2+Z7FYWJq2L8zas5reIhDZNohWS/rbgX7bXLgQqvtWMot6vZ+ktX06olIA5sY9
jn/sy8VGnzDxzQSrqsMZDB/DN5KR/lztV58G4gze3XSlFYzVw43Ad7mx7riNIn0t0RLo1SRhwY+I
v5lsdhrpZu03YPGZFL3uKyuOHdDnY1Tv4Gj9MfQDzOwZClHSsA4hsrOCwf56bERS8MSH56L1xtEC
H6lAtMDWzKimCl6PLflxO5riBqFBNOip6trGzsdLSeb8m6frJVHh3sJP3l+r1sPgXs0AFL0f/GBT
5XU7sk3u1VFDpQEqeBZzdgkKQLWojkV17s3I+rYv9P9Imk5llr2ch4AU6lCotQwfXECMCCe9vKRu
dKTzBiEmH/nEqQnUH2KzhA1dtGBdCFb2e/TSusIyf4jw2k3c/Z0xcyHkEMs6qTEfZ7bmhfqY6Zgu
fvXuowzVq66EO5HG5XDrFVsvRCaMfXIZ0Q3aKL5l8Lb0M+SrkBR1k2pH74jewrj9mlqo2wfrASDM
SlQgcFApkbKFyVA+zfEkrakNB4KQ6RqCO2jxjvU33Ml4AQQhgkVJHjYNalKPRVXbSBWJpndfk7MA
1CgYE98CHJdjCfTIc101hpuButPhTCoifccEw/Y7vnxn3zxpShWzn8qRV9knzNkuzy+C0OoGgzqj
iVz+DYkB5QOiuDRcK7GkgILH5E7u/D+Eyz2WuZe/zNxCIluOLC+oAkBTAqqdIJlXupoQOTXnK5mH
xERxgUYdRJrth3R798yYh0R0PPAeBWKwFzOhTIFYsT03It6Y1Yn/KoYSdWnaTjpF3shPYBC/0yAN
6C62zNYQx5F0m3MDcDZsb3o8r5g+heaWy5fA8NOCe/yAvWqFbWB7g16HDwH5syN8E47T6C+/hUWv
fRTGzj3EYzN19dS6T7TWcAkXD/58GGL5VN6HQH8ujpAigVg7A/qZoee0rp91N/MRpTkK6UBPG0Dh
kZ/no9UmjVQxRkG6N2AtZMrZ7H8318tA+NaYwl8bLuFxUuz6KITpmKZPsTtYihcoTEmeSMdmuqsO
1HB7ESPw+Hdb8C3pcUKGrWTjXXz+E/O0ljEzvY7B95We1HD4qaPP0TtUZ4Edi4eVe4IKbsuQr5ZB
yQYKAWFdbus7uTykQj2vG1xjZGpmeVDFpxdYtY2511jyOwz/PAG8mfquaH7DU+sAzyeBX/u0Uc4L
s9MG7Ita5RoRx63A05Apg/louQLiBT8axfJ2m2c4x1RTiooW57bFmnu5YR+3THhrEg3Kf3/GtxET
LyL55S0vj9flBpHjM/GYxpwlsK0/+8ChxM3acGTLmLXiywds26zrEVR+Vs49Dd+VBvboh7ooOvGz
sTGHikWrQlCogAe/8SeUbm4erF7eDHVnCjY/LDLfZGpSMGx8cdxTcqvBSFbq/RrzIk/YxhRobFOv
974Q074K140QLR1Zx8NUsLYXueoa7jwDhnRDLrDXAwBq7hYdawmrwyRqCJoZFF5560vTY59FnWGi
72TAJYC5YpYM1d2IhJytkwiPydR/05MAU3ZgMs+Q+YeDY3j632bqHOyb4+V5v1/Go7kIRz48Sy01
SrtorAfl9fQ/KRBHPAjR3A/k6SL4WYU4X1Y6XLR12lHd2Y6c8jUw7v3hmmbhhijdpMK/Tp1SE0Yh
C/UyZgPWnAMX7jmWJCs7uK7IgDg1z3rfHWVsb65VLiGZquLJTi8oY1GzkVAV9m8RR4EaC1J9CNQ3
LXT/Xz8Nb+DMer1TjNxm5b+FLjhl0ZQPDsjXy1Si+QtaWAhlP+4uKTnyLc/4pFUvqyuw+m1Xwlks
20ve6546KBDR8U/EpP8pdIjuGRfmugrF4YvMxQixRCw/ZH3V0EGV4dB0I1g+2+uUwHnmYk8oe2JD
qPDbXLprGzNh6xzg9VIXe2a+YE52NZKcgy5KgKTY3jDndxI4UknAa9N51HB1Mg2PNk+7VYchKkxp
yGJHyBQniw04UfkbrvwPeO5AAaprCM+lNVje+oTvkar9UQNg9Yn/JHRN0wK8cp9JxD6u/iurheUs
Swb+szOAsJSDU3TeJcT/+JFWptSThcVv8qf5tySjFur7bfJmgtWFjNkgHpqYDAR4tWM1Hw9dgw3g
7lC7rG/iZhDz91xhhrbq2GbCqyRAW1kgDAhCFRAik7NKkYCI+R+hceid0i9Z5yeGk2Jfqmiz7Sio
ahAhubAVBEI7hBQX8nAnkYEW4DJC0uFD/ODNxeI5nyvCT84WSru2yDtTtapez3tKdYpuY9oq7gJp
SDmNlFydFKEh5bIVD/FFJ+i93+WArt37UVXMn01jRGICUzO67MaqQsrOoIlCnPVbwAqI38N57A3b
gqyP2GLdZJkdztUl+KbRkmhQl0FDEppBrind+NCtUnlVtkMcN5FuDKHfi0AoNi/x0k9pFuNCMEui
tjGYyuh0Ey5qA89sy27CXfDOiOEIvDvyOkICXjlqVJS1gqt+U0kFh5/QTEVKYhERlqOgFQ+RIC7e
CWhgtGI5TpcRNPnA5STdpfRTCLwMUReP5WEwHbETkQwz/Sz3q9dk+gYNKR4oM9iIZJnqVeixXwMi
VEf2ZqGlR3vUvYdZjf2Yzb/2xHIg5CfpUuwjDAajWahJaab5Wid3KygOz1klPNAy0OHXqLJszmcs
agVU/z4ufslGX19+VjaxXk+YhDDz4gQtmgLaXDDxxoh8Dd+b8FTGwcwxp8aVT0ZUQMA1QehpGnpT
UM2koqT18dzSBY+WBVbEu8s6Vm8cVJeFzTVf1omjmT72zyxi9NhCUT+v+J64+bwEgwRuhDcuOykV
6yhQeJMoGzAbOABDwJgUjAJyGvDgPsAEdjYrJnsHbFtpKofYsBk5evesBGuBerQwwBaL/I9OjQyN
RiobIvJUAWmHC29BfY2k+SZqLtc/b4aHWwKXyQtgoGKjd6sELIzHy4gBD9tSGYeY15VVeTaWfk96
M30SCaHbX7HekMJ498Xz+DADV+lLK+YR0A0hHgFACjDfrxAT98BwBCngfj2h/rqma/6OQSdRu6ts
LN3KzqyVlpm9fUJPTg9ypGdedoGBQ8arBJTLBEL3xyqKRiHzZSyblfFCnWGQXfrUr71XtQGvfQ6V
Ife+G82LdbR3GPBCmQSn0NCBKDaZYk4bARR24ino2ctl6DQZJuT6mthk1ypPKwXEp/Rm5O1775Kf
/tEMz6YuyBqT76vq9Qu6U6WkXlihSY4l/nzIp/YllNXHhIpbfOCwHEJSFGM2kibbgVG5lVeT1jtx
6A+6iYE2F2jufOKG49w5cl5kWBS1Zm95z+cPNdaKHu4BiDNvZCUKkitZwWTuE2f+qjJ4FB1OyRdE
esrp86MIV8wduzCG6FO+3I/ogYGUiGEseqtOH1u5mLAdVfG7rUFwNlXDtH/PWZbNP0W1A06yh6YQ
sVQ0v7CvO8+tDHm1IqnSBXemlOAQc4sIacqplV/gyJ2fwcktoBSXgzNzF+9iaxjlxc3RaHAPcFRA
7oJXMsKiato2PmbZ/1fK7OZ6Uh1B5GLxHMLQIzk9NXjXQY/u9NeKkWiiCcxFkQzntfExn0Hi1mvh
9vouE5iLH+jm0jpxNs2i9TtuTAvMtVN4TuBDLEwqhVjEhPfwny3lus5v4xtvojZ6B2ICcUhhEhrq
vQaGR6hAYS07DhDwoOXIs4TquM8+u5OnHn5uWVohYxBC0irBwWZWJZzXhj5zSc6iKQ1F0rm2fY9Q
/mOGSIft1B6XAKQCk2Vv87RE6PgD0FPFQNA7xR7kNFha5gq8M22dgM59LOFKUYdLezHwCLVSdp3S
BhkP8/DZ6WfcjZDlYkiv7qWdNL0ASuOIqxVa4hlW26fNUDemBfQq3yk6CKh3iVBJYESYr4+irD7E
Oe51xQOyw6mU/LrvKqnfABJUknooRqo0yEIXejMLf/LeqO6N4praoMxGLZFPHE3qsfzUkQsbd8/s
4ZdIigW03i0Y9nF7de+PHqs7TcN34yIIxewJQjoDZGnHEaqaEOmlVT07ahWP+rb3flTl83DS9vmZ
+wdRekLXcM6ExwjAMQZS2Oi5G4ujzCYZrTQUCe7BrZakdKRruE6I6cRKoK1exnOWs8Z1H3TU83Ky
QNpHSCnqt4tm3ZNHYLd8gq88Nx7UDLDQn+aj42eMwDNdXibnv/uwQse1H3GNDQ7E2lVfbMxStrzg
a8dv+EsmWJVaXbIsDsBl7J7JAfhdd3bED1ohKuLfBXTYQQ3RJ79yRcW0HyOHnNBCwA29EqGWAqK4
J8ZWDOlp7fBy+n0dtA4s4r3J5icYYaQDiUVC87aRsHTy/CCdQb7fXexAHPDhjXVmOf2wr/D0+U9F
g+ObqcnvwJdPROBF2tf7Oy4CpxK7hmUr/bfYDBBUdhUGYtF3ff8jTbUIoyzXnKu//9QxBo1NZiME
I3aKxjQT7ldW0kg1MDvGQU6jtqMRCUdWHOsQ3i9kkgqv3NvAGLSN5KDdHHgDZt6YX4Nyafyo8khP
Lue1ja6etHwhBPomvb7NQp72RyUmwCVnqeQnRzqRViyKw9YJk3pNQLjfmOP2MfgU+ucWgT+e2j1R
TaThELHujf4VJr+AVdmHeW00rjhlb4r2zB4twGah8HRIBB4EXpR2Q/2uRnow07dVJBjq4XCq/7le
IVFFpVCrsrCtVY9SKT4UmwG8Np487FJ497+Dl+gvaJ7Hz4jEUwfLyGG6calV4pdEpLc6h9HLUfLO
26kuzNu8lzR7PDBKkwHVYGuZcYQ3+eUUQFcjyavlDiZKISSk4mpx9t4F8vXy+iX7MtOAuElGyOV9
fuqkbqOjJCHV0EWQpthGNQRwSXfZFT8k3OMrhcDkl/3PoXWqYz+wrsHzx/lDslUaRojOM04BaJpE
+F9EQjG+cNDJsQhspU5N7WdMtvYK5RWsxOFUs4pz12UvItqBk1TfMKoNvGeHDt4MDYuS+smMeoGL
3/HraSb9CatF6roEFyjJfo3+xP9rLp+qGWQtM52VounQ5gX8VeiN+UmfzSTRLQ2Cy2Q2XKzoTF9r
Go3tT2W9Xz1uwCNz7UHDCc5+ecdS1JljkGVEx/N+KxDQpHxk1OKdmwPJ0qxbX6y0ZJnquEJ3+mgZ
OG4E4fxtUNPa5Y0Qrq089UfYwPNp21HlRDRGLMU9R1LFN40XM88g3huxlD8QhnLQp4WODC1kCfYH
m8fYyjn41rAx+Ay0sPS8VMYGboGPIUZO/UaWrxBTvye7edkW+0JNM3tmNASdiyq3UAnf+A3p+Bzg
OBgkqWwHWc2zFkZ97NwXlZSssAkoEKeY5MPBGKB5bxZwnARl8CE9FUgzuhC+T1DrfJBnyhFXlvtN
FD6g4fadMmBkesZZAW7cmGYpWm7OUM8qZMffjQWBCPnlKM9LQUo49n6TwxZEAOJI2Zouk2qqWwdB
FT/iPeVxmQ3vAsr1I22tCKPEVpwMsrgdBCOzLEpxa6s689sWTikbRzgTBgfUDcJZyMJqCjEB3jhS
pC0lmV8Ldm3UnitEmWMWn2O7YLOiJ4nFMR3/NYACg19FWB80E2jvc5l5lfhj4AOyCfqHciHwordI
u9YgSizxLO8H8xz8D/krakYJn+okUyva9954Y6uhPnJqd8aGALX9Dt9Mv313RF8kvyGefsnhnWXY
aX3uYbhu/Eyb0JEDxcy7f7rvTRONBLo5thuzSprLtRvLehp06JC82a3ug2y0sMwOBib/W3pO9p/H
z73kjQp+t80QfIbqms+tTE4LGMrX1jRxnOTPKEo0BGHUm/yKPn53GaZoWauNCSIPv3R6l3ap11FX
feAVzIu+oBKnxjfDdDP0Z0eBA2AAI5gu0A8stv0mdTmwCjtmi4v6ou5N3YP0dzel6RGo2iHeLfxu
wvKbaHB5l4hWvRY3gVL/P33p3oFkVI3GgXGScYL31iY2pG4hWv967Iz2KVXic7WLTSNajN8JWqmq
j0TnWLKSWY/mR8rUYpIpYShtOxxIRB+8SurNnM0YKinH/9+stYULePmlMrqfPJ7IJn3ussXwRzKD
7+QxGUNS95LGEap62qwUZrKi8Vu2+YuT49w7oUetDkHMamfN5JkxQEoe4TLR9lGFvDT7nddN1oA9
rw9tUp6zj5SKHYZxqWmK5aIbKPEdeYCg9xNHIh5lQzdyp0muG392FpnoMFXRk58FDOFDgQouPsVM
mzwU6jBliaky4QNc59rY9bIRqAepSw6s5pjVsQisZei0afYThuCZtjGI6DxuReMGVzVp4zFPziH9
hYHyDj3JeuRpbfdbtGdP5K0mCqBzWxdS7PgubCbA9Bd/c6VUwxZvkk8jRUMYHhnv+nRdk9zrYKrU
TLRwpDEvNdlSveFwwmDhko0Qrtp/vUjPFCR1ktm7b7bftnJM+4hT4Rj4ze9DsJiRCqUIUk9Lfd+x
/BhDJRF1Nx4kO/iC0xBf3BirSjgF/JNACHaFdVbIc9wfzNSZQNDX8MjdSY1LdO4IKGIKo1p5/sHc
KvobKsJlIx4rIDEFzSoR5uKIW0CLVXG62OVAdexj5dTHU5K0sRdkjnXYjmhNbEirhdKu1letYwGS
aGEj/qxQt+fP7KR9WBYhwHaxCTH5vQBK18/3PpO84z8YEDfFAJD9FQeWY3yAXx5iNzSJteqUBhzn
/CvIIw5M2tqaXdSjUr+tFlbemBK2l5ZB2RYZFGu1OvxYpiCHvimyUdpfzVBVkyXpyYB/IDN1g/QH
8PIAi6O77qNx3ap/vjfgxpFsS8/7gsZi9yjBPpXyDgyfWZt40wOYLaHzfuhvJZjUpA3cjWGbHri3
iKxNC1SGF14h3880NnKJVrYEo1Q9PQsvoO5prqlLlsogSezTRX/ylYqRW3x2pbTWRWrWsm4g9rsp
Ck2cmdFgWTyDFsx2lB3MDcbZkTB1iJinH5ywN/9Z3ol9I7doSKrh778IejtVRyPc7LZkeaKLNv9+
bblXB3LYA3vF+uBY2wOkff5jstUHPzA0o4HvENxlZbbePOoiywRipAPzWwNT0tPzAkPgYyFgyx4J
pD9ploYHx1yAMTA+aXWbBWN2eR3Txt5DyThR+GFT5ONuvT4dIALDijeFwrU25NiMHPNKKe+QHgDY
nVb2lDx/L/iYnH3Io/swyAsaisCXE07QW5y2L+ETyfnY6f9FYRulXSak0KjLcZKCSCffZEIvIZdf
eqFtuYEVtGaV45fFnfQGnBE9TC9PSGZ0aQV0axNhz2vRTx7we7tG/CImQR+SdNZKn5G3Lng1xctB
ZkjrqwsLUvvoKdgbNAY9Xlq5KMuiBLkgofpBVB3PP52Q6JzKR+9+3oVrtBAZCnfRGZwk8PW7ZuK+
qUTPX2ZmILvnj6xXcw2nlDmp/IXoWpBKL1vgUYG5a58vaevLNPRtQf8VrHP2z/hYeArLb9u/w+9f
kWd+KA/BJTJblVGuQ2m7/zM2PQpEmRR8uEwJgOGU8ejG0KCjt4KtvCur7Kw2wXta7EKJ/vAPBQRX
JB6hSfj1SdlO6HMEPmCT5opwIE/x8Yng39URqUUJE7Qez0zO7IjeemWo+cxvrgOphP0rFdx+15Uz
bXdJeec/9K/3naQT+J6g5UKOz0wzg8xUTq8i6dwlPy6D9OQHvNgl3TkA2dBx9tMqieOpVNCSJOXM
zjEhpD4TFqh8qCisgnSTWnEiKP8k0PpOnuCrvq7N1htPVXIySBi6pPvMCBM7dEkSsf8zbjac3xmH
IjN/o5MxVj3Jpam9l5zJ4GStqvaHAjJxT54WJMUPooOPqQgwfVFpLI6tP5sOgA14E18w7vNRChat
scn8lCR8H/f7LUGsdP5i6vsz157/lYRca7bosC0cTvF0rmOHvQQbQ38gaVcgnf6Cqky+8px0Y6oE
RVi7l5pREVLzZAbodaywKpWkSiXgo8vFKYriWRsxgUcQdqnzWu3IsI9fqhi6sB185KgOyfTF6NB1
paWUBkW/G3HaZkEoxIIqqkBzZ1gq/68kHa71bWCESF3pvcXwe3reUJ7klUPwnGXM2uFYpLCltwkn
nGdKBbYLMN/9JOxXjh3HLCBHZiscVIwf5YHNxwzZFg+lDe2Cyjbgr8AfNSU1ia/eJDGMMG7oT8K4
z9WC20Si0JeqUi8QjvMF7yqYIsaKYtG0fDwzAuw0FsBHR8alDwX7NcNxqjqGadN1mGZaNSLoYXUR
fBQd6GpMj76wraW5C4YdJPWVacC/VdzdFVQOztLkBKLN2Fi7SDZKPQ1Nzja79LcDJ+Mk7V0STgbL
odtB2I1Uzjk0A5ePZ4XBFvYn4D7+jHYS1/WZR83Qbs8PmubXvnEQsZdyVVTuXSEEBo3wa7G47ks9
8akTfdl5RebrAVZEqSB2nSCdtZFR/pPbwS0Oejv0HuXOMB/cdwzjicLqKx6HMn5LqD9Dx9i321PR
SF1b+3ENTmTUG1+Ou7EzU8wj2VHFRkuDSiKGZQauky6Tk+rVvRfJKz7YDlQW4t6lvDXkmZdX14su
DzZtA5YJMr4oi+81YiRW8EGwXBmys6sKwr1m7UzN3sKCo3SfFXyvzAtgQLnUVvcGEbV6VxfyJX67
I0RrZuVfNyxdq30qFZWAshWYY4RZRn3fDakocFokU5jHAFvvV+WF+4SwZfwj/T98rZf4/7eZzTd9
l2mX560aoGbFVKILGtdPAbUeiCnnSYreWqkPwedWOJ26dCRq1OxcaKv3N7NNNzipTcN8LRXhjmyA
09VF10osDKJcKzwAH41Q14/BrUn6aEQyVJqFBuyBAqp9rAzQeOeaqOs7RND+l3TVkUTInKBzvvM5
0MxdKUV8or37q6074ysM9tHJPO608D8zemtcCfiIPBQEeAjzmZqidL3WWwAo9XjuR8gnCeCgVXqe
pBiVpUqWho8kEcPEEWNPN8JfGZNw1ZlKQAzlogxkfotPDZFcxOWbSKGTDUyYRN+SV9RW5cNyHWXf
5lj0+Bng/pYsDEtFmIsXPtb5WZzHz8vJl+0Tr96C6SOcm/ltc4SqF87vtCuEqFnulKDvYiFU6ZbH
aaaLnPgHoU5K/52EICkM++LXnuedDM1VttnLY4Ox5GuFg4B4lGAhqDTt5GE2achT6GEZ2a4cIuI7
8OqQp6+c9NrQxVsmuzM472Y7NrykxJnJVXh+Xy68D+XZOFHTP2VcBT8ZWdgiuBJk/7fdxgkZ+GfV
qBVsfRdKp/DI2U6UV1LCF0qt1T1/ADPcHXdhZ41qjJUOEd+NJVILZkZU0XZ0qhdtQR2AzdBjmvZQ
GvvuBVxo5k0/mCmHbuuz3uIrhDzZNCOpqqxlJNcHKDz3+pMdA5jZjpLhMuJH8Kx5pupzzEmN0Ky8
WmiJz+TPOmeQUy9MQlzMP+pDzIn5vTZ59vRZk10U6il1Q+aRxOyQr+3I3qRUxvd5KDfFppdNVl+w
I4VXOgFHb2C9VtAogXYpMhk3cS1h1p1fTbNxdytv2dGVE1o+j2VNco3rkbrukmoaB2Yqe5thxtB9
Buwj53DyKab1IcH3h4OTxlm5eU53PsqPz6RNg9Ax0jyE5UFdiIzBwW+q18y37LXdX3euf+JIIe/Y
E1245TOfXePWi+sE5LzTEXGMZQ9WOuo8Y8vLyFiytqJJNh29SrjcPoGdn1gNCSBHIGdFrcvCCSzR
fU+8OTKAx3D7O4kIcZpwd6xdLqqKYXaursLIn7YEr1p4RV+rPJ7+9aJ/Yiot0GcEEsehI5B3csnh
It5MLpxvXs0hH8AzSyn6M81XgGiNcKg3VmZGYOkJ12ivNcz6x7k9IRzT/kTCOH6u/cUuyO7pSjB9
YfsSobiMWuwJms3OaC0JSgablm8eEYAuEXolvPGej/K4fTlyraFUilX/ZoLe7ixpAD5CnEtoPuUt
ZpdRBOEthe11A4a+uN1OUXy8Y23VaIRTXk20PWAKE21iQ5IzBXsndzjPeoRtIp69QgMADimkZRe5
bA0riTm5ka4MDCt77e7tlloNaWdL228EIltlCGvF5TLgbmx2HgsLC3jovkyEDUcTOgRsZPXTcHwI
QN+lBr9h2O3gBRCxPd3gGuphfW85CAxqUjB2PWhQ+14LF4xKxiNkNNdBkc2GX40pm1ZG4ri3Wnqq
/VBB2UIoyiI2aDfXqeiwLQz3G7jsca2W3xmwcONyClB/9qWB26P74+R5bpL4JhQmDVfEIxqVVL3X
A73DybaOjOphz98E1Lz/oCKszNy5IWlYZs7tLzL1GTWD0c1LAadOTPnMeCJ6KReE+jfpZpIvkMKQ
4w69Y9H5NgpFd+LQaXaeBthT9oNoPyOfwv+PNqO3/7JYKWKJvTcaYTI1xEDIGdg8xrsFVI8tleTG
+lWtlejIADB0Zb7KnmNoRWD5l5+PQ//HDhWnW1MINAVdo48E+sGCio2yh3/YGpr6P2edgGrjW6ds
t6tVeRaeSjp+wOBpKPhhUa0kitJHZWM144RaO0vKKdpur/idT7MQwEHs+vnwH+U2IXNb3T11jTQP
H8yE1VVwM5yxUsScguGW6f4CjXaQejJAw7I88fkcpSG1OdDy+27x3ZzKfDREyUN0Cjf8z1XO0273
7JwukvG0Zw62m+46ZmIrJ1/zJDeK07tRV+k72xmqO6T2aaSZoKRMbKRpASBlglBm+kzcAMBjyhXi
sILKxtJpU3OitC7BIHGEpHXDrvjpJqeLdcH18dJv6Uruik+hZYB3Jh9ywjYo6TZsSgV16Mzo9zwi
1FM3ZcuBIX3Y4//U0G/trJS63BQwjux2I0hgJBx0zcG9kIDN9dlFuPPLxLQDAvzmvA7oGXTzHCZI
4SuYY/jqvc20cRlzXGDVo4R5Y/V+do5H2VVsNTwBDV+Erb0lI3xW60XTTpkDqm7edfI1nXdpTGxQ
fscFxfOopx7BQrlpTTMq6z7PsTs6FxVFB2XXC+E4janSRJQE6ofPqhMgfdSRYb2MbBr+wDOafVvN
gFBWjO+zoWbrDvnZCXS7aEtUCg1tgOlw0WTOeaAAcYi03174py0LGdp+4RVpBUNEHENVRJqeSRUy
2xUEGlSd+q6icmlgTJZ4r1VMs6PxP4sg5ua/6PMGst4Ra7Xyh4zg/5UfLBaWK2yti9lLCj1CmhNU
Vh81nWuwuDZJLE9WC/A1ZW1znGIDYMnRY5kHa24uBD3IN5lNV3syXHkF6jrqdWSbn/MCvZuqIyL5
mKN7Gn/LRSL99cGmqUISztTQ/6avJVMKnFrm98KQVuoCoQTW+uWNi409uDLXUdHcomJD2YX+jiou
OmVvX4cGCxbRUMxyTj48S8z6rz32sBb7EBtESkeZcde5uGPLdbOitnqQ/kFZumPmUO32T73FxeJt
R+q5Nf1aTeZYnXqPxObsCrceBqgnWEuiWj29f+Lk1R6fxxHom94gWZfylYKTpsK7+zgsgtHj71Lz
hzdbQSpFNMFP9pdEBhLxiOkvcXjYECJuF+b0G/2WkX8cqBzrbZMbjCW7QQJ7Qvovatg/MGSi7BxS
wwesr6rzZw53wdhhjN7yiHgbnplmO9Qp8Zh7GfhNgvlIqw4ds8XizBqNG8DYLtIyk7QmlEITGumY
3MsE3Kqi19m+9TI7XXj2WO0K1pbYc9JQCbw3Qyeod6DDt0j+Rbjk8Y3CRY3bh2oz3nPLehuWJQJo
dGFJEDNC7VaXQdgBMFOCIxpa6QgTaaBR/SPJ+ITsrajx5MiRCwqfpYfwZnxn4An8/e8UcheLBpuH
ozWIEPsWW5yE/Y66PzS/fGT1joBkEdUWaQ3+pKYYQ9JQhOT6xJ3xB6rbA4EjGAyN40Y7MJNSGgP9
uyf8FKbP/P8fs0ExvI/3h2j2fD6YWJj7giS4BpEicANggSKqpHKRSEWp4TAY7WFoowK3KSGiI/9y
MILgPMW3VsRY96FiQ/n5zHxOB5qi65Wj4bXUcMKKo2zh2PSpcKZS1usNz39g8Uhzlfh3rtMKHaYQ
y8P83tKeuxcdDDS0sxp/plH2uRmrmjO5Tz0yuIYODmRVmG71icpkR37AUqCgEZ3VVMgLMU6uwJJi
6i+JfmTBVOw67LNTqgVqS0HSoMqxPDw8lTxv97aeZoYqNW3ssoBxUBRCaCIw4HS6ei9sodVFggws
WtGnME97yba6z0da/dKHEZLpi9b+xqRxeHmtB80USGQWk0JJCelKVyGZjsChrFS0T37cAJX4FYr/
7OVntlKX3P5h+SbJ6pjmlRR7grh+01gaCfu90nfwAvLAphFEFQLjbDfRgJPKrOA2Vp/3PZlG3FW9
feqJDqS7SdeNdL3vR1ZhUdKaoA3RypPJTXq/tEkmthxLMShi1/jL7vrBUmzZtUiJDvYFLNfy4iYl
lamlHatgxLHGS+GFL5aB0N+r5XQKGOd6Zq12jxVlm1jR16Z5OlzWn0YWnWxWsYGuZtTF00eZ2JFx
jqr8kVjqVb7WByfYFufzLsf85odLQIof0c4oqQ9muS9Yjao9xcugcgisjIhHXBKhHNrHWo8vpjdk
5xKq70C74d8lGEqG69Gjexfs6QWhIt6l4W3HyexF/ljA6lTVMvX9kyol05OAbwS4zEQwcqZYKmhv
RxvSIFCzMYdhTQn/bpa4qkVB8grbflQIl6ivuDXybeNEfgnsCLdjrwzvSfMf1Ke4coMMrxXJvSNb
VXQA+Fyz45u+2y7DvOpKuaFDeEpeHnD2/B9O43PMmslYe5OFmGW5qW/3Nv+ppEhO8mB9DUJKnqIR
43NB+ZMwCgZvQFROoI9GMkbLX+wEEhLSODD5POsL6RglHHgwwVA9EqR55WcHG67xwcpNLsX/lDGQ
U8zFbEgoXzVVm2UpKputasEn/RQWv/T1NIxWK+WZz6DHPGtt6m38LniUq2dUkcs8Qq5ByS5sZQZa
FUZHQAFRjRY5KeHDXdEjCaN6DA2wlsktPVytj60K55BNsg6sbAiuPvnBsScw0nXBo3OOYyoxcfhH
D40Wu6PkcVdmfb6W3oQzqiKLdm2zAmfRu1g+jvX9sjskJuUPo8KthBp3e09EyndKrdg3n8geqxet
QiXb1p0xXe65ArmvxPlmcshPDf55g02OfuRBZkK7SogtVV+qyvgH6wtuzr2O//sd1cBZkPbGmc+0
28rVoc9A3PvhpI8r2B/TUCjmyKy6UjRaJd7CANfc0FoZvbiUipjN3o5yAdeFYQHem6XR2yiOK8e6
uSk1X8d+uycNb3xNcYEHz5dLe5y3BtzKTtRRH9ERAFzpAiZ84cRAE7qYUlpMwNJZGjJ2HZ9cPX1h
jwQmoaopWmmz8TcTOvB75y/8cdIA6+PYLLbeYqJ3EVMCDUFyVMSnYn1HXf47VLI2tqBe0RZXXA5B
DONd3pWERVfS/N47BdOSYeatTneU8VhxlNaYUZFd+Agx4gEFZ3Yfp/AzrzTCT+bl075FSH8kcvxi
401/ICvIKCSc1TNHkcMzB6YN/2TuoKvnLzgtc3qxdAGO2bVTmCDgUuzCk/YI8zjmq/5kY200EM9Z
59BUgTKbaMRXgQ77hKRDY/lgRx4ML8wwktk02FiwlDUbqGy6AMLjZwfGXMfOuUbkRJZXIfdXNRUd
Etqs2wcQvniU6jknmOCWgBYhAVhOaz2Wuyqki1nByOQ3x2kqO5FwyfepVsjH5QznxzxxG0LMotBH
azVIpWoDlvdZoI30jhFLNG7QbXusBnAw0uXV89pFuGwxNKDkmrtuyVXStB41+su+h/gvDtbjXnGv
xfAPHyQxaJgqgc+aqdAXX7AMre5LBxb1nJL9w8/tu0B7YBIEPWTsLMKOllt+VI4wpK3vBGv66pZ5
1IVNNYoRuQ6RaI5KEV4NOpbV2I5bAcU9oTPjSjcKIwYpHHm7MbL5yJbt7SjswMjQCjkChrtwgba3
bsGeGUxB244SzMEZxcj1V0R5y8640fZHHz7y7Zlp70BTNyoMn0C8xbTKFyeQ7q0a54ikYSHDmsAr
JVpmJrjgSb6VjqvcssXb1iLrcgvZT+oSMHdfr/xZrd6KOpsN7M9U7C/d/i2vKMkIXJZXT6veEh5b
wWIXhAV6ZNxL/EbqINo/jQd3s3eLuMYJhRxzeI20NdRNNfeaelbYf+3nT9Ir/97osQCZkRR9wLcz
4Y3B7yvFxySL2UUv4gcA8r4iqGW03OUaCvSBOlCWqTrmuaaEomJQJkye0b6FQ93OJDl8Y9P/wpw+
gopzTrENF3TDSI+U25IulOj03v0l8sxBBdXGl4E6gWqEB1SgJ+5sgPpBdpRbDyWz264pnkgBaIMz
EmvN2wUwapiYpBuoPSMfFayyhvNExcERQ0zDhiBpaB/EcWVH9t+DeMsCIwox3KzKpcwRbLQ0xRux
tWgP+2qz/rcig1t1pDfDbabZnlh4JCAj8bRMl0Cmu0IWs8g/61FZS1sxskCzLh9Zh1pbM7AOhy3Q
OPVy87oPkRaKjxNC/kKoxB5wnonT7AMprZ27SqQrh21pygPclomZhBWsWQYQ+ke8k0q921WrE/Mp
92D1orHH9No82zK+Wz3p1CTGis6ooPoXQXsrkBSMtw4M7w59rbONBjUAA5/JNV69AI5ip5fh5o7o
Mu9BKz6D8IPJOC52AW/JHjvR3RvFqYcSqVqGMJZWTw4X2p/3qTmtcPKrPrkzjFlkO4UrI5N2kKhL
A8iH4qNBuZ2YJO7bwCLKNT2D1b/JU+cAO3NIwqoujrTZoJJ5einGviiUC107p2iBX6OiG4TcHoPb
Io8O77jFquoi5I8oENwi3hZvwdrG9hPYgf+efp+1JIIDNivPDmv3AP/+3GeeXi0A0+ZI1ghXri99
cl9SWOeUcylhV9LpH5wNwGECUDvN152MkElf/Z54+cIe6WE0CGomAAhThqcWjLE0y6a77fTteviO
YK3FzGvG8xQNrbOZG20k3h81Hwde/tlY1sNmNjy71q4/nWdYc9O/Mw0rWIAluvzMzgUBQzTr7g+Q
xFyIbYnLcVdM8/hOXNSrAzCo5f1hem0WBT7gnJyRNokYOL1ci/XrDx9r80X7FjUulup3Z0odiTEf
ZX+hYf1GSu/aBffP10Z7szq14CV2vP9xpowH672J/HTahvdPWKEfwCbl4yV6ldKizImLbPCFFuqY
WPs5AdhAbE9KZ0TbyzGHWrtcxjln0LnV3fF+hcnMLCOlLxIYYiItVm114QRAsLe2DPB8uipTR3Tu
5SQ6+yWlY0LvhZ76xljlhVV5dRJkTtcJeBr469YwVPVzManMYdZu3sIflAQM8idMjRc8lV0KLk37
2DDbFs/AsPV6vtA5xHgZimBCeOFsdVOpPsqSxeoyqgNZYRI3uGxMYdEJY6FyEwRNsj1bRNuffruo
0F3zft+gJK6dAYj4DdC8o9gG1bRCAks+5t7CohWXlz60Vn9c2W/5vIisB0fAri8eOuLwCu9rXWsx
29P+7OyUje1NfDiJ7L//nsxpgCjn8mjsgJDxNMqTtz8H4OEK0UvfVH/c6Al/ox6Vf9m8i6Q0NZoo
Duh4Usot1pu4YxygGZS3kc9lQqpeUY6+FsNXtWAt/4JvDsmFXcYvJyvtTDTZGya2FvoDbOWzMch8
qWhodABKo6/iNVbj76vec8JQz4RPNbqrJKhcKjgv62iboq11C7VrM1MW6FeGQIPa2Ljn0lh2mGJR
j514mmO2bakzjbCAg0hQoychHSvVuUVo23BLijH0pj0PtFm5l2xv02f3hY1yA1/ROl7iQXXnSGRp
Ap+n65f9I03I99jO8kg2GnRebhP7E0WpqKH/SnLfS0U35lADP2YepO2v7MAAhUuvBjI4yij4UxlJ
4yiXrW6JncIPj1vQwjLTSz80FNHkk1cEIVFC6PBaVfsSCEj1FArlofIVPhucYi9YRFaSDsDuPkqM
JdvV3Wt1r2zuVtAMlbXtzWNExCe8WQOWIeZ7KiaL3d/T4MggAhQo44l67HBz8GyEbj5dxqVIgVD3
qtoaOLhCdNjpb5azFxbVPzJtFXvCYhfdURyXmOYTUNsGZOKb36WCw5hbK67wzj1m7DrULiIctOSb
PK2pMTDTBmOvBqQjuHyc73fFxjqe5UlRMP5PA0Z0Kb1WzF3f1z/VZkoQQf+zuYmVq+bpC+wDBg9y
A2OD2T035UpbPPjd3THiZ56sB4nbLFivTqWDOoLLphwoPqbc+MPvNs9T/pXxEp/Q4i12Cb+L3zgI
nzyM4BSI5/TscBF8InP/s6JrAnbPl5pDZ2LTYgun6qk7Besz8SQtBvcmyIigjezrstHqUp9snzls
JJSPTy3u/FvB/7tMvbPezE5k7AhbwdGpFbveWW426jWhcD8N2MjQRyiK7liklRrac0fNy9H9hCRA
v4B9Msv7xvQPTRn39QPViWa7PGiSBL72FdDLi1gUxb7+KcZ1bB+i5nSamu/hjr65EekBgbKAEXjf
3xMSshhjBW2+xzHl8XUkA0jscY/GfGFvQ2qbV1UinO0Kn2qO/A+R6ck5cT+YPK5PYUZII6j7KxER
1uTHFacxGAduNZF0Nah6g/5ahQMc8OM6I7x4Jskq5HyN5uhzGb5zZUxvtec/39GaGAjgYw/ZdsY7
QC1eqVAAhfHdM2UOAlsAYd3TulO75lTysA6dXGxt31TKDMrQmVLEoIJID0HFB+Gts5M2HDuMjCpS
9mpqC5m8qTPlgWmWbqyPfOWk+irqg9fXCCR2i4HvRWw2A4B3gBOEAEblwro/ee38YwMcWtXGzu1g
LaL6NcY7mfcrleaZeDKhy+gLZJ+nWAHWm2A2+RBjaN87r1hMzpCqQ83eR8Svt+jY/nfJ7buqbBRh
K+VRtIhoZopeU7LbelF2fW2EwOdlW6E/AZY76/5qHh3AvNfTkLoOjV/h9R3PWoSVeCjk3Ze9RXL8
8BSa2R1ULKBgQSgHenmrf1jvmlLCxbR9i3JWgvwXhVyGklBlaH/Xk1ryofvpTMq2h7vgmf592J+3
HxZ/kOPbHwrulV6lh/hfCh+o+LKm9hp7pLBBtcmo3qvur+DNWZkfoc17bzdYpcTTuh9tz+7Z4mbi
EsHmgw2ZEoULO9PbB8MI86B4UgnLuixzdcQlv+6cBGQvYqiXSpBSuCFwO6Pzm/L/U5c8oScIGk2U
s8k8Vtsj24XcgN4an6HL95/PCBrIU5+RIcxBBoUbfOKu0bvAUdxftw/geNaEg+6Tme2SXZVCJ8Y1
HdohIE2JokWR8OGtxhdacL80LE3YL14ItIVzPZ6r88EcF7glCayChHYac8aTuIspcrE7pT+zSqp7
7oCuaPY5e8nQ7xd+JLqf4e+quJs4/pZBl767PDzzJom8HiBHcKedCK+28jQZuKqwDgiv1FNaFJMu
IjR69IbgCC0yyu4zbSoQgzoHhjORqrQTa7Vvaw0JeJFT1QgT4jjlEqGAS1X8Hvti334C6GJrWQB8
LulLfvBCroFZyIYpOT7NI29BMOOEoOzmLspse5Bz+3SAM3bMmtzI3gpKVFARFxmNOeoH6inFsBnv
DTa4GOoW2pJNgrz7V8Dk7tr34Pn6rhk5QHDXDnfn9HGGPtAGYGLHCwajA+nQGFZEStTDFgYRakD2
8sVUNa0uSAebTIJKhOXQwba2nTUUctMBkWpqLmVJKmDLTWTIzz2fg6tlRWvVOiU82Ek7xsgtImiH
O2JTWrOsYPqOilBbJmNEedAT90l2A2d/UBUIhxMqSVM7TxAhqlb80CCxh4+e3ExzvkveT0uVWAID
ycY4xdf2Zuu+eTGLhWmXQrIiQ7ZLWLMR70/rimIUO6WhfzpVAEDURSLgDG3RrrtKOJu/vtdjGiFq
/pkCEZMr5+IF9xuKzG1TgOhG1lnV00yh1ggw9RHn6su9dUtAzb0ICgS8JHQKCJ7tFBhb9ES98sA9
T5mP60ys780hA5Xy6r4KdhYYI/7WLybnoNBDTgDMgMVAW3lVmJYNpFubM/Wyfvtbq+V2HRaoh+Du
h5tx0IVlwxzGdi8352VPwThO/A0gKD39l5LM5pgd3V28LVzL2q9fqJxL5Rkj1DVOCf9yctLPrGqU
yQRFRrJBXwzKZwNJ8LSOjZhlYZIR2LVlDBYXsE66YHAS99jpICoc6k8craePjkUFPuSrOPknV+x0
INhqc5dh65hCOIMVav5Gmzn5xNyOjmhjRfKiqEGrarmXJ9hBzqhIbep5duOExWfwQa1TKUfMnRv9
D0tych+/Q5vpfBz3OtXIRI1TMa6jdmv2Fi4ImfdNxeRV5zD/9aCgPsp48zjNMpnJsqTMZ6OMuZyT
OjNxacqJTBEH03lvDLwIabwJPT/OIjNerTuSp2ZF+0oCpDmvZo7wrrHo4I4vqC3SabziQ6pP3JXB
pKv22ZRr3pSW+YFZArTDyQTX8ervL2M3YtjcRWdGrfJNLqFq34yhRJyg3NJTEmwcCkh9QmR2mrS2
qNoGCadPkjYa16qXXo3PKFd307qCRRmiSJDAeaZaJUPJe2NIwpZFEtNxeJmjGSIpwNDJPmzXJDZq
7jAZIMDhQkexPoaSGUCZU0/2PcsMBNI8ZijSx/oO1A71h2qGDVBU3eD5xb98eaT/MKZAeuMqmU9o
NINZr/E8D8Mg40QBwSR1Sh4NDfLmd6hpxaYYraNIw/yn10QO0DiqZXzxvcer/JCVpY4Qab7wVvkt
gQc5kqvq1jkdIrymGw3RlJJiik/g0k1/l7BEhOCnAyWoLwKDD+VUvOC9/8uA4pxu0MDJLTsq/RV3
qpq4/ub7nt8nzwHNZjv9U0HmtJgCbIIsc6u/fD+W8hFDvAggKuA2EJXzAqhvChH2TReh0aoevtAO
SALCQi1I6pDQ+NXxhElIw3/oyaGp1cyWw9l8BvDMPbBUpP297rT/k8/sgO+JI3McM9/yq60P43Zs
koGD6SlsVLUByEZFjweeEjC2caug1qHHjoZm+/r2OxKB8bbKM0iTwm2H14qtkyQpocIO27aktQpP
wngmDNVMqzsYMkZIWJxe3HwYDtVmuSy8PNASMX4XWIr6fotUOYGSkP1EZJiCihjSXj53qvtRf+P0
svAnkVu3ipMmxzcLOMWUQjNB0X1DuQv7xvOyofBk843MyMWYkJXfXZQVF8H5lO0IbZ+IPMejchyn
Tgq65sLRwgpeawaGwKBioe/iY6cxajAB+iNkRIxkI25aHzbtCiBoUyU2ibkX3KsBRcSwRA1rKWo3
P91zOd0G24d9gU+d2xYtqlRiDAO1ASAMBDhwEeBbBTluyFfjBW8QND4caHzLNGmV9j+jGR8H/Rm1
wB1Cf4rj1ibpQQmcTmEZGHk9hPQyMPlmHxbOl9Thi9uNegfJja52edA1x5CRm3Q/fYGQZrnDW4Bc
I+I6JrR/+Uekt8FncdmZFf6qYzA/12ddQlfu4iyrYyn/ZS2aClAz3+l1iUgx6Xc2hIPiHeIgYmhg
LfzDwTivfUCRlThHb9jDN3P5O48JlgX5A1EQpFGVo4J6a+11iVr+tMBaTK8xcum9ppTqOMPGQRcf
f+X2LFLRiJ9DVK3U3dbXHtsYzGGs31eNdETYlswVGC7MqJQX+/VPNbvTbEohzP2jKW2ZK3EaC6Yx
W4Im2TbipuAOIY1BUzHVAFieaUjjA0eOCXAMOrt9OsDW36o7cCffcJgUuYv+zqPrvsR9G9TZaBJA
rqfviEgeKgsfqGzyPe7esfz7UiZnzjNqUlHpfkaQx3oZUt8EMfu6KWmihAK6o758ebs7m/Utv9Ps
QO3RFs/sKIBVcPJVuWsPxX8wWkCjqiqpYrmlKo+0hY8aShYHtjxf5Bw2SMu5/Ztlfxx4FmGTR/34
Xsay1yYyjG5kEEUs0k7XhoA3NhE2E3WBrH4+C9kSurcbeq65bk0CHfviBVZfG24ruFifjyy/fETw
XysvDHpsXM0izLYambTIw+YQcwd1GEz7pOjjQbaEbi/Q6Jmtg9oHFJ0jzUvKIjbvgSka6qfsklh3
pPnp5k4kp81OzyviDyu+7mVagAe3VKP1MtYrS4T8tOGCtesYsr6i4dALSW991SnA5OoiWKIhxbN0
MRLDl4X7ihsX/91nh4LMizuEusXPsoLn9hHn/X9gaOSLZbMGbuKJ+eFxxbnQOQP9QLGV3cJDfwqO
gg+93tixC013E2YVGRd7PCqoutEzZuJWACp4iuP1UdYmaafO44nnGzeQUHxuQay3tSObf7A4WaEv
nr8U9kmG8iMYUFeIzCkVNFufqzlUp42HqsbLMvOHkzwK6W2B3CJeenK5OOE1jPIYc5RmVnR5ZltN
oIh54/xiY5mZrMDiPY4rdpLgpFc+PG+IyNcL17RKJOXJJqFWW4aOJwZRDJfmNX2Iv3Wf9W+CLB8y
+ruTsK8s5H2FTHUc6htJR6SmXFY+4jBRjRTsDAhyfU4ZzjJRcoZWvaid19u2WSk/aynWSM6rBlbx
edcl3mVCiSkDp6+Ec/f3Oy4IW9vrIuWfXxtmJZlX7qwwlcs2yuQWDO1qMxWfBvn7AZTS9aBLQhT0
RfFUDKEGqHH4szsZcCIQQcnoGVe6tdMKywkcFFcwnvvGfBpW9fB8Jn/ZAV+ZU5IOZcaQ5keBCDGS
W4XJAdORewVKdidjX2GsSxK9xkaPcuvbmyB0gWBADP/8mK+yEU8qSn+0XmczpBqBgdeT76MNCUAv
DehQ4LA6fqZf26Sxw3l2dRRd/Y6KfqmbGcv3MI9/ICbTmTgBxBB6w873qEh0MMZ4x/gpvCgXnuk2
AKMhXOSFWzra67PFjD/yPcTuvMijIrNr60h5c5qvsR4qJnQVafhxwjE7RGodW0tokFOF2fKbznz4
jkpjLIs1tjbA8IuwAUnLC65dFI01B/uTv1OiGim1zje64BMPF5huHWezXlQDRpQCXANFVnUQmo32
2d9CDGY1lh3AaGZEOWSlSQD+Zrz01cHhEwqDuyRNFvxkhgZpnuaACzX2/M/x8CWFnJsvXpVw0pRs
nu/a9GsLgT+6rg5LZ/dBNK4W+9IdRzSN8WHPNJq4SD4+ehwWCZKDao9Iy5Cjt48Gv0ofzdPsS9dH
TxnXwkkjKsrfyvd4jAKCmVcVs3fbxV0oHIE156RBW+vIwLZwtN/Bb+sxDB9i9nEUMc8uspL+LW/x
AI7QkovTlX3va6nRQsTe3M0CNaV6FCITnFOU4xwFH9dRevnXR4aM9iSQiZ5gxSmjFg0rAUhgwYO1
Hs5G0X+HT9e54u09ebCnWfS+Jf48/SrrHNSTjSBXh+gzaix49R2prYmc1TMt/u22gihll+AoNHE4
iOTIHJnN29RGz0QWYXGDDeig+hbyW7DbiNFSh1Q5nVD/6LyQTUf2z4sbw8t+aVyx7m3fpIAJPNXZ
q1gOQjEfgTSEaLWQqGA8tZzumNag8cjI9XQWfhGhisIfsNxHd+a+LOVDDLDC9SUH+RBJmRwJ7K9x
tR2lYPTJBdoaH3d9jL6kzUVh+1MRzSAHXeUOMh0dBxxSsQRGKUBzgBnhZZ/8IWrMTNhVK4eiseO4
caHDyrGX6cgQRPe89C7Uw/9dOE8+OTUrfoi1XUBPDhVWoQlFP3BD8LkcuwSUUxGMbmNJCC/wc+Wq
MPrCLK1lqyq2gd1awD4wtK16SOydmQtWjyupgdxKADAEd7JqSLd5TkhF4H7j7r4qx9oO5GTNjMsb
sYso1anZTRYL+mWjImJENXoSYqltEuZRy9+xeDGR34z5Z8Q/NxpXr36UabDM2MDU0py6ZtMr104/
R9SXRu6yYQEB2g/Ii1U/4K0JmtHHlTEe0DFNJu6l+EI8A2u0a0EIGoI/fNcTdOt+QVgsojiKn1Cm
SmGzTzIhY6oQf4/CPn1OWMV80HLyBMSStpv5/ctr2lfUGyO55ILWoy4gSpGwYgLMsJ3gzyUq8zxh
R1OBSKNJf0xllFMJW84B92nVteGvsF1vV3xB9+hdsqtXS7cV+KtlNXiY15g3I1hw9lPRxwhXY71Y
WE+FDbXDghyn+T7U0TStGvUib0KfLn9CGedr9RKD8zESMlzblFfXznVOD1BkXSSptf+oeuKHD3zY
+J4AxV4l5YArWQMoF/jM0KAFZGIvCWQ4EIAINAj8P8Dq54Tpstcq4bp2xO0qiAb3lCMST+IU6ps8
DBSndo0O92Mm+oyORzaeAqr7z7e0NHFXh4RjOdOWbZ4ryaqLow2BxbW5XBBSxEKBOgOzAujBibgd
i2iRAJINtmIvBCpfeynGGl7kc/Vg/Q1/VaDoPawXt0HOzIA+vTAFt1AIr4oVFSa2E2dCZw15v00/
KddsXIJ+MaqZSkUhFa9RbmL08zaIzEsrw625Tx1TIQIbAGbFfDrss7VHgD37rVvDwbQmqfuJwQqy
7SAM+Te6/iFzm5L5YbGPSGXYfiRMH88Q5ZGN5y4HxMDiqdtwOAsSoxT6PEbwqJelHBPZq/ehC3Mr
XT/ESC2BMVqkBIkeQnNTeDNVKm5fR0f3FBaDtORrTXOy8vxS6BgT60Xx29/w5e9rgllDA6UqAcIp
uWqdd711yvv3gCz/F6DVYLYhD31Ywa+AOkUfq6uJW13ERRl0n4wriruSX5pvhRF9AL8v5o7XOMIW
eG36wZQ07mtKZtQAfDqEB7fwjOudnpR3eW+n1pmU6VTRoYmzn8kulh8Tqs3DcaJ03DDffNqHRZIV
PQjQipcMkKt0/aBYatj1Pee8jKGh1pNiNe+ArwwciJSPVTBliLa7IV7T0mWCHnL/5a47GRaOO95x
IW6C7w5d/2q33t2GgvRAU2a4a2cPSrK58LZK3WRsf3QNneZetgtXhsAkYmqO3WlBIB6ispyN3Du9
Xrg9EgFqmHldQ4OCVfIds4n2FKb1+woJ6W4ODa6W+NkTg+K9TlHVS2Efkzh20H1eZntcV0XNA3Jg
UE1TszGlbRYd1lrDokizUuvcKbFla41JdWS88FHub6s3Y4Bbh/wepeTj0TAnD/CHBMh6GPbv1kpO
ikQ5b8rbJHgW8IolMw0//cvW6kvfg20pHb7+FDkVVYVtJcKLf1lgrFv1M2oKtZV+kDz/mzYz21H3
kjMBOFjxLpuNuUj8EgAI1DMfjwWwXx4PGbRxYqARk1E5mcA2CZ2NQ8Kg6Ez7/VQxVkVoYEtgBk6f
5nPKHPLMd0c13It/mPorM93AHjE9MFXk/K2MZBmvTC/YO14of8jfqJ4/5RVlnFTgjmu/ZPHcSXwb
aMA+Bd0H2diBvrHalx9g8+lEwqf2hk5Tp6ACVCNhmlSm64sF+/DSdvUad62bmvMB1npjhZ1XImA9
ou+Elss9x56ukcIGrSEhSKBfdVuBVNcuCWR7LGfe2hswmSpIOuVjbMb0VTTDyQQBzaWDEuVIWYE9
d8KVBHa4HvmOpZhNFHPieMsDETmpwTdZ0yxh6unviLYuSwD//PmKGAOAW4yBT9EER8uQwGbD61BF
pHjUDTD7SjI+xUCBHNKbFruFzrMW5cPDzcIsqb1jE+Zm6IoknVmWzBaFoRdai0GHM70kudiVrmcZ
EpIVHsiFzeuGGJ8VTRQR0fx46zGWbVEaZKuvIzLone80udyJDNYERbVH8XcJRBGRbCj2/8A2+QKQ
j2tk8kUyhqI8RF4qHRJUZdK/M6pnHzqfBtbTzUBPXXSan2gM0to14toTW7bvDDXSm1HKvZEdV+12
RV+yvy3pGb1sI4GcWz/OBhLqvI6gmVzh0QgPqxtPWT6adY0suAnG7nrr5ddYocOw4Dg7Sz7lHgOx
SCEzVsJqywt6zbcfjtWGd2NVYdQz9idMsy7xcvnrAbFCoAeSHG/se9HiT1ptaNEsDWckW/buxvUn
PeGvlsD8ShIP07YhJ4KeWiJi1MIwchsEU0LbrNiHls5ybZETyoA9d0ns6ZJhIABZKzay3AE6udNH
VFrQ0hf0kQVtpuTUZLwIysrELiAeIZvHFeZY4t1COSJ9S2cMQ+PHa9G6IXnq6S4g/19XypJYgjTx
xhmpFRJVPu18ciRWIme3wuFa1q9asCG5pb7z1h8lzJHVrscBEq5vpllZPXeWiTCYExR2/OpdhkXD
Sk4OFzUveDiSMTWO88mYwiK6pcJGINNd7AfkBK/nmzXdAVone/Y9us9EdaaDPflsblzvVv5UwmFT
Qqp0Fni+oX/0HbkDOONsf4/viq7428fUZTr1Ucp1ea7Gh80EP7WQecir9gwPDKU7dxiDDm1pgSLR
Fn/GNnVdh0UkOhIB0eVtz4p6sQJJj4Ge77jlc7SRZHzuYQxgMlQG96MlcWzs9dY/ORvgWFU5Dxxa
XjoOC7pXiMFCdvbJxheaqG1xbl5mST2sUXNoV/DaqMHHcwr5q11RhLLPEG4TvHRK1I023TOa8JuY
N8BsMPq8jslGD8sLf8j+e7zPdThql4lPwz6JVKPWAIRER9OW6YlSSwGke9ZeciPlZbzU0EtNk4h8
7dGyN2uFJlPWE4qaaOle7oWqLHDYj/A1ariz/LdYN2C56T7KLUEOTyeDEw5WbrN+gkrSkSAR8kC8
1x7xySgu+q3A2SkDZ48wQzB4BWzlTB6KwZlzWqFl7/htXj061D4he3a/fKFuVOCoWzUQmWvicG6D
Lv1OGALxETZxly99E0/XfGjcFuY0mmChgIGWARPrBCvwzEFUAxsj7S5YSUYWuKlH9be1GJYHFwEl
XzxRXkwHl31fT2LhWG2U8I2EkrWMlHnZPqH2tb4qkk58yHk/Tf0ahTNHGzbQT62TNGJi5JtX3Y+p
gpduxSlKlwUQjbDJBV6UtAnUKJ9EnUnJUx31UMREL555qNq27LxZKd1XMDof6FzelzNR0RrrZVfb
uGz5kG8K5sx9/aE6jj+IMyFdaqD6XmTli+Mz02et7UOPJRV689iKnU/EMeWyicFvl/2ZvZiRCbN7
+L+lks/m5nCXjZQtGzaHyUKE6iBn9MLZK3tzhQDRR1eM9tWlQaGBc3U2ESIoOHlOdtDq2pAMbITV
OojLvHqk14xskV0NEEo4RfI3VGBbeE2JvCl9QEXTMzIKjbXYDCyEcaf90Zr53TY4OXiQN1FWoBOl
DvbcjnPeAARQzjWHiRhGfahiU3O05QAlyIxOAcO8W5oBCNMRG8p/vbe6a4+YNQO9IESXDgvlDhJo
IwD+ykH7JfQ7TKYx1Np3XyYbMcrWf3Oxrk+cykNYkU8mXIP0vU5knqiD2p90jmpNEfqCu+fAU7b7
7EL/OJ/qA9XymDD6OQR7LRXUX3xVScxg/dST7VwY+YP1PrGGzyr66/CzPi1a9wIDeDltJr6EiSnA
ofL+jc3OogzPmpmYBX2u7F7mJKOG6l08G+//g00jQKs4YgYP3LY0x02E3GSJ3ClKctG2UYJJRson
o2dARCEUBovt+ydTFIqDD695krvs26+GWxwofBOmfhMoQ4CRKnduwJd2Xuo8c3z52uWUIFHymf0+
uYh10khpPFwH96La7M9//f3Ww6Vk0i0Pg9ns+OZY0lx49Ucqq9Wozgg4BpE2n8CehddmBKW276Wp
F+7Jzh8fWihYhV/eh8m5hcp3SWIBKMTm8le7P8LDpb6M0jtZ6IvPpI9gXE8U/RHVJ9PCox4BtoOB
pTJJ4N0qnwJOW2OkAgvEVQt5VfGUvfi7cu1FMuWrhPTj03gvq0CfVIqcovDKFz6+4L3CGQ7V+pqZ
LfChqEWyil+o4ti6yt+Gc0Wtmor2GIwfEXPRkPt9LqMVFREZHeqRtXn9tWoDRJRK16+dD48O8CHd
yjWh8NwJAkHtg88pUiHHjeWxQHV92XMNU9201ll0KWUhTvlJzmfRq9EoKEPPIu6hqCI3AUF64V0q
gDPU5IseceTW58VXElIdjmVCQNUYKc5vFQKMO1n9atyPZ6bGHPA94hi49PHiYUvOR6uLmc47ejVF
CwzKu/bzsJAWD7ceOwOHvf2LF2Ef95MBfY715cDL9UUyQdTyGcmYrsrcKfqj6v/JicFPLhlhOaQR
ifSE4Av3UXr4EtE/yNifblkhYXXicIKv037UfUyOQdiaPuPKsZ9jeomnXt+3p+dsBamN+hVlnHeM
Jyn+38YQrx7w47WImyZQzUJqwnQ5Op79ghcqKpWUQnxxL++ixMLdP0PbuLqtClTbLejVzSielUuC
SdlupbL0L6xP7mr5L1fOh3GxeD+5G3tkEpg+mRCC0oYkGByI1yrECCy3Uj54kJtlZ2sup8J7l9Bf
VnQxqJ5O4NXr6Y8HmOw+8Ldya6osh7fMmXSjvJ2b6KdayqgDS6Ory+SUsMCW3hgtclNsoFCrRYT2
WRn9wsP6xnTrlyhcmKBebpUG2yiLzlI51EoNXZ5xq+wq6Vppj4gb4tFWnp+ac4aysb8011FgYiXZ
WzcDda45n/7Tlo8CpOud77yS7X0Kw0w4kzK9/AnW4oxao8MH00CR9zCoJGfMkPnaJt51AxzTcbzM
AdPWUi5NPr8vR/7Olo2n6zLoX1zYemwuDcueSZqwTGhr/nWBZfoKwZfilpEOMkWK33nXTaKcy19u
BODQdHxznEpD4VXcx2IqDJry5eyYan0HwswTD5BTJYhUOQaNsmLXJ23xkhm6Wke7TjUw1jlNYd/P
k9KRzptsPYmInJGd6q9nWMeSaCqpiJAuE05ko6/gk2uE7kNKDJ/nawYaMPtFDB+i4qBmsPrz8Yht
F2gB5ZoMTB1ear6LYILnI6mI88AUjJc/IW3KlPYjLLBY1wcI4quGM2XOrkk/afmlAzQY/d+Jrevq
97VkeNGH4ZjSj4tm8TpzP1DHsFv0Gz9Hz/DyPkunBXPKiPqGnGDAd/uYKS/VdahkkQ8ADc3+NxbN
1Rr4IcBzgzOuuxxKuuGWL5hcog+cB60SqPLHiDF2B0mRyNn42gb71OALycs0m32PNodFLjcNLr5M
eeCsp9cxsSQF9NXPx1zBtix7u0x5aU3i22+LbOsHo57u0rsoeRxwpzj34SbvNrkaXxTPPMGnIe+Z
UyWKor0AFOH6vBp1REq9F4xK4Y8PTiyYNokeaOQJEvg1bGonqyMU02VyqfJbFLOy2BKyelo8gEGt
EHbzcLdGfouJslcKsTL3Z+hLUlQV8YLZn01eAqdDoY3x+0ZV45YBf14sikbGvaX9XJPzyhhC1Uc2
kjJBbkVjfD+L2A7GFEh+VRu4t1vpgV4GiJcI31vwv44aKWtOrwqoqOifMILtImD+uTqvaD8LPnQ0
yP/FfPI+gpjlnnvD2LC0LmAFvjwJ82ZYOacnX4nzxGaf0EAnTd+BeooHe7BRF8AsLRrDX9JVwcwI
3nteQK7aqgfUDAdtgcCgcvEBQ6y0mJjnc6Ijlvo5fmnyDFKXEvShqCZ1T/vC4qg6HrWLtfX/IwHd
0tyfbjyJtWM/qrCk4H9rMXtwavHcIJ2E71UA+MqARKeaPbzvfntoTC9TaOOVVxcHBwWmRkknfW/X
z2bGrmU9ylExR2ucYutCLDvA+JzcsDhOo/kcaxWNkG4eSJto6WUl4fDah6vNqI812hlZ9W9r60zG
UwuToyD8AQwX4SCBt2Lqr7jgw0gT3Zswrwd5qpvNwhs2M9d3g81aXcUqrutI9nRIhKLPPZ8T6jRA
5lvNa6aYv1gRpzEssHQPWsA849raE3ezBkhH29ijTcTAsUaSLhrruo7niUiF2ugDD8c7tzk7+jlz
qogHYMI+LvE/aXeHRAPD7kC2/hT6idj/G/GwBqSoS/Rucv7lsq1UfLQJLyHKdEPs27meUu4emo6Y
GRorWvCOkGItv7j/Jo38Z/l+nPxg0AjdChvCcK1NK7ioo3wm4eZJNlh+OhFeqHnGPHhfSyIhwwER
IViJOtDvSvi70HaQ9k6rFVTMk5k2RgE1XtiVetrWYuOjAQjAiLOc6WBgqkRLy3eRCQvMnJ0hBEmp
GThP2xeWb7bc9NE8Wp5goxAsIjWdTE0sY6wShqUDBVszdlOOxSYo4B46ADYcCuHS/RcY2jyRVXi0
xLj9vq55aTU9JBCUqJzBtgX4gihy7TI9OjM19p5I6kELUvkJwQ9awgtfLyyuHH2OeBEZ/p7g/079
PVyvKr7fodXjSy2q4POq89qAawIK5nxHg0Y4eaSaNJ4sX6R08xIXfq5f7aiiRBeNLN1umdV2xXDZ
ViqIMwJJGlUyJjRMG6b/+WcI43FPcQ5S70aiwvMCWIls8OqGrqG62y4rMOvWGHHTYDhLlfPeKfiS
K1+cWF+dl68c/7EzKAz8/eqSrm/t0U3xO/TY5+kFea62TmJUFP6IaXL47EbWvXNEmkr1bFGSrXzG
5RL2ciJ0UhJcEA4qcJ1Aa2Mf+33XpiL+9gz2hsL0c4oRYJ/VkpCOcnl6TGnQfcMXXFNWDFK/pFkp
vAYuU5Cn50WjFwIHexKB9hc3qcnKD3AHQc3LY5MWeGWW0UL8YBdYVMKywTj03w5Ds8oi0qfD8DgB
MAZQmznMDohXSoAz4T49GBaN8aGnu2YAqcl8SVBDkBJX0QZkDLNXMj3+FNUnXx+eC9DJIeB4eomC
lD/4uckhWCzSIx98iWg4U65/wy6WdQmZcx436cEkE5JmoXnwwDiUBYyKmvImF8jSzdXrE6inHzZC
nZu8RSRcVqoQuXBTsvC7DGdfPHVYNPWJGXusLoPTcdr8cg1kQoJdvIFZTGjnFSk+3TkmQoCfqSTD
TsgIyXjvSwQwZmJWCh7Sy2aCSw3LaT/m0udeKNGQpzXvq55azimW95P+aFX5NiAFTBrPs/iByZ4Y
dW1GWw1gDkR3wEhEcziCqm1LbUwoNQCsR6VN/qQWl70ktJkZQ/SY3i4NCm3YX6sAoCwXl34YrrIH
ZlVv0wXPnah7WtAMRxzFsj9R/JcqZc9l0/Y0EINrOKV91lmkOk+LNFrhVR5V6evWqrgSkL/UJm+o
CAXRO4uXDKtHtynuVA+oQLq2e0wsx6Ly7b79rRtpf2aunqaUALLRNfUOuWArdkXGGKuEDwJERWDx
keDokuN4xLcpjYtsSnA5PrvZGv8Gemc6rPLW2t3htQLArQqy7JbyNWNugUT2wWOkYX6SXqGv8SYe
b7d6R78FK7uBPQkXXHbRrN7xfgy3b1zuk68s9Dklx2ZG8fng0PLlYorheWOp2XAMkU29+iho5w8A
3rVdFFRLuao0XD0fEwt8RBHrnvbFCJ5JL0CR/fdWZ16Qtm24qMwWKoUYGKgNhMHrLDQG8MEEmnZ6
cC1LE9KOLrtbpMT7YjiyZz9de1zo1rWE/CefC0FxCb6I3oAdJMFYF2Dbpi+4K1wY3LHSXpFC7iAe
KmrG/C3zWQ+6UKqMxfDL24+JBeiHg4LaSxaLeZ0fcZf1+tzn+wuOPf/69zdrNhHRvnDUWaNpzU7O
NtGZdTuQKIvy52ARM2dcO9NlnOnjGz6Lr05MxsxwAW9u/Yu3BC+uamd5KcYEtpbHV1xoEbuDYBfm
qfmLW7cAqmTcVzzwuA8FXKfRvrbND3PW7Vs9/cm8XkAIZjQutsTMJ0M4+0Lk6oA2/DZ7sMrhljWy
jv4bj9qX6bejOsCdBpHxJoCABke7Dps8TSz3uSjGPjeOI84RcElddmjYK+igjZJipBPaKhaj3Cdy
iAazfwpJ9CJFhJcpdAJoWmoQusJfAYKU7jd6+LSdWe5BP/JG3yYgHYE4+A9uo+3o8MMmAc22JLV3
lXz7sZzezKeOd96m5gi6qQ2C1F0uMMaes6ztpf+HF/51SIl8T11xBjmKUvnnbDtTGrtT/EUkmjED
fS+NO8P4nijLRJlC+qggHHuwIv+cIzFKuCUQd/Boi3tYG3vON57MG4QWAWwQrdaujVW2RS1sphI1
vvUpu+/3g5YzjxId3yeQOlV36dlCvEtmI92W4mTaWbgXJIJ8z9keSp/sVkdfQwtQkMqUEQ/thfYE
WRVvg2f3NX2KCCyqJMqwNVQz/4hyRVjR9pIdw4XiARgMbRbgySIaVy9stUNepT99z2YLg/VhiJt+
/OTbn05RGeFPbgiebboTlLooNZljfL1l2S4+tNUnDDda2kgq5C8Xg2wHhqumBnA8Mlxqt8hNqABd
LE8wo54l8bVv6JYSAJVAa6Ho4D/9m+7B/SMbcERleLW4UaOeOtV2j4+TVOVyFMdSFhGe3uibuV88
00qFbToJX9bexISP6zb5zCfvI42RsZjcGF4qM242P5PyjYl+81OVECN/NgGvXfBKUekdxhooSSvT
u9zI4TDEAjky5bPpu8pNOPSYweC2FySgu1ezaYwjcYtXoi7SwBkKBoX91JGqybCm7qQhnP8tUPAB
m3B/flg2sb4eRjIXmDyMRleEGKIYkIlOkxG+hCfXCMcmsCIsFSc0QVwZro1c0S3VjJzgr76dAAmB
Qh9lH3GSNXmQQDI758gk1H+CcCMJUUIsLgFafvtSlKUyJZ3HMH8mpeM8/X7SpnA2kfx299X0PJB8
SjpsEoWn8BwMKELbGXAV95m3HDsPeBfrMZ8/tr0Or/FEm+vci5JKKpGMqdG1TF5Xc+9oTFDONR7W
2GNoWB0W1b7Lvx68F3fdEjc4WJUDxXK+zMhsOczzNoO98oERaihOfEk2ezFerB+fezVljCFM7VDQ
lDH9zmrA23BSTDWY/K0nMMRCUAeT+TsEMj5Pry+NzrpNXk4rcuLpRZQXxoSy2PrV4Fos6x9ld2n5
VbLBb9fTFhXUit1zhq+e4TBCZtWVDgf3akyWJi8ggRw2C36H48XoS7SAstPzqUPCFYR3VJM/fy/K
bKMh0cyWG0iMS9/uBKw0Ca91BgXNTJmlNN7OmNRz+Iqzp4Wd2aYUt12hwJ6+JTiiyOWmsINEt5Km
fhk/wm1ZxEJCutpdZEFLkrM0MX0bzHrXO0vaHPsMrdecBvylwNSG+lc9oUzRQW9H24/z4Zhau++7
zTx4Ka+5zIMxylztZFE5PFpXYpRikCzTzjXhvMxcZIEu3iZ6E7xRJodYKnARd9UVtiQv0VoMLtZc
NDCpbVF7qbvfwRJgKCbDXQAOMZxe6VICHsBZe75oeQ9uPp5BdsPKISrvOtn5RyqUHJpEIQXL1rBZ
QuCGvgROb/CCR3BWzBZ6RFlNz1mcO3+2k8EAlJydT/jknNGm3IOCqYUYp2BbW4H3VE7w8LETSJEw
AGKeCzHB2Ioy7Rn6DbvxCvbQ642mldDyWyMlrWD+WyWM8m7aEVh4HUBjufzkP824hl3ISygP0wFG
3g6YgEC+wkfyzYP/7nxGDTGRMQxaI3RcxqgoB9j5oGwe9TElVgNhTa4SJCLQ4g2Vgxr2PEplNrQb
C2z0WzVQl5xzp029RMZEclU2od9QkGhC9CK+oyaB1mfbS2zAhb76R41Px3/+B/I4zDzcigSO99/b
DOUizxFkSRIZOarCbVpHDMCzxzWLMjw46VJc7jLYeYHf2AhNNO2cvrDPWn2VrjF/ioABnJu/BXes
ywIPKmaBi2AgXZH/BetN5zGeUHe2AIv2+m+ZvECYLxAeEXjMcrZrMHLsplKivQ+tOwLQb/TviAaV
Nbr8W7T1NeONhwc5lt3tkt8KUvXZGkdeJUn4NZdwwbivQPoQCfm1XG9Xd4vB+Vyw0FIOfH4bAPXJ
Xjscb/x1KXCkoR5074ToCUxWrIRDY3q63HkiiTfE5UNW/GBis8Azy0K9sGn1lQLrpilAJuqiY+Rh
2cUB8+NakgKK/rczGll8610J1lr5g/fCu+AdCNK91YZVf+usB72l7Rt0drKWm7bIYdSVuCqpHXjG
B85kpcAdbuwfHYqmVsRpfrJylhbHNm1v2uiCUW+16QZqPXsWtUKajgandA0KPfGbm5bGxERcurms
b2RI51fuoUG00+EqngEEJmKjVdCcEkdwqjTQLs1iXGhdy28tvhm5HqSV12KVNCQ5KRftYP57ODec
dCnfw6DKUUF6eDH5z7QkKU1eryERsu7Tq2Fr9e7e0d2OfcPXJmgRTVuLPjc10GvPRkCyid85n8V9
4epRW0iMQ1ITKvKUxtWvh63V/vcv1ElxslzHp/aMaAMwOc1R21XESORrABoSBkqPfega+NRlmzWK
P6xSkFhKcbwvLCLkaxbQ0eOIcqCPebO6qKRzqvfY5uMtSLiQ2j1MAyS0uYBVU0Gz2mctI34k3oO8
DWMAgT8k3oXYO5L8ON/Bbr+7CguobS7/FOeXeY9pg3IN3CMs8YJZyZqGnddNfgkeMUFO6fxlIakF
oWtRYEdSazROrFtlLjCyT8U76UjxtX5oCc+ff1GTeKvFtW5wNYp9eVtUHNAk68M/4/9yLtejrYcp
izDnAFjvvh2aR2tGpjiFhPMjNyaVT8GUi2O9k5T01qGLQj3jfcbRzIOwaWMd+gxoA9p3lJiVROBO
WeLUe3vPMIj0sHKJlCtqx6w7467YcQnHjHUQewkxqMdO8imjBaEX4ECOK+QM/leFYgPgX7Ws1b18
gTZmW4cQ9v+G+gTcPMeseoHF9XtYtykRB3QvU6GwQ2O476JxRm9znuqMV8+02G3a/e83ToLwAlcF
s+zNz2K9aOhwwcU2J2zdDuCYTDfB68kysAP3uJJwfkkMaLQ2yhplWzO251GeL8Kzyn9X9dCmhdOb
hLFr3qzKwW41oz8uhzE6Y3AnpJsPELhKw81MrD601jysYGJC9jNEGHoXek0N2wB42SXFair7VZ7g
ROxoVMT1XzVWCQK4pBB/Rcc/NdjXWWhaAIOQVV19jsC/2B2IBInuH9g+nJnijMSieTV+3+pVmr63
StojXQevifl4tFw/6mBnnPz43XPvErPCCb6yzwJAzcY/wHHi+M8igOgzCLIQA4YcWhvDIhdUHv4y
VgLJtD/Ogjw8A65IoQzR16eOg+57pAejEfuwoPxmFqkk9f/LdcMeCYB5waOfkPX7mROsDb+wK24F
df9QRNxzYLrT3OsQLi5uFc6SWOHeRt+bm3jiOQoJUkWxgPTnu1FLcVDaWSEk08iK8KC/EkRMoY55
fGFjKmotVomlsHXv8g+SoW5WOZbqACT2Mkv9ePHgcCenrXQFwjVAWgfANpPgNKJEbIWptOoxx4Yu
3A3rOs4+nQGOsPdpKXLV/XATXHz+8aT4GUs1vzskqr9dX7ptkm7286o0CRvPLuNliocA+AKxjlQV
YI3T/drh0ru6AZHojs6Iw/e5ukLXZl258ZzTVsg4+LHNgtlMp8U423cLOLWMxdt8kPI3VzDgxHvp
ML1HOixYPCmFYg1Eklg+1BVgd4stIJjvL0XIsShFNguoM/2ETpi0R4FOV88HQxmGMVUeBVrFuJ+t
yXU6A9IP3+1FarUhserWU3Jw2oxoJn7FaFUuD3PtqLN2NhUoqqHF+K90K+eok1WCHdtm6EqCogXu
wca/oZZvJfAkQuu1J4QhWCgXk4PotiUkeDaMdEo4+TuQ+6cZ2JreJX88uU6Ahcep6ZH+DUGwlI8Y
LNDOF74hnYhuAa7+rIp+zBcz2DKw7V9+eySPb4g7t/WudqZeIexvlNwAYPJen5xS85AX/NfIdkqh
8+GAhPoHTXSjtquZqMN3QWPVWsGKyUiv5cpLCPTSEPueKg5or+4OFKIkaMveDytVQSvOj1yh/psa
qdH0K9z9F5wGSF7EFu3kXpFwU9ICaMfSwDc5Y9mUOZez/RlixMo0wtlb8d1yH93X6grlLTHitF9V
haWokPz6iI7NKO2bnbv7MtRsREzwJgv4nfu3fvyHQcuEynqk7AFhifT7iHEXBpeTfwGLt6JPP6Wt
l78PS3oILT6k6vZLzK/x1ojphPw7Q3OkUijLp7U1NRKSkOtYebqtdjeV1HIYgOEdBHP+YrdpCPJX
yU/HuKHoHBe2enyYzsMwD5Vb3M82m/xNspCoArby4MTyTqD32xtfhSdW2mq8BdIGHzV8WXdemQae
IfJInM+/xXfaqNNQ6FWxBFVdj9/ZNejyjegF2kisaQKTjcHjgDjZcBJ0Apn7mA/G68OLVr/xNN0X
Kd3k3JgOGVqDdxTGiV3P6yeYH2CfQpftfhumXGcpuQMp+h6e4gmBjduToqsR5F7Iv70/iF3UQIut
dFpwehiEnIB91pVwiBflcgdtCz4EEIHH8bGyxBGOPLzAHwPzbZubJ6w+cyDz6Kimkg8epW3IE8n1
FvM0aNg2XHlPwPgn74T3zHqlcSna9WHB4OSjfjAFC32If4dP5IJE1htjYHh+FUcBs6l5+8xrjqjy
qw9Vv9Eb1MlaWXK8r55huU5zYaVWPiH33RUfOK4cf6X96cdZDcAPg8e2DZoJPwt6iRL/RP0iCEyw
jPMBDudH0bgPy0J1Lg+Px7jNDJxZsdAOT1qCJpVTu4RcpPj/TQXfuaoTG1tsEARgAElJ5CAIfNuQ
viD3m/IxKk8eVNmrl6flyI3flPac3VYQrof87rtwJiIi+zh7fG9mS7JwbSOp6gu/UriTUelAguVq
/88JaYnq1VsBw8E3N2Teb/flKfnBngdAJZim+kkLusqBpF4IHI36JOVLxAkq3bPCJ3ZKNtGG2CFg
XEa7hzs8oPIw3f3+FyPYAk51IyUaM+WV8u+JDNKVi7GAnN1oE9M/9iAvahUM1d9sRNSWB6lytJ1k
WGJNF4uOR7ElsKqSvaxx3TTKg9I8cffXFrJDXSqxCiEjW+FJdKxzUVhp25/gn1E1zRdCytX2Oesh
S3u+AwOCsdA9V/A4cDJ1gMESgVOn6Hz3ou/gCf4Slo2cEsJBoc6r7zpXuItJqoNcpax0XJJIj8gC
pGz+3ru3xhB+4Zlq9XNRXpAPm+ktMl+/usA4StWpbVDD+ql2sv8MfOS0QVGnLqUCAVvG+X7jclCZ
wQPaHlN7mkTcuSx/6mZHFQXg9JUzAVjBZqfJknyi/f9Gq9mUUxjP6sM37X8UYn2fDWWlGU5YMDaD
+Jk4A79x70m5oib9YlnxWxEmIiW/Wp7iA8gvieEHOHrLHfiQ1Unq8WfTaVwZXHJ7pZ6H0VaOkl5d
ZiToWIp2ouKWRop3PwoZv1Cz2g/1QQsGdqvPsa0f0q36/rjfeumXVaHJdWgHTYEJpYfeSw0GC43p
Zjj2kO4e0uM0PnnTMModrVMs+5JVAaYQNrc1ng5OMy2STK+7S/iBlOqzgDKH/3r6dib4K/TczneU
hH6sX+pNPGi6tIDd92jN56DsDf6T28lMoOFcKpFWS3QErb61OiogtLW7d7djBuoS7viuBC+iAYM4
MgdVKOh99pX8A/s0a9qHBqXxU4pIC3VFLgy8uTUHwTC8IEi9OxueZaefru5JDLIidPbw9TRXEIix
TiRKE8EmWPvbuzXMaK1EvD9rEtEI8IEhWIG2c+oPCskBVWbV+D3LaQeOV8oDZ2faaAX9F1zutHcJ
NC0uxjlJC6hPkbxILdgAV3+5qPH1QsM5mEKk1ltig5T5rvMUY4ASi13QtrtoAWtHDhaNA6Mux7eo
3Cmc1mLom882ttwhRTizZ+lGE5QKok5cIBuCpTkmnaz4upiGA5LIsKn1Hm+XwpImgpDoIvWpWKav
nOmqClIqwez86msVSrZrY25wLKZ1CvDKSNgxsWWa22UXzHbGL63qTqADWBe8Q3hoeEjuvUfgZVHd
1CZfxJbE+o372NY4wzXO+tEqEsh4+dyIsNBLlcngahSAF3xNw3P1+0yGCRlv3x6W/mJAswTs9jxG
+rsQ020CLa76nnMKWl2MZDz4ZQu/svURTEP+qDL3ow6Mamy38TUSG23vh5TTuMUCPFkC00/dOadH
3BDIYh8VHQf5Jx3lqd1KbCUiCt2sj8qeRleJOXNgzcbso+OyJ+DEgGKmhuUF2mFzEumQbsrjUhcb
N5chwJOYdGX6r+MFvppiOd/Q0A99pdfSIjmj5FOAa5pV9RL2zj/r4XSDhl884nCGh+D1+ChbDM8o
jc9qgqA1T2U2AamqtjI2FpAGCAi1ri+Rp9hSpja0MqoEVvb1hr65HXosP82vIF9oGRTT2NUDfzGN
ZV80IbS1pbXto0EyP0giAd3SHXMSW3tp24NUJuneGEruPjBwZ0ZHoZ3cOztgm48pzXd9BaYJDskR
JoIm3rOHnnMfV8z9jrU0iwMiEjvFZRQYPbZctAIsiVGeHx3+8T8uc1vMQWBShr0FrA4cLjbzzXPI
fS3nRCZrc+fU/UkEMyklmgEun119TyKwbRwNP26ap1G9GSNXHfOdkwHPKGQdjU9wVMBjRqvlHG5P
STkcWqGOzvdgIW5dItTIq6oxpRre3FMEZo63GFg8BzqXhsWtshrydmjldXJfF6Ji9AraHdcTHRgs
bn0fGOi/ni3IQ4Zl096GJtAQAoZMaicKs4MWhLQ/AOKIBTi8I6vzZVQDnvjJA4LoV1FjbK4aflX3
DbVapl608jFGS+ahRM+VMkT0TexjTW9Jb6XBUNCdoxMlB9E5fVx9gESp5UTSxLLOVoPpMXocVKs3
zPCzId9ejknzGIUsRjcI8qraOrKFZPzMw5YaqyBx99MtDlYBaoek8p4VHbGSVcvmi95UwPE8+lCm
5aCTdXO6LpXzHX7UmfNyBjM8/vZXJROq4K2bMWeC+gzODirolad2xQ9sMkHkt2YZQ2Cal1v/Y563
Ii9jXxukNznteAUrFmtdT6zQ9cY5h782TIvWCmizD9RiersUXGGOo1EsyuqWhaVyv3t08sAEetaP
UWWz3hiUT1DNPNwJ3W+2Ndv9P5BTKw1gjqWDirR6/HXda+hy6Xj8qNMxsY/lw4e9ouWxasMU941f
bFzC4hkcUOcVewPimS6T2KD05jxZgO9DAujMVliEE5Yf34lVgukFKxwQW5wd5z1M0mt8djjNSeIn
QXRY0d9bOdmR28TU4kNdqVdm0QoGjt2MzO+C7/JV24HDZaAX5NSor7We5Fi0LRCksccVZyk287xk
vKasQXFdpPCATUibbxvSb4mT4qxaD4E0ISB6eMgpxVCbtrh/ml4P5fBF5j5nDid4CUjPWio8/+pY
yqr70TekLKEXHgYW9lcKEFa2Lf/IlcBrzurN322PlrroCDcY881dUfeZ/JttjXatYwDYzi/PijCf
Af+Ck01aIrFbsmCWxsrp25+gHIVcNPuQrX6Et1RouNsZbkakKZ+NLCbo40ZaQ85HasOzxO6L+33S
xG9M9Oa+Zlrr7M19/2UcgR+LuxmN5fWAHs/NqtSJhlZ1wIOO7ACuwemK7iMqpxlmAjEskYnfgFDV
Xun712ftOOkRgWJLMcPgBSd1MgGLYTd2L3h5G0QyEOM8ZS0QZnUDunbNX2n/SFiYVvRvguAFoSci
jVVUTnPBJ0lRprS7twEmKSEmQ+FfchEVQ+wpjp5pzZU49tL8mIYkembksyUehyYrVL3T4IKl7O03
3Y5ZelAJhmkNmAA+Y5B2+C78+earUQJEi67A+gfA+9MGCNISfPE+4Afgbz+VOf7wy8KaDECy4MQl
k2UxI/eYXdtRib2OFuRx6bi2KjBJex9yNusSJikjkF6Cl2mcwmiSlqFk58BVRy4e1UVO/IPRNiRM
RXOXzP1b7Tgpa/zB9/E1Vj29zKiUhWLANLcfPvWlVBZpfAJRBX6Sr1Ql4F6Ux9e7i95dS+SiuGUQ
pmQUNyLKgJNkMruXlVKgoYnkHDQQJea9/A4HSfOGFWlzDY52iU/uIDxWKkn6raJLLw/q2aq8cBKH
G5//oFK7tKLWqRv1yqUNaW65has6fj6wIKsAQkM3qv6qw3l8dsCQPOPaiptKLVt32uCKBSaT3V5t
55hDaE2EOMDWQtxD2cKGKGNP0Hi42Pv9cVGau1NoZy4kCL5KgrYse/s9xI0Uy3AVgccyl29roX88
OVTBy5ds1DV3AQCmkhgCpuE46Slr4lLVUKy3AXf1kC+rYZJwYAb7fdt+pF+o+D9MeOovHj5srtvw
gmq/KAM2153LMjTcyO+8z+kZ+0Dh0qgoPz867QVCXoqp27XLzezjjLUvZZer6cHF5wHqp/PUyHVV
KOpjTo3KE23k69xEbPm9XFTrTl8I0HYf6a9FpM6XJQRr3sHoX3pRBtt41k9je8KdCQI3G/kvUD+A
UzFhaibghZDbkBweitbOE7WqHrdQbdT1nXkk5+TOLMZ0qsccMecIpsg6cEaEbFmAhzXBYmHADRC/
EFcBEOzeAr+fqiBfxpit85UnXH6IdNMMl6cgoCoV+QwOUR20YLhipjTtVdwVdZcxdGNyQmAVVsOI
CT+GN273xlnw6jGXvVZDuZeT8V4DI7295ITtQzJKthtGgpX0TjCQwFJj2nQw5giFTC6L3z1b3le3
xKSxagAOKGBhelPdOOjatXV6XwP2o7luum2qIBJsPdvu2F3KUyRYfHRlqC6Iw5JtVdJubXIlEKRx
o5WC8C1cfeyZ6o3m9kqPOYk47HYI1q81X8uwai4taz01ijEDP1Zn9OpCZViTfpT/PVhdGroiWUlQ
eOpbVyK4ViOC391VuTXiGB4upVJ3LiTu/eM5WqztEwimI0hB8kEIxSsWakJSx7qBdfcvVA8Jne7x
duhRBWLWRGrakuqXig6h/eFY2gZK3sqCGi7a0mcws4MhBbpoUj3/xZV/7NEaxAbx4UMOIZtxoLLH
irj0nxKsWhpPHovv9oekXLRo6YrctddkewNMc0ecFBxqsUtMb254h5fg+Rd9RroUrjlw9jEEkncm
kSPXLPof2FhOaEe7WSADkMtrojld2dHnTT1/lI2VtxWBYJzt7c/LylIL9rQJl856CFw2lxyzhipW
DlJw8TQ6I5cbUFaVIGHnGexv3H4wZBP+XkwTE9NQUSp9AqHLzeWeZ9WX+X/ZbGx6AH9561Dwyz/f
P5uIzgaVZZKGX/3IWCbs9qyk0rvQhHWp6zmUgwyEmRWwfqQIocR29yESFNMIoxsslSltVXjLNtWW
AGNKuDNpuebTMocd9r+uB8zQ3YONAnD05vbAuSykE2HP126l9YZkDT3gBrhcRr86bLQ8W9qLmWWj
domWRZBKQ18oxXSZfz3T9LtgmL4Ljf+1Vv1TXfz4mdlrCJ913oV8OUMuDTWQ2tGxfChdBnwlxTh+
LFrHQ/qb7Eave0KxkZ48ZIQyokkfyV3gDGzvxejr3CldZ2MJ9x0ziRcyqnu1Kxg5xDJurarpBZ7C
6MDg/odAyOiTdUqsF5yXc20OiZAqpuaqWsoZSEQnefC6TNDt76eYxnXVDZRsqM0GyRc8BsIouy21
M1U3mfHXtRGO+Qeo3nue1GF3TMYZ2F2wy+VFDT1D9PMIbla2knkVu5l+8NjtpmG74WtWAv9CKYqb
2Bk6ecmENJ5jVEUyEjQYHzdhrEd1Axhi6Ct5Z9NqqZQ/bX02mrTDlJmwrTpggfPkvbG+zyxeNwgS
v+1zYfSMddkz2zDRpHuGqba0d+lgiSZLefDLP7EcT2d9cSV3I4/cJYTaJwykHYPvu4rwPyDi7p45
iFSLc7ezVYyUBVuqBB3VLuTySOL0rcFTm05LlY9Hvp7UXFHhj4ds3UAwBjRVGkT/sbjFYFeOJz2U
Zl0XuP2GSNksntHL73DNV61dV1eHsqOhXMlVnCxxsBBH1VqkqLAtTK4gZHJV3FPxCIUaW9Y35MRq
7vjx9LNJNQs+Av6S4Z4QLPeVE1d4j2bItTThmQ/g7k529pV7/kXb9TCBYmJcPHMOc1EgDusjIewF
gVvFHTsROprBAl67e7FLEXgnt4gQI+KuwHEtgJ8Rg2H8mjnzmRXcVc07qV697hc/G37Rt/Si9m4C
r/OIm1qLpjibNfc97f3pC7cyc3galy5BBo4w/qIhbFqJ/1iIk/e7CFn1XVRyzl8RmvvM1iAg9lw/
YMJqoqq7uCtEhgBpGQ3qElFzkRR2JU7dxc/DVrXvsg8weRicjwg7myoYhOcUjE4TWbqzYoaODE91
GITBb+RX4sMgQlJPQkA5+9Kt48pTX8ZieJ9e5P9w+566SMLuW4Sr+/Ku3eCWlYRo2L1eyyotxnfh
fgyfzKU56KrHyy3Nv65uus4DKXb5POEKGGOMm1BvW6TrzjcSy0U8rzEqV9Ac/2c2k9wWStXz10nF
rlVzBmx/cYZZkIRImizkv9RIDFdrPU4dTUjyo4aBmRWYENfZ2jIkS4HkGpr+FUTHNgGsGqHOd9JA
ymkKfhgmEGIjZmXU5vpiE3RIuONd3+emOHGD1nXmh6pgGzYqofq2GpMSJPuJcLsYusiejL79kJzn
VgSJZhQWEZqlGck7aQwKQCj6yDCB8Aols7jNLLC9h4Tsf51ZwWVADdM47TS7B89wL7vUDsrFCEBN
mO9sdXJHmh9o8Y1VFKhyedcTen1SgVAEjhiF7I/XLqlVxu3X83GjIEq0jZ8jJdcbW0Ntdhvcf2Yx
XJL80QRcjgkT+mGAuQw0JXiCm3+PU89+ltgzQgVyFS7xS6DXSWJjzrZdAYxbEi07CBDWB9By+fE6
8uhBV/ALahKfJ5mAzC9/j1BKU0xhHUg+eDoK4/12Ne4/Rz7mMk+gdiNZK/PRk2ePwqq/leYKhCNu
zvyozFFBl6Sw48ITGo8wE7AlJJJWOmxrDij8mxZBAJumXo7NpiYBEqq23VfenUz6xkMa69wdskud
/0eGCGvsvmeOojKYopx/qaRHd6kueJD4WhXTBPiM0n8NQYjQ0MgnPwmi6sWgOGfNwtQYxI4c8uaG
7w/uvgrqgli2sA/Th6TgsuupwyRSfdSu2QXvrln0srmEcfueMiPg/k7NRUB7nlLpXyiWpIvOzW39
pHovJ9WlgXzFSjKHwrvzDsXx+cq9fu9qjaA5jr+iIo1NzV/9MzZYu5h9fsV/QxcVplg0YqJn9JPX
a2TB8r7ihzeO/vTrMpryrQVy7gaGPo3siQgSaNoOqTQVqW7KKQeDFzHuf3rbaQ0zjAQCwgtd8KAx
b+5dmgXxmOGYbLH9MFuf0n3Ddwi5MDp8555UejP+a5Vm68OuTGOSKt56IaeS2T8OMTr7SLUHBFYW
aRMIz0lJ5WgO/SL3JioD4tjf5smvyTytw6p6+XYTSHkIrqGt6qlRrnNbJmL+vL8t2+42vDsYdS7r
i4cJ1S1EoS7EBrT+z3M9R9C3JCE8rklwjMSWS5wQGhSqacf1hXy/PnJClJLnIwMQPGvvUqcf/SlP
YjvbHE5uYkPF/IIJ5K3rBCY+vXq6W4LwxzYAC10PT4XkhY/jKjqd3/aRXz63j3Lry/8+TDJUmEdS
uYLuvKJ+NjpF/+prAgp0s2EVZYDp9n/YCyAhdQyNIHVfPGm5HN1I4D+j0otxHFBbbWhTox5OAmWx
pC40jeAUWFkIJhc1Ftjnbe5pP4bzRzbEJDY6wVJckpuw0kJtcEA0m0Iepb61vH84Z+HBHmKuS9uN
XhHTW88gMsQOGzTPio0HQRqW7XNDGrdE1KKGPuuGoQUpFvK3WFihfquqtf7a2XZ/2osTG3EoumQT
2t+liLyrLbMA3JWEnyw02VguHbfEjlXt2Y3tCNx9Ng1xnE2n/Dn0Z/dnks7wPMOIUNJDv2MxI3AZ
fami6lPgXrcWbnM+BG3euQmosjrzmwAAGmGha2c6OLyTfcmk0kA67lQyZ/IxyJpgKrWRCuUaV+/k
RtonIfUXtW25YYsmAvrdxM/3xw6AK7kgIaa0PF11Pm6yS4Q9m3HRI4qeDVCbEYhO+EMXFUuBtAsW
+HFaEne/TT2RtZLQQxZeb84VT3wn2sn1yl832dDBFO3KcDckvO2vTt5IpN1OATNU5CK4fJWrXdJ7
viobKN/04luogTgxRWGUu13LNZptNfVnZR/8e/dvDemDddSzCGscOFc99wWWTygZG1f9mpO5akCn
DTnmmgsGz+QqrwCr1uF/VNOP1QyUmCOYmezQUPhwMcNmMHh8anN4z5yvJLGQXMQqnkQudq9LeQLU
vi+KRZmrsfgLV3/sGL3xqvPikgaZd264f0OsWhMrNnftk/gj/qeH3hmLPdcxY8ZwjwiLVuIaHNu1
pXjcftg2E9yQeENkZ26YUGBXtJLNpU9JhF6pl0N2I5FgrBpY5CUJnBf54kc8QiFDdVpJw7ho7fAr
JxnB4tcdmDdT4A9WNBBp/dvr4H1pASI6+ro7fFjIztI7ZjacdbUBSaKvQzdwOqLCkypsVVGq74Go
I4nmlungEuEASqpsaJPKJNRM78jXvfPHj7qHtRcvf0RraITgpKzoZwgV8z4WcnB46cXUCSgXQ7dA
owtrrs0tEvfr40O7t/23zonQ0wyXOa80ZACZNT8yVdlGfvrJgtNMhfNRbhsJbBwsKtvSdL3OG0zW
lI99iHKg5jxb77SgTyibAjtEH1N98vUXpLGQE9OByrS5Z50aevOTvg1DUDNYePnk5QXbya3AXIJE
jhKBALPB+1+bBOVa72fVOnBeKdGvqXnhxuq4mlRAPV4JFfCrFszm8Ds5Ko2Wtsd/SO28IkxzCpog
tV74g8PDwc4yCHth8XKGF/MkHhF1+gDYYSS+YVjHsKnmURYyR/JEdY3vWyC7hwfC44gTnuCWbP8b
RBsebdq+HZARjC2ZUODfGVL3zxukEt7YtuoyIcmLaozkz1EPz2XBObxOvwQhWd30Ne3SozJV8151
GvVgXfk0tZ/UnLCTGSX4Rf0L7yMrlbGP1wepWle5noZWbhS4xa3wvvprjoZPHlWVqm3SCx24DhA5
ds75e5LFd1e5iegusd+MuvwE+g7ReJcF/MaoKrTYCnHpqdKNd+2V8kHR2VhmzqzIBaamP+hVcHsX
uFr8EJpOUlD+PdzIE/kdfNzWSjF5tErC2v6GQ8M+/Lhm6rkY/ZZ55zR8W1TNU75KGGdElgPRRyhG
wqYU2o7VBRXEKuwC+IMnc6jCy3AGaWjZ/wP0tSDSBfHvLSmF/4FEXNlW+1auFk1yLqLbD1kXvJIi
OHwiKUgFriEwWdKRnV4w4Q1QHOigqY3Evt/iqKo0FaCiLxQ1VYQdoVlkNJ7rOQL/XIFdJm9tLTvW
LOAgq2GXB6lW4jg6+pRCIQ+tyEavxGjqHEt7L+igk1nMA1Jnc+vEOzeOHSAvCW2sexCYSybHYkpX
VB9dGwZEXFOaWPCTPrYUOXK0e737ntm4LNuuU7ITF7rLg1ctdz4kEhon6Dd5pl9CKHREY+AssYx5
wwl0S/4E4bM8+qybaVMy1qV5EYGiesCZ6f+z5ITq60cKYYZwrwZCqc/Z1JpVDiqhPAbIac+KnV/Y
PdaLFjmtG2pFZQBtl3U0jESTTtZlOGA70IAANj7CbF7bzj02edTV6mdfTqk4NBChD095pdUFJbnI
MyVSs0mYwlJ49t4N6tF58fsb0c/MhgEOUOcnjrcQMEAyfptVvDqOXrqKOGBDSkhl+DDy/aBipVwB
jvWl7IX6bOOR1/gjSz2sjUAP/0UL96djhnztfWCqJCYeAbxPDw+0Lftfov6om1eXh4vzw0+6lvEb
+shns8ypdcT/jMgj66hxRGEUiEGtPGItzXOhiVHWuDoYqZ5T5NaJj8bdgdUWtd6DD40rJWdb8Q/+
GTSXLDhcdQFzV/gGFsPYRCuKK4+pf1LC/WmwYp8SFHhqJXjIMW9/YHaOXc2eLl3vg7T+fo2+AzYM
Nz0uP3JmXss/0i1Y2THY/wdOfsKXR/u6CatgZzEEWvJmSz9SJOe1pNedmrXwFE4nKUBY8gVd1xR5
dsQKCERGP5LcFr5QUSAqRT8TajdCJAKhmVOMvuvHZnstCA/q8MrWwaKJRQRtPoNYZ2RlvzIW8FUR
RFfAcsRJMfsW84Tz3s1dqxfkryo6kE8BHgaeDahLkdJfICBSgjyH+RIYYU1lynbF0XxyZPscua1N
FiiEkHJ2qYzoKcgrM2Cyx9iFg9ODi6a4BDYVQjt3x8eofN6xOkAsMHFRkqk2zZjr7xtvVY+hbypM
BJC1M4EWcr/ITvUz9h1ZAsRhTuSSO5t9oUSOfVuLhGhZDbtTcW0bdhwqgV3wVz2TnaUbJ9QTkUoc
hQOZeZ2SLAPVbPLugrGPlwqd2bMpCB2b8rMWX4VNae+bZGATkMxjkg+i/Hh7W7sdQEyVKNsf0Nxv
BqPlYkVbWaLHoCBP3ByMBIMWJ90N7GMrtYjynNbIC+TL+HvBtPtR09rsegCSlKKt7joMOWhDQGv7
FqTWHhGl/CMvAArJj6yqmA2FzU5jly5s4a49lGQoI3UOTTEqcVkicYD6GVWcf7D8WgK8uFRFKQVQ
Q7/zrJeDCWBBikwfI0H7HMHTwvoUwXI6JfCix2g9FLTiYD3q6esX7BlFJTyZsXVopEJnPsWGfTKA
zCzqFzA6LXEAdU+zp0prIeZdKP9nfK/RZDeSwTTFWUH0vNnoqdfNuPDi4h1f8nhgazC9tsDrWzjx
qfLPQcuMAzzx5r1brqb/B7g2M7ifWsnYBeikd1R576EHUKv0OT5JGeATNaNGgBFHDr9zJ7aDpagC
t0U9+DoR76OMKeHhOvvCNsgDXpNDRV5zHPoO+6g4dzJK8slFWMuK3/UfKVZtjk/AzHXPbcNdDb6v
tvBe3km2KcN0iL+0HlgF+NT9wcqknM0hzqjszQYcRgH02Nb15Okofphd00l2Dp5U2dNBiAKXuTFf
8zOtGeYYFByZSWF9uDFx5mgJiuUfmC2mrkd+DjcgiXWRVCcALnv++/PIvh4k6/nfOClyG9awQySv
Q8wm3g3aZhO/qwXWFoI13sREdZ3MUX4EaPYpKDOjhHLXXgVdD+zZ9b808SWUGqYYmo8oSvtXgBIO
gxyHhHaSf75RRlFiqNqNZYGRod8y39yNiNYuZQ4apcXk0qMo5mQkqVZzwmEsrlhNHRti5umCK6t8
dkU3pnwsbmCfZar+B0J0zGMOstHoKwcz0RPTXLYBQ7uOQUGvcVUbGKj3ZI8HCyljlA2eUbn30YeA
YNMuF0lQa83YZAfhx+kqfLIubKKXnQxO0kbJTuxuoCm8VXPmkKHJnjLy8ZQsOCkqxiswLj+TFTel
0hQ/TXDb3iCp8UZWrTcVCLFG3Vevi1l1AB2gMXdwsp7ABkN2ago2vjgnEJUxsGgqjyQcW861mwCA
+uvpUbwQrJhq0qe1e2mEpTpaw0UfanVNizmwDuXStGJZakHnK+cw4wJBn5u+9pjM76/2ym8aqSAI
Puki85ng3JMb8fKj/0vTKPmCa9XW6zRPfBlm/g83b2SE5cozbsaNSB4WSubx6dn89VPe57q7KBkp
vWJW6clcOPJlvFpaySOo3oX/wPZuR4a1SHyLyYtOKsnIGPuNQit6zR0tarkx1oJ19ww5aSKcUH9a
h9AQcA2FcqySY/Ng4afnxSqivzOAdHd/EZ+p4tCoKHT0Qei2r8RLolKN0G2GArOTc6Ti+e6yfhXO
tVsJQEzY52GIzSFGEBRMT+XZFBVPsd6W58QATxG/vRsqbZtI+t/1FOheS024ovY5QdR9oGl7sOfT
f05mdzGERbkOJ/zKvxgCQ6ikQ/cuhBFXY/V+zYXsaQTsBt2v7MvG2xeRsGn5/9W65nau0dL40YNF
IaskkGPC0HTLibZLAJBsxZY7PcdfimBA0tjKFPT5CqOMjdzbV5vLVa2u87fQ8e0pDDK/HeBRIvsU
Y2nklsHs8R8mD5V68shn0TP84MmDtvfrZXrQoFyMO9WcF83G86oVTdOJBjZmDDiGfq38d8uUU79j
7DpOVF/mdQ1X0cY+BHLKbrq24CH4eD+uw2sV0k37z7M1vlN9MJ1BtxdAqKMtgdcqdGqaX9tEeQKL
2M+y2uWKAvxsbmdKEJdPaQl8LLr6uXWsZd+zP93ROH9ewm3rIJgj9QKpHTOMP//3P9Dx6R3Imw9Z
S9jKqZ3o3/jaEl6vU4XGLpGjhBcbk3Zf5TQWgK3qcQnJTeyaA1KnYvy32nMDqehlqgwu5himXWhU
JnBNc3Zn7lon4YWAFpKoIW7aXlgLU0e2FiEQnaoySSO20qTds9pt8XcanaKghON4TNh1ol5cXxFZ
Pm9DSfj0ELjQfqCHzA4wceCGW4o4PmGVEqbzlE1+TCTak66z6OtDXCPF9bh2T8msXjz14bUYcoCi
t3n06g3XMeuOLvZVBTe1F0+1lkk0q7zxfcI9JJLuofVK6WpjOG8F4JD8PxzuXcEAWGHN8TzwRHfe
IUVL4eYUaY3GseIFwwJYqOTb514aYcErN5EXofpbwJ6N3gFduGNt5dmS2t0thJIfRaDeBXBwcX8O
37jzPyU38EbhShAN4i7GUIabMKF1UAqgK1x6aZFsuhX9Y849xwisURQsbWY8Hdy0gfDYa8QMx/xh
/VwlpasrhBCdRA9F19i+yG4N4McDB9CQjG4TIkELp5PUOnJsNIwY1cP9OuRrA3AFmHe5cbbHZZl3
3hhNAtz5UPvIDM0UW5MoD8j1lSGDY7amey3lvlUPyVnJ6Ph64aKuEkZmJfKU6uX0u8hysMYBECgn
0nAVDOr6N2wmQeGVfWLkxd4ZWzFCsMB77feNTK6MzFXf2KZVnlg+skdCv8jBjMXza6UMl5nqCHr7
bxn+AQEi/rpKnrS3/FJMxm2v+mJe79Q1r17Zru6QclbM37aSQ6oDI0CMl58ceAt3C6cCJVCqKl+V
9z9NF0P9E4FIvtukEAowUqLO+mNG5UlXzzvu+gsxgxT2VJDlZ5xmQfzjCKxPVbbNGbdgw4toxBVl
f6z/fLOqBL/PvFIg2R92578/Gq/sz0Pb8ipjo0DxxicCMphz1xeEGvCY7VyYcQTWt8W8653dhiMa
sYINn35NcZQeoIfWoDrmRLzL7AYCXmMQ8SchQyx2C1Yk17his62wZ5pjNCfTnsVnsjKGQhQpic6p
0SY7vFwAPWKdTPE0LERcc08WDqPNrh2wRA/q9byCsGso5LXN5+p8IPRVIFChtoItrmT4DOV5YyS0
TIXrI9YM45E9sbRbslG5vCQsfY+Rjb2unOTGKUumHxgOam8J+TwBi66uHa9jR8CKoFAonc37tY78
WNSvrhFwqJV+ekx5+zrYiKJH8G/pA4mDwbHFtFX2yMAmW7+qjcYXv1prz7Q3xciG2bDXp/KWKaDR
JYg0z9Y6QBM8wq0ngPzHvMF/18Mr9+WhFlqxw2QxgKpWSMdsrhGwF959ZpHNHs/ySBRv3Is7wAVW
cAatNnoCJS5OogfU1nhRG++bikW4yW2xsoh0rS0+Y1BkYaZYnPNdx1kFTzUqFBGxdFAUm7iKHgmv
jLl9E4nzvaPqWsgH3DG04CVW6hNxwxKNvFXQelWCGkSRpMHcIi2FAr5oOVbZabHLQmO2zYuch1G5
jw/pnbWlLhRqA2UycUarDx9haH1rUcu0LwdTWf35og6QN9CC2ZgsoPruxzJWmxuCNs8NHV01RRp3
HkffBct22fxtGg+vLoUt0hjEU+c+Q/7Ts0cVtGwpqkinZKPtcFo+LtW5uCQhfjfJwUkD77dhr5eL
Inzlf17iIVcCtdDuR4IoCs8YFFfCfdPxhCur+IHnrRbd7Mup6hlvamDhCPBeUacswvXpuSDYBHmY
qShK9EKN+fp+tEYsQVNbvqrSZRLh/g7gb6jv90UYv0Hx+jJsUHNxEGXxyNrqtK4WZNpM4BKKWxfG
lVKil6ZbPkH4yTKXZey73GskBhSJ9lqhSw1JI0ui0jNyJCgduy/7PUvSJ2WXmhhno229irRtCAI2
WgNzfAcCY9IEPUAE7wrfhyJ0EDNALNTwUPlboTpMwZFqD8JjK9pyG5x8NR7gW2oWNbSmYN4PFVzy
v6YxAH6vfqSNgDYJi3gmi9DjecuQFiS4q4HLrqEe3az/v9KUDiH3m5AukiY+Ny2IrlIs1GSMqOwR
h4HkjAVdwxfZlhBdPEy/wi7TO1NuehT9eU45ZCX9GEHHGoVwKPOnMlMAZQcI61dX/5MKJx5O/R4E
6ime+o/ObAbKY30VCA4miVFHay6GbUd/ZBpqPCoKcLP6mq1PB2/lfKkGvHRKeUyeop9U0nL1/SoF
JQCqzAK6bNUfwNAIWJQrJ6OV6FdBOUiZkccma0PptsT9ry3bm4j4PLKpco9VRbY50zQ614l3DDft
tZRomt89PX2Q9QKNq7f5Sa2IU1yeTEKFGbOagQvE5ZAlWf90YH+dbOJPGAQK0jZNBpswTsrk0nah
HOiwGlkhMDb1N8e3VIqqd34gkLC8oogDCmsMkaIhKwm8JzNR0KAgoKnJXdu3YX8No0koN2+cuWon
+EC0PzY+2gf95ARimh7t++afayT1bhf8epfvjgAOzLi1oIxEUTPHwgd/IqSFJMeOGALmRxD4AdKG
slRT1eXgzTo7vdOFVbNKsfae+X4P5arIKdf1V57pz7iE70IeogMAWmwZ1RXrze0RuCKYtpTTIB+s
Y12cUK+Txc2G8/sYkCcztKhAUxfCW+4dpzgBWJ//1CDEzJCkGqYINXa6Bcm4cpNiVBmJzfPhX7U2
V1Ohwml0WRAG6Yz5VTe4wbVwKeTr0UsBvfMB0+OudLVM3NaXAhHudek24nUqGWIu+ZKgXMqjQNlQ
Lk0WKl3ydnjUq8jTRyMiWUn+8dQENhZdDd29hHTwXArlMIklnejT6RsFi2zxGwovYpNQqI0zD4ZY
+qEFu34IR4bfATxGMt4o5oCnEjEcXlsfmD8vNyWruWoewKTHvdfQ0EkS79rhgx5fvAedppZiNOHP
f65p52ZGFMaiu9Ik22YWwXh08kh/tlMS2rNkwKc/1u22lzQn9BzGnYUkLUqU2dH9I5hrt8dlr9Ce
eZCInZFPvvNbNEQigL8b5NYLgpEO1pEH403ygX/7eND/bOeSS7/EyQ+J1zdNFAlLms/raJhb5RJ9
/FpNvdpkrOiaAD4MfpUs5tEWiYsgPHFECreH+G98VbiR0DUEeldB5mh35Pjn4GTtNoQ8/NG871zu
Z5vB55ZjNIFIy2CARDMLTKWpMLmZiT4bKWyraCBmqtGnvutHcdca5UqSRK1OVtd7Gbvb6rCIrigb
Lynw2de0Huec0nAwJTUR+ZclEK4JTLucTm9zOh4unmXGkH1VyKsH2yNUodEaTCkRXrasgYVZ8nMC
8E6YJPHWyAtydgrKET3wMLgq+450aloTYAMaSsUoD8beCSSmLrexcc9oR/SYaTCXrGLe6JS7BLhi
RNZHh8CD7GQsTEbXovA2S5G8u0gFoJwtdct0IjzWDv6PR4tw2/bPCKioF9Z6laP6g40AffymNRRZ
nYSaDRILVB8J9HjB1qGrPHCSFrvGNG7KpVzERKXHPQLqb7WBE0tBaLxvEIIuZOmW1ez9Wz0IsZEF
yMnlu9H8AzlmitC7cDpspEV72FxL/vxXLw70JOZGx+ra6/clzj6ZasqGonaH/B15FK8NKn9sUl0f
roq7bSo8/nBGdq1r91z1BxRN6zVlPzmUVRN7Gs9LxEUQfnFeLKdMUolnMWNArrLrcONnirUr5zR8
m49xhKQR6CznwZzGtzeZYkdiaOH1isR/B5W/PhjEumJuOFYGuNg2xOI9bgym40YwcvaH9+6/5mYb
q1x/Sf+xhmaEn5F+61Ii78yStlsc8tsDpozOkzJzN/7AZ/FSbCZzX7QHQVcq5pA3gq1oS5ljTDMe
h6kvHKqlpyBxwFDUKxoX4u6fthJ7hkIkl9APBpOKSA4P0rh77/mgQlNHtQmV3rcna4c2m+f8pOOt
/1raKKCcWpnYeqmZGOsh9e9KaR6Dp1NJmOFWiI2OzdNv3+1Oi1wT1LfRRru3TzxVlHR1P+CKGFxo
m92JenzD/ZSDMsR9WbMo8wijkfxWmTc6umQ496TMHxuY0N4ardGEzyoL5gH1ULjZwAZq6G8Fxt1X
LfvlXqbK2MvwK8zu4u1ilvbVbyDJ7S7aTuTT5nASvPe368S90B4hGv8wLIEZD6fiRoplte0tIs9I
LvQIC0iinTuKNJovZuGKusxSYgBA9U5KHXVbG9dGp5o5YkxIZlRf2+8KElC/bdrhg5rZpKhpIQEt
vJ1C16gFlabOr1SQrb7DVN70hpExtb0aESra/dwwi6dyhbyu1nWk+Nw83WTFpvdeZdeqDyYgMGyL
k4cLAEcj2UhL4dLeDKiwThTrpO8DxNeUcQLB3z9c+FWWUa/0pDvyX2VbOIHanzB7etsyLEWeYBr+
RsxS4LORN9nCeQtGw9eWQYjPW/CV/RUa573Ebr4rT4WdSxFqX+lTE14vmi3tU8fu2ZmRmj1toM5D
64F4M7bOpOmoMh5T8E1Af2uyQI/0GWslBlZC7rRjYpmuEUCRoWXWjhsa6MZcDY+mw66ZTXwaLWpT
YoTiMtUyuCv3kb9/esZ9KbwWI43qG6WuYR9MS8mtPrLuLe3RnKDfOnCza64yxSzmweacGAYfqxnH
7+nKkoccMJ49zJiaBuFQlsIYtrOxp3oxt7JrXBkBNhiKhiE333XL2lQsi3hF7jHxznAeThcL19iB
zbkQAo6f+Ag6w4ziYoPhOyD6uzmMqwl7dYEXOreIeB0T7oY7dnzYxPsQwtx6V0B9WOwIjPEZpu+P
Ou1Y41dJV9Dlapf7iRsifgeBB+OP/30Ix5XRE7IQhNFDVSEi9I6LiS8k3nAhrXj389k2evo2dGHT
8mOMYflwF8p+5ybScPDYcjnJOnOqbSxfy9TaLWzLEqIaiUAQpqEM4on0zD7gaWkef8QO4VpNetLW
Aswl4Dl2uUBWbQ7Hdlqbt8lVe7elpbQhzB5DPhMo6NW0jZe+ekziYbBwyfnAnD4UqgpAX90fygEF
txtaT76+Bh+PlgH3160xi8sJcMXCWwi8HA5+BWe/PgGev9rei7fjOdD4/x3uFTt+szi0zdpc6SbR
0bQdduNoml4EcBQIeEvwjKaqb2T0qhBMpGe4fz6XpcsSH8p31LUKuUBvsvVcdgwGAiqgLBZB95xJ
O3RgoeJ/Lz4/XZZfhrI7wCRnt/KfeNV8jZP1rwaX0akaY/Rtg39eoqAoH+3zSeBOY//3gS5FHlY0
ITtWpoF7SlrmFSO7Sx9/nn1hx0/R15aq1n4lH9gqlYY2bhg49l1sIhcTV/kbP03TB/w1XttNZPor
3TAtRRS+/m4VEY4UfabmcVBTKQNAD3Fm63XPeGY/s0zaTnGpDDgBXV8g9vxvcYrP/rSUre5dvSqu
qUAjP+kRhQKerkZzt7PeOmvicYwdk/AD7bigSWGmQ99ReUSMPYUvrkz77Ck19jh4d700gyUtQBY7
luoR4dZFtpZZRipcZHdAdS6Zcl3jl/ZIstMABF4Ad0/BUPDKOS23KW6LRxo7Rs/sYpRnMnyOPu+r
QrlBFCLBTqJYCJO493+v1Z/HE1vysRqxy0NVuXr6H4IFmL3loUS05XDYIfoRbjXlOLOgrcJpwfgS
BLp1D6g6TLILSNWzIN3pzdFUCjYK7VLprm/lbbYOoTCncA6Nsc6MlUMIl3f6tfXFDYl8mCzVHK+I
UH38fHwNbTKtBz4MIDiB3ri53fFwpMtDnK8HVeAZBus6pKss2kfPW5CmbcOZl7gYYzlfYcYmU7AM
TQZCO/1Ob28NrVgbkAIRyrY0rbolclYuHSPUhJp9jgiJvgGPvbMDdpCW8UJGElxjUb6frWNfX8mA
SRzMI26Ekd+PY0oyH9IUhy9pNPhYgJZ29b5JkFaLVwkb77kcFJyyR4qOHj7TCLLi7j75mZYtuzfL
hoQfc6av8ZRlWpfghVqkzPtWAZ4uj5+C7tRXb0BBlhjggW790dAiRezA6ifPidM0kb3/xHNL27ag
IK2O2HMZnQIaOoqFZ9cF6Uu+JqKOt9xtdC6oO55YlB7izAD0dBUl71wBTjqlYS52nLl7KDTvAyMD
IIfXj1lmDjkFcqE+CVsR1X7pOFSE6vTPqMQmYfkAG/VMcTJS90OI1XfWb8U/R/Nz8NI9Wfpl45wm
/daWZLyp6RPz/OpVajXiOnROQL9Tr6F3yg/uhmwjlspMuPNqtw6V2tCDbhucXei+gQuMuWQaUHe9
RqKc2eNiYLkyE+LDjdCtLelGWZMq7d+UIgC7aj4WLT/eVojQkeHQVLABDGXNMdCQ0ZyIeBFeqOEA
+dFUki2vd+mr1r6sBPyzNIbxIP64mRmDjCKW/mAsmt8jvnG7v/LyzmkZ5aK+K0jPz31iZWd/2pPm
qbxZUEJW1cGlN0hz+FncHTjIIK4Xf0P9AJiVa+B7AGkvuBUpLiGAF6KZ3ET5JcLNDaF2+g1PxzE1
DYCXwnVewk2EjWuOeFdtpu0VVAGDx3+CrWMvtgAX23st9gYHljLGpDSlWXtAlAXl3mh183ETlg+3
X55z76bm1nlihClFEHwVpml8WXTt0OhgN4/3/ZBR/DrcjPX5C/gyczlZOpM/fdW5GyCSaiblQII2
WdtEnPhKenatQwT1azk4xUq/0NTcnS6t1GJ7SGzYtcVDSYpmYnr8Bww6yCHnlh32aYFRJQUpfj/p
OdXrqMlNWe0ahn8l2b7rGnkaZw4iFb17yKw/LlVupQcCpeonm1WwxE7o8K7mbK74aEgfEBfyU8Sk
IvOW+2toUq/zGXxHC8tiMOAKREj1U+sBdehY0VtnyL4pnwho5BX0p8lorkvNnLx3cMxiE8R1WZOc
jvuYZ8S777fGSEvdWZU7IMl5jjIfksiFjDx8jCeUrNeAtCDt8E0zEZ6jHHjsZ2AC4fb9vQ0gJTzv
czzPgYwqAExCWfdL/tXVeYGlf55SIpz9EEZUa3wnfR8huNezampmYnYYK8/kFf2IO1ILWmT2u3fB
GEDq4yAN3opj4/ZrFrpOFhjXy75pdtK8g6tNSuqRVMfcykpe/btjDqeiyqKdGLwUjeuM6ZGcisBX
L1gXi0rz0REBlSZWj21PWoDFkyGboGYkj27gMtkE8oh1LvsUz8sBo8pc6Le813bOemuDVAXm+rhr
3CPlDd9jpu9CKU0eA/cFH+2zBLd28VvbIGwe2eb2YhsdIS/KpYI8+axcSAIvAqEBlaMwHF3Fq+Wj
ZfghogQWZu1PWec/kF2E2L4u6PLSKBxJWTUJC/gfqunOwCFwbPyIcipbvWpjbDn9TSpiPhMB/w2q
SFjWMY2CVTBlVqLB3ivOWwAUCLlTc9JUJsXExEHP8v9xlo95xeKz2WHDLr0ETCs79mC5btxmvYNN
ObihqWsVlenxC8TVO66RBzU2mei2z5c/ASCuScn8Ne8kvcWD2JK5K+DFySZR7+qMcRE4iHGQ1vDZ
425efUszPENtGhzQBhHlD5bEbFeZHwtwHsy2tntghUSF2z+kzbhqDKPMOt+vCBp9A1sCA2dOKa4x
Jrn7oLOVdX9GV2aUJk5fRNVf/rCJuHFCMZstJMwfNkEdremB0CTRDauijqcvbnZKQ5mRxoVVGrOU
BCRSstl5p8bsQ3kFA8GkvXL+2U7eH9nWxD6N9jO813Iil1tMPJw4he9jmU5VLVPhuSixk9H7CgcS
F9gsW8G++OalhfKVXSJd5vumLyjKON5GqyFGFgcfyShF5gz8h8gas91VvkS9Iu/m+auleEQCmEAa
n49kETFZFBMpDv6t48RQQPoqqKZxGByxpI8yQbOrbNMEwY5g41ll3Yftg6WW6upPm++Tvc0Ek0+7
W19Vg+XsZL+jzgqUDkZjXRlGFnjWCXQpXxqiUFNVFQPLCnw/YbMymwukEUbRwsiA86yhKPyVwECJ
ejluNxLw3AkMuuMFMXumu8BGLNk1svUiBe18FtZ1yMKMzIt2BJfIbEGFBwB/3MCWAgIO5RFXZjk7
Lpxo9wrO93TwArHqGPxjyO/Y8AUzlXRlVyaqf5iRKw8bW0bm8OuX6Wszcb1yo4YwfDdXOL4LcWR6
Qxdl9TAuD4s1MNDgSapbu3dZnHnNHrPuGstHIfYjcTs0RBSs9lmOUJ2rE3OnLaq4puybeSwh/5oG
go++TrWOfQJB81EV1V5UAJz00FYWE/CNjxPq7+dXaiB4C8wKmlZxWL70IIfks6BZCm3Wy/i3Ck+2
a1PdewZH26xEFpiyr9jOeMzMlqC+Sufb+IVCIKJ4XyV9jZqcs9Sshsjx/u1ID79ZAArJqbyVZMja
CQYoR4qhN4ZDnIAFADF5RgbjGWNPgd3bM7Jj+A2JVfOeU1yxNtAulgTaSFmwWzjmz5Qo1VsgixUH
bGZuEsIvD8rNZGgdLkYRY4wiIKua2QnMqhaQuO+doisRw2mQ1ZOna5IXlzBKPwslZG4f66HS+tcp
DCW17hhBOragXXmgP03ZfKd/dI4Tvhqt8WNuyXcG1ZfENsqj5N0SPUCuex49iNL24Pg3PhhoY6XZ
D9lFaalqAW/WRcbLGMmyon82NTu8KOW3C0LiHS3nTb4P88GLHksTKAFIzx0a53uFEd8ec5JCzp7t
1Eufbdr8m0zdQ3isRII0nnIrUg5c223WHS43XYTyc8MQcuLS9qAbq/2Kc1FU0PwkEf7Si1UpvNXI
0yudyofCY6lGRytw7b667dF9vNHvn3RAcsiNmD8FLtq3TN7p599nuXbgWRSnxYQELbMXeAmQXUsi
Bq1jCIPFUaH/DsQZZh18S8b9FxxOdz7cOpc4adX20s3O+WDHSCq8TpSccNzCpEzGBAr9Ewv0TKiX
R7u7haclNRnXZlw9BLPAtEcmqAWTslM2KSfnxnNISMRV6usJcDOKi4KZ1K/LKrarZsveBrWVzmlq
8dcxqn/N+aPYZaQxwEu1mcFtHUIxuNS+dSnu9NyWVlspsfrYJPm2Z65PSx9ilb9kIDIF29Drxkih
Cove4k+M6XsbPjzQUGZTa6pr2a9hGoa9hXsKBkUStlFOMljHiVLBsD71w7b2P3bGLMfv3PmHu/B6
aeNqjDT1GOpTWxwwh2A7Hjehl3b3f+MktJL/VHdXiJACfBWqufps/+g4Y1djNbMGuvBoBAuQ+pfU
CbSw3szOWt+BNX4+V233/yVnp/7WcZ1PT8l1aFxs48AJquD7K0Ub3O9Vmxh1yoc3xgS1o5+io9a2
QmbBmUlfoeRwDSfY4AqsT2LbfM52L1Ss3VkQ3pItv6nffdbvpVhNBDRmK1miX39Rpbg6ksXUpuuB
1n8tmSDeQK+BzbyrEHCoOSOeWSgM0O0AyxPiN8PVm+y92a8JHwJxKUli+HZkVk/MIisF5R3sJN8M
788rgXqbKy0nid7ugJ61irzDyIPpwkpqgqrNoOqI2ne8ktZrEzfGurZo07bXQCpLWbPSxzzypbft
vx3FnESWbrCsR1/WrL+tCNFthn3Asnbf9L1IxyORgcFqcVVEDfW4P1z8cok6OUyAVo/oTyytw2gp
tYxll1ReQT0zK5EknU49cvAnIa+g9Jmb4HT2Kq77jtuBeApzaXzTZiAfpEu8EkysuLAbh3dLyPvI
1KGoVw3JwzGpTAICFhanLZkZItkBo5zOQvKA3VTAgIC0basNWF6U2WPG95JvaSE1R8zmJjo3V9yp
pJiz+9GL8HtMo8J3cnjRIGGvKTslUqua2+qc8AgoIjiBxVEKv/VXg+IwY4IzQsf+vvcqbyN+e9G8
wUBIes0ew5MC2SC48rFlFrrVh3tPOaJ4Q4GQU8CwmfN05ZEksNzUCp2XI6garfuGxjAEHJrv5Eef
UKnn6Nc+EQzngUrxza3TtVrzEUOgOi75ges+qnH5kmHvktrYm5unsr0d8DTfQ7vLamLidJUUg5uC
Nh7s8jimBc8QpG1VmVHD2B6YoP4f64MCywY9LffqkzUKr0/re8JeKi15xlx4BpvzZDPlZda0Zxts
WEzGx7Cn2JuX0NUHxHfJ+WQufGsJrNUOjOtTOiS+q3z7m8CsikDppPHpEJV6Bj6OTb3RvCDemA8v
lL99LtQXH1rhZwngfn5qm+blN6L38NrT9VuXMa9Pwq93S1PvklduVmUh/gXlQjcqTFJTOQXYYF4J
GK1ECHjO1M/3WZAGkXwz7l9IWLz5MPzHTLVt+zrtHZFq0WIQOW7BLSnZyqsCfKlXGO49nNUco7Ry
BVS59lKTJeSdh2Duae3Ga4FtxM9LwgE704HMtmJsg7x60EYqMTOUc0nhf6YbjLHXa24gwd+wduIU
uehsnisYKjbQWJ66/NJcze4jc0KP/S6SufPcLSvxznVKkNfDLlVusZzsRGHVfXg0O7KVYdoFI/Co
ptGrLusL4iJAFz7+3tosn08i07nvpyf2/ql4nHJ4T9Dj2hdkEuvwM9nKSCLhO57bMV7a5FpY4DKe
sFjnUEGrQBeA9L1tv1SAq1i4oa2C1C/2in3IdgoTe/IyrNYmLZ6qx7RVI8PsHnhzjU1keLj1KoBO
fBS9LXR07jRksCxSW6NCxf+c1gp2b/jCRS6zk85z4PkWdET9bDJFizbybbSKYY7Lg0if+slnpoPM
rWvXTsUXHQGS+FK9XfTwC5+dfcfmnNjWzQTlEu1LnKGXAsVWbATmXXLkACO5lzb8j38mIslYqCsd
l8aXArztb19iawYLSGna5LJ7RZgbr9tWAlX/H4nFrIlLFByLU+C3LoCsWWVi/ox+ygbjwaJlnBpz
3RoV17RY/5gWpL8hsZmXb/NuCf259rsfGJIrc5UWXp5zTfGE5o1cKIKbInvDVR7UzN+wOnKeAJUu
d8qFrsGnw2cZsEJsGpU+yBarPpoavuPAOnSR70JiGOTWNgwzbMVPsvh6lWXmOYWE5s8fOoJkUFNx
DtDKBoef9rcJlzVx8wmzsRSyStbVd7Yc34F2vBz4DIAtyGUzTjk9S56gHGxs/8UtvV2XVfVAgsNC
tpTjcZLvadMl17EzaakxwmFdbmjgpZQiFq8wgWviRUXPlTeQREeoX/iTqSViqi5bwJ71PX9dxmjX
RdyAgRlLvhBH/MrSJr+e46hs50F+BSVIrdScfgZ9bsaGRdtih5OXMFQcwuoPNqvRERS0xTuKNYq1
6P/zzfn2UPzQztkXmFRy4oyXRDvP+rqJTZEHuc7xRY+37+C0v0RI2RoLehhLyEtqHhd5BUZSOfS6
JYw8Inkk4fOmx56NeoVzUFm+V4Hw0cSapL1yYCGLzKFwOEXl/PB81Yv14wsvfF5GLOXf9pT8uU8c
f/XIuqNSQflu0359WVkFctbQ8jzfLZ/42rO1AlSMsWPj/SU6NAQbEPlCyuaj1y1bePsINydpfuPO
bDq5C3sg6iYrYNjhRv+WNP2RYYx+m2uLL5U4t1uRbq9TXdAceY1b71Qo4XrNKPNm+5FpZ5pskke1
3HJ7xo+GNBbdUblSBYZ+fJ16o8IwabMiHw/RIlZkkDAnaIpYatiTAPIQmZR7qpwO3EEVeuCmOrKY
XZdXcbnsLskan62eumzPJ9WCuBXpqRCzaSe+6c1ZYKimvrMWZUxYjOu1wYY+xOgjRA44j2VEVlXK
JgPVrePgcTtBhFkw7D4BXPetyVwkbpc5fHTqGncIM8dVhM5r1crDGMUjnjzLZEEOcxYnAzwSKbb5
EV0kMtt1RTaoM0fzhuPGYzOQEg8hNIhV1BPnCETPl9p0JAwjMR7CtSSCjPDjZnq6PY/u5AnAObHE
V96NP2Ib/qLGfcwbK3EXvJF7Dhha1+nbaek26pq5wIqixcqaKxGiLschg5Qo1j4ZqX62Wi5eXJmn
L/O/Jw6A2idhVluSBx5aB/Kilvd0lIhAZnWLKdE77ylXD1QK83DCK91viH2CzGrQwGCXVMk6ic/J
aqs2c23XVIE76ia+2uSsk0LXLvzXCzlvzGxvarAC0EuV+x1LYpWAwfal05020VP/EntaQqQkUWqU
RZeb6GDU2/9TQDDxZm7F8i+JTkSS+mn/xs5lLcbx/3EwDvxY/CMPrUkZevpVOzpk37cR494STNKN
TH4RIME+/HZVjzwrMua2dD7liGgMwteZpu0uDd8xU+2GhV8rFmEsSdpraw9KrAh/uRnTYDxCUDku
vLvbiF1e/ixPeb7zdB4CN53XG7E6JEAdiDXGzKqUUfD71pConecCv6laKXeYCLhIa+K38j2Cm+UD
BkhfbKo93hv41PkSccklV7aVmtxzkkfJwiDtA61xJHUpA/GsH2/GuHC5Ufnx3GRkAIQ2Y9oX6qTb
eJY11GquRQtqtKw7s2P7jsVoF2dhpH8DkDtsRULb8kEHdhXavblxMdBHggFJ8wvImIxI9iWDSaNb
8E0u+2rH2+f6YaLd9bPrhxXGRfwWPPHpwVkLU8cZxuPk9xPNQ8Crhjews34c2f5YlW6gfKFvteaX
EkXij/UzcbQ3jrndoiGmVxln0IWoTWUhwxUhRi2JkrYjKMLtP7T4AQELgWbEAHyT2pOlRgxyJ5ac
Y/oGG1Mbejg5kizB0HdsRCJ7p1yZ0cfEc7hx75vHMruW+TCe40lpx5412xRiwRvp7vGWIHMQL95h
IQTZZ+5ifP4oNGHsm1OguxPgWjlYZxZxucSqTrs1pQyngO80icM140lwBvz6Rp8LM8X0i07T6ftO
8RTZSti7NohWTu4uJTVQWuPoFs/A0qe+4e/lnV0GpC1n/1Gh1enomaPaKrXFiEqVcq3a65wgFUa3
qqawGEpFyPzuwId3jPuXnFZ96tk00/SmiAXgk3XcLwHWET+dFnOja1c6eh3un7sluxji141tVQb5
Shkt2VZ9f8MSYAmy0x7dBpv6ltFF5h1SIFa8DvjbAvnXdSjFPzNa3xXYpEFDhJYxJ6P4Xtv8KPUx
Y/sNs2DJIQqJG2EImys54LYqnkgbesLYN7vVD60Wk+u9pxRRbfsERsQHLIT4vaRXTY+LfRiVTZiu
1CHQm9wetMBHOs34jRKf701ky+J4USh9xIEiqXV4ta7NIIIYfio0nFwvIvT0WE3kGKIVhiZ16yRU
cDBzt8DUaNu1mHFfWWnNr5MpxlTtcfAG1lzHZKsdF+ycmRT/B1KUY+Jcl/BnKkEnhFfLVjyyOKw8
5p5OhgmPZi6aArpDvVzNZ9OEVtOA3dMURDy+bzkSS0Sus14AprJGNWcxM+Kgz53osr9RjJ/MjIv1
MoH/otZ4PMnV/wxB7vTx1aCw5MxNvfU97GU3SMyw3sMRuERlIcrPF8/s3mxC2ZYXxnYbZpDEVAM6
XkxYpq0ILEJb7NW0cXwfSsmxPbXZ3H8DaTJpEWTUi1M//EbDQEIM+/fVWZ5KODq+P6Xq0x0cnYrk
EEnvkriz0ct9qEcD6kgclMrX4NqDbINjZWA5v+X3jlai3O5S9gz3nTOgLfdfsazGZgEnY9PYYtkh
dy0AnUzDmbeCgpMFznUoAD1kwzpPsiOhwPYBdolLPCHRjnW4IhlfdnIDlLEKthOS+rcV31ceTNlo
7PgN8W3fgNVRBWnP7oom7ySOHy4EgxbEvtAQh7LekB+SURoJfMiSg2lpQA0mZu3iOU/3RfZ9MlMK
Jc62YatdXT5ceTwgvT4zDo1CM/M9MsTW5eClkmnLhN9wqnEAIWUTsboEX16eH0mjf1t5qX/U5L1K
VMx57RvDAVxQ3/gZLJz7OLo1h3NoAv9Y+RESUDEi/RkwdUtG7R55uuYCPD1GCd/Jk6rTDyVTOH3r
yVfKZjGdUwL2e0I6ymbpjdDhfka3IC9jjQlI/jDSUd86F/swVVVhmAtZIzWphCpmJbwoxQBL/TIa
TJtSC56rCRclBCMmoRnpAuJ3t2KjxLzZ/mGolhebCJI64As8kPrKdR+1F67fnr/FHGB4hvjVqFYv
rCm8YJBqjJF3IfO6QZlfn4YSt4yTfOD6D+H8WTjX/nrZAyuN2hFj/MMKcNIZ92iwonCvV/l61/K2
ZFuVZ385e9rmMdNmCx0tr3QPzKxx6W7/eCYj3kGvHL3J3kwhjd5JYlTvGC4NnVaEuAzfzqBveHkQ
02/p+I7PDkrsHi0veAh37yrwxdGVa7DXxqP3RaTzEieVcrm9c6EE1ItFMcNV3RE2cXofh8rJCmNq
s+KwJRu4fsYcs+HC/pLuF6N3eGo9/ns6gAKFQH2s6JrzBWuFiUXqNopVeeDuONXtnbrXA9Chqh6w
73GI4tUFpQkhANZRuC3CBDVy3xc9cWpFeRouvWTZKFxJGOBycIULxeergXMSUvoDqHvimEhGLLXw
LfdgMrKgfztbINLk4MMbVvh0fVi8XDtleXVMa23AnSgzS72siyazBmYruRmgEyF1FCvBR15vJj5s
RpA3zI0hgrCUQ4btnrfIePGNvl1wAs0zGWKnjiQn3TGN6d+6eahMFT3vCxpTKv9uV7jy1MEu049i
2KpqB1SWA+MXoLkWrekWckUJJtvdPc6RjwqHFtrjYhBIpZk7SW99+3DZZhjQY73R8WEtaZiBnXuw
otCgMXLLy5ItMD3GGstar28thUo5lVSzG/Z4EKnXhTSEau1FqcacntlxqVFIj5YYhVRNAHQrMhdm
AhVuUTvIVCmMa4S/FPsGwyWE325cYnApexgGosVJn5LyyCEXk9T7clhjF7w5hGh7amVQ+bX/UwS9
o4SCsEh6w79WATRxGEWOVgIt1fX8q1OjsLqoWIJedQEkue+H/pzakRBY7A7ROfuBFJ+Beoo+AkDu
tEB2mU+iGrTfeLkFcm3SfpDqbHLOAPVBOPcjLr8lHsKprlwr1WbAFRpurowepTaBMX9vMBP9xrRS
Thi/4j+xOM16Cirbmq8hGR5kxZjkFeJW22KbGQ1ytu6qlygRuOUx1SBFKZ1hGhHyEJy74S7iEtp6
UCEVRVwbEFTlUieLCfYyr9hznjEblSQJ/GC8Ad3ZxMDdpB5MDmN3myDY8mleoCysJVyyJmerUgHP
/em1xyspib8zKBJaxkYIrA3F8yNXm09snhtxRIFmiCbc00spNij4tXFo8boQ2amEiU3au9OUMv5r
SaQ+b9EZ5b6KVKff+LpwQrSmiQWuIiicpp/sJtfBEKH3uiA0k7cp89i3knPyzw4TCozQbUOeluqG
18XGSOZPwFvXR6+4fvaQzx3ws05jn1b/pOKyoVmvAXtPwge6dlWX6Vgh6VqysjypqpbwNkfehxPF
zGkYBYwGbVKpDeqlWpIxB6xNRY4EEBS18Fa0QxD5ZvlnMWRN2wNzJEVAM11xkLZQ14NyMzUFeYGn
TO+waLRxHupeFeT86nVTFOzy03ViXDVTvkzx8tET1lDKEIxSkaacolvcRfdg73vk6HsYf5Qg+Y5F
X47JSLj9XDaKnI1mJ7Ha7/l22azIybz7Ii3cay5iiEN44dLjAMIagqXGb7n/Xl9qfplrF4ynnID1
1ba11LGi7lDQM/3srBAbr+/vurmjKPN4PAOx8KaW16a1q7WWgJBQA+VuCffYGjbjhuXaxAaNmTTo
WIiidkMWpVNr0F8byL1Z1OTV8xl6+XrDqNXsAbmWAd2wuUKhAODYJ8AC0Ec8HypnwxTH3B1lc8tG
qZw/FiX0cOEqnuQcFyruFqW/O/UFzTZwEROW0EDupW0nOWMTl3Z7tIdLsmIkzA5D6E5SeDWx0pYw
pZNZW1OA3yl9Q4U8eTPsyyHLiVO/Ea+RzGj552lNJdjNjY9GRBiX1QvqUgMCvfUYd41akYQ8fW09
mnGp/6szbB4Ffr+7DflrgbIKqWjTjkeiZvg4UPcvo5My2bNk6/oMfOjDQMczL8NXLDQPp9qqxpJg
II32D/9F2teD75IXgp5Rlpms/y7W1DxpN64W+Nt+xHD6qryyn2b82azYTsKELHq+8i8rhA2bb8+i
SRLscxG39ox1jV0T/pdMqViDzW0sbPOiTT7YhR953Yvvzm/SuTSkitOaahTAGVY51yZvFL51rGSL
cBV+gJ8UgNtNn8mQTlQ9wMd/BHihFbfqwLNvp60Uo6K5Ho8VWsnPFp0fI0lo0i3FwjcItqTmm8Ns
yeYJ6d4vzuNf6QMHnAqD3XBFbaDUUF41CIro2eyXNR4u+6QwkyzNqqXAj8qIuQkMtbL8KFsUg2OO
VL8/VOJj+K0FfGqICK369aE8TS54uvbSfFkFHyqUVyyyHJLWitnMqUYMnn28JKrdl78nsKlWd9EI
waI2kEynV55U50dBUzamJDKCuGOTZ30xN92lU89rHXqeCKoL02rhF6SG+jyjxeIr/f8d+RvXRYen
6SRNeRg95AcNPqpT7HO35Ph7YuHQrGXuCKgWicSohfrj/9PSFtaDHaGwl+/v7HmF486+wZHzBgdK
FLffVx7CCA8514W1U5T7/f1WrI93bBoVSZlNHusdR4iNJeikFmRzqNWRlNsijPkO/fENv+znUv9A
cM297v2TKpS4vem9ouxRK02gYFkdPXmlSyb9giQc7VEBfhaecKmr6c8QihGtJo3+MnAX0iodjw4I
Pmass//MCYPfvDiBoImOCfVYeVRvTDohveFCjffxTumjBHZKbm90EA9fHuG1JS5ueFsKnR7rHf8P
jPKVQWh7ja48i7AyrrMRQSHrP9ALIKQhKTYqlf+de0YEDK0mGEbi3uAGKmPFiFG5Neas942Vugyz
+MLDrtnZzfnJ9f4YMkx/4+GwBXU4quRdaO3WIENgo3wDA2CyAywgp2X3c/yqIii8OAYPehEb6ttT
hrJMeZmtsknUAm9l/INYJOTrgafP0gmSs1VeZkR7n8hO1jXqOX/fvnwUdxmnaT45tJ8QLEoxKMWK
cn439QM9quc0uOKlOZ+wm567/QgUvsJb7QdOfSlUiPp1qDZ0aaC7xl4y399VTHvDcWsKwn4JZIlN
Uf7tMz2nwNG1q7gPSsaz6vV6xlUzg5hXJ+pEiQOG6QwfhBVW2pdcCqCR9e/vdTXRjmomKvRGYvNr
OsL4wMGuUtSb+oPuZ6JEyyDZZ1JyputOy+NG9HaVDV4h9G840NOkBmBMi0wi9ObmviF3eW5rMCSH
+8EDofA8YkMmXZNBLhTxgEXhGPA0KzJVmeQurVNesOnrQERLTBeXGqu/TS6Z/DU0wWPgZ5zcO9HC
lWbuBo0q8PqoHvLm/DU49OGlbq0m+sPdmsgPltz5pRfK+DmKeXzLSxnJQ+4KwhjjSyRLMLOB6iW6
Wcm4ADDsExmVfvmxL7Uqmf0HMYP+zDX5Hv+RLFkRtDQx8TonJR7Qi62w8t/RqnWLTrAV7ZoNHMgc
f/F4wXvjIhg2jzVkNpz6KQc9rkOtUtfMwZkRKwih7Q1tOVwnJIMTmwBewvU04XZA1OOPffLPZg8L
Waec/zR5yRZm8xuxcvoqjYYJJnQ2DF1rhj9GHFVOwcUvUt3OgGI0NVlbYoWupEreXc1iwjVOyGCG
jUhI334ufK7ggCPQTM52nGPBduwnWMPRWPYNVbqOL8681GUmvswLMXEIVEPI0FkcZveG4pLyQ1Rk
h6vlediQ52kEGvZOrMjU1HQ/ONKd69luAWbe6lgoBjPVcxrmHOZTZR7P7w/td416os2lofC4aCMV
m4e4j8FetWLYoM/5mHvcfijHzSIgEYfzY/ya61l3a8YwZBu5vGjQHni1OefvTp1Vp5fK9eja67Sa
oHwdcHAwAFzHhuMW1J3KZDR/reLO/N6GxAqWdmpvjuNDayF++m8ZVwKRf+KOKBc46tJe3ee/nqHb
eTmXbSrhGkp8KGS+PNqKSxocEEDF4IXvz+pgb7OC8X89yBLvm3inNSgHewC3d++jec50sDa1GjUX
wb5DZQhqyrc5+V8sYm7WS3s/J7e0l+tT2u0WVReD7O06yaBRHBtfPB6hS8GezTLcQPCl68z5JR69
BBioKTnwnBAMPF5/DXHSJsgQWE0sXAQeBcQ6FmYuZ4a+wYzbO9idwCIr2fEx0rs5path+x/N6GE1
oXSXfHBtwpp6oht8khKaYj/UWi/Lr5q+mzfCxpFozyZnEE58ackpM5M93EWd7GYa44y8tw3DR3Zy
p2F857OGEPkLEpP00loxqWFryNoopKlHNAd7zNckbsmO3MZnvB9hJQz1Xs2mAX5WExhcQ/gUpFH/
ZzfFgeO5SMDi+QIjJDHR3P6HDvaUd8MhXzX97gPaX+fPRkn8iKXIJ9zgT8iuqrilQUj/29ZpJ711
iuOhy9zaYOLNVuoWthX1sQMGwKqFSa+Wrp+o5JvJN1ulb0nWhwzcshjHx3hXPY34pg6y867ncRRY
iB2X26hd1WXIzJAcRaqCr0nkq3vRBKT0SB54tk1IUzfRzO9zzo/GpzmaUED8656uycYRSQ5nClgd
BGgxd28rmYCd8GwqyCnw9sWQhGGVo5L+X8Wu6PmoAp+Ho5w2nDCphoQ/A5o9xyT5vR1qUHkae/QQ
oah/9bCSEodkgAS1CyoXpw7prJzl1M34zMJu6qvm3ZQc/zWoYl6YuW0GHfty2tjLXuARh6r2Jglw
QHw8PuI3yugcmzojzZlNMQxwqFXP5E9hbgK+J3Dj8tC0YCJT4C4JG+FoFpdriSxxw3eNcxOpH48C
tqRhxaybiQ5wPSdYr3JAN5jSX0FxtbMgamWJCY4SwK9lMfXrKBI6jPF9XPQBHSj5S+0c9XtqoSxQ
l9cB58/nJbwqwiBl8ZZ2atnT64ZvBuwzfezPYfm5yD/VACiicsROIAj+7lxgj1pt/5x+6KbrAHGs
c8V+X1gdTR/UnXUwvpZGQn577plU2tLsiGGqvGsLT9DQsR5VvJ0z6w3rs3zNY5129GmrsAR5I3eq
raN118UdPYJCt29ewYxx41b0hytiOga0J6Tbu0xEWnjHgOInGWWJ4vdxy08c7ladt5Y5Hae/6kc2
3XNnG5t99GZRTnihKzO+aHq52TJUbktr/jZk1W9gdrCDeXcbQMqw4z0qSGDv3sUKH6/paBaiJ+aA
fVDKjBy/yXEhRntg1sg/fFaBSJ3TmNB0Ql6hm93rwoVcYZIUcxhQx/TA6EM5BI19wKSwE8dY7eVp
uEujtoYXqT09PHKqeQlc3JPM5SdAmJAxOnacKoGywBLl3qfmHF2kLivh3OHMDbrzn1QARZ046dlL
Jq11OOuoONCQijFV0273ZZducSu29Fn1V2FXMMKaK1eZuUnCYkUTbt9Yalm/WihuVyQG68n0Zdzh
qG7nuUAUkz0i25P/bVd01f9fFP9qLBencz2w5uMdHE1NzdnpudkEGg6Vqwo3feCptj4S0FWqb7Nc
EnPaGfdOCayygPrsLVcJxMu6xs3Ripf3rksG55r1Mvzph3DimQWdvOnDXQnGnHkMrbinN+59SQh7
D+ALxXrobaPUHd1TTZc3mBGq2giFIn/KmVykz/qzc9HJHfWjoQ687wjJfmHQlE7fcBGEy6jcw5z1
gB2/NjnaX6nzV5fM78bdPnTK1qHPkYYjbD0C9w6XP6SYHpGlp0usn1Tw5E8vd5AIu+A3cNJ15WWX
2LddZmPNkX4wBfwUhtwUWIqWrn4Pi2eHYEr48JGkojrI1ta7udUVXWOIl4himYkHx6K9LZgySlRx
clU9zWH8/ZoP4W6ixtCoWqScEtMnLNKk5IAVAQ6xxuaqL+nlgIxyw8ZkNh3E/lthyXXRw5oTDq0d
uPhzn+c+j+gzrwNSEmJDlDX3GfHkVY/1BDAKxfjXUlXnQ5KoumsyLHyGNHAwRvLk8FuyOnwzgUS8
295lLQIWetokOWsGzAFcIaREHivC0nS+wOt+etG1i/msTzuZQdir7tdGt0buQKiloGRln4NcA0uu
UPC4hVPMdk9MnKeIqw4qjR0Lt02nJidUqaDpkEVDb84JSMnWtR8zhZmxj53HET9giGVbHLdiu8wu
UzEjinYG7xS/wlPEtx4xwBTmBRW5KngRP5W7K5aOdw5DVAJvd5d/RtxJ7GSeakDt9cZDccUPZrnA
Gu1F9TiUXef9SYr6QGiId2ISPE/NRkYnExHL9KhKY8vQOQ8fojZQ4FVFTCOYpU6AkGvHZlmRnrMQ
xmPAY8qSt77k78M17dx23eP7oes8LVEU19qZP588tQqrMCStRFrMmMNz+MSdQz07SvNMB5+I06iL
BVDe8BR7NI23pQxjEoaMpERpz2ua7ibNP5rXI19hPmtLP8afQJbEQMr9L5piyhQXypW8fWrbJV/2
ZSCW67bSSbw4lRkCX83Jvz8pOl3t0ODvR4baNmjby1FOdJ3c13X3xmTrtaAERkRJKF7sDYwp3seL
Tlmac1EhDafDXTDkGiLilYT52UEcCpwJVA9+nt0vSKUTkZGoYM2iqW1nXTOgY5F/GterKZQGdcQL
A+f+T/ZxEJG4bGZSkkz7JZ3pkEzmX1Rw4b2yaouEPH37ndxxbNjKK+Dx5omQkk2rSBuwGu+FQIvE
o8WCB3SfscRwVX3ShDxCDaBh2J2Dd9PrJKf2TXsVqswA1MX/7MXTws5QHIJ4HREyZ5CYHc6QLMIm
GFA23ir+bU0oTFTekNz8zt86PYZni3+eEabjNmcxvGtdRmjZ70wplzqJ+SeV6AXWQhtvYiESLeU3
60i8Zc8JddCSX8W0oPKWIpUyLpCA2H3etmJSbr110dsts4+epvzatTIyoAzo0Dtv7E6+NOZe8JWg
d42EvOzviZz0k12V7sIC6Aan5AaezfVKjNToaVG2s/NuXTyXBBIEyg6d9dR/2k9GodwZsFXlDp5k
HXFO9yTYrobE3q9gWRwzP8tnwWOGOROUJL1/zQmW/tGW+d0LFeliwXq5xRrfKq7/B9j1xeDqTCrd
vwlxw6lupJe85Q1n7i4a/sh091Uyt/LXjw08SwRqKruro57fTnyRtfL5K1i5NqM4+taBz3Kf8LIm
jy5HY0ga+iqfnrKf29yKdncDmswK3CIqwt2+nfk8OBTw2bEAF+4aLjhtc2Ho+/zLV2CU6w5KTTGG
HHp3EMzHlj3sZd5tyi/3709cUtXCuE7WG52Yo2hDiHcNMcnGx3tkz+yxOZEgBNBgk5qg4CNcKxLp
Cq4lJAnZfMeyjx/phY+ki3mSltAsgHIjMMfBgCOgZr3ZySMv/xgW1HAewqpl4XGrFUo8wCC0qFk6
o3xsEoAcX62K4j1l0s+DNT64dd1TxeTpyx+vGdh3+v0n8C4kB9zRrKBE/emq4/93xIiqL6kWoTOW
Y12hLCaPxPwLf5jLmu1PgNXH4kuh7p+7Vxhgc86fEuxLlfNmBgbJqLJDV0bkWkRe0oEZxwzHz0Zr
OOywaXkfSZbdhnKJnog5Qg/XxepL81T46orATpH84s5OPMoqDtlV1Jzg+jA0a/Y//ZZ1X0XPGlUC
cg+/1ip1o0TAXxEE/C4MyEJ2iUM6CuVh+HdGuUhoN+0ypVrkghkwdMThPLLNYQrEY1o/prCrpyzJ
W/1GE5T7pJZWrmcHc/ry1Va83op54bEoQ/MxdH8g/A2xuiacfB9ex6JVJCYDu91vBjBSBGN3Es18
s+Z1sDoikVn7514rkrpSLSQVPmA5CbJEESF1TiJ229YVDcETgBaW1Yb5S5XWfHFXf10G3GOK4dro
5QQUnfTseG2C/iMkAzJPu8ZnCBsS/CbLRoMNcAWm6DnKuJeIG5gyZ1s5h2N5GHSCbv/rZDjYHCH9
DCqFf4FBc1ojYiDkg3J8A7s/zyVDyTx1lZzOjE5acPJ7bE8cNs7Ey3cblB1bqXeOR5Yzrqt/Wav3
Gc4Kkw7Bc2iXvUcQTDN/tNY7hsaeTYK4gaoZ8KQCh50oc60hGuu2seRcX46pA92Myl+T/tz9iYug
f/9NUEmoqa5taRcvkmnZTB6IQucex9Xo526erPfst22p5ASJUwL/xkBB9907iuCSU7Io1RgEFDfD
DVVUHyimDzVZcyZyH4nEPIu+efyIneVLBRcemu2mnfJzuIAvg1GV6xVI0Uo/U+WnN/I4nUtpRB2V
bpoJRVqU2n3QJrPNY9IB3hFdj+tqAKn6QM//1x0YAsMQapxch8SgCdVX/PBfN2SUi5IzOBb6FkBa
flyJgY896Xe2RbvvC7ExiWBNNXRHGBUa6vFTUwffX9Ak+/l3y/Bdzkfbas6lWLbXVSStwnhveM/J
ExdHCauJx1rarnskzkg6EicQtvRU7o6ISXilxh0JicZVgVu1yoig8ESrDJsgfNIOa7EZdu8xp1MF
ZZN0LFJWSBPhfQSSGNbpmJh2Ama+ilvmz5I14ifij6Dnb4WjgcF28EHXx7IIHgyasGQBsGFGI8sw
GNqb6Lezm2Luqguoaxs1DFDKMVixII9E8ZhoS1cJy+UbcLN5kCk/I47ptT/0qlM3tJhj0Bhc8fd1
6TCUiJD4blAQEVIKBh5r0wQDOb7H78QQnkJWMjtFPjaFiItaNQI4NJvLueHo4rGypgVz5uafXUZP
E4aBpoDj85krUSbU27s8Jnktt5UQfX3Mq3W0wH4cWUql8MhpywMFeYbMKVsGRszXLm5v9gTjqpwC
i4/cHtYfI5u/ciM9DuMi/Su8wNb4uEBu/2eUEZuPZf0eAZazqiBg+o6h2e/65o9QgPwRNzYMU7X0
puGXXTVSrFn5N8ZO0s51Pc/jgJVawXXPURH7lgPuGaX01sohAPl9Ku0PLFHX4wDdqg/lk1Yp3kEY
Y5JvM+NhumDpShsw8NP+uCOQPFn5EqH3uYWqunIjc5BXuWvFsl/eoq1Cbgic1208Xa6qeWeTwmbD
kM0sXLNMV9YNUDW9snJfP45cgUO1XZujgIV4bTwaSe3SXRUWORrGomz470f6uBrO8OECXh9yo3gF
wmh+99XXQLlBonCmlu44CRRdWHixOuKP5CEmre+FpPJiOXZOhY+EmtxQUiHcnxfHOAK8ci+0WVUZ
y/+UMnQ/JfFx7u1eifYEDz9Eu9BUIop6c6DtGQsmlgxUDFJSjKzPs58k4RznJ9plhu2mg8HNWJc4
vumstLAkZ8Tr2mDK52qVBxH2KmWG7iGPJKiPq1TFhGfEOBhZPbaTyLwr41gS8Mv2x1gLLhE0vqSE
S5UeWaElarT1Xso6K+FN15VnfilyOoi1LFgONlKwJo3+3vpmSxTT3b7xz+3aCV7iSRGvafRzOJAR
9oktLedINjYzqZhzDTwvSSft9cxrpca5IlV/Yi7QXS9yl6V/dx8Kv54iXNaH6t9THLia1gs18jXn
wR1NjNIsJGKRfcIwkK1Ftfnm4mxzxMk7ETI9cqqKbN+Kyr6uiTokNGtnaqf6r012VVUb6iH7g2pm
jxjlJSIRnE/m1zw7sCvtm7y5tzbjBPRBd5zVpLqPA0D1fO7VTQRBN25odxcSWGOlmpMcIPWgFG5K
zvBIxtGt5Ko46PwaJfhGJ3kmtQtJWlsHQUWEPpZEuGYuyKU5uE7MIpU2KU7Hb8eQqlVGL69hWy/i
IWDTXixUZq1+vxdfNuhYJKiPP5cXwGOgAGppleC4qI2Oe42u2OWpU9NjyLsBxH7vweIdd6SbmgQ4
WD08h4em+hmW1tZunJda8lWH2aluCarsAYeRhSjmgHWMsNm6hFwF16EY8AIoBTtg71FXmRea0Tfv
6+NsIEQu0TC6sNeDjA4qyo66NV6ng7dyX2iNflGM78ZIkWqtI9WiCvklTqD+jqDGFbGYvGmY6UV+
HLvT6F+obCAuBkkuh9DBE/BxVhVYPLNZu3t3lSehsOrkU9VDN+gE+J5F+wY23wXciDtgO6OzmLXH
QFNQ8cE5/fHW7zUJl5eHa1hZ/wLizPT0eDgvr24Gx2o5Bkcovqv7CajJDT14XalMN0hu3d3QQ/5/
8WEndWtru6Jw+Vd0yk3IKTfUD06rlzHSySrzzHkoRmSuW/87YPBEokqVHY5Dc+jaoQS7qJfyGhZC
wbmmvrHqx2rGSd2zMou9dVwtlIs0Z/yZMmtNTBreg2RUWeY23VLivxQTlyg/A/om7X2e1CHR0O1+
u+segQu2Nyhw/gSZfcbMw5xRexI9kJIu4pVAWg1/itV3slkSL+eOFq7fgW8QcNKgi9fvo/oLpK/N
/gsuMfH+ewoIZb9W4b2tiAqV5L9PPiCWo5X5lcO19hOqm9J+6Ndo9rKBcTRrnqcuwvngMEX61J/4
LDUovCPNrD34AKJjvdpYDCEZ3IU6pbjnSu8k0HlrzAIuNDKW2slg8YzjkJDmzsHClTmwVjOVtGRm
UMgkAqDeGbjt0GY+C0qXi3RzoO24eS5UpW3dVl4Q8rcGY/eH0E7535yi9/owK1aig46F8K4SrPrn
b6xTKjN95BbZlrtwc2Iqi/8DyS1PgqeEDP8IohvQeqzw3L/siI3Ct9Mn6aHUbtuBpVPWb66XSXhv
dcsNs8L53ArLP+NanH+B+BS/0v+WmdGqzuhSzQAWOrMkiIesP8mxASvg4ii2Eee1vDtOjMqdc608
Hw9f5IyxfhQN6toPpYtTQKpXtj6bZdEnzAMXQ1KWU+jco1+oSskYoq+ES6xwdYR7X9tEC1zx5Apa
4h6gDVqJPr56na7kkuw3TL70jOE6EszHgmaU0LvvPbQdXg6QccNbTnHtB5uGU18zEG0bghULHG0a
QN2++caycMn0jFJsGB+pi/CAmPKyAQx/74kEX+sTyF03PWUdl1yYp+c2X/393LlYnYfAqIrR8pQ+
0hKng6HIfGoEAfyLeGrdRwZ40xv4T1+RiF6YXbdqbysfMnVPHOaSXfAqAgLYenAjk8pt528YFW8u
EMq+YUoI33CzR6RXspuQR5XC7tz83IURkg4wdQO9Pi09P6zCqktKMUPPRou38MR1hAwlAgIRsAGu
HrnTQZ7wSINqLcCKqLjl33NphmIdRKbMhoexLAsow/1iv3UTZb83MLUMWYs5oI2EF54qEabnjKUM
FPfGAhpnPDsDbZc+0m3HNKravGk3hLP/299xPvorxaQaJTTePrF8QAiZAIBKQwcOlt1XZ+j0hKDa
yXUQ6+BfWK0TeCYT4lNVc5lsQFxsXr480OWBJXh9V55ymldEcex4NVmnO6GOV2J2TkzoNEMMLS5V
J9THWVXBlPIGwgD6cCwpSpO3SCNqnPymF4Y7I1Mw1LWm1EozvRMPzXMLxUyeud/ymOscL3YguWSU
IWGP3Ng7OwooIQgTMSHCODcN+1i9sOVoFVHVKBMR7WeiCP8MReStudYp7jBXqjA/+1Ax262r/q6k
WM+/Jpn3OStQgtJTTu43beDvRX4D7ad7PgvQQcMsWn4w+Csyw9YF1e2cOgUh0iPg2pHHTeD/QzDM
uKxmsx4cEWT2doaPELcn7UDV9+NlcvBNCWDNWiZFd4U6gSVrS/23QbAVh5ORs0YYBe1pG4mMG+oL
q/u1zWd+yfvppeYnIxwAfkC1u+Cl/gV0T+jlFHTXCSmWbhNl+6u28rkELW9CclJA2kLr4HsO0sYO
gG3jogRtqram9o7GF/wa6WPNG7PF10Y9xywnVpMNFbYYtoUOXhVBxRXXkY91TzHEL2I8oyMoBvxP
DRqLegI3Z36khSQVw71nAacR3jdCX0t26gphyNGaSDrTwQ9yjK0EMTM8fXLFOwgyi4Q7EPEExQBr
QkgXmvhYJla3MisolQm0ep+WvexpqXKnA2X5BDezrn+W0jXAyn5sDxzRgaGoQTdnTFT60w+/RFYy
unHtmzayTyjE7iIbkUbfTLPYkbMAjJtHt1xlO39zJ2WPJQQ1bSBmddxMf2hkaBVJwEay8hQ4v/jk
ikv3TDe6WV5g+zGoqYRNNHR6dAT3V46JjSW+ct1szqQWV8Ps2JrUcIvonkpfuuhHvfKaubNO9AF6
xaB/ydf2kYSmdA2MGeAKOsbRASOa443wm9eWFmu3nYwPNE46tLT3NBZ5t1zz33to+lgTglB66kVZ
sT9eZVasEFtcMil2bcFxdxsllymXe+Xe1cc1/jrIP1uSK844lPJKgXGX+1u0trEsOIHBddWKYlvl
j7LvBzVnVlwL0RmSXm2Of/FWqqvojS0SYB8JcKYsjZYt/gN36eLyRutaz6Ky3XFFNINbY/8aMll8
A5zRml+dcUjIuQrHBVuFyh8Cde1P6QHKk/oYxTBwxih5XaWL7ZoziSZa3pIqQJVkmMMSqKOR11ag
FsSn0eRSWTq5dElLdntGRACsXHExOv9vgRdpJ5Ul7tMLeNUdRwxu8eE17bhwEQJy2r6gKU8JpQ9V
PdMTZUuRfTxbyIBDwtFA3irNO0K4W8zcDoLDEAl5EvPPCITKpB0hcQ6wLnlKtoaW4x/Q99857YWJ
Hs9+UoLrBTVBrvNekSlwgXL2PPlJZRKxaKJb5pZso6Ue+lLUwcJxvoy3Hp/y9dbwgp1d99W1w3mA
YRFcEIePdzzR6D8lkZxw9vpY7THCqzVIpgxr29hmHCqnCCg/Z8D1T+s8X8cuuHpg1joEo+sxvgX2
ss37LnUEAYd9n5WvAoBuAz4JspPeozISwNsCKGGjVWXQ2RP6brBmouzm0ruJCub9cLKvhg92k76v
QeAYwu9dgRmiT6I65Y/L6uptt0gS+TYYIbICfK96vuIOp7g4aiaVKorQKh+QrzSbcgaMd3f1LE/6
EK2Gz6sWe8/chKc7ZhLjBZ3cprWvKtR+KyDc4xgJyfr61ZuW2snYMHz2iw/8z7IqawI+oe+EZ4O9
0oySkw8XwQVw2gy59ZveR29Wvd2qp0MoK81MJqZCXkuZ5MsD25nc9gJq4+70akFELlvGuCF3zjls
uLRYXbPW25vKBJp7ayJEPJqEat463X8IGbWCrJ/wOJkfQw5/mlEl+KwODAMf7x2f5CxY9cK8f9MD
pnjVjAaWPOSb9sIefiRVyQ2aiXZ+c3QdBDSqcwP6ts2WUyULjSEO3Ju8lAb8KOQ/LRvqBw8fnHY3
X2QWpRf2Anfi8ERoDo1Lyk8x9971M//dMYRIgMuMUFhb5FXLuz4psTLrPGpFhJy+/94z3koHHi4C
SkdUY/0jeI9mGiOmcstKrehYXubo7ZXAGmLHuTxN2lFGEFqRtNJXFbyuv/Dsu+5WMx18AdwanQXB
f8MaYy3Ae91o36kppDMeZA2/1u4rpUHQcqe31CIDZERl92fuhOJyf+3nOSh84eIImHAZcaR4w2Fn
g+dOgYQzf492+PokeAAlCmpjvSXXFKmwtyN6l3aEvUWjvj48Wdo93s2aKAO8CO9gv2emK9N4aQFF
n3RndpfWJiowfTKaX2FiZuFpCrbtW/TMjoB4GOeYCK6GWsj/jIvQqJI/iULZNp/F3VNSH0/PqPqk
VuQ/GxYECkS7KcDfHyGJpMy7TuiXlG+Darv5OAIKCOMVhY7FO4axlfKrHDQEQvzJyPhhgbC+oDMs
8uC7QVkAdsyP11iahzmH4NQUFeMPQdBC7naH5QIHAJodc/h0yE0i3Qhv7D+2QdwA0r0PODZr2/Jc
h0cicGQDUORrnNlT9gMDo9LnkoyLURahG4Ah0gAoLrSLmlZdoUKDZl4N3GVLJkc3KcD6ybyHLWz0
fh2pbGjfEtpaQBvd984Tgh66zKzzCVBBfp3oLizpGlPvS7g9FBPysGszLdxt6oq82YfBKxkgVyEl
ntH/44vmBoqzHLrTH9MArgtUkBUJFzynzArFeDThXpVX/7xrQohRX/jGQcf5xiVwKD9SNnHkJMUc
w6U7dEg724WbEl9uATetVYLmBS1qOzBZ6Tp7AfaXrYOFL6QOY9OnNHJXq1y063fcb9gl5LVCxb8X
mfoMIe198i5chmZE5h7su6nz77PgHFqRzwRbRqGXp5KBw4cuNz+hdlcRQ6xQBtJHNIkRpwcFt4Lx
qEF9ajObrbU5HNrK9GZF2jDLzlm9JoeLbcTVw6U5y15g4jT+b8RT/FSXICSkDhEeBPeFCFUBCOEc
cnwjWKK695tT0ebP5jyfnwkn6MA07v7ePumPA9mSL5RwqO31doYB937ncnXBXL1zDTABMZ3P8VKD
eXHcPwaW3hZqgATjEkJg4jerDbaNYWnKo5El8kyV4yUDFWkr3+/0y2jDm6c+h4O2jIyTeo7hOfnH
EPZZsmZHdanPLqBjpRa3oQQ6+NvlxvnMPx0tsiLvq1Ju4E01N54Q910Jd+6fejyKfNtRUtH2UDuw
G3GysPlH8ebNA7Jh0/MgwuINmDFVX+59NFEiPfklhN/gkWhXn2OA8r/Uro6dMYPXWmRxcDwErq4i
nFsd9N6EBiIWps+LXLO3qGVmHtcv9Kir1m9FI0EmFDKCAzTjTIGi9wohP+BzE3CH+7VCLvucZ6lX
BEYMI2YlVz29bbV2xLukhYAlDJzyTIaY27eo5N55/6LwCeErBl8k4i/Rhzt0n59IV5bv68SFoaoJ
A8gblRtS83AiLHPNnH2E6qND7jt4X2fTxS1vKGuJ1MpeB/TdfthyTO6GtdXgnPu2yoccKGSVYY5J
6cnAhngpUut7bj7gfA+Q8Hhnq8O6P7GXR9HAma7yz9u2mSj64ZU2589fOu285HEBaq/MSB6o3ed5
1JGDhTOxvDxR0G/lYA6t1MoWf3df16Fabi5N3AZ902jZnJvYopYYPXTgMbHH3/nB+Q1Tb+90fwTz
1Pn2mJir4nQLez5smsFd8nwbiInIp+jHaIRX/qmG/h0Q3kvpHDiS28qIT9jrqkRiqMgWUw23bQ/5
iIBDeknSObsLH5clID7CruyklBsX6OtYxptv4QBlxxoM7UhacFi8Rtb8ocgbZmR8AXdDc5O1ABjC
5cWIsgkVbodnxJXVvg2AbNYX2vsSzm2iT+am2kpsbmADLnx26byfAcqwt92hgGa4sG0sp7IUTcWm
djSgww6YNxQjimxc5/z3CSRyYCyeHrqwRBoNL225bLJBu/UD+sZlJZWTv4tvFhfBSmJ4Nghx+Ltr
fjBzT1VVXWnUi/UwMkXIJAarTLs5e79yyaD+ss8w1q4nVsEYi9wsG8ywW1Dth4d2Opj+JuJLVUV/
76CTYr8zrXWjLazqh4Qe4zwc4gr08o0BDbv3P5RARVn/DD1cBhS91/mBx5tv9TGHj2l5OUOJpjoV
dX7yYO5kOb5TIO4MGIePfGhHYbRyF+RbxZi41akKOnLy3UVbF0zghJt/Gg8r2ahceeVolN+qvhjH
s64nOpxJrMPxT/Ol6P9eXh7NPLmlGOx2mJm/2U6IuCyC34koz7l1rMxZiPUEYw2MaBT3OeP0t7pt
MlUZ+9CXRmEH4zhkjS+L8+oX9BJIcrBCBktK16r64xW1lEXf1Y9lNVf58Qtv8E9T5nUIrXbb+s5r
WhvmFLQqUQUoafoKxzOK73f9HTo5brvvo7ZyaJyyZOe8xen2sbBB7pVCsu2D89DUY2U/iKIiUpca
QMhOjAZC44fC2PglmNxFRrGBIxzqhF8VfhAzSsfAip4WRx/fg3NfDUcPiKekK/OQp3kGTwmkH92h
XrUeszCzZVqrphfsxIzbMLpaTgKSnwrXzl/4tGGWt7oEjcDR3Mbhta/gaTKdPJsNeFWedWD1cXtC
iAdwGgKavIGOC7izZ85KrFiqi08NMnvGkdlmr+1RnIFzRxK7Zu08U6jHNRPBfxTuIjLkauMQJg1x
I0fKJQURUZALy9TyLrI+bpH/duxEe3YXs//Umqty6DkM1KkWr+Ebc6fxg3xSKndmPoNmR6RvZAOg
nC3QEItKUDVKTLZ2jnXF9aeHgj2Vc25KM8Ga2JF4eZTxcS1e/MtxmrRh5DCg7D5Dh/9AL/oeB6DQ
FO8LJuqhUtJ3FPvOB/mPqpYKn8j0WCkM1FFZm3yBvHm9Vuq6IsZ+sOHlTWTndPS0tugLFd2d10fS
VbM0gpGl5CQe2+tHF66EwbRbKNJfBJIs+wCDyOhKATcrIyMpQdp4QcjL6g99LlisvC19xJHVDi/t
gtEK4mFfyYD2VkIPkwIRP4NiEGCD24Nqbmt8q9BDazMmo94h14JhxhylFMDiIzXayPElWYObQnOj
ZFnEVEewktdalhoTWfMEUT5NElqSGG0aUy/fyhWPkcdWKg4+o4clr2CIgayvUnJ5Ho+a2N1fqcQR
8E0/Xp53NAp78+rWxwXlGUy71CK+KURutgpCtrH+C915JkBVyhJhX49GckfMrs9gA6hqkIbyk5Wa
j9K+UwvgujUkzYk6jRvBoa1Mm18GEcJVKbqlIKIF7Y5luuP4x5cc/77xIUq8/lo8jjCPcGpDVzrk
ySIMRQ4kWBJl/Y55sy6JUYO46J1NNIIkIfcCQNCgEw8RwSmLFX17aqVqbfO0JGIX27mPBJcLy7WU
GFI1VjmSyntHFHexeWguFYFZr60XFaB4pES9gQ86IuLFWmqfvOqfm0V9FbZoHGkeT3XzKIfAOrKf
M2mMOV7rycLhY7ioDIolxPUVKWk2we6NeNrxxf8hYvI1PeqISnE7I34e1MKmJ1M4Saqgf6oeOZ6e
RzO2BRKFc/nU3F8x2trrV3AzYpC1dID6pWlWCZd9DFkmGzmSn964vxwgsjlFtBHAstkFiZWTd3ZV
NFmVjtCgZLFDonfiMUu+HMnPg5c7l7E4iVzEoAUxoSFXLjkFud4r4Jn5koe0kBtiE1TppvyIXkE/
F+pTYA/IqEeky5M9u+CBZK7mmSj27PzhOpBIUXPFV+02CJRuoLP9lgnCZ3I1rOqR9FhgiiDZF04T
hoz6cNmz4odfAVg7FYLaDiv3L2m/dI35mOQMsWXyMyRP+BATOGRmt1kiI6WLNzTGu6Bl8HwF6MHH
0oXfWXuo5shAdqjBOV9cDfryrk/qu3w60IXGATbd0yPgMyeZfwts8rIANr9sIQJbJUARYopSOSYW
lN3P+w0EKDiqMxMJfQ3QVtDyqXpOJM6e+QuSceU+9wEq517rjLLT1DPAsAclwRqai8gEH6KVejti
HB8T8Q4PQhM9wKRZr4pPDGRqsza7mIa3idhSE/Wb6MAUzFqOJjzOFUMoMp749JCh7v2SawhQbbOd
+1wYJs2mC5TAWYzv/5da7snxnlMyR4Hyljhe3GiCOiO1noQvWcXRHNUBRx5O5sNhWFnnWkqg9geR
EbPCAGsWvpfozFHiMsdUHIyPKZnhFVTXR68i1PbpbF0iTq2mmjQINJPk+MR3HpXByXUGB9SMPiXv
uWke+3k4XmRkyQb0wmtlSy4oDuW4UdJi2wWB9HfEUJO2AUABHHCMo3UALC5DubHQkMjyPrrZan3E
MPdGv7LucQ/yUNRL37Mm+paV8zG1+A9Z3E4vtzqRov6Jjdg1QNZrdYdfPQUaBwiN+9tkYnrWNOJU
HLx0dqRDWtEADOUfgf6IrZtSv2MsocEgQC9yqPGG21ZITyJulmBN039tjNQwWGdpZKP++0LePiH4
j3QQxm9P6YhWKLwHDe7w9P01EwTRPiW7QWPXINxi8zh3wBJ1E4Q8nbRdNAPy4XilW20PuAa3qetS
l9Ae8XIxDH952EIc54q5ARBDJ1Aye33Ygl7voWGgeIZR7kjJHpYTB+TcbJhltn6l5ENILK+cG6t8
CT+/HBsNQpJbgWnrBm3+OqKcp3pbIIrocVwrxf2hUVA0x9PMBjU1uDSqcYJozYvxymwJqLCPNjGu
9gYIvMkTVweCFmYYm2OuvIxEd0bA+L026nyq8ywgkNv49C3XqkjM4Lto6GUeDBNNB6EwmRVhaCM5
nc/k7eT60WJC7Tw/yNXWDXu0zpis72MPrv7pEkuFOIiMb+uDVFA/YYShtodpaqJNlMJuojphE9z0
Gvy6kbV1573C4C9TivBQg2pGjfyp2njd1BZwLw6KSsaSHB5mo6Om1tt+ZmB/5Lc+9zck7O5+IIMf
KzwurLn9P0Q3CjJiI2+u79APDoFhAaXKKMrJZ1j+Q7bDeGgHplLX8zrSHqK1byAPvqZwQSVkC4Ja
6TqTpcpJNEadajByZWwDgi+5kQ/9gW7i8drNnYRHpqKNs2O1lKiBaoMGjdUs5FHTyAamjKItRHKE
duvUlJPN3VqHvpVhx+tl45iNaq8WtIUeu+Gpt7H7GHHiDFfC52sQ5H6ielrNdS7Jj/hI6l3OmvxJ
gjbdxGDCAW2sKGc4Fw+V5m17bTPVxFv1E12ljK1kEaJvKhLjUWHSqb0t59ERiu/0nWiD3fpop0hJ
C2lO/QATc3Sgyj7UqB+SWaO3jiIR+j6VIf6sSYyY2YkIxGPlncvFfbwEgwNAeevIRu3pQHoBrce+
GpoY6WEP5EkS26vdft51mdbIPdCRvkjb74F/3H8pGyWHsBgPe7rxFXT+7P67lMnF/iwvUVKhy4KV
up+56y2i6DAb+Hiw+8xOGeVk7xnem1jLljLuMPf9f3vXDq5xjdyo4VeOPNCH5MOMYeM2c038La1Z
9/ua5F2NhSns7YkPgFRC7DIQGX9flbzb5cWKFhVsS2md+cVlGNT+vuRUXSDtFmBeBYQTBPh2maB+
DtQrVMVLFu0dMJx20dvLw7NgtK7S1QHMCpVn6sUQwhyT3IBwo9MsdNVOju09XeR71rYQKBEIKcIq
NJvsu0rjkGK6uhmwsP5el8l71VmmeHOpu9kqQofCQtWEdrtWSzbbnJPyuETpesyjtod1cNJnBuUr
YXArVzCUTwP0ctZQiuERsagwAxbtkvkOAfX8JPys4Jj26PbtIcWK/7SYsFwOUQXhI19cqDOSFxLC
Asi27C5gr/YOHsvHK6fOJJI/fuEfHfDGB5ZvQTx3xE7Ib+bKwbWetThj1EywKHxSiIc/y9CSEoRI
EptQwsbAgvCtjdnrLhvD0o4ykNGYV9xYKGiAR77EDJqTMldyMLwcZddQsIRws400UEJcPIAXlVTY
PR9HTWtkgQE09PZ7mOkTE9fnZ6y2Mb4EcK8oI068V5kRbBLn9gOHLCnodPjzM9ohbXWcoP8kdUU9
LCjUHMK4Db0OI1JwJ7hRoVzNdecYWrgu66a9EQZ3v+Zrh5BpYo5FSVuVyGrcSczEDO0ySR8Ti8lB
yL/M7MFBoNcCJrshXcRDpuSpXVPK5/Xk0TLsgAp6D2P6872YmXK8WYL8p9q+co2Qrbbn3hNXCRJN
IkOdbf4FcvOer24612UwdIimivoubVY7meO+QDUhqy9/iQyqWdgEf4Bzr2hWXEhA7srzne+/+3ba
tbH4TAl3f76Gvy7mB+W8/bCH3vs+Vau9mdpkk76d71+Q6iL6aIgDhxi9tDnRFJAnDTOb+uN4pN8j
GIXFQgl6R5tzftnCt8PjNt4a3q8QnHSOP8pRefKo55lxnxJkftBXkJHgz3tEWYuBmOuGfirsJbo6
P1Pp09oddEbPxzItabrAO16yx26+rqFnYFKOmpMFTvprN81k8Wbemw+w752URulDgHRmT7yvjrE8
1zqBXrtzkma7r1sLZ6QcrOcMjkfqUOmpeex4S3mOUdV8ELyrpiAURD+iKK4iJJKcYvh1bOlUogGn
lGfy2maM+D7llrp1zuU0dOhMMR184QlbY/FEJtb0ky/siYorB/4W58CCVHKZdeCtJtlZWXasglPe
fhGYFBHNHlArrcM80uUt7GpsMjmV78Rb0Jyrg08BHmp2lrAPM5VHck6vtgimfjT4cSnD42mgpXV6
jOsNWzvyalqKXOog2nBNxZTd8xtpPYYcKRblh3Z/RCDPqajRiXy78dOVkI3N6+rtBUbVTvA78KGC
NiEkaT1KKIYN2dFi1GGzAd2RB+HArDCrJ7MLk5S3sP5cD1jdG6ey63NHcHB8cwXGJvaA4qZMHlMF
hMHZ8AnMoVH6oaJvIj9bl4luW4oQZL63Rhtux55+i6P9zsS7p288xtUbBzD1QR5sRnE8o137ZSoA
uEUzA2N7UfYDqfm66R9JORNVEsE0Jk4BgCfN76lo1lggwaH6U+XCOPagY09pDYU/Me6LZKjbIs9C
g7vkVjn3JZ9cSf4sbpQBYdpKLiq58UwCWetU9KM5648GnLJYYEUYjWxsIkMo3lzb6fq09a62Tnwf
rZc1OFBOL6nJQF5VfG55cMvcaAFwODIb1m2WQHge26ezf/t5AA1tTKN7oztSSI3/QvfYd7puznZ6
ecenKH2qE0EPwEYenZxd7wLY67NoGlN7lLyZB1VP9rfdkIJGYolvaGPs9m00OVuGm4L24eE+q9vl
rBZ8nX5Sg0M8Dbre55KIGCVvu5r4mvGkG0lhQMTP6yG0/jpyoVGiomDiG/Ca8BhKz/YIqTFO2B5I
/iAzImOOKaDYEch1wRyfGZoU3+YscCcojIEyqZlIA1GTnu+URj5ez3YjiM1Aoa0NCtsc6kO7+MzP
LlR3PiJkIKRD086mrwdlwTuctxbxtdejer/NXLlUycQkqj4dVrSy/veFBpMmyvMfOeaFq5HWuUHh
PDpq7TLzGfgEQ9vtoN6uYMWBnpr4+JmwjFpTNgVRs8S90LgGLHh9iB9zBuNfPH8qV8mJxS4Euh0l
8Y9bUMTPrYKsliyS/4AjZnoOHN9JFiyhcZ4vksLPZBOEa8nir5PmCR8Gk+ugQqsRWi3CbG6Bjej5
KpGib/OQ21mwWG8ZEN4qjQdesTU4lQ/cKOSQFA83cZ7H6BOb+cEWYNwAgPPO7uH32gsowO6xgVFq
TUuYjx03/j5QojBcYFfGAMUDqc4RH8UWI3OZVjLA3z+ZPrmid6V04Wm163JQtYot8hq0CS9ShdSM
e8sYgHPrkEbsqswF+sucm2uJg37FlQhow5bS9o9cyNNXBWzpDT8bbZe9LL2fUaAVBx3R8wBQdBY+
/+p4RB3sIV3+A1bzhT+IuMYO/lTuuTDWZfM9hVwlldwdBzkGMUyA/AOMQZbrJ33D9BQGLEw6vGww
V7Tw90zIxpYGrwGemFUfKTB0cUOOH4n4Tk/GJaTy3syNIXQQVtZjRx2mA21AeuYEF1irmmNd7lwV
w5uP3yxAtf1GVnIxJ6Xpp3fgS4zyE40eKvB6TGLncl5t49ZDOXAOG68P5BAkyTCykVigjTmTKv4q
nc4ZZOxR813SlmHan5ialM5gRlCR/WMz783rkO8P3tjk5ArfguJfBsHFnVsT4ZW4Vn5qt6TZevg3
wBp/kwpbC0waAHqc7H+7fOoU+g0E9Py2UqikhCV6Ns31KwNGEIZouaUUevbS1Q3OaJouU3BUCbnG
WK86Uft7BKlZWDWK2X1Zdz/vn3vCWt7O3IjkYw7SWdxRHRA55xWqNOaC8EVQuj0RycZlZdYbjUJ3
UrqW3HKs3ChP6InHgNnfUg8hblGNpGmGR6/qrF/6LTb4Zb8YmcmcWJhrGaYQ4rY5eQfIEBmdXpiT
R9pAjFDlSeHdr8biF91d/fZjJR4KdQqj0UaUzWPYybLlFFR4jf02YUHpyIzOA/3zsEr6Go85IdYo
OEulPR4/Qa065rKdFHnIh/nwks6+HHcKROVusHyUttXdNI6RPAYuWre3EQPNzNpospTeCCR5dmXu
0SteTT6v64hmEzlv/LIe6rNvBmxdBvToglyIRM55wW5mBj654Cj0j/LSzWut46/AM7s50BPMjRmX
y44ONeCsSz+mXFMjNRmCg6kONZoUJmQKKypHEWrsMJ1VZ530YzQBp5dmJcjGU8JYZ8AhWCWpP0k7
hzicq5wlMlx7x0EIR7HDazmGaWumTmCSr0DOFvz0uoKVwjVGyzplMYl2pu9dc4BPvdfTtviXa3Vh
MsMzCSOW+eWcoWlazpaI9L9s+FY/iQKOBwQL+90jh/IBK7wY0QA3daubnJRoNXVDPylPKYvMpP/P
u+55Nm33GYuD9nW+tj2bsXg9gErljKWi/bdROSmzY1JmtpWLmndQ/9eY5dDNvq86NrJ1Dq0vEltB
RM2NrtUjL+/CN6GZTC/V3GBXwLA1XDvkm64JAVX4bGgXcF4B+w2Gt5HKwT852q5QNwaIKiX9wz/V
uiJrAxSpR5X/jBa0RGH8Ecbu0h1bcJ41gz9cOO+HU/jH0MGPDqnLNEZ2XDmUG1qEc1GUBtUKHlqh
YZSjDMTIoFBkmh9yqUcbImtJ1lN31YkGmId+iwLhM2JaKvvlVKIpSXmGTtkzlHEtdiXC4K26B8/t
0X50VmJoO9gKpGXDLV1q5bnP8CB1w3xRSXD9Z3xMfoTqCyQzoAc8gBvC3aF7t0cYwoy3A01iP/dm
S1sIhqQk+ueRiyuqaeY/3r/bAbKhEyJvl/v/czCFl8rwrWc1dvUMUV1EOVDCdiLyiNxIC/wdLXi7
PZhRXh6iJiTs+FtBcitceYJHOG9AscZRPr6CG1QGxEA8uCJLG6k2v7Gw5tl6iAALeVslaqgbRmzG
6Hg+npy/gUSeyhFi6VIuyrmLS5dc5p3adeRq6hKgh7S+fgaVQvHGLw45aMmN5lczAZqWQLznaSmr
dZHeeyZdo7zDzS8IW6lAGcZC1LPp9QpPDv1tBk+XYoawI+BK9a/76wqmzsYchtxlkGnegexafPKZ
I6NOuHXJuAN14+p8uHXz0KJ14gtSRnLZn+0lUEZxLipVrn2Y6POO84o62fSmbQDhlPP8tOp8NhHA
JwCuTsj6mIbcm5H5eOI6FRoyEoEK9tptl1AvKvqHh58eyLE23LTNVaBFNyxGfjea2+ukqDVW9nx0
gBeC43F6wDuyv2jHDgD+2HOJkmoQUC4Xcj5Xmx7bMH7x7Qb0i6/NCtASFSkPxK7Ubs5DmsmWjQP/
kkgm+pc/0UgwOCYvtmFUFZea+51n+ZcVFot71Ri0ia+DxfWqcPnO58FLrfYYsW2H4H7bGq8eMzoF
7Bs24u6hAvZfAH00yScM5E4asA6mJmcVB5mVZaCtbUAh2B73ZbwZvpGMYLYDSBtgDTfpclKr9Bi6
JyAaGIgfI7Sh9kWTWMn6oLLMgotwzmno9jWQrmSfQg8/KvPdhM4OUrm9I/fSB7n8VP5geJoYN6Lv
qUTlmmwc+gcN9teHnK+5ZrNkc47HrhiJ5hxRgCDCuZGqA+uassQD/00Cji3sqA6hmH/saEZvzhpI
YKzdh3S7thzQLJ/NxCij/P0MUfATl70JiArCWfkVjr0X5xVShSXuJWpTxVRrQdQlmdGVZw4cLQRK
ED5AOQrnERcTthX5A7F9oc6nCeVMvRUn9LJ5bSCIA71LX3z5Yh5IQV+TOUqs9neAwt/raBvuWcuI
PKJyA1oa/1RRETPNtoUhJD/8+icMuM9Ei75o2wP9tA98VXul9bt/tyJsb8gKaQWnIDD2cE2vIgZ4
TjiMV+8KmmTrCjQWPJSQtNR6vHct1YBnZwQqQVrX7vcWY0hHc1nlx7LPsWGE7mRB92P0Vh+Jkfs4
SUzT33+R6EVcpHE/P9B0NBmxkP1abRNTg4UcQ3SPdk69573EM8LY1dQir1ste9GUnzD74TprL47D
hJ2TP1AAda7Yjm/2lHIp8V7iPwZKgIMNUrII29YQnHtct1BmxUXkB5ti8NYnLwHCLTFB3jtd07kC
sz1NccyIvAAedLxa1SJQNRzgau+DvJkdgrx67Ncg4KjrXg6gOpCpNpGNjYQM0/aAomviRyKSfFl0
L1VuUdRrbbTji3ndzs/roekZZxblwut1b4vPKqwdFjIi1JIAg/bJqfV5YRggcPW+sBSkRPkor0Ug
/+wlA9QjOMXoAY+lpb0ZNaBHTe4tiutGTnQpd3NlMelWiSqSpLblHiCvqkMzob2PfTINquXee4B1
OavRRkWG1KskwkiGsmY3egpooc3Q7gXaIowftdZiaRxPV+K9zAFCvmBo/42n2bSFFp5qCF4UH0ok
6xvac8M9FPeJylbngqddD2NmuyMKJ3fL9A7WHnbMgr8x9JNUsaPWMfYkc2z+Xx+xML4kOz8b+LGU
pp0yg6w7ZWetGx3m+FsTQ6jL6tNWtN+dt1/3t4TWiSpek6OsTTfA8BuD6FTXQjSJsLbQMtKocXlq
YK89D1QmFn7cOCzmDeHuPlnwYHGLteD05Wp2+YLptv+vVhHicsCtHfxsm1PiWikxsSwjnHFOX6fN
8v+vQjaPMfKEcfbF03+zv279aotXGfK3iWHAqxjdgHhB/URUiOgi3gis+C2dMYGi7QSEryqZXPB9
+oOCUVEBq0l1xu1h5nuLqwekRLBTjmRr2l2KXWG0Oap8xa0Rlq3gaKW3wFE5HJ21n+YpsiiUUDur
/lTz4POj36YakdkkbNPUKJeSteqj3jKK4vqr/JJ9Z3L5Rz5h4QQ6DFpEWgTpnMooyVyNBy8WkLlb
FKYF9GQq8t2VhH+WURoy9bXcsOiyqejIuZTkoakNi+mxTXTDZ39eHBLMJHTBaf3jnfUoeRXMD6VF
f70bWLRu7rM6C+OiCQ84dRsFWPuTVqFYv+wjt7Fw3cQGK3HFppB+4Cn/pMcNtmzF7To9tKE1JdPJ
ahOf0UL7IFfC9lb6EVNeONe1Xo+cAFMNn1KcfJ9XgqVr4AsxwgmqIRo/X9QfE1uE9yyCihfe1SDo
R0vLYxq0i9gamddYRi1QrM+M4rZor080SFG9cMKLOEECw0hjAB6pr8rJ5Ita5lTmpt+fiN3UfByB
maiv2bkOog4YJKBmHU0kSk2HYFc6/V4DTUFvg2SKrYMp4F0KOIO5A/yg8zcpkPm0ZlPihRP/zBNG
YdGHrzDgSwTXcFjrxE1tEFz5wcNdaD28PuSPwO45mFCUbl3pHTGNidaYjOEmqbVNQkBj26cql+7m
mDwz/SRdS4gwwDl0wiK85PpiPRDywIHUcl+eae6kd1YXFo/AGbVFH0W2k8/OAs9akRWlA5R+BS/R
JKQh0DPdjlvbFN0bATkTQB0dUkOeJVB2s9MluNYPlKf4I4QcKTmmSqy1a6VpN7n4bdE9IfW2ViDY
lPFI6uWGlCzm7VQ3PgoUJ2hHdWzTREV58QJPWQ7Yi5IND2D3Q/AxoYSevPdyRcFaxqJwrtqIkPb1
WT+YdQ2UzpN+l3lvVS9seQLfrsZ85Vb2MDuAQZJpMg3T/ns9c75Wwd/miU9Eruv5TsGayYVrSxXr
hClGA/P0W0D7VJXDFJekchqJ40Cj2of5UtyGVmn1RDvAEXJABv4Z/f2xG3nN7dr6iwP02BYe4h2c
Lv23jRLkGVILuYyDfcbrPuCShIKetsL1xLfkzEFU4SKBQfQ9N2OteT7pbXsQPqdIY90dldJqHOvk
LIX9gFCyyB/Sp76daKLPiYTYZMb7L9nGos31Q0+l6l9uAqRY175vYZXC1D+hZcf2b9pxZXGD0bFr
dp2gFWLLj0kIuKdSyNlyICFFsAFXNfFb1NNp1b9YvnrEciG2nbuNt7qwN+UtS7X9IiAcLQALhX78
LnhRnvb8daGSQVJ5uy2vVoWGomgIwBUuF0YP3wskqYKzKgrmst+ORRRTvXIJFYYwZ7ujxSe+/FyJ
HR0zemFUIhnsSn9wOOsmf5LbJppBkvAgo33HHfUtpwjL3d2N90Qul3f0Psqmo2ecLBfY7sJeahvh
1b3JSfMm7JM3DLxfWw5j8IEP91QGHR7EbjGlncR1g86jlUjytGkMZRjHzfvylyFldtMhLbmApzy1
uyfPh1lZSdTluX3iNA+KheGbf3zlSfhRoL36u2ROXIkEhqNDS67oyseuj5N33zAFv2u1kCJQWCgK
ccdNMv/o3Oqo9kAytNvHpmDv2FlB4dvH0EkNFYHpictoaqSZnsMSDeJR7S/Zjm91R0qZWFFEECHK
zfX1YM+Z+2enZnBKEF29xY8zN5YoSQHaf0aYlQDsvGmm0ZALoHbg8haNsYnUKMPTIZ+YyC5HijDr
hVXRhP+DFLzzD5ancUoAojdg70cCo4b0fR/lCTaoaB02MuhvIFowjOfDDH2dCdr3QYBONQuVvRmY
S4V6kGTSVAyPTcY2aoa9M5rz91rnij9z25X7ybSJbDyjYRdF7A5L2ITBjamnshUFISq5AsoUYl2s
Z0cqjTuCVgiucOOBU+eSG7MB/6/2tW+J8QhXmYmdnpJmLlYm1W7EcsmgCIlsRr0ZC+UBXsSdNBID
GElVI8N/2buItJhbqN8NKqbTzzXYVXptX0L39lHkocyjSSliSEcKDEnJrirRov2mg2t8k6aYnpJn
bxCDC55n+TxilGEY/WPgPD6RJxhqqdNrjQ0/E4Mo7dOpSrqmgC2yOpJYeJRwjA0OwLznfS6VEr63
/4rIokasVn60t+3QZ8CgQ2j/WxVKOWps2qou1/Ai/dtveE0+2Qmkbs1MFaIHDPCLumXdM5Ljph41
A56PRD+Z7Jtg2XnwsoyYCRbbwwlhSHyOAAf8Oo4k+Yj1wZAcCkZAxRn3wYuMfhYvsBFepq6WfzF9
pPyg18HOjAyxTRBzz36XJz7ziN8h8zHNNzhv7zqt3mitydkK+P9J7cw8iPPJb+h/WeAfbibbTiWi
s6eTJiuIOP9YzFYcV6Vr1ikLWbM+gQUkJnUq9fG9v0pd80xgqJj1rCYcpy3B5lis608m0I8C//Lh
7GeOeHdmst2V2NQMtSZUhi9TwPUKF/+7Iv5imXdAanLAqrs8p+xoiiuOEHFKPn0PyxIwAtxM9rw4
DKfCPEEo/VC4MAyv9gbGoS5zyrjVU9XRvd9Y5BFX8TljjmnbC75mB+YYBKpeLpNH1nEeM7izbfLu
4EchFe63lJqPj2AOdTey9doUOPiaU2WIrAO2UcOqyEh7pgtIDLA0m3xNds7Lmj1Rn4//0558Lkch
XoTjZO0V9YX5hjcZeqe7QbpcnTpRhTY7cB5m8lcBpS0MliFSe0JfA3ZVuKlRTIoUfwVUeUe5HBfA
7kDemJTWYk8PntiIlD9HWPs9+NqIQ5IQnpjnPOluAd6f93VjRN70YyKAFPgDuILEsB8kZRj09jBx
t9qljjq3DP8SKOdXv63ro1ytM1W74fxBqTW4YjzW0BwTnnB5xdaxe3jq29u8DsrPhYR11vib+Wdn
UiPLVQovxs59dW3nIkKVL7dTEmevXqCSbRndBHofHwh1qbqpcDZmdvPyV9VFFEjXqbxjWHbFfwpS
kDGitXfDj6Qdl/Mi6nZLyztX7OgrrEfQie+TWUcRzuX/xjJbyE/0jAK2Z9cDRkUjv7gUcO2hp62N
hkzS9DYA+pBir7hdFV3oNY+z+zwZpUWSCkkuxi0oy2jXD1IZywQ9MDuiJckcVH/1r9R7u2n5kBn+
4UdRugFHE9kcCRHEDcrO6SEccEewGWYd3Zq+9miNkdOyIYz5CQydSAE5eX8lbU75aIz9O9GjO1cM
Gfq6qMdLnTVGvJQaSTuIOEUWTHp2fuuPvxG52+GNR0BaXpGZD8kWrtzmQllT/OTbnQ8WIVaRx8jJ
DKC5uJ8kKzSeCzwPjEuo82GDm1ED4/lqM/IVPp2/qcOJ1PMiTDBXHBJXS5U6+SdfnufgLyBhFErA
L6XtdvtV5kpLjT4jcARk9GqVjFzzwshplml+Oy/KaXeyk8gCCIbKxaE9ihu5jSgLwrG+h45nB8ow
ymBD9bscshR+3EgasBEkXHvRF29CF8Fxe5MwgbsuPHnDbpcP9lxjgbfh+fQCPR+PBCr2krHhYlm2
hrmqYGSp8igDS7M1IRbzL+IlPkmSYMICI2wCFHHlwKyNJ9hN4eTNQeYNvto0Cjq+TnYP39WbNN2t
nvmrmAXgkd2jRBLcRSzRTqphQs6VryViJd5W8kMOfXiBkUKTjQlhhEZCa6L6L3fcsL9FTs2awCbI
GauMhMiSiwl6yw9teMGkiF+yQE0l8dJnan6qn44hs3/85MALgD274PCVvg/9bfvf87sz702MW8ok
cDJdLhx1zrwzKPRmx1TNMafcoPsUM9z0wtj/2HafVo5m8i6Hd2LrkRFburR7Jd7MBElafVgifhI+
23dlniIAPUevICjzX7UO0FBSnSdXTESCtpEr4JW6VILp8ChC1wV8vaY5/3PPCbWt2ynZobv/O6pd
CszD+zKx4bYMdXpi6HTL9bDL3Y3RbKJWzK1wEQ4sEknDkGlhu+amV70UUgyFBgKu+6JfjXrwr3+p
KbRw5G8pjgJ57OA38iuzMdj+ODMEZdxasZluneQtV0B8VwPMW0voBVadO7Fvj8ihhtldIMp8EpMm
d+vfSwIFO8w23imcNuOjC0T+F1J92QNx2mUk7ykZOtlFLFBOJgTjeXWl+aJtzyHkXe3F26uQUjmo
rSsJS7nHjvvjSL9DOuJH5s9Ubn3pV5BnkB7mYdrw1Fty5ykEDE4o7zeGBVqX8e6dC2bpAQY8oNj/
1TMR9wtsuW1Nx4qMWYJZNV0VzCIoJREtEiO7zTghtqo3EX12/zL+rFBH4+75z3lNQDMREwKNDPaz
8kvST+iluULm8Sxqc8MjpaDkPL/YK+wnXpKSBgJ5WGZQ6TvOmPYzPr8JvZDOCrjt2Mc5iw++KVmM
M0O5c1hT9j1Xdzw0YprCqLfRtwg0eFbKZPGQQk40P6QfIMQTIi1jyu7ndFTs8X+2skMhY57+6k/C
OQyPnyu0ChwnY+SpLKjbV7bgqZxBpROtEW6LIPFOeWwJSGWOp/UAO3syfW2RjGFzAQsTmnRM+7GO
xOAn6w91pwii5j8QYgInRyCuCe/Wei1tQZWeylKtK+MSbUK+5Is63MjQm9Gnb2qnGrcnA/oc2BnV
dNAjg5wtic4XbHL7AH6LY9h9Pk94xblGbaGBs7h4L4khnnplLDyy38zWfBMsC5gVETDSShiHtBNo
pKhmu1ms+wM7mr8pzRfb8mHiEAbfDqB94vtwS9IUSj/8iscGXHlUQvGLCImoWKPbNeJ3WwHqyipF
J/UBpXi5bqrm+T0NcyV6NMMrIZcYEcJ5YZHlXUeQtwC2SIa5AZtidzelKNT9bZf0CGevlFG0hZ16
SHOzYPoVzdrJ1w0kUR146HT1Zd8Hz8i9/m20JsSUsjiBpT1+7HZSCNAjKOYiCHb4ONYXXiv16D6r
WwF2tDi693OwewoMhew4OV2L47ygTuOvSPKAIxox9AbQAO/5yMma0id5D87Ie3lNi1d+V/EkNvlm
3mTGrcxRKFMHcZ/d9Ljg/lddwnG02m3RBY44f/bw1OZ67s1DJwLqX8Q3dr8X/6lnBDJTtG1X1RQZ
QXY+4aoLGfIbvBQVRDdPghLm4Uni3YheVHF3FDjs4OZOWTALrclC7NpgNNHwpImDXG9K2EdvfUpc
a63c0+9hKXXaX2G4Xes9y6pL8+nADxRwRxh9bFty6l2o3uygic0CR10WRm8xAMYuK2aSMiHDe+OC
LrF68LpakKSOWGhATwu4GzUlwHPgLQ/SUQTuzzVWzjEZUl91RuSz+WHQR+Ejz5IsWyv/TbL9SrDU
3WPvbzuVADLIcGEcu9DlXsy47DvG6WzKtxs+cmsWUA33BfQbNixBLOs67RAAIYYzpOQ+s/wqjwb5
JCFvfRfZLsCxd8wad0gZGcew/S2/oPBfZhnBlx5FTWhewkZ0ZmFGaA358fxLVMMYHWdk7bTKqcQW
5prjx1TKJy/4KGUfSxUotI/3Qu7lQ+gRmj8pjyN8gYHvRdw1xW95JAo70DbN84PtnDxB8U/fMWzb
63iw3u5SWPgWGemkMJsIHkwGxKE387j0CJHDo+4PsufGpaI1ALqxAALfJAIfLGJ1dJmg+9yPg78K
zqi/GfW4arETeBNnPHWvXFdnv25LRl3kAxzxQDx5RHpLc4s/GuB47K6U4sJN3Ou/YO/N8wmaciTY
rkyf16CF9eOgNfPmQ+LlXDDWYhiCo1HIQ8OhecBx3yO5vKjnkcDENgMopU/rKKqxN106AjXPfxub
jnH2c2lp/qKm6r8aVfl1YyITMFwNJS/cg0SCl67GqO/dA6eZeatCr02A4jWjExAGNPWPGmS+iLAK
qK9CyOp8FH8N88I2HzYAwCP09PZgYhQVb5KB7qAO/V7wnatTWqfl9vt88jTHTFalb2Uui1rH5BBG
9mEAZVD6Xi41w/5xCX50ow2Tyd0eaY198m3EePhY8icCxNPokANvt2t7XhbNgJ2Lk0ffomx63UW2
6bEDM2qpXDGJvzSjWABk+j+HbdU8b1yoYt9IGxR7UfVPg5LDQyk/B6Ut3qZfwUlTokkDqEe2KsY3
lQm65GFIgy/JUTzQxG/nreBUobUHC2p/A9oDuqWGZl9u6XIBNh1NyVU9nnjgdi0ptOoOXtI5JioF
SW4fLvvJpZV/8ZINdPDz4DItXBvVHsqmNqDQSn8VN87jEQf4401n6tpwCKcJBCWsGRqV/s/4Y2Hv
kvoSkm0UKX8+FebsQmmrGv22u8bJCrxURUQLt66yLZ0yxspDSKx3ANutApKwNycUDTtQAPEdyOdm
4K32aTON4CMIDxXSenYOsLAVJ3y3IckTYxfk8+s5Z/GDCxINfBLx5EwRD50V1v2H1H7rOOvG5SiM
70I2rAC22aZGBSfPvqx2kJYLhJhj9GFOKj5eIXtUY3IDmIHwW8XYsewGAB5/El5+926ujtw0KPsz
r8QTCsz70JzKaFVkE/R6nr2VfCAY4Ack1/YoB+VJ2j5oKRihWNBAVJMtq8HKXFEE6qslyYNFmYtm
d9Ojla6UUe379XTUx2bFc4QNM94XF6YkQRKsjPKr/yRVeOtVFwZXu1O9H3bbM59QP9s0SbgfuNxk
jX98Ik3T0p/jrWon6eXtSMM88ueZSY0Sb5q14958GZC85OWiMUOjwpWzopm/PzbiF0ugw+ecx9ub
znjWiU+gud9TAI5Kra0csIhcvELh4hFMM/xiA2LN9HBwA2ws+IcdOhCwG8QhccaSC4Cs46+3R+jE
mQzGMK6wX0BpmC10pA3/T9pBxxxvF/IktXTKFP9VFhbmB0jDkZAG3pqacCp6r09ISBD5m/FBIDfM
EvuF0wzAwjjoGSYMi9zjAIiiIXXryULtDSK0jRuWBBwZMLGKmtSyjQo46YRq5Qi12xnhT3KAt9I/
BLXocEmu/u/Dzg4kloOHeLE4VTO/LaSE30obUPXsENUyw6G0qxAjR0BCOmxI4py0c2zOEDDLSEkJ
U2rcA5gT0/tf0MX6c1H74nhuS3NHZH/3lVNQtGmAC4X+47xa6gAmj5T+YIjLNegjW4fiTYxrnVTG
Gp9DPv/ml3lgtytfffgbeoNqrJWBGdY1b8hNXr+RgLPhta3P+QE4kyEzEHKuTsTVgT3o35dNb8cS
wirBTsdoVdcAm2EDfKKq9O7MYpnPN+BRceUflTA5HMpyzNnN/htGpq8MgW/WmjQHYcA6Pj8gp+sZ
WNJyyLiac/N/J2MJDgy40Sa2RlxREHiadN7pL7Zu5Ly1Ks4eSPkFmYJ+0V6orvHcsl3fL9ukdkVJ
y8qFm+EHIhaB0HEDiPF2TkM7x3Zy7CPcm1syHmpe8VVUOpW3dZjlyCflwxBBtev17NHhinJo4iCC
+nUfzV0OHhD45yALnlNrpPIXUbbZIF2yNdGkIwD7RIw0mHb0oex8H8IyXA3f3SFCS3v188RUfvkR
KcfzzrEm/5ats2VO7MHZKjgkSrX/DWOvWQ/yqa7LOiekcOJ+9xd85ZOolrPshHBRvzCme5IQ6Q0k
VpZF4mktZa9ePQhqkdAdggBhIRMjyIYSbO3P6V5eUsglevXSCwA8jdRoDOpmsyFN/4KotUo7kmDS
fnHP8qbbBUhxDvlgU8KPQgNnp1lVCza5YuNwlRhKKUQNVY8IhDu1FG7AP5MVjwBrlkBi5Nhzbaay
f4niH1+QwOUt48yqrAkct/TzhziyyjXmI3nvaTTglK407JtOJlL/UHJ3xohZfD00zqfz45mBjsrb
tBz87YwUZU7cNZue8jkVSGwt/zzfTcdViFQwHvg78a80jIWypWuqIVKdrD8svXKvVaZmSZ81LKYT
j+497Icn7cYb9DPfqfWevYlATGjcv0TZr+b15WLQsunk3rsTYhsTaVYkbQdio4q9XwA3fVVAEbz2
EjF4+O47V2yPpUjtXeNo9Spx3E6YJr5ZEX7doTlQQk5ETJ/ibx8oExCKQ9JKyq1iWkiekec3SDO3
uZ92wq62B5k6AVpBD2g/QahYMSi+YbovuI046nVJNHLWHmMN4A6RMlAmb3wAGiqL4x7xD1tYk51v
NpNVNbG7jCtZkSgg2hnOeII6Cx1XS5Umgs7QwFLaDWvZqy4IjLHuCfyamzqaT8PH18JtwVc+buBO
oOd6NfQNu+/KH34PxgevsNV2xjal1w778umTUVG9dd6+xk8Uee79TFFXsbWKnKdkDpucqyKvZgnJ
OIL4DDCuMpsQPTrkrn8FFowqzd7BmVJ+ptjMeSnpr4YmgKVHbGd+0zoRA7EpASuJ4HvQYBsg5/kO
rgpRQa30wGZo+uiKjuQRSe/YazM8CSKU02RWuUNsmuPXotoYPuKkESHXCO5ypdyetEI6f8iuSfeu
afCYyGWBPvFl0wNMLg42iiKxnLvQv7sx19RH+qpAdGk9GsQjUp3MOTuukRUcgXoM3SC670LaCrZj
Ss4fZIxzMNXIkT39Gbm2V4UDSPd0DktSPhcwIrppfmOzk6pxxGP8ORxJsWJ8RiG5ScMckNi1G10J
9dhU9vqz8pcd8l5YUqO8CLO2i2PH2tuX22hUBogQYJCZrQK/D/wt1iIEfcpiMJ8S7F1DQAEzxgUX
4KPsxpZG10SughhZjssdlcSiXNBntztkZA5Cw2xS0dLkLP7H3nShueOZW6szd7MO0u+l01ert79n
UrkTcTDp+CgNJrfup6/KSuzFh1SSE1zNnmwXJ3yExSRwcqGDrNHauNyOf8g/4FElMH6daNimAlCE
hC5ZmVrrfiXvDc8K9gDnyACr2hLEnQPKrunIOdfMQAVagril/FRCv4sB9yxVcVH0tR0wb8Oq3zes
a1GRvh3A2JNnAmm1Kl6gbde9/ordNAEkvfNVdgFdD0k6/+MkvmJ8gtcMGJOxgiZtB8XySL7gjam9
kVL9YrUuSs1/KYPYK0VeB7h+jSunQfiWGm1jyc0YJBwyinbv5yb3gL7xL9OF0bT/wDcMgtjhS3zu
BCfaT+ltF9f6Bs9U2tJvyL+ub0xOvQ45zgsPS6ufBwD5Hce18wK9JiolwcPvYvF2itewQ9lXVB2A
DlhdJiXxgtVa+V9umgAtxvf50SckGn03m3jDr7jOqkrnBLXWsBSyp5bItcwMHlLHB6IP3vV4Fb3J
Tg57dR4B+gLN7UAXsMj2PcsnmRFQr99ICgVhX0p0McU0bOl/l8K7gpZvYbkyROjf/08Bdpihi6OY
73HfLa2ctvaUCPJDYrG6PMxfOnDiN6JhsrGMhrYXTSUezuI5c7NyVlYDOmkRVT5u77TY+USM+SAa
RzPDbbr0GbCuQ5R8EF9sAE4cnaGyYObBxQsDu6j1Lwy+3E/SrPoCgBvqZBqWZVW5zjRKny8FKN90
EC04ZgzmTmwTSFhxIOCsvxzX68jd84ZNHWQu0pz3fGYAyHKqPAe12yJXL1vi9Q3TEOeiP7B9stKL
EpueciIipvNUykPxxEUvgaFoPlAcZdpEaGQuyXTgGnhgQJ3N56g1+2MeXfNjCinCB8pdAgO4IEc4
KPFKwRP7E8F9zAZNezWUnl0dCGrITMpe7BCqxvQ8R10UO7qlbItsEkIN9w/Sf/aRIUeLiZBKl8KI
uLIn+YFUoNEpuEk+c67jlz8LlhsW+vyBrHZE+q/0Pk64A0v5j7pRuDFTmmB/ii7gv8eHnaguRiys
op4zjv/nyWQc90f6ryR8UIgggvNAP7X2ETi1DOQfLyQsJm5nHikUhBPAglM0u/e410lRAsk6HCaw
xqCa8GtRbM2UnX+rn8uMFcELTvkDiuc3dty/GZFmpn1Mh5xwOQyMZPaGixlPUpkUeZoBOW++RgJT
d7WEq+3a6plma1MzIihX86O4imfMXeWeE84MEsm1f7VD1tNAwePqQ7Ro6ym4t+mloJ2/aX6vy0J3
tUduPom/P7QN11ldBI0ZnzqHsIzD5MFe5FNIgHzPeUwEhL/x31bP/uLFOla7tkOPrHJB8VOy/aYK
CohXBLA2Qaj7VRtzFYS7U6kn9RP/JQJ72niUkW7s1KbsRMy0CUqDSf2vec/YxEeVklF9DWevP5L9
mOZKlPwJur05UU7wz8oIj/XVY9ENnrN3igXE+d58dxBtS3XVSIX96T9E00EgPWbFq7glT77teHFF
v+HAIyIKWPZNSzLxcM61seVQKiP4WMeq8teHxIMxqmbAJYH5bgPyQr6CHsSZiMuwCklv7wKF7wAG
5pgI9wbNx06RMzMogwV7Xruv15Ux1HUs9Me2NxuNz22L4GVu62TEe66SGUWT4R9Sehc8Fq4KGdoR
Xmgk9YgwFGNoQisMcuKQI4PXGBoM8OVl8L069s86CO8hj6AR9k+FafoKaJTil1pdl8cB7Iw7BWQm
sWTlec9HH62eLr6yhDhdzNB6uCcFGxnMQdb9jPlArQNscNy7f3ZdnKTiBZsmCFGvcMsZY7K5vXTC
ejyoCDp9STYawF+3Oe+klGd0Snk/Qe1AYmdVPLx4mRRA05NGtRl3hNrhjUOdP9hbQhazZEFtBpu1
DGSmqW8I3ODjX2+SsEfEUoaUX0rY0iEdLKMXpXC18w2ZuDmGxbzAiavPmDD8e123wb8o+7iZ6aQ/
nY+u10sddrI0PhTk8jnshw1LbXCgYGSydjDHmMTvTRdLG2keAePHbRJSMtIDXzSuRhMqr7KjBzlP
NIn2zokL+2BVGHioUifUKbqS8gfucwy5FZc4qED7YohPCb07io10n0kG1wBlW/VxSyTPQsCi+z/h
QzBkiwrWZ69zP1nw40r5k9EnWySZyCsREz2jtKJlDQ7tJwT6VlY0mwiskneZiFzo+TVXLiadW6wv
C2HaWBqYO9iBP6VRovf5darfNDAapmz3IALQjMU3eDHev2YOCFfa/4z3+jXvT5xHLTuYTFksZZu+
j0EnZugoB7l35nh6sI/cCRQU3mEq4lUdEMZ3eUqIMzeN0AxzBN6WLjaYMv3Zh+3q0kGsumCBXTp9
Jb7HfEuIQfdpLy2H88KmltZr6GyAgyGGxhkEF2Fy8o3jCXY1drUS2ULG9EQXPwRLoN/FJTtNN5M5
6+UqTQcqckDz/c73T4UtJCYZ+vPDnbZL/WfsQV6RYHW8zwc+KxGj8PHwNQ5AUKiPTJ+HwopuWHQz
Ow5sl7u64sivVkXrlBJ2e7bn7qzAibXhlSLgbJDc//Bs5wtixoViNdk3IfmrngeIqjBfvjeIvihZ
Ixgv8VqL8kwusELvjTBVYsBp8f38oYXAoElI2javgg3y0BhgORyKEvFqN45KA1pzDbcdEt5FSKJt
WAcrdNer+iwyT6ncrdqx8Lj/rl+xKuKn3DDGKLtIHM4A/5jPcZavWTQUYsZRnPMhxEKNvFh1EQp6
Rh+Q7KKc+/gDkq30qi6DO9EQyZEYlxdTa9Nr211bocHDaSGA7/Pmpv8h1IkKZROFpZUFLpXHslEq
uEb5ivKrOAr3sd3VFewYtuJJlYo2CUk86PsZ2hW1abJuCuhiljDAIwwa8sNi5ukpXoRufmM8lUp1
ZGvBMQpHkZUUNhPf9Wf7hOXQfi8vgL8o3+FX7+BRy0cjZSPonW20Sp+MbZl2UXLGnuwl7b/TYdeS
mck5BjbU+harQ9L5J0U0keS5+9FUOTAY8t7oVT8yGTD3eOxVhshwWEKrpQSSVZJuvPqHUyN+psjn
tMnLjlVLe3mda5jEdMMSm9aSs+6XSeVC37rKd/P0rNtniY0umogo8HqP8fFLeV9l2NJwh1K5TYRY
t1Oui7tpNYDaPcC8ZIJPRP0IvHsDLWavUTrFa8G8qnLfDzM2UJqlsw8wsGMaqH54I+fB6jAN1rMW
1whxRzMYF0XXqslPwHsBouY1QyJVt5CH7efQ9T7PtT7hvmxOeNW1LW3iAqWKEHQrpyMf7iR6If8b
VKCJokAIssIWDayriQQkRm3bcZ1QoDGBNV4S+KFAu/q6ne1Zn+fHphg8Uda7JasAeAlPIcBeYvZ2
tzoUDoRCbrWsI2VvLDGj1wZrPPPsBCllzmzDXU7YJ8LK+hV6M3ExbcXF/IlksII2VCJO463/k7kJ
6pOM4CrFukjxrCsQ0nGzbWZg3Cq+TrEAyRBePI0lgpMG3fqfzjxY49GpUlUPyWUbnvBYo8r+bOUs
4p3XhpUF8XzqwObSDuLoO8efAP8YkhxqYYskRcgFjGXn0s+c9qDQnkiFRR9qdqqeuU5NdSzXnrC4
VwtHyWMi6BbkqqyGMQTJjpwg5EkpWNpTXGU3GcMtDhgoXpnHBxNAt59HJYPhOMCBOxlMYDGgD7YI
MeuwVsIdUY3oEUjZDB+/XOnIg5AhN8zthBma6k78w8gcHprZ/7QWZrRMsB2zuM8LsOjN+5Os0qVb
+cEt90jjJAR7tNU0Y3esnEjqq2zSm/zuXnY8IZKUGwFZjNnK6me4oB9fBaL1V3otdixAz0oLEfTD
1xCDp1PtaLNuPzwBOzCdnYX+3wPnGCG44xKTPMREeZiGESexnuW8iUCYL66yhmusgRG62ovaqwGW
hpb+BCk3KRhtg8o74dJUA22iKVoHRdzxnC3lQTN3NRJRLupVD2peglUq2fZW5iuvX40oz3X26Va1
gGkX9GTBDTWyS+/+DHfhzUGw7gh+2hamE5TwauQ8CtpUvrD00ImAhrDEeQtT6s6lYP4pllPDHpNU
7yy6GbVzHsnrVNZQln74eMUh/br/9j8McppARSpzPpvsmZP03vuR/zCbbTWTsPOuhORK9b5aRFxs
gNQ5SPQc8aVp8ABdYyLjcwPPLFlmtS7k3C5Agxnt/0e1aopSJPRjIJS0kjAkmVw6puLOX6nnkJ7u
9BNxvRzwjY6o/1rYHekhDdYcp5f5N60UrIEZoTqdjrzpkwsYd0B50FojJXYas8hgmf0iaFBqBGzz
hpiEOG2JhBElywh2SQA72QCda/JEhL0k88ZtgNTz9ym88fO4QkfSNQSP/OqzPaSGhY6Z3watfsR0
ZivmnDlaGI24NCBhQSlS7Q7S/3fKMBXoMuBqEjyi8AecnRFF65KfBpHrsrI7w5Bmu1kal0lANP8/
xrgknykGGsNmziEBbmmwueRe4sTYGoBdV6UPGUyX3BVI0AqlRz/+QfE3v6zdZOVzrZKziDxKQmhS
omKwsDLprk2ZXU3cKZpqsC2GPXrIFut8nN+MVjW9UDxLu/8gg6wJ+TUQdeuMUgUJ37JDEX2PYhy1
YVILYrUEe0NYMT/U4c7FE9kCKaL2u2QRSjqXtkZWT5M4v6VnG+1CSuP1qEyc46v1NnH2mO+XW6eR
qhuZuS+vkyWj//9Y0caHB0OjkZdw/Qe8G0AiCbKPf4A/GWWndWP9Qndkl7qzSdsRqRKvu2a3OjKe
IKGUL4iacIrNHDfGRncqSGYQNQre6Hzpl38TDbj76JsvDI1UITDpNrFpu8tSH3WXBNocTEqKjBXA
1x5M52tpZvZ/piW8zWY6CCRC6+2xl+1lTXHEqU53ecGNlAAib574Mm2UPHVsujhmvvSBJHTZDmHn
cBO1O11YEPrY2iH704MCDnGdPr3kCoOxG8IXNjeMmzkSW2QpZxieAm0igXCtw4NAYzMVN4f+dMJA
iuDFubE361WzExhRwHm5Irbk5mklnRrdsplzlV6UWzzxfDS1uaDdN/tJCWNZIxvOQeEfYlo0+PCq
OFXEiKy1Ri2srCPiy8cf8zWc3aAGOgQx016v2zB4BHish+VhO674iURKG+TqPsNud+fZQqHu70Tz
nxZRAJXkl2MmtdPvJOBwx9y6M4d7xExxQEVSCEZGt/R4kqfiiAAP7UOPXh/FyE9VzO2i4M+L7Wlz
0OKIASgiSDXnPFK+ccZMjbFT8amEI5miaBwk2tTBHxmpjCDr0cueQY+yJr4o0+329l0x3LIjmv8m
skRU86RydE/gX4Qy3Je58z1uz8bVl6sbyVseZIeIRh9Dq+XDjr56IU5l1ZiImHEjPdvAQcOcSjtN
2BZZc0offlPSEmtGSWJr34Hja9LmPoPhS0hHnt3KNghzx/djWGTEHsCdM7SV0w0Qh8PuCxJjqbHY
0D6hWHkjKh/qWZrc0BgtXjgik17tyqhnZK4bTPoC15tRqCZAFKEQ11FkwR6WEiFruOuy+UnMmphE
M7Gvzsz8QrrqbtPlNIhnjCVzu8v/BsNUgTNSp/a6ZjwQyPXqbKrpPdMS9Kk4PAch80WUmzn6zf1A
mV6BnaGn/bEAP39vorKssMd50vEeDIJXdrqU4pV/72R6H04XE90ZI97TbLnBuX8olhAk9qXwnXwY
VzTSl2yl0Ra5FQxPyYq1dbb6oiEt64fh09YOKc5jrEIqNtaa2EdSnQpZCOVzeTUH7MgOFyc2faeB
VR78gkVGMU948bL7118S4X/Qc+tCc521U9mKVwGPjtGS4MkLMjOYX7dh7bArO66DV2DDoubUL+iC
nxv+JXAU2ADuRKpCkBhJNcEC+2RBXlEoF+6GgL1sdGPJU7/t++zsjRSKMz2CcMfNHJ/av/C9Gn8n
hTdHEGjKFoB4Awpq6PdzL6tyE++GFR70H6oeLTQEFkD8Ng5OoYrG3QMReqRECPbT/fMTZLrYcTyy
a4pmaFbHteCFjLUwk8LCtt/ocmZOxHFOQWu46W3t4+Zc4vWATF13admRcr5cWm0a611/X33em1/7
NtXrHEn1hAF0gXmUqlKMlCO/3AtDYk/f4W1lPD3W0K3dr3eOnb0avN9jOtJJe9UxxaRcGj8huwrJ
/YxdghEkDNF33SaRKdqAAccOF+EnBLI/qmBuvB01olebxa545wdfsheDKm7cmicPKahYriYIJELC
ceLZKPIvL2PpJkGn6ZR19FLSZvwfBOkGY5VYFK1nL+ehJ5ZHb6Ow31oZ9wy8Psnh6qCvTJQ942zE
WOYi27KYalvg0U2NKRaf30nbUkVp5TWkx1nSH6QzpuasedEKnheHlGDF1+9LkzKNp1j2aP+UdFUL
LQZIBdChFC4tmM2sIJA5iKqKIqYZquKXLLt4CdCBOVWcyqbUoFXqjIPGEx40I3Cm3dkwDBMLHi5G
xll/cYV495dLOGYjlu4hTm7HKFuhRYIAEbKEQUbCS7JXLFgl1zoWZkhz9SZtfBBZMeiZhmnsuQtL
sHHJFiWEri5lNyq1+3Gp0Ejx4ei/JaPT2N52bsnohntd3tEmeQZKIJlU02iF8fffkCxXy6Zvojqz
ru80MB8v8NdUa2ElyiiXU6XUYXSdvuHX05YvGVvmJNYgrdnvfDE7KMNspxkBVKiFXT92lGyr/azZ
qYCcB91Cfoxkvin9k+fea6jG+oSn6BrBLfTpEU1DyvauNkafyEI2X9Gf0xLu0dfDRJa92hiIEGD8
Gel1cENRRB//ISzav5wkZcJ7rTapvPdUpShaMqCvkVwuAk89js6k4W5/+iyccPecLBPqzWLBai4q
w/opgny46dVMBY1mEzdsaE/a17QgUtg0Sor/rOCJWlo3GwwgXCQoHhD/qx6MPv11EjgcIFvOGD+m
rTvDq0JP/B338ikkK6ePf6giGnBasYJxftTRSE0S17eQuIIq8Dt+PY67uv/SEXc5ShcZMaBCOv83
ic1+PsWHTs698NOX4geh+Tc2mRigOT196l7o3w/Sye5o076ju39JQQk8dLQ00+cy6nc9z0qiwldp
tGPAtfE7KAtDimVUeh/n+8Vw2QF/J3zm4FO7kzHGNM2VDN6JirzwyNBmL+w7sgMInLdbFaN2xIqB
csUYjhK6YsMgz5EcZWknJ8f6Qg5g1rm5NuDnE8szajAkfOeR2IRbpRJ7ZGcHeCvOcsHv0kgNw45L
Em40fY8ArIzB8CQm+wQTC/9KZo0wFLPymchOlUY9B4jmsm27MkaP1p+CJAJ1wbybTWCPlFsYSMkT
QP9kKzReMEwX8Cd5fgaCmE7aBIy0Zfgv26bvK5dFB2ukWk++AzcK6YqjaOND2F9l37eKCJRk6laa
CmdweAl+HZpAdK0VEfZceh6pgOWQfpXMNipgxO8kOkz0d23O7o6uXIvuz2t0KE/k8U+Tcm8j81+i
haDxweWOEFRMF7DEJN3g0ddWTNg5AzZJ6PGR5aclDsmpzlX0r7ym9s9yCejEnODXw1R2epmyegYM
xrTynrtH9JW0o4qjWtxfnA99XzSdqaHIoN7iMWJt99T1Lhtr4y2wNJ0jgjYYMeRR5UAQOTgDUEj0
DNfSSbON+FWI8mpkdzfTRGpt1WSKpmvSdgEVqT6vgpvclqNEXake5nJIc/AaqtKTGKdnTDQD0pIs
AxeF1eviEWlrO0tiEx99VzVJBCXAfoJBZM0z7q54YxBZD5qD8L0HzzVzgfg9NHUDZmZLwiFBrCZY
YIo9pa5tLgOvcyEIKxmbxVqURi6tXyWAMu6w8XQW0WkVry5zKd8W7/ef0nOCeZmj/yRY2wv8gzSc
YQKSBQ4i6uTaOKbjqw/JNJb7C7T432GJOaD+JhmAVip0ezfcsW5a7KNOwmbVBXwQUIzN9Jkyp3Ax
LwvukRI26M7q6xfJfGQnngutR5EDt/ui2/nm4mtKjSveZwBkt2nRjUyxrhdSk4XEuUJ9UtRutvg6
DvDa5dI/STILyeL1wKdcykcBmboEToyDYz3ocjWDo1TJBSr7Sz1piRbm8tULPz8uMnn/lzcq8gNk
ohp33dbwQVqIFSbQsV/b+/AEj8e+tP8drAb93/yndg1SGA6NbbdIpgQwJ0XEdFQBxhd6WS6gb77D
CCAxzzR045CdF4SzKCrH+dw4o8PvUcv2KCg313TUYTCVBRrbJYzrGX6gZbTJ+L/dE0hLDoQmQaAT
Izdg1pGJIsQiZ/c1K9owM0J0Bt/9JkL7QhFa7eevC1Ub1v7MPzV3XGYGIaEFzMINmFonKZpGheiZ
OUSRdseOiGHKoqFR3KTjmarAN4HDEGOlicrW6Ud3OS/GLyel3RV6bd3xF4eOcs0WH/J6CTyBA9uc
j2/uzKjVhlUsoR8jGpqfFYDV/zgkt8guEhAh8QiY1qKfySj//ErF5BsnXqHje+VwtAeb/RVOKpj4
sP9M3Wj/boX+VaKwZORJEuJsDWuKuTLKNXfJp2kcZPv36Q+nqUZ+prNoum/XGmX//EAqBcS4oHhu
B5YFDrV1JVldBvxWvWg1+vQ35qNoXppsb2OzFfWVxvlUTl0eDcF1gNERWVoVTVSouA1N1SugjIme
EADd9odGlvbDfjM4gk12qevGZypXjJCG/AelZt78P/TQhNzZt/SybE77+TmKJoRN/Gdg8ZTclmOi
CUqWyXhNuMNSY5d0SM7mnaPL1Ldh/Qq5a2epthyaJaDO+GmgMRmO54iK6t1buK7etSyePLTYWGJB
YXZBy/8bHjH1LIniQs1kBibEopxzrJjRw5IoWErHjrqCa4pkvINQu5Km1DTjdY45hYTTKEQGZaHU
0rd1agCoY/2uG1efDdg9TDHE/Of9SD/5ibNEqYptK5hRLv0uLKTCHHiulwAZNUkdweQ6iA4c4VtH
AhoMmlVHvTGuQI5bDeUtM/4HGxr4+hmSbqzplStO1dFvgRb0DI4QgVMVGm1ZGZeoglsGg7iz0+ze
xWhAgwo8BetldivT7hyJH73rcoX1hV/z/Jt+GVC6glx7AxhuvLf5i4KvS2NMlda6P8Xsc8CB3eT9
knR0LmdmoXUWMvo2dJf/x4RWnSXn/av7vsKe6VcmJy9vrqBxplBLJbK+0uQz9ySsfkN6ZUvHbbcz
dF9gUGRnJQCpyRQvCmSavD2+mEdMXy/pg2mwUGFqtZu8hzQc/VFq+m3UV3uyNWAUq6NRnzwwhesz
aJS8N1oNASUqWbg7DLYq8yo14iZzqsp9h2xTY8jwPWLwEiWflqZVEHYcuvP/yDMcn9ljHpaCgSN/
fSrTQj1uJT0p9iice120OUNKZolW6r7iHkLBvVg8ySV+cHIMeevXGLpgZ+NqTZpsQmbvEpfx1KpR
NkVs2kxl6MQniGqQrygiNLM+TG3NXUmiuxX1ezh6j5ePGrLXrMnLtCG8/FN5SOQRhT/G5PpEaGbg
ClOOQv+wCbaCv144PZZkAa3a8t1i3LdbdTLAKi3ZxpTMRgA60c1BPN4Q6w7Q4OP1X3iPTy4qfc5L
CKMx3i89oNhzY4einmnGCMQ/ZzSPJZWkZHLhWeGBKL0rBUEvQZuLhdk/HuNG1gdcZtE/4eGo4mU/
0ZQWlUdCZubpJKtUvUSMxJ6sApx9f/P6L6WT/bfp2sJ45EhoK3jGabNu/OvDni633SrvuSlAs5Tp
AAkKkwawlPgZaU0zbxGHhKL9DuKVui45/dSiD5eiH7TONpclvQvokGkjmTMGcOm2jLJMbypZcCxG
pGWIsyHHqZzORyGD3+/1TXYDgOtiE/KZ8Za9esLuvYN9TLvRYbJhgEbKmXKqfUOYIv0mQdXgPIdR
hSKjF9LOblu3U0pZKHPl9iV2Hb2C/wJNlYxNx9R8BJD7v0HalOx0EZ+SNXsuHrkolX70Q0SxH+DV
FeQsMb6vbrMauOfrUuBMAdkKv4qIfulcKk3HGbZ9iftAXK0UIRyoM+BrDUu9EX/EnB8sRXP32O5M
d/ZEk8GOOJVVACwd1FPEfh4JOHIev05ztIJjRKiwx1EZ+lGGONhqc0M/ORDT+r8KSgwjz8m15dGJ
RnDQJMzyjcPpO6pwjA1vYgIWV6VEGHnl0dJKGKd8tqIhvDFCEEXmGQqeRaLxqANZ2zerf+j62KvA
uktW5Fgk8PEZZ/2hKFIxApRCVCVlQ06WLEsEgVDlhXp68L6iBA8tGNRh+nzLSsxaCRAOFxNtbJJQ
Q13LV36kmqk1wfsk0dxVDre4KDdVhPekj1F7sBbg88ip29pvk3Zsn4e0fAw8vZVduK8QQgyKw1ym
0jX0Oak3wRioM7SW2UXwMPc8KfUyc4zvXkHMSkawisj567M9OYieonkCD5JA7zhQsW/wOfC5Nd+v
lnMhrOMKQlClBJcVV7uZrwBZCNhw6Y2dOTVI5uJO9txVy75iOaPwn1ZRh/yDMP2E934lrUie4YKo
Ze3++bnuvnh+cr2bcJOMQanWbz5CLvNMnMQ8kVs2N+cCk+qJRhwnbluc0n9TYFJYQMmQ2SK0Dx18
/4CNAHXjj3AKQ5hm9RT+OFjrG+ff6b1lgsHaPS8NYtC02V2T4xm3pNNtCI09a8hA8RXRHcGf8hn5
QZwZeVhtbIWgfKyuxq6qkECFQcoSknqCYh/LSsYlkmMr/mdl1wzRRFxWYxOlgtTem0NEJ51aorsG
aflgpGwBnQmo6HY18ak+PJeZUu7RExeFGKmrp//x0VVfXlZPn2ThXhH18ds73BajWLU+Aw5RGJca
KV5JdXOaXARY285/+BxtrIbi6kyUhcnYxvJDfIYPbLv7fyWWiNVJy4LKe7ka7jxmO2H/O6v8OT7C
vasTW/Qbw87iij3X8gD5ddwHbaWpr1kWQ4KHEW+oc5YnTnFtMfnuy2PUB6IRt0grE3JsokbuQtpy
FtjjYiJkfB9k/7cR1Vl3sqhsnpF3l5zudPwdxZBbWiOnwwV7+UCedeSiR8hD+aWcVgmKiNgLMJst
xjdIh+QRlL+WUAqWeUoJjNYz+TLXwTVvy7NX/3t7QxAf0tQv5bVYU14XNgLW85/MKuJe93itPUL5
lIylYbHIxzNIsi5pftpK22LmsAuD8YNGrnFjIETUFGEc90jhJfymQ/osY8bPOyYB6cW3yUFqDsl2
BgWo1zJuUG+PJWRAxhBdoOGvO6XtmYJ4lNxej0T5+cJ3v0Ejto75j2A00O7p4Q6XLv8vgNVnKTaO
36wFgs9iMMjWDSFLoGLY7EFcxQVrpSbq1NvAxKLhr1sTmPdCVBREQU2vNec0uMlhKtp5REe3Hq3L
csDj2Idx3tR4zFX/kSfsYjHXk9UEwhmVHOTi7fC5q5evOnnEmTiGeYPfvk9Ts68Lu6KIF/5SP+TU
AjL/KRNoIl13Iv7w4AsjQwwvS0FKrAYOKezgjldfbJEjzsMPgNFPRaGdzhvue544rrbULMrtV34g
LMo0uQZc4zMeWkBiRp9DpXvOpPJrJMGOLynGL9rpkCKNW9MMP0fJFDxyhPOS+XUf2uosNP3f8mUw
SK3eie+Eiw+o806bA0h4hDNsiacdMtcbQFtUquLDResLFfl7Tjd37xkvfxFFgZoySLkm0XBtfFW1
14twvsKMgaWtDznXbygXCg/aRTcEYEjF9Vei4JCEFSB0t57Qg6u1Mt+hzMgK/lLtF1VUDd/e57cw
ei9JG781Dsyb293s3t3L3IO/rCG0LpyhL7MAqn5+jliOMkV4myVaJ0kYblj1IjHA08K6xo0xc7ns
dJyQft4UrxC1CIcGt6QSYHQjP7t1bBLN+e3cceqaxUgBR9clgAI4eupV9W3J6+/sPWrq2EOq/ngF
YbN5zbuNTb0Ve4P/ob42Nuyfob3b1D0U93u+wNRQZmKqn4zKGxUSnc4T4Zo9KNui5e7Hk6tEgW7g
BnVGPp7UujJygyQO5Xzw+1D7+s74dTahnlDh7FywiUYTocizUUPByUkaOXH9e7uCpt0S8zeGQSbI
9zxoNH2/ZQeyJjjS6jjOWztt/WMyR97507A/G7mBVuAayZGbb+ixM6fX4I0AvkWigoSMgxaEIlaw
Fq9WPA7svJ7ZmCXu1kD2A5PBWIEC1fvAXPF8R2oFcb+IPcl5GOKOgMoyzWd8rBU97Wg3Xs01+Jwx
rl3XROoRPJ9T4e1tVTYP2ujT4N86H1H82EXMlXw5Pz0sSBRyFBnttk0gSs0YtcVQ1r4kNk5Q+rgi
23fmFLVS+gmjb7pdEt+B+0bv0IxEXPlLzWqAQeuIFUoya6UKaoJOD8H5HWMkxh9QiVp52TBcD2yL
pf0/RLU0hZPnw8JvbfdER+Og0kIuHgG27Lv5Fx5U56q8VGX7y18bZ4VxEC/aJ3xXvQ7XL0FKr/EN
4K3GTKg4xn6lTMg4edX2HL0aQpjqVjbWXkONKTrgeRvAf61fzGMPDbxoB+gOtbDO5pgpsyQeQuyU
fZqXIF8TOmOpGbhDfnHwidyCfxajsWPOM9Ydcd8oBKwWySGjgqnq8WEsN6HNA4pjh1xEuN0ERgQz
DtD91BJnj+x5WbzcG6wP09ip3MlIjo6QCEqGqqsxy6bNUzJ32kQ8BA6uqT4ej0iaYROTsNEX0246
CpR7NKQXBNoIdrJhts8F3CJp5mow1nA6ULDy+V6R5Pi25rPoFI1Wdu+IAmKIRKeXUMI5hMXM5dgb
0L2OxJ2jFEBqHEtrsV4Ot5GqFaRI/bvH+HX93E2jA8iJh+Ju4uQBA8ofxNbsjhNUC1r3NTndQR+4
jBYZR7E9elw80K5Q4LL8A6yURW/Vd+u7ndKXurGQYBjt+coZsPTKtd5cG6yuiLWrvjm5C4dHbW2y
R24Kf4+n6u0VMhqSbN6j7BGTezW4Ax+LtXhXjpvRPAPCRmTFKJUNzdnDxA/TyNofuuSDuBeChnpj
k4JRNlKMijY9NK9Ftj2nN1zqhESvq9vY/DSYYEACOQbN81okmW0eHxGkAbrsnNIQiig17PT5Cjgu
ZlW+V6f3LI/xZkH1nT9lVZBwCp37XABemi1JBGDSTSxZ2ou58sp5WZNHhA/JNpIvgteTHLNVQyQO
N6AEdpVjGK+u7qazzc48nCGjpVJ5Q6SHh23A9KNjOxFdSdISQX3iB09Tedbqpai2LK1La8wM+f+n
fapWGV76pFKvx71bCpATmBTyHhqgWAQVzq6924lPVVqgH7OiIGsv09MaePzoE79LOxxAOWfAF60z
X3Ivnkb9CCimxALDkeSorS17cSVGQNZkdkxfoE8K5b264295+p1xwI5/M6VsZ95pi4Kuz6wJt3UR
plDzzn4BwdLZzyc5uZ+bnR1wbZph7IHeZNXRghYHJSHBC9XKggjGfAuQtHU5MRRveWlhlrQgjdOa
5GCN2GHVzoHxirfJgj3+q9szEmrYPb63yc9ovmd5k4fCpT56EznDYw9/gGSjX1sVS577/RfIJQqm
muXmlwvPIVdDKz30Nifem0zyZ/7DFwgx/SrRnqcIws2ok6s9dWBBlhtbyMmwVQFro30EW/slUfkv
1E+GKACPX+XXNbZn9lXW+As7LsuayhqfoW2XY3d7/OaI8Djb9uUQNjZou87+wv1Ew9O+UMU6qNfR
jREFj6L7tu6K2uXJ8KN0c6izZYSrlRExB4V0mdGdK3VEJSRkNf4UcPfIWXaupWIyr0Mj5/JKUg1R
o9DwiRggai6Fewm49GkSjEtmkkBJJcwDRdeT9pH29Cy+VZOSv98sqgL3WtOE4BZJmXQ+9IxiUlbX
8KmmqV5Wwrgm149HTYFNzSMu1zaNWIh+AAme/K9vvuDrztjNj+STAkYFtTrTV3VeppOcSKVRcuCt
YJ1D4yWL7rxhsQe/xmibyyTdolaOGPhFvcvadLfKtpquPbVGd9XQFP9rJOwU08oF5XOn0SH7ExF2
vB8fp+mAayBTdITsc/3qlZFHNmn3WjUdCEIfP+8K3ApuySyk/n3COAgH+E96rjKTz4bbq5kLAgkY
Ff1JJsgfb1Pe42wMy2WA0fDSk34B8OqIqPHdM9wl+oJsYD0reRk8Rs9Wqv2IWKu2GFBDkrIKqPg4
AsdMPSTQRv6bwsjHiUZj3m2wP2RO/9MEJ6MvTLBwpvibRFoGx4GUXZIeWtcAinRmijkuOE2Ecj+F
hJN7c+zCLULAsa/FPo0CIn00UB5sYnc8Q5t2D8vtObn1D/2wlnd8PxD0ZesljixOHi9XAZdfgClC
ZKv3HHGFdD6H9WoQ37v/0hQDcHVOyJGw0bXUQA2AUq0k3OOB+ci8P3MkftURfdWSXB1eGRrfiZzB
MTwooZubOMv+LR6Dk63v2XCwfAgcJy/rLIbikI3hsPAzZZMDcj/Bemb9H08U/hPi7rECyv92UoOU
wanwQAxA8F+SpEhxxK1ML42bcPWggiGn85m0kb1HijZmsN9A4vKRK+8bFDyOC9KvqFYrOP2DtXLf
bOnNbsOtXyj67vCzOJ3AUiwnB8C9a+Aw2kdFo1kg+c/SEgXC1u1CsRBqF/dhm0SozBaCKRhOjw8K
WrwfsAricntn8VbgYyhyGko/pxSyAEnPZPmNTpluvQs/LEPSidmY10ACrFEzaXUfr1WwkSCsPi6i
h+KH4akopSoyk/1GExlW4gzjEgiBCSXHJzWEpaeO5n+OnTTysNdsvzOvLYUQFHVx9zaNSNC/s8Kw
zUqh93NI940kfQKS+MeOOmQiD0n0i7AepbKhQTpc2mCN34OI/g3Ljg4qJWJG7Adpos2Cd2A/4oun
5yZ/pcS8lFFgK/pFxGQlHmrM1vCGwhyMPH5S54BgrJNFDg87Uk6+iXYdG2dKZ+fdrMPk4mecwTZ5
o8qfbx3A6D7I382BcoEPAa2kHpAJzUhjaT2A1coS3iwAoaf5yueHeL1BPJpw17E1ODyga1pdYVJb
aAWEGk6VJUfDK0tHDykOJBCzxmDiTKeiYTp+i17iOwr6B5eRHsWlI+bP1G8yTVkN6Kp8F/pcyxPE
YXN5XiNO/y8gGQBxdPLF9grxFoD1a+WztCpWeRtf9CSR6X/h6AGoglCC7/8CErIwFOwZR6zKIFjh
w0K4fdWkAbOdoCpzWvFbVMr1TCcEurIvvUcTlq2AcKEHafLIsia5H4SRpBSaxndArjYsbAVQ3vhx
19t2HWBA5A1maqpyJhhQnFagrEBBXBtYJUxm9kVaJbbYk6iNFEQlRNwsiJkVM5B3z/qth8wUNZUv
RyeaBUGYjb4kksm+7rKqo/rdTCTyhpNBzeNeJGx0mFHvj7cClvL1SBZ7FYI3wYqwuueewrydYHh8
apkhnpLgLhx83M+Nh4OxnNZNMn7PrhFfFOw794WDnIyPDXyV3qRAmyM2TQl/TYcZv+yXS/HmqGQm
8p9LDvCHX1I7y735a41cAZwZuagv9w+AHPtJyQ3kjwV9rx1ldwTzwT8j2CmBlr/HGIv3+fsLMA6y
pX5CUYONIjFw/6dEjg2eiGDhOoad+cUtxa0Goj6EnzOvMxOI3pJFuJHgrSU6YDODQUuzdQ0GvFgv
vmithiWZWSp87kzhCfPoVHO27HBY1bFk6YI/1Xr9gXdj0KWib1RhH5PR0HZlPBCBr/oO8Rbyqlo+
KHp49nhMyJyMm9WnuwQXhfytqTS6+HHBaUCvmoCzmEtBVaabuvMzyxc2TpaZbD6vRNHvXHTFkZei
qL3JS+oKANi0wMVD7PX42FFZa61DPteNSzj6j9IiwJq8/hc2S5359jR07FAh7T4nYpnDZ1N0i4cy
h+VbsGsKCbdFr+xus/sgzskryNfJb365ocJDkmga4OpeElISM3/zsNqApzH5qwvsWCCB3noiAX7O
Jv+qUAJTGwLMFeDbanHTXfo/oaTJIeVnmgzejJl9waRFE4JKvo7RAXvxloQsMEYxiaiZck9uRt4/
9nr+5lXQCDZSNs9kw5NiWzZEcB1MHa0c2QeujTTOa5vEUtvyPZ2fO6G5BsDAcJbM88yykTUfxcE0
LCwkFS8jqFEdSh2bxQlc4+GlyCrqCP2B2upM0JaXPjXQOsYlrV8zAIk/oozPL7CGOvV/NKteslo4
/qCKC6yoe5l4JT1J5QgrARCSdqEP6KPAZ2giGJd571LlLsvtyF0tpsEcBAsgtrZDLuMqjNDbk6JW
6ggxVP49jJtmCnNAnAu1mxVOj3VlfVPQaKnhJEYxevvF5mK+G9wlt3/R9Cx1Njl3xivMZ2qYaYTN
jbBU3JKN4AuGM3jH5wfQSyyXrLgekPX6b9U6jmkxxH52KxarGkRPJus1LoVrh1eqq8AcXU1tLbMW
/N9i3gwAb4dS3J4f83vmsQgJW1rpfqNnZrSnsNSIx+jeY7XzV6Mf/zl+rACqQenT6bKn3OzoKY/k
SlVAQIirDS6VlBKTY80gK7Gm5v7em0U58cbbnWc0cL4+nk905egqdAkO83MDW5dKbMieOUx6NKMh
pKYKcRW84QLyscnsM3SPI8kRR6ZtIzVjIv7Hy6K6ttAHVQrb9VtSEdu2Y5FDKYlduymT32paOAwP
i+lSjpPT52RvDsmqqXacShdWo/80NlXDB9gLwYSe8Khb+JU56Iq3yOIhoLA9K7wOfbt/GFakB62y
AQU7QCnlP9f1bWuF8Be2Z8dlQStfDAtT+A97v5v3/Tu9nv2m6zNKa4MwZ8K4uSwJzgR3onKN2d2i
1mxu1CEeo74iDKSn/f00Kc573OIG//SdpwRaahlqPgniLdMeWYeRVwxCOgNVzu8t/B1EWZmVw4yA
bD1JWM4NHfaME78H1TD8UFvOdH44kMJelpD48j2+qsY+rsg2byQHHMwYQds32g2ojDQHEge1M/QT
7S1DCov0EUiANurMTJBNHTwxWKIdDs2f7hK7qVS/CciohsYbH/R4nD/vMQ3s9JHjwgJSUtcHq5Ag
nayZOCWm7U28og3t1/CfDm9QIJ1siqUwZbY5uA6SOdI6/Ddx9/xyOHLNN0KI/eDBLzIXZ5XhRF3C
XrUGWlRmXiqbPZ8nUumNNkwpng==
`pragma protect end_protected
