// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:57 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KOlEvsDmP0rucR7lqpn1YRIl9UrT5MBfukXUq4IDPcBx68nXBAhV4N1kfvUlfObP
MLHJBYGtdA3JlzIPETLoTZnKDozvbYxC8M2hpfGkjIrGN/ML6a/2gaBk9yZ6On+7
MCdW95fXvWStzQCN2zJlxScfupY7639hBzgZX2HN8dw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7120)
bTOiY9P8kAq7MlLfB/zspzs7lNdJtXpa+fmvjQnB7FLtuH00H9hyPuJqm8FO6kDR
XqmNWTwZAFNQZBJLevlQ5xk2OUeCVV1guDcygpMXm6/lCs57cS36+yqbMmybQVK6
NCJUw9Ga6190kdWhR72995L52UUdtPUxAa5560YB+DluQnvZutOKIxtQ6ZQHAcTm
11UF6IQrVml2EOvI42rxdYscD7NN46fVkFQGsaNK0XyQnCu98uvxTSmh8q3qIpvw
JjOsHQJHZEwjNm7ZFydsXjUjbE4uZP03z9tbu2a2CjJ8seoqbPFFMB92K0qZ9yYD
IxIzJlwbVc18I79fP1y3lb8n+at2ng771E1jLHYEJTwZdezvDYliRBAb8tvc1pHC
PpFIofZV4xJVIaytzVu550EecATlhFBkwJTFQWqS+q9AEIPeyXNElVEeocPsaDf1
Hf3k6/RSg+S3YKMYr8PE5B+6fPwTWY8PrmI9ao0ve2Ci7YYn2+BzhCwvOIdG1ek5
bJLhF7N1+eQYFeKT80Zhbn8gWkQPZahNRdR7acRyrqh00mdGQDHYzYZeYa5uSRDc
Vq3ihBVBYywqdWIpjigXa1Q11grj6+CjCZMKUP5dksjEuNMsrpyac4Eetdf8vFvr
2LhwwImYg3RvviLfkggJZOfSUZ15xSboGs8W5gPbkqyGRQH9PzI7gfijyM0wVzjv
9NgPhOyZynN5dlQ3icnM6OfZtmzDnjn+lN0asq1BXoebu0/UdxaDi3s1EDWCcjN+
X5bKHXLaGvjgAZMG3KqmvYWcOgRX4WBr6hZxZAjEceXirqz1aGEnmmoIvGtpM1pf
qx2V9lJxXrjEqFKj3UxV3V0MymlDwg0xCKW9eqcPVhYQMBDZlgqHhVimdc35sybq
NKu3WdZ7vZQoD7BfykkyNVet4vKUSuhqPrIhrVHtx5MQ76mHWeQqH2aY54v0sP13
RaPFuFG4We2ggtdl4QcHwTHVWavu2lMK6awoAaSpKKB/4zapLSu9BRUl7OUQqJL3
LCP+fNYD6tD7thihwiMaL1aG4MMR8IjM5KzTzIMXKQ9lOeDwEpUmBlyy07M85n2f
rOPWhKgLVtUzHCgsA48Nf7C/TxJ0PcB9XDdsneCcXcmuAL9XNHG2YQ3MG/mByYQ3
vvYtAPkyEUh76YYkOObpDHxb5gqIss2c/UTiVL3fMuaG3bx1K9ZUDOzGolNTxSZm
S6HzrUnSCXo2IWzqyx2FM7ZuH3zPPPlnbaj3pQtbGCCT6Sq9wpEr9gxHdQa1hjTo
BN76963r6eJygrAwj4wt98O/pZOIiE0U3KBzVCWiuZCmWA+5MujmdTguSuRZcago
qcGbCJhR88T+zLY2M1zTvwCYZxBHFiWvjh2R+SKnoUKZDMVta8pmbv/NFgwRQK7g
B8dSxIJdYLsJT/uuBif9/ViR8+9qerQfMNxj6Ptglvcmzvosszsdtl6wAPZU6B+p
c9u8fgJbS50qXuJTGzO6tywxgUoCAhmsHjoybwH0bj1F/mzyhWpkwODG3hSq/hbP
kBFHovvwVH8u3DhmtqCo+KEG/7W/B8Gy6opuYzgz2wV2DVfEYi67Y0idJOkmKaBU
kE4ztua3nnlfbOIXQBSVlW53aINgWpfZCZ2YSAB5yrXw9ADswqPHceZUNo8nMqjL
jcUgvJRv466xX9RLqXMh5ZqaEywTGNUJQ94uqG82gtDYvB4RGUuGK2sMrfu0HM8p
XJIiRzpOUxGebpcTIcpwZuskzyELOgMt/GhKVH7SK4XicMEVH5ucqUEFxaYFovUp
NnIe4btBsldT4O0vuNA6sYs/BINC0nD6cSLSx0n3S9peR5Xb9YqFeKBuL5zxIvyJ
mdwPGOAGpmkk28NzSWsHq6X5QWTL1f89c04G6c0GKCDTx+IQek1Jufb66/cnUxk3
LinHcgIvA4ga5ZUZFuS4eJ1vvKIRAQpm/092noqvmOm9m4UBAL7f1HDfiZ3ILgzw
AyaPAIG0AyS43hCTcBTMyJtq2gQWCdJ4UUhcAx9sntni4iQrCSjJra2rxWE/8wpJ
PDCqZc+F7HhLqOD8UUss4YsInlue+fH+uaWC4LmtXkEk2smaydwW8lE8AMW7RKXI
ipssbQwusDrF6utAqsqJZoaOPT2MAO+fV7dvPPb2QRQQt1L+5m5FWt5y3WYTKMjY
UHOplQQNX4fPgG9PNwjFuMkyPvS5gvrpTShlWaSbHjBU62xqJIhJtLJyX7fDc3dB
VYaW7t/6NGw9/imXAel47YOzD3TT7y7BeKiSCkUHwIIBlh50bwSoN1D2RZ3uAHNb
Yz4FhCdEeTPnu4RigtV1YP+Ehck2fbpbe/TdkEOABwzhQuFD6vWYRnCHQggpC7J4
UXcdKi+hB8KtKead/TkZI5FeNz0VtGitzH+6yc3wsfqzfPwqR9j4uvStfUAHF4PI
7cKcKPxin7n2fpaYLW1qyXIZ7A+bwXgDwQccm6grCfGJbVSL/2uaThJGTkrgMSBW
TpooujBhbPqbJRfCGJfyzVcJUTms+rJ//uIyBd4aM/al0kvK9B/vd1OltbTpRxId
hCWtAsp4FsLyRHp1fW3u77AD/QtznGQMkWqS+uQ0/HpiqSv1A/vtePD3G0KjYZ2u
50GdZqZWiNEDOtVpV3oUfJ4opE61+Y+yhnsdhiRS2ZfVOBExwIFunYU0HTwoeHpw
oGWVfTFroWKwjv2GalYLEms70GbgOhAc2WP7D3tP6Tb47NMRAg7Y67VpmNeNiWcQ
fM+O7vxBBlI2CVGJI0Erf1B1ooZQrdqOezgsqZr2NKEefior4qSzWa3ccMDxhTnV
ZRyEi/OB8m6noMgXjGAN4aG99Y88KKg2wktAH2NoMPqHLGHmw8Hl+MDVC0O3fCsm
a+TqcgGUkIiFrBvM/79cPFaUbbcRQoZnzN+SrhEZTd1EAAyqmKwq6xc7oR2X5OWs
+OR435Z9/sma2Za7xN/CXU6skawmnsAA/KTpimWNXlylqWs1NnwfsXayUy0uZR4+
cB11gdHOQWIz+igKuke1fYrUMA64kgMLs0El2B9InWfy36eKz76lUbLzDTjD37YX
og6vmVvY81HCXoqprVqTgtkbHVjjE001hs2R2OUTfYNPgW8UXLe/9o494ZpbOeUF
hwD+iY7rgPXYaaBQo1Pn1ct6mo9MWkUAjUjIF1dXU3T0ZY0cFZO7/Qwj/yxPG71B
UkNPZXNSaBYCWRMOrr0CEgmaZzj9KfexU5Ui5ce/l84tO2fkn0aCDv1ysBqm+uFx
++8NGrUpzkedIopeAdlnLE+q2CBIv2YP5R0NYN1BEClMPmDTLzUSly8t5IA4SCbU
4S0AJpesPVfh/J62lhlqmCvAOVtwGhCk697cZwfevIzzOSSb6qMvX3Lo6QoAIVeA
THAyz2EETN4+w1soB3FoPqp/vChOZY4FKhwbl2bDtIIMMMDZapS2txHcKY3ajZx+
xjtT4TGqBiM6i6GPSIGD103QzQBlqi3UHudD1FGPCsNl9UqcaQn0wnuXsjWMJbkK
AEZJjAyEXkQjySJWa2X93vWaIJ1F9C7pCEzAC04v+sWFK2V8wMsk5Ax6ALueckc9
UOaTScQVoqpJMsu3KWYYBSF2qmGJhTO6uGBkk9jrjZHZJszz0rFo8gfbp/GdyUMu
GvBt3aqJWmjoU4Y6Aq1ljgIwBBUHBYzEp0E6TyV4yrJM0RyJqjJBk3oSdVDDzSbw
gqvKg502tw1VL1KmoVd2gw+BKacYvhhMAfZmLvpDxUJ3k3QSoizWRPoIf3SZ8wPM
fG1uzDePEbHwFYTEqQde6AVJGVWo0l66rsyQXyCY/gcmJ8+5uj6QFepty1vtgKnv
cjPlik/AldLmrjZzr+EJEUkk8Yl5y3/H5OgFlZxxUPLBlHjfPOtNEald9g60Ivj4
vcKA/4ySHK65o8nC8abCrQ/evxJZwyYjtGtISiD+ZKanB8vOJ9Rv9ixrQK23AS//
LaBEYC2fcxWkTQj/mQJvm7btgRzH4DOZJO/w/JyZwCBds0SBlaPcN83CgAnK2Rre
zL6giDcV/KX0jx39Cp399FwQu7Si8nBs7lQVTa5Z23qdvYyEGWcONgoMdONjZ/zv
MDfIIYqAAG2zRo41n08l1P2k9LlPIL+Fbg8MckaC/MsOExw/mqdi2WuJTGxbFugv
VuqVr7KhWY78tZjR1EhagWGM1s4r1COneLoorvJgypE4bwlmdh/447odminN5CZs
CFQNsY93XYh2qO0JrYr47py3BDOUsZa4ukQUHQeyVfO4GU0wPKipJdzbp8HDZ9cZ
mRPrXuqujvZSabMFhH7dZ7RJGLoCGBIYbM1/6giDX9+aTXdbLGFc4zdRRng8GOca
FmevAMY+lHIr0fOjyvbdu+uw6pQSCJENbdDMznDQCsqi7Fr6JfzjFWF8ShvOIsii
YCgtzUVnmFaehE6NtRuZqsQ7/MvNxz1hJI5rCtZLYNVPCM64dBqDFbsRGxtCPdpI
LERS/ZPdIB1kk5MHIF5t6etuDmAaewZyi2DT64fRyDL2NZ5DIf0dEfs1A6jlA8uQ
MbOAa+w8EKBI37cmPOcsc+1qji7BFS3fqdyAVGSpCAKop/faxHigXD5C7BWU/ICz
0kV0BpjVEeRpS9CLRYWdMG7o1ADWRUxFsR6tWAeyUUhQPj2o+tb4XWI7YekTWQvv
GbQRRGR8Bme56Lo3tqueFyhoAgngSlAnZV3x9C8Xu9MZLv/rZbTHo9+jvB2vvbCa
S6N6aBp2O83CM7GmMSZtJspNz0RXyyIo1APaIKLeOHyKpfR4j4hFepdesIMyDZE1
IIgQMUZZOLWruZx5JsTrOb9yX4nBys/xmxRmghKq2e0bh6aQWm4viC9rMbfC9Wx0
0Yf/5xRgHTXgpJZ+/2ZytT4Vs4+iT6WGf3vrZTNz3Fmo28lSphepXN1GUN9Djcb6
+749ETLR+kf6zZLI0OE9Ddam+A+u2U/kL38Ph5mzgYo01rrAl8pRzlvLiYHJvo+I
jrTRtLBwnGX9wtzxTMoTqUFxs7c1fy3LYrmybiwCRaX2okRbpDK17ap9jZDnG0LZ
xdLdFSoV1IlDwXfmq5KVoP2TxEMMphcspAoOQdJI52KKxF0b9w0uVvX8jzbExawf
mVldfGzDtlVVZSGOIyatBFkripTCvMnqoqjc3aj4PIscqNOYmnNfSWqbqFQOjWkT
iLJQHNnZfVMF1C9rTiSlao1lxvTfdW6RtXvIq3HFevM2wUP2qJJU2Wr86/zrT96x
e+WUuuUWG8jCUvhAl1MnRntck4BDI+xGX1KQhNqt5CN5pGtHDkw98Z+Wrw1QayXP
CdwbPlei6u2CMA7snMTO1Ut9+tE4+t8H4qoa2nTRAAqTZru3htb/YxeCe26ReHZT
uCzUkNv7blsamtki+V9A0tIAJ+WiCn6G2MSgEZ4CKgTBrsJ7e0B9eBTxbRGrYSnm
pQMLYiWHqbQ6juCJDF9waYoptoKBTonHub9srkWafVLfRnC+3dpbVt1j8WL5/P8i
eKICg29y1lxh8T5THHq7uVQnPKiHZ2dL2IbxSB6AzhQihqYZWW4KGhqFpw3Wb2Ny
4KgLf/FIVv6m3CE3prD81IFu/0OhAYaHDyhTcSl/+FbW+7ogP0dCyZT5OJ7vPtH/
coFUgepQcWfpFQ43iKMUwwUUa1+dMC4GFNG1gxqAfwUV7Nx8qdZAJ0b1fDsJwLIJ
WTPCqoZnk8UCXEXqNUbhDQXe3R8vBlVq67y3fMnp+kHr3AGi4ZbEkiJlw4ReoqCw
NkDnLYlwgIakDc0MRaWLE5ulTBr6ez7kjeqNfSkzQtN5aA29bOsIj/lrtAGTm7U6
nbPvNd+e/I88Ea7nGKOsDDJtrcFkhnPO4dW2ZOOqYIvVhakD+wDq7v9wAG07B0Jk
WN2OgYxJTEhbwOIKZw5bfZUnOciQtGO+xFVxuZ8gk9UEQinoLCf9kzuXa5OSOP1d
r4GtxbT2o/uYFi6Ronu52SXxHkZSjgB/Pw3M8Gi4WcgOLlmrAJ06grB5GwEgbUEL
NaGVnOHlVE//Qrerx/cE4dVJO97bgJP0gLCxi5s3YLc9chNx+YnFkTh+UapkGmh0
1Zj3bqQfRI0n4tz5Rt1qBIsawO21gHmFB+Z1s4zwpDZH+iBOkg0LaqlY+RJpwEAK
WDBTF2LAzK2ZGC50CvD4s/EEv9sSrX/ax2bpV50Td6HhssUcY0FSRWmlOV2THvPY
/rh5mtUCUSIU254x4Dl7AHS01h1KT8OBdKB6xTd/CwMSBoNP+U0wMg2teGNtVUzM
vQL7FRSXJDVABSQ2ERF3mLIGH6diGKRX0DGV2tuLbQvPO0varx7+4drLZMrXICRY
/g9rHFq0o8TmrxUJqFnnVXdeuvDEnHPYZMNoHl9WJKAmp1zGUUwVRBmsxMy/4cU2
uoTLeNsFLQb9ugO2N1R0uw3PDrjvTTFZ51M4kw2ldkp3SJAgVLFdGoYVS70AxpoR
/EqEQtbHfgNH83hatgFeScWAEwNHb4WrpI97y8pjYyvpCYNvvnMRUb0hNH2xTDwe
pkxilu+S6S7skshh4wncDLgVdA/Q4C2YerNfoFpznl2z1OrC5efTfjTF/JSyMGCM
dakN5TB3XmLet4cs2w1nNA5Lah9WB5+5csEXz8SLStNLOzscSVg06jeueaRiD2u9
lbXMi+JR3RfhRD6V7mkAExyBnSfaSoaUNCOIzW7Py7u4eLPK+mA62uWZz3lgGbfP
O6T+l+GH7WiD/xt5+ITvcy1u2P/C+NbITejEvIPVDzeQmz6K6r/xG6psOsyoqWuu
QXZm+TF3lL9mOsqBIXWTYdblO1Lvv1b/WKQdge4lEzA7pH955A3H2vC65cUK/yhj
BKXIxjU/Y2nlYQ2SMGz9IPdWKN0Bjl3Vu1p0QuIbdpoLM6o30v6WVqFnoqL3mksI
hP0p3rddApGiJ6hoHXki6WnMh6jluXBaB6MBOlvzPWwcoYEzEluZRzv3bWfbLB3b
ox2BfA80CKE32o6ybtFXS0Zd+jt+2tyhSW7xNSk7TFjXMCf4Ed6SZHtBXPPiBwyn
hVCUTLEZAiDw+o9X3g2PZ+0FPBQfB1r34gFvCljQdYS64fcsxyVjmilBUNywZJ6o
sOkHeMNaenYKFh4r0UzK6ZtopGh+RIHRGpz7YBIxMGqsUrra0V1UZjSwLlRXQkt6
/gjAseGB89hDepZ1aM4/L0Y3ibswjODLB8gFawKVZT2ZoXQltbkJBRoRsnRBrmTp
dAnM8mMbgh5bSBCOkDWWR5NJn2aMYLHUPSY/q1jDtJiqPgOMndbOCsTaUEhgbVvy
lmgRUKE5grhX5GRzF4Zx8L0AFnInwyR3s/j4rl+C+YE7buoCksm9TDmSQJqmJlgI
aJtM77PUYERY9hm5K5Q4J38oSzXKxioa8W5Ch8BpRvOSVX3ULz6oX41dEGXJp0VA
cFAUkvl4jIjUPliKuIwMdjYPYpMLv8yV6W8chXvSFDXh39xBx+bSBYOp5fIiyVNU
lvKWdw6nU+20wz72rncaniH8jO52PIG3pyvrZcJQFlTY1l9awmiQoSC+m5HVAQhj
9k32F1k5alQZNjPDQXoYOtMthc5o2KurvX566U6dyoHYnxLSica1TcCgY89K+858
j60dYit+RWVPUAWFLEV9nndQGt6BwbvE6UZ1qiNpjGxLIO4hB3nDbKCC3udkm2Rk
Da2JsJIT7TmW1MeSE1ThQfHBqaO90m4TLOUrt4A6QhYbMAt+M/TxT3e3any7KaXU
y5Fa8jtsjFUPpydljHAPCtthhAj6gOXpWv+VRK2hbTu4pDI8CaecACzjzTt/vEew
ut70CFfJxmUGmWC2jtkCZUpmD6vztUSVo7zRFykL3cjEjGJc4PGjdY6k8thzhORi
FgVte4UZilALnZkJtr0wVeqUOoxSVkm5EDoIcsnbLapTch3qPKHqLP1ffRrJ/Y7K
hVryNacKfSi2P9HQQZ5p9auxTRUjxi1XosycE3p2R8KauhbVxYspYWH2OHWtccNS
XWxcCXGQ9funss5ud0jGCi8QkBw+U4S3BnId7zPdSCG7d9I5TmTdA0T4Gyfg94Hx
LK7QK+/gVWpncrcsk0dVe2zaJcrQtZIc7n6ZhzVyEWtmKkcAjN+zWMBcNk2s7TC1
eB6NIXf0jT4FjZgpZqLqah0gKE0feM9rDWL508IZO6UAWTqSVTlkcLq54p1B/Lka
Jr8WFgFLxgkkqR4inQsOrE+m+yyXd6Fa2pPVFr00bMBhewXMg8PXULEEz6xKUkVR
Zk/DUkH5tithyl2lZSv0dxBaByeyM3+nbkmGxs9yWy2F5eoY+I3CgZgCzrFYpZ3i
od2AeK/S8lP5zjOCbPm69Wxvzh9GO5XlG282MfftPNlrrv5ZTlv6Tjm2/iB7Ejfd
DgN+cSkzfLw7E0XCrId4dnzp9iLvux9dVWCcI+l3Fznwd7o8tnCJWLh+8Dv5R0D+
S3vfXAlHJacASd9sTistCJ51rDFKt67txATIb5THDB72vjzyvE+vR+wH9y7ZxrPn
lDTAPVe85PV0njeJuncjlJ1qqeHqrYUWUaTFFzKvQ22dTh0HSs4fu7+hW+Haq7bd
jH50aoBascGl6An+Oz00XSRh2tx2d3v/5CEWHig/OJzekJf+OZ58Qfj3Mb3LlNmb
xXGOu8Sk2dzJHtXK7Smf3rfbTD1DT6wSVbH7Y+iVoV0iIauqPyry1fheOcPNkbYc
uSJAmDQWvf5h0xkun7PvEL8H40PEVJq6VBXJvH7dBF2Qr/YXJQODMlzij9qE0YCY
gytcrQKws87PAELGxoF8Jq8xlAftPwnkVkLQ1BIfg9f06FWw7+g5aT2fn1cKa6pm
N9Mz3xUeok62WSGXm9j2qqOvD6DYlwrGSkA3UdbmjzomAbAhJjecC1lr/aclGT2u
Of9sLFZGhidCQ8qf9jSwBItgeQ/FgrfDmYBkEaWiNNY5a8cP+DpcaI1zGlhwH+ZH
97syjicgavnbByMVMmDsaS0FkjswxiAzX7qc8IeAE2K52FjuNkipGGb5etjrXkbf
+zCCp50Mul/UljgJpOrKNm4jU8XEiBgeuS/kDYB+KKmioQI5WdG0Cts45A4SCzxi
aP0FnzcFVxzDJRprAI/Zyh81xE/2bK78JWf7lUJQoOTrxQQTVC4jAoshoUWorSrB
+5UICYi3g6P1CTlGE8SwKNrTRJmBtPQ2ZnGjtEOxTpuA4MPROePtl8ObuHaBFJkX
HYxxnmyORwdfKiRPQ0ZUzxcTn97G8mVHbvhA1NOEsu/OCJGQzjUow4TRrVDAE6Mb
AJBllENNRaOTe9I5900lU4L3yUW+CD5uQ8RH2lJCvBNreYozEQZ107o5l0TOu3a4
u3Dp0w6SuxpKxi07d15WhzMeFvcD49Z/GnVbfDgmw1YzV+CDO96eICLVXjYRVJ58
duoJzDEE4A1RgPlEGvTNhxpxVR1bFFDV9KQmAKVReH4SuNgR6zoLAwejcGkOf/bP
HhUH7Tr5R0WMsyTkOpW8dw==
`pragma protect end_protected
