// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t9WA2hlW/vcolCuK/qY7ioaykaIFlpwecU6pEnmdO9frSjpGfULKMDyo8pDnmr8q
olwsd1idWmi0906iF6utLbD9vKSY/QOm5gS5/GvIZAcElubhXl4kVOAm7v0deZu8
BfutRNVdBoyyxVdArFrCitr1cadDiNThCyaOcor9dWE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34128)
gZwOtsPioCaaeop76hzessygDK6iLMCEJcYva8mwdwK3w30f70dDY/VCgmJp9Mpi
7PQFKzsgxD7IwCrPpsa74IvOEJHlcUllpEQv7HWjEFrf8lUVlifetpD6UimKF7yt
i2XLiWQI9UV7DTFTnxmahFtswP1lRSvgDSIcquy/fZap+5z4Zg3P4ZKQMV8umbQB
Uu5xDevW59jO6csHUwiPuU/lR1Y94R+dfXshkhDIaDZFBhUdh5D/MfemfauCyDGw
nQLb106bxPkLV06gfHr/O9Au8M0E5iCQ9/+U9hzZf4YEIG0kY2dEAfvfd041i1Js
ooT8509rqx1HA+WE0pxGMGy7ykSra4Nk1GgYCYCsK7RiulalpOukxJWB3b2nENRJ
HevkD+2qtLUepIOOeaHO+4Z4QMCiRaRI6TQj5q4KVPVezxYU5490Pamxzq0b2lAr
dg7eorSEiSUCLdILL657tAKUmC6SHe0BCViNiUGzD279oLqZRry33DnsSYd6t+hT
sVRXdXCk6pb456rbLbLB75DlcB9PAu8QvEsRBKr5uUIY4SwJ506NUcNtrwsRGzbG
SzipsG4bSAR6jn5aQYghfwdPD7u1wzFF6FixPZfzl6Yg7Dr+EQe5OGdGcy8FZcue
URQREpEYD277c3fHJjCFVj+gTZKbqhr+sX8vXrYVk74SHvlaJlNIDiOdufFJ4XPg
vgYuQTwDCcNjb/0Gij4GKAlSQ24rJWExL9y8rtUMJF57AUTIrCPXyF9BE+QhA8Lo
2qN92yPSDLYUXKyDSERXc01z80VXOYOyo5Y2ReRitwid7fOSIR1r8EW7UXB+Vfyt
NlZwYE0Z5nebar5M+CM/vNOnlYUZkwffG0vSf/C1I6faWFbLh6leJ/IuzWPpJJzf
BoZfNqgViGwkF3s1gNc8nrwEg05eGbQ3ZGw6IXkdrK3fE7dmD6uz+ZVvW8u42uvJ
4PBjA5vATvgQC1HTV9472wL8TJcSO3iTS4+9kP6FbXgO3xPbhku8szvJTORL3sEs
SfJ+Co5KUv7U4zWnciqMpDw4LljGrJ6IExG8yhT8EqMtJaaUSWdAXDaBvRZ8mkMF
J1B2/XJEh9WFUsf8J5KMmbKp7+PThWhyLAopM2qSucNALWujlIHzlLmr+ClwvVuh
jbqHemHIrn9gmEwzJYEo55eWyMV4V7X/BLkEqEzJtfb1ENBhc/vU2mQr9OZQ1GtW
+/CwVbk+MvHHE0sYRSyIz9kiSw5tiFae5ACfegZtS2xp/NMOTBBct3GPHSOC00wX
FUBSBEAYWINv97X9eq2v9iHzg5lNsO+Q9CGmDxnrPE/EeoudsSqaIg+wnaizMJkg
+aq7hx3u8APQbWDN78qmee8Q7upHQDqoieaCNnyKKj24FmC8tCX8kilDST98C06n
jncqnqlCzYvMYXgCj72sCbyoQDI1uqJ33D2t/cR32wB3ppTID6I5fKYz/GdB+r1V
hJbUjtCdrC/Jk5ctjFqu95g0Qr+MdGJl6yTIuCHO3iraYHHDacG2oTh5bo3JbXko
ntIkwmvycKt0B6Qaj7IxL6VHEmO+TSupR0KIeR6qL46zkhgSK5GPdiGgpUA5/Ibz
iggl2yjQsze9ZE+7RpdI4/tadMUHZShyUTc1xdAGkS1B7oUhJt930C1qZVrs7V0n
3dU6SovUrigFgY0cm6DTd/72CLB3XVqnM847VxI2tb5HLwMCiCGThw4eRRtXXrlK
Yfb17Dq8BB4wCtqzlmd2VZi0VlBNg7ZthBsTBMtHEBvsH4BdHBMjpR0+s4iCUMp5
6MNT0HQvbxN/IOrGaMuNXS8/q2dFmKqvoGjhwNOHEnJUf3fPJKre3GgwB1oRU7Nq
uYmAEyJ8cvRZ+RctfeuGHc6q4bDxA0EUjk9qZAZdaxK6DjE44QZ2u1LFWmQb0u1Y
KXseKRXxJLdnJ9t94jgSgYBjtxw3yYOUBF5b38+8avjOEyvMuDLIzdRPrfbDEJRS
hWmbPBc8DN/Wq/LdEntkSc1whbCAfuEBquAdum5N4T5FDWjDg6poR111SIUsGSMI
hJL4rDMILtzfTrNtMnuAhIQCkr63sDKaEIGByRf/qT9dg9eANdFsna2/Mxdb7c/M
bjly/Gq101nkejfMktWl8At9sp1YWGNKMUELt9o45MGlfyPReJvQXS/7P/yxhnVK
yhLP1AlMPkengILT4Zeb+Gez0hz+Pp+nHIh7bipcaGNqiD7LdmwDlHOyFpoyqRQG
qned3BnuLMpoTlII5h7dMabDqgdut7IEzPQNGgTo0Dqt80APyLQ1k/lPR3kB5IlP
RX00OJLnDsACk/im2+C/ypMbJci0kj6bwWBId1Ix/CoD4oz/pw1tSPnxJa0ptA3H
fFHoQnfTiL1c0UANgvBI2VND9to7z4vGz31/AjTJ8+GC00YI0bEyuVYrZIcdY5i+
XDZ0gzoBxO/ZsH8fF2YGsepm51SeK0wzvP6Bh36y376GilGl7ON5sexNH0oBMIg/
RMTxZH5MDIgGlLloH1Ak/akJInF4urweMw90XIxRIDjR6CR9p16r9h6R9IxKzF4M
AytDwKFDLT1lM9rQ7YQ7aQmTHyYlBgeOHRKEK/5Cv9JIA/zuA60/2gfiGOmFpstw
eJ+DZV6UkfirxFjwrFVPXV1qE/NgnsDSlxZ6KJ8tTdn37Offx/XiI0FwnAa8JZmw
DH50gqKVPJaXuYni0kyOsdfPeXa8bxlOuO0ZZKLlxuK5JZwmjHsupBFn9xMNVgko
zfxRS5ennD4VhcHTs/H8j8r+vf2Fj1rHN7hokKA4xg2jAGKze0Abn0xeK3ZA2aFN
0HwPhrJ1W/NKosoUXTLpS3QYduP9OqKNz9gLJJrzEc/FntFWdWtF8YVn/pGiBclH
wuwliPgzWWh+8lqeHd6f0Kr9RQfv8XGGbi5zZqlrFK/3ul4cC4YgqWXZTs1ET0nG
Syw++8lGtYe9/UMfUnJ4o5HANns2AQEUDvUUterZLC0ZHJB4ln7mr+8RggKc9zwY
BNCF5I9ZZk4ikX/0FX4nqcz39h5icBfOhiQRGfM5i7tcXbTcC85xL88ivtYyFmxa
5jY+Vx5wyrlpoBxSFc962Qzny3voCSFiRM079eaVMZsX3jTdDd52ujTMNKXsqmu/
J4DHJ4WciqV4AstkqYdnDwmJjkkVMuqkguYI2JYdWOL7NIDSzeMYzq3t8BIvWSbU
S/W/bwYalCUIamYGHwTWbmSuKBAHK2vUCFJ5+lIeeCHrmu8MhIzSZ/7iYdBnwaGn
eUd7W/jRrpJSk6G5zVsBwjJ5Q6AlxCA19bmzVtXykCP0NlxUmNN9tmlMl3snfr/E
RbMriYtUx63ohmvFHKLShefiIY5LrywPkgrROL4tDb4fLzdfbecItDqN3g3ZIWNQ
0ykF8d7HOKsIAfb5WSvOyRLjLJVeeaQRscEUCKPuYaJq5pFyN74S8iK6neVkEWik
7L+vjawYSFUL6Ze3+fzjr0SvfcpoVMHEZEFZ99NoimGl28fm0XhVicTh7mbUHSPI
Var4dx7Bx6nm89bpNYFfmPEriIGzGr3tbVhwl6jo9LveN01yxmbzc8picUBY51R8
3guXUX4GmqMzG8oDyMFrwVWBz6Ck+lP5Uz6vLLHyMQFUEmM+9E9+MMMQ7bWK6ZZh
ipm/N+qEVdZMNI70pAFOswDZ8Z9y5fOVB1lucbEJNNJrPloXtsJGBUrXasAeC5w2
KXJtNescT6rrMKH+6HDWjj1PcPojvFjpgNvNPm4LsdR86Rd7XdTjgbUnO2Rnx46z
2ncpvL9BfGF8fCznvHnNTmz2gSZCZqhmoH2SuV9Y2akrsCeQ7BdbKGakgveY1jSd
HiadbeaKB3VLpzcFQ4pN/Jv7uLanTE2GYsApP0OI/eB7QbmR7QE62M+bPiyGX0VX
dYw+As069P/i07cBUX8z6OLfpftLJ4L1WMcnkOj4C+/Z/3vVLphna55/BB8oIG6n
K/1LcbaLkV3TCbLeumtpKrxZ5q/6yv0anB2NOFJduv1KpeXPi+qM6RuDCec+ENJy
PgtzHi7FMeWYWPm8f6bx12WLqVxF3wEE91UYZBvl5wuFiFUVRzK4WrsRth/biDPQ
xKGLqOaT49C0z+0ExNGB6uaEFIWKCHggpbOyo9kNNj1eDSaznLbXPMbadK6csSLt
8oCjvVBADV/yy6ArQNHTIwZLEY5joMrSwvHVXj9Vw7xv7JxuX/xEfql1bUppNIr0
f6VVwYVrRUbaYyZh0BtO3H5nGPtMbnH71yT9D/prne5QQlbxlJsklJU7bwBIz+Wv
6LiWk4CCVnUKTO2VSiMDIETKK33/bUJuPE86Yx0wCS6g38ztFZF+i5oEbmUEkHDl
D+xouzVHLbqHngktNnDxSLcykvyptCSFxn1XcwAuc/tCtWHuGZxWhVmIDsMiXyzi
NMSH12OK7ttVTVQAuJE38ifEgNS/Gx9j/5oyckslC4FtCfIIAy7CKljWWiG0uFDb
3Qdx2H5c5PxdQYLUmSgROsXe3bgVXMvv4FCgrc0RhxKO+mxkmW75VhNNv/5D7G/a
9ZrOG1+duTj3rgeo0gn3aAk50bQO2z5Lwvmnr/deXsWx8oMVRbMnkBY1BGpEyf5f
NASheCQTY69CNkSeGvGLPU6YECcB0BphmNCrT2CqRw/pkiWswgdFlKs0EEAwzVdT
/LB7CQtsm1VqF4Hzvv2f9A7tfAlyWEsQFgIhQ7ovMtJ3qkvoRwv2o7jKsAsjko79
aJzPJHWy1xWHeEaHxdmzkZhlapCj6eN4g4pNrU9WzdshMaLSgt/cDY0dqP78Slk9
6xLgSaBJ1yjhRrQHrOPmTtihh2Jy8b+9QuKVHABD43Sv8qpOQ05NVT8KFLEGUQf4
qVkDC5LwUy19+IYn7jV9P6kZNsUDeWDXHky7yXP0BUIY1rPiSIO2NlVAZBiHRngc
oOHGh/OvI+sWPovsUCxW/uo0jU6WcL2ZtlKNqfjEdaMaPwDV+k8XNLDZUm/I3Dfy
AQO/UL7dQUgO2Jp4SBDFnvRE+cCPnwkSP3m8AJKokgT5cpAPNfv8Nb0d+kUS/jtQ
NLLTJs7TuXvdFM9ovG0cyqDmOZoRwFfgwecfLKRkl2g17J5INmGBYkkQFOSnjc4P
JBtrNtWsP/pN4NB6ahuEdthGVcuWHB0dPxw5gPRMYP0VxYrT8uz34YliB9K9//DO
mYfAuJXqSmMwQIvVsBq73mpCtpWxUuugeXFMVyBjUquadz1sX5s8ouZnXusinWhb
54Yg9/YN2vhlQBoDROOlpnV858yii7m59NNmlydT1KR73WCS6d23fQTPadOtSrGC
4DhwYRLNg85dwz4o3cETbZsLgJEdtrAK27qaPLqQCnThXPHrKgp2aGmdxjZcqXmS
aDvoVduD7iCje7Pf9yAfRzevP6FGg5oFdMFP2SUgaoA89me7/YeX/mEQrW8wb+JI
LajKrYQsvrMxm8/VAwKQWWy5HNsC598OGx1xARcCKDiYCW67m1fw0Rej+I0nY5Jq
CqiS1EUoBTnvfTZ75KcL4e5+xF5FYiH7e0HOi5q5hViQmz36bLJMMgctnXEB9z/L
Uuxtxttz29/7rOwzot8upPIieJQJR20OVkXjpWTS7zSbkSRNx2tU2XiYClb9pfn/
Y/UWS5dGahM/Wzt+ZrHvv75XdJTlgPyiV0wdXsi8sib+oKiUP0HZnwEyKiJ7U08Z
cYqMD2gdBQSYlFzS0TWialVHWMNRlAI5q+7uBotylIxrQGQIIAR8qc6VNNmXJPVG
tCfUPDDBxGyCcaN5ANvUijgHCSWqveOe/6B0nfDjuB7q78M9qVampHy7SiErDkYu
Z8WR1+gs+CW8PpZcf7LUvXh5K4LaD1QKxcvmsm4FI8cjtAwFdEygl9N0n4xpIqaI
SQWHpeOrdH5Ma74sn+ZMMkADOumtcVPHwGjxzddVQfulroqdxt8snRppA+TRGf23
U+xfdPYZNNVNpNEusVMN1emMmzColkn5TvSBTAYWCbxFNrx5lvKTgREF+STwTavu
nhUW/SpqAAg7gmmNLa6mWszzhNPoSNfls5S78o/ZpX3XK7k3I72CjBm5wujlXv/z
KMz0i1Kj7h1hqaaECCU2+q7pt02xas7SxHPw8JgEKRzbmd8ZsRBIoisggO/XE4ub
beGWXJLbWKAg//hLuhrv8m/Xy14ObGbXwSykcbuD/K8l//eIByZa7uKs39UBhHYR
ZG5ubCvwxk0Ojk0jZ6reJW6h9jGGQzpQlZ+b7f0uNgODJncNizAR/0alkBnQHQrm
iiZ1NntYwQbEjHxw/iw/814UfR6AF41TCktD7lwgKK+y4JyFLWPk6qbuCXl33oFu
zJNiSQ/FRlsHFxppVxxnuYXRW7KlR5srMR0RXOQkrRWYOFI+757aFerY8kRpsa54
tO07/JoDfoPeSbQVT/9d7rzVrmdKAx5ut7t8LSx2gSdh3nmPI/+mF1NNyJedzPzj
ulah/MixUPvkgpJvlodQsWwHWXXYf0mZ8dVjc2DqVkeXS66hzYe9U89dIhVOHgxo
D9CUVArPXJ05GKbVFp3pNfsM4NEfMPN3lPmM1v6fDZ+lW34sdyS68W0aK5G2V9O7
YoJw3XTBQW6JbmVyNmiZr6D32u8Du4ilGh97NVZXe0oiNfuuFNDpsr6L/7BtkmEM
UJEcFNqJqvCltjx/2qkjNBEJ4pvdQhxLaIrhJdSIwRtu9+rYwVjm411p1L0sHZwL
q2Kqlsge+ai1Y5+FVRcv+5iT920nb37J4APfJQQTs1CWXVsMtGGedkABrdNjDJ0B
4gXhjeUkyuPUhI9yIZeqYL5iiNhVFQk5WrXepp6t2km/GkJKieKnpkU9w2qt560O
srWLi7AwLhKxIBt2AVnjI9VQPz9ANqrRErODZNz9LZ9kXZgW8UeVtFcjbIQBkdUz
rLZR2csDcR6hKbdRu3LwIecwp3/rJanPR8mi25+XVqtg0/xZZEEJTO7d3X92bojb
O70Tj8pW6VkVufd6QFtfrQmxM41XHlCZSRDhNtY43GsvTYSIjQEkPIyn3UoqfDfD
FeoRe+NgNaojvdUAIaOmxb22AP0lZohrRe6I1WR7nZvhxSj0MfOI0xFePBfoLwM0
umr52FK4q3Gf3Tc3ag//+7nqksNigJb/I9ui65dIjCoarTsDgMFS8COEPMfFu7Yc
NkGdy0JbKxvez0K/elrHMo1eHMS+rV5v9tD/Dedu+xk7paDMiw+RvAHjP088yoj5
eg3p7o5B3Ss62W3Tqrh7pKSgfTJBF2CMP4iex56OofTKG3gftE/HEUZS1uIB9BhW
CRHCNDHUJW6n0JTy1ofJJNLhgQtTxPkSJSQ5gqaJlMcjd2tHkRUDQ2dQaYoayZvY
SfXPzIQSzo5pcCkEbEMzOQCMq9fpNFhSWR16DNXs/WkONj/cv0SODdsDBe5hU/ZL
JSsSFgHDlCHX7l6dOLFXSew8wfpwrHncAPJUODvlTXZfwbcsoKaBKQb0xvaUmbqy
x+WAejEJ/z1UOUfxKM60koM4eGGDYFX1HFEZrooIHlxxHr6wh/aJSMx/zLYQcDGD
onKnFd/ZaF/JWFIOg9DJwLKZlFWj0VPfNxFQgoDLwGZBqVQMOAh3DpNBJwM8a7IP
f2K9uavXLBZTMP0mQCJe5LtAJI0rGS5SACgMHbii1IYPsGbhAQ7iOXHgLgDXRAE/
rZNsa89t1hKsuV3/BPo5HXaB79xb8pB59jC2VgnBR+lDiQDW/zoTWSMO8ksz8dn4
FHmsGYY7vX+SgvSIa8bTAyddHLNhmJ69g3dZTmgWQ//KJURsc4c4iwE4Q0qaGfAH
LrllZQb4FbXm1c5ttXOAjCVFzCIRzNbLdypvclZ725ZSQ0MZ9eOC1bEnQQj/Ke5q
IOek8VtNIsTuIb7X0bWuOKaaP/IYYDaqydh/0dFtnjwg+4zwYD1erKa3T0UoZ1sw
KKC2pjn7nuFgkUNX9yIUUbnD88NOvWCCXO6gsAt3q9t4fuRMDsNBJNvgCT5n++1K
sdM+epx30HqHpx1uEmUL0LBPFU+mwgY5dSFBqhe5tms4qjGqDF3Erzcn+y+Jl3KW
S89PG2OhCubOILsurwcZlGg/ZV2O+kBuyXFHPVD4L6WSjiku6//67+i1HZuqa/42
TjaxffeOd+RAVoVrwpFKTs18bR/pxcJVlVDGMw7ApJn6vaqxpZn+DhgwysMh2qPQ
5Cpavnp4O50AZhVJvFEkSCrn3MMCdhlhESeg0bDyFG8txNTEGRf2n7gXvqDL7jVX
2vzvXfisgxZhltbBPBJiCzzJMxC0KAnykc+nQix9ucXYyCHen9bb4IS3sZgCWz9E
P2jWrwR04X/BQHpCO1xPCordhhCmlhhEJpcGfoySHEgC6WzP0VW0/w12yrieDfla
UeqEP5SeYcYTLMXdWdb8duc7iqzgXu3QKHqCPg31+wZPtt3d8gAj9CPFxXIgfv9q
Vrc4G/yZevTn+lccCYsYZR9M3qb6Ow3pR/6ORdrhECOoqP2Rw5nG5Gb5NeCZy10o
ryzoBfvmFL7AZ4gWRIt5hMAzo/LEWytSG67ot/cfoP77LsLGY7H59N5u9NftTAe0
RsP1lKHX+GCYeSA0FldsZ1S45mHQ/+Isg4Af3jOOPg4ODiq5tvLnlT1uJ86gVpy6
36YdZgD12YE4ew/QyBWXsu07sETa9j7UBJjKNwrIDB5niKXpusFG7TAJSkB54IK9
e7AIxM3Vsi+E4PsHRNHec0mH6t2WSASyKoSdXcX+8P3SooLtZOnL2rB3Ksz8WjLZ
pAtD/2nnIWWxQ6O26HOVQt5F8iUqc3/PM/gkTUL5MO7RlpM6UhEx9vWaawuwnXte
3LlqVGD7YWU4MNeiCRAe0oPqdZjO8QX7EXgnMO5hxmWhP/alf1/gEG2Opabd/7qh
kiOc7l+C+JDrtksHwPWxI/BSecGL0Vr/OMYIrQpFJlJcopRxhCFOR9yZWNH2jmPR
dhIZ5l54Xw/LVUivI5VmIK2Ncm+RO/J948cK8V6Ryja/F4/WS+u62WBe6O8EYGfA
QqzC8zkvRPOQpC51SEQZAw7V2zP5HAC/pzw947PutbP0upqNHZS+B5KrOU3nLzO1
DfQKOxVT+MteIf2SssMvyPJUCZo+VgERUMlbnJFxuiH7Mm8e8nwe7Szm7BU2vY0T
Zxt11gn3HoC0DAJSbkYUNfhPnyKT8ECVfPAahy6xKw7n78nzfyYVi3T6lS25mAdr
WMwud4bx7zxZRZvkKNYV542M1Ec9RJYZ/MRxUIsdlSs8K20q8UhYEIwFmVUpA/zQ
jjm3SK5yV+a82qlVYickS18m4shTejtqeTqq0zyq0anrrKPzuq80STGqRpyFoK7h
8AKm2PzV5fJIfz2QaKWCHP5uEQEvi7JjkXeFPTNrdjtnyiqGdMpTpI/uGN1YdQyk
yNN6GdirxeHyxwc/IcIbpwvH7lwcgya0+oaqIXkMrTL6zdQ8+7HIvWA7PSzuOWwF
eJsBglNShtQJoFMJZaL0nv36qcQrgAEMxwEE8Knt3t6JsdgsDM9UydDmieJtnkwy
zBEO/UmGNMy0+16L14gd1MigY+65skRDe8VNr0LJRKV2vr8JyXBoZId9FvGiUD8P
bFU5aHQ3D2I4KXzaOCpjFQNpnGADC/wedMY7hspvdE1yFN49sUSKZvz2vzFghyyl
QTKADap1Eevq5Z+L/+Tf7I4CvN3ndYBktgQlbULNRJ7dVV2tRpamEtJ3iY8Er+GS
5b0wM+Cl29VM9es6RqQo294RepN/iMJx3GuSrNkoJgICQafrJC3TWgegrvqEunSx
9WmjL4vYxq/GhHp+mpDkud0wI2ukC18+LzBNoqi5Ydx2HdhbNl0pd+EQUs0Ozi4Q
PAWF0+0tobmUAEroIYrKCUoaMyCKDmBD1qyDDXvToVcqZuEi7HMzPxmKf96txc6B
nuHxFWdIRsquqSDG/0dE5QsI/vAYd7XSDRPFMHwm0r90w8X5+mmIsZ75vNsuKpTj
y2ZIMdpjouZbNs+fPvgLN/SYKJwNCw4qBcwvuE1dcXjDN9c7n3N5pE8PO5NPjpXy
ERGBfufka9MWwrZg7ur1mL8qOG/rzdKBEVNtrDt05kkM1IpYizK29mlbEC/FksYA
8mWzNGjzd8d2tc3CxMFExtZOvevRoymJ2p5n6mnKtMJEKmbt8oKnvBp43QSI40FR
9fOuFGtgh/dZF/462Sv2MDIqe2+gqx5z2uhk533/kxYIsKFtHS0s47Tz33EJg3RF
HnDFChv7B7TX03SsbMPWUajNGeBhbsesjMGGS844yWj6MR310FVZATWXfB+g5F69
Y+W6gIdV60eUurT6w5XCwC3JQDsLslc8v5VmRZ7+Zj4feVuUz0dobwNphVdP05kz
LdOo6Y0w4WV3jWkryb5oYnbnZG0DoeH4u2Re9yOPXGHsLZ6X3xS+c1Ofq9Rg2SlU
fvaOvx49KjFThVkUqNtcLUuMryVS0N9xnxEPcgR8A1c2scRgNZDMjEgDw8+JxM+q
Ac4d4FG3pQs5oThMr5AQSRI4aNVhIJF2r+FqQ3dJSiMd314hi6Zgfyb2ci1kqmc/
9KZNDGttx1NsB8uKvSwshWDbNGi+cZMZiU9A3R6vveO0V2pxaFhWWYni2S+QhNbS
o/VEssoWyO8Lf7QVw43wguvvRGrSayPikIrGKmrJhUOwfr4JnWcUUk6nvxWYC30J
3JXsopPQNc3wuY2iamxZE4emkZiG+tIIkT9kh1EJjnRxRzaB6ZqDdAknZqrJ0l3s
RpqYpBTriW7H3jxQZOVeFDMJoOG01Rg1V1KV5BPnPRoaPx6Qoxkg/qdvzDpBLohJ
PT+nHYHRab3hfg4jfkyfVKyG6V+MRO/zc8WKG/4G/d0LeI8Kc+FscsA9xt01xLY3
2zDKYAhqd8rXMjrfNaXXvYQXQ/aExeOplXNSPlMv2xIgwNw6SLUgCwwRmZ8Mag2e
sQbAOS3XEQ9vir2iWwbB/HKLEKvAsS2KOX73ybH+7GQQE4ghn9cCFX5oGZwlJ+sS
tC5G7jmPrNqOAhOX/BQkY4BbmIOcFWtSbGVYOl5ysxkEOa45VQQ/kp7Yi6syODcW
tHVvy/rNFI7sAysQ+SlTGHfqVIcnS+zGkd/EdxJF6daVv3e9RNltrmmU331avskF
USklQPuKeVBF22F6vqwzNNeLTjjd3qq8nwKz26nTDCtzgVtosmdtx3EcXFRuZ69G
sh84v8/8dFgVNVuqjjzlWNw5kiZkhWRC2bIdNPQ9qknKiE/geB597F5YnAXYD239
oOSnubq+Yjqz5unlkjvuLVdQujSH8jthZRLJEF3ZCAwrO6xeoQ187V0RUIZNyjWJ
wZP2nFIvYaIgxO8MT8JtzNPY2V79H+rfyFWP74Mxj+twrsHNmyyt07dE5IHSuoZb
eNDlrckuDIcS0+G1j6DP0Gjl0pB5w2pBewhw6G0hym00FmW9qijsLnbDhfziMtkD
PsehlZvt6uJml8tgZ30+Y81nl3UJCwtPx5KEb6NMLC2HuwIA0XxXDHzW8hKR/fff
ATKEH8xW9AhJClTLB18xHMt09CsFXRZPBThMtaj0owSKasH19rYVCP+/vjDwKgeJ
0QOPNMTfisKDd2ouDAfZk2YMU6N74MCTx16bzTnePdBHWHKPl3ikxhNKTjNsxZ/Z
foziRT9EOL4YuWBzR0FC60dXveoBq97aZCuBQF7uGDHglWh20EQvHam5sv+2TlRt
MTsY+2yDVb1MVGBxD9ymqaJfRFvWKvDkE+EMxrq+QfUjdT26eVqZy5RRQN2kMFHP
xZ4yNK/BA5UA9Kt68/w8K5/JrBYMTASdi5Qa23Pn1nvI0dgDk6ao+HXfPOtyav2Q
VRwV3SIyj1P+HlPRxuxT0NnNxkkVAKJxb00sl+bFAaYx1xVjDoXSbOj1MzpaFt1a
csTtAN8M1LFxEbXEskZzXAbfJeDEen/XEJSTAum59w4Q9iZoY7D/fEROChfL3fBU
U7d/o84npoCLEOaAd8R906hFV9SaPMsiZgCmi6kn1E7iDlRsHeoM89ATxgmrpzcI
+jmwDRlHv+iOdKeO2GQ+eyuKb+7/SdyQZOY42rGftaug6y0rnrUaQRus/wIQq+gX
PsaoVRjk1waPHBDVpPt7dOQRQ+CR0wnY8yoLXXUadoHJ4OgL7Hb6wfsubEpAqb0q
mp6OtVEPLOrYepDpo1uRK0uaiJp0at3+cMMjnPM1zNGyZqjO8OQNTUmorvR0w9uL
K4G+UzSNmxjzU3dHqrtXKq8WNXu6eDTXwzPa0jMI5crqWJVo5UVzRn9JAz2rc59r
tHce/jv0Utt/gMGb+quQ0ei8IzE5hv44bPHMfwOdTG1NxU3XYKONqW1JSc0g77NS
/psBqsvyZV0C3ZKMd1ZNI4prJGvyGtUYs5tNFUKDhkrxI/G5I8mpn8RgCQvZ3fHH
KhjR1qUAdjCEdIzQiRKe0Fd3V2ZEWKLCOOX5TiMJUqlolthKImy8q1yYEUSkOC5x
tYergx7yJKS4nzeOSJyKQhIBi4Y3cyiFWs3GvFjWYLHxU1cnRPIWgdbx3PPAcU1T
VXK1L33ZhojonDk9ZdxkGW1LCoeWbv0Yiv2PSgeN9VEndirt1LnEqHp4SQ8Sw4cZ
wAxhLlM5vKQCTHVq1WuoCD4N9uTfRtb75A1vFoNcw7NjZvVpfjRhwUvUQs2G/0fn
cK8HEZHSwRiVkDpBo+aQ8Wx+TftAPksSDOLxP1r5kdHhzHdKV0pwkHJWrfMJnLqG
KvNy+M0a+zd1ZD1c8NkKkRnP5MvPOspKSrzxsHASqcs8yUrOMOM+qtup0PrEI0YW
KJti34/V7SWfaN4owpLaSjrN5V7ShJ+a5/y6HshTwZPZ8aLvvID+XaI4USz9+Uy0
ozmFAltFW5IhRDJ+UtYhg2Miqt2xS80k8G0k0eaIsdkiu9KYhIxGyzyaTnAb67Fr
KRGYuDn/doorkwg2SnGQS9DEapVraKKiiiMpbpvs19Z93OlZcTRWE7uWV9H61Qu2
5271BWh/5AQiuyuqsZu6FQc1rgXIoISqTsjpLJDuMFDdNqwQ7o5ErbSMHUEeJ129
h1P8xSgoMy8p3UKZD0nD94s7x0zD3FCra2WbxS//Zb4CaWkNZOjfdWk7Kq94bycY
Bp6Xl8kN2DZIvz5te5J8CkJa2tbBhViIU0ec/AuBUy6iy5GiSANsCWEdLWqL8vJk
/HAn937FWNQNIcuO2TSYikUPFyZXyZbeQefKArkn8HeK1OGz/3JW6Od/uHi4gdxK
awvvk/C5YrCNIpghmryFos3AzWZrPa4SO+3qcYpncoR/en5pVAhTa+PClWRv75RG
z6kU9u9OqMPMz+Fk99Zr4UeCCVHXkfnHxDLnfOOuZ079qaqAt7rlEpjl0PDL1uV7
t2JJ7fXoJlsIUXwvs6SHvobBPyFd6/pV0u6CRN7RcumYRz5BFBL+DLNWuBdnvTaA
tOOFdhmrGis9EhrnSla1QA/j4a9f+on6gpDq5IXsMZIdjUME4ZMcEuLTw0DxTzYA
ndHJ6VYiddPhq5DeU+uoKKHs9w1GctwYinqY64HZ2GY4oJROAu4V0xNcbOv2umVO
KXJlFyaFGHK+4cTS+1Sp/abESi3zFAPamcWSekVmESEtca/aW/z218DvOiSLdM2s
pvevwG552NL6wvboGL10PMYv0W0NpnbyLZ0uJ+SlpOVT7AniiC7zsRE1ZW5eQ0JC
E1zXy9XdEZdzRqsmfzDlK88Vwzl4krPIfqnU4901twqXS1Rii/STAuKE4uJLXo/e
g1a4M7bz+JPpnIoA/WcpiLen9EtmlJ3ivLr3iv5jXQQTpRZlHIEcKQmkkSE2SLhu
qd1l2mhGgIPHT87VAw9zVWOPS8Y1VMjuzALuU11it9hIsvDIvChulIVahtfZW0+L
jvvA59QqPx7xwaOoCriyC2ST15CBd+mWcIsQz/IULspEt38MPXzKeMfoKPDYAhYT
YLLCQChlx3EMBdPRl9pWC8EtsRPT+VHjY2k+FrvUiO3vcUfwIE2AOoA1hD1E1YVN
3M0z3a8Gpw6mT268HZBGnvW0+AOGLg5F9n+VkcuZpRuMv/p0AeudYn6y+2EOARAQ
VewYl74mqhXYnJINJ7Asl5h5gWuurz2saE54yAr9FEO0jC4mYc88E/F6TzB8VgFu
v6hc3QPyGNN5N/rucPCTkUkpKA3tHlhZoPV7IHMjrfyYEsEtKPVQLdwclMEZOtKa
N1JOmIX23yGrnVpYNwwY17XZ8aXz/8zQEJShtDLjBkgJEM8QtHtdu+fIpFpm3ZKL
hw2vETYmfn5H0imuio4V+x74jXAEd4faRSA5ZlVv/BFMHkGc1AZal/KQDOk/C7bF
LVyDvP3l03eWSL9N/WKbwSCSx7YhzMufp7wqsdz1nFGdkYstGaAqlDFRmt42uMlb
yg6vZ9IgyGolybh9ZXG8qp/dK42F8Q+sDXe/ORYZ9zpqfCs+hnUT8lG9SL/pB752
q+mSuhuj/uLBeANrz+t3615cWODetQhk/rXFqpzoESyW47AqYVFkNvN1FkvVy7ye
yWYbYWIxdF9joohGiRfvIR6IH77GQ5j6+ouF/TCleT7Sovzz2pm8cdo+RhPGqcnj
S8yaViHxcEjvFwTSc5UWIJX9R3GJ3BXeGuLRmW1pTqvVtYcVwVM1l5/LrOIIDZk9
wjFDiwnBgGsuxYCSrNvtgXnbAVsPh2LWZZkWTM5uEz1yF82tELMA108QzcwTX9G6
WgONYbAzDyFppc3RZfsGcrmuiXALJPiHaEPSudiw8P58gbBG6du8d61hICBSjAT5
cUQv6h828KxnlbU478CzkjCccnoBV1naagHTyJgkWVRKuDvvj3df9RZ+hu+Kfpux
HhtQ6T2svWOVOPPNqFeyLXNZWYG5i9rfvbl3JsKs/V0Bdzyon00aFBXiWYwCK3N4
y+D1kWRW36W5J0QhBPdvEmD4BQFP/d6l7PmNWxXg0ilnWc8zqgu6AtvLcBMOSn0z
nTGwIdOmSwg9wzK9tu7UKcSG4V/fdlDK7lJaAla0cb5xWBCl8c9jYBBfBRxecmlA
HhO+xJeFl1mW87VF6iv51LTLlWmc7GzWWEAMk3AX0OXe9RtLRGjwqvUQ0/MifYVe
zBru4lXWk5a4dKTmePzPE7Vn6ZA4sRYriRHRuuwp5m3R/J0voAme1ofnDX6ESIgU
Gv9lpSG2DNL8zxLyaRlpnGrkD33ye+uo4zdNt4h6Ds4uisGtjBZVGaTMph7yxzlS
BBhgRQeH47UVJca/EiV0p6R02F80CGXOKnV3FN3Jnzz9p7O8x4kLwbnsj2BkLAgk
LS/IY9gNpdqOrUZViFBsK+oQRg+gj8mRdrJTzk3m+nY1Yb5rtY1aLNeXcsAIgoIu
cdAo0jak/VA3o+LxfpZsUd8gtKGEY/xzS+UjzcyGhNrySJ+lWWYMt5e1Zj8TtBnd
hJ2INbn5W/z9Noh3RJfR14euKQ9nKvOUfOHJmJaNXPB64zYxQhbNZtex2HKGECLb
H1cM4B1SFsr3cwKXahkfoVs20hBFMEl/QhDv0vjeLvjHtjST+yAiO0fgYpxBPpTQ
f1UG4jhfY7zk6w33KnVjWD8j2BptTpxsHy2mVKvoB0XGnaaXKMKdWpGrODhaxqoR
j3cHSRIaI8FR0jcdy3s6Q3/6bag5Fbx1bOxT8nZqJbDIDIThD2OgFZsTtDTSIx9d
H4pV4GOsFcMopeuCbMwxkNFsalVYVxGilX2HJSfi+5f/8cg1wTCBddVb16htgUEb
T7VaXIcMItI9dD8fGTqVnbXfGktikJ+pFjSxdXLttS7gbRqFG+p2gCtrSoiCZ/RA
2+N/WNLcYwujVbmQKcS2wE3AJejzIthaKlK8k44tlcWpLinST4/hAvFXBa2Oo2oZ
+X7k6tJI5ZlzwK++9IOSatoHKAWeZqgPHvKKBZKtuhCqCK7HFxa1JvC1VvxReidI
6NZe7hIAx0tAcYopzZjNgsCB3dtQqg/eUe9h4RFWzgpMkn1lU99j0QmbKJEyXeDb
uMxZvGq9vHk7KNUmYzrwluZIYqDZmj00z0EOClluwk1rWhI01jxfbFI/wAbG8yrt
EDMBhdcOpxmJzBzq4je6WnpYMvGZ3Tftuwe4uyGWn5tI8FEm+qrF7GWwxNe1AlER
DPy6GW7xHhFiGVkpCHVWd7ZheLQL97LYJx3JXzjWgqdyMhB+hYlFxDWuTj81qmwA
opOv5HfPEKwWQY1dVsd0gcZsXR/iYxWKkwpDiR5IsDmuFK8yK2Cz87e64c2GKoKf
krMc1FYXNTJT4enqScyU5Tmr291LVyTzq1zIhBNy0kauXHq8+0ebrDlWOlRp7WuG
+19SzcXAJuTBhFzDb4OlgqUpD09yczV4GwokFZ43vDCbkdsxDOP5XEvZly1C5Cen
MMKW7efL5YOj+HS+odf9ElM3yatxF9MJeoOmx04nvWY0E0kDuEM+qXuceJu3LWpr
brLAz+/xD3onNYpOPhFzeCBX4aBxLFaUP4NhqB6Vi+Ru3Cq15l3G+XdrkvxkJkcw
MIG9+BMC+XG1+FUM5f3CEQ3yK/Kpj1xY3w+118NKZSOOHnOaoxEHsXJQNEY9eBm9
qf0yeSsWALvtfQc/rQIzp/5OzhrfVi9stcvs86en7lBlcVPC/RdxNKo9QLr6dF3/
KMDCSIva8FGpiRuQyQke9y32OngOXmlH29lMQftCTGwdDNxCVoVnvHuqe8v2WBeL
RKRX3/9zjZQLXUva2EXGgyhqNrvhriCnDYZ/zXMIwEE65DPbSeblOen1cprvbXi1
NLbcJem9zvwPfrc540gXhfb1Q8oo9BldKhl/hMhIU5ESwmiVsxd9YBDFaJHxVnl8
NAdP9EOmgiiLZkVNTGFR5CFrtPUkKfsPgWZPUpUbgBOMnASfHP62cLmj/zKcsCLm
/EuWiywWRk2NkglKmuVBnGHfQNj5tYwoeEVTLUf+u7DYNa6MuVdWoQuPfTdtGWlL
CnE2DPClp9gcI4OalvtzLAQGv5NvzW7bfcNFiUyngJcGbAazHYtGU0faTAH9i75w
ia+RBPlSjmCPWWOUWudoD21RXcbYBu2PBkE60YxXgCTr5e1bspj613uk4DeM6AlH
DTy8sDjd0Grgj68ZtrPaH7Juh0nDpEtnRgMNV/EBkCt/jDfKQeaLNNJkmGKldyHU
vAPFZdI6p9P5ZTkykEyW1R4zk1hys2/VTx1Y8l2AcUHJdZvyFSXJDHjnsYx9huL4
+rj3niCFQt6ZqaD0lXty3VWAlCTVVpdSBdqqYMFfwCEXsGRxkD5z6O1WGVUJP4jq
TNqjkJYZKUyafW52JLlrG9c9UyEb+qHMwFN0aQZrcrq4c0nF0lpsVt+XkgtazHv6
7yqka/ROZXCKxzHaZzT66IBKMpmKFTGlZreamk99qvSpeefzKDpNMA3qwrqAI0/w
t9EWS9HmbvdHFe3EacVLcsw+8Q58YPLBc4Zg+SgkCYEF/l5JGvfX7h588taM1mKd
yAe3sJuPQZNp3vNTn0z9rg5OPgj/w3mrBL9hKS7VAsBucs0opd5OtcJiUbeWZWhz
1xH0m6L9uisd2j0hcfCE3mAZDTRFRO++S7tEdoB0Kgb2TeYrl8M4BJLW4taV/AJQ
CZs+S2NjZyeXYh4KGB4H4/TBTjWvbmbCxA1hbnFOPv7vrkWZNzCBcK0Ak8FmtllA
NnHEogaOe/iOtjCOy/TxJM5m2NvoTIx0/LhJ1UXcR7iTLb/qjHhZwGLCij9WMXGy
VhK9AoHsIHRIRuCiWFIm7XJsktIRPeAFitj2wvuOk2rfDSt24JQU+ZeSNGEiO3oo
3gmDeUtaEu5d2lu7Vjlbng/9VaOjH8CeeU7nl3vlK/GVCByzr+IEI7KqjVFSBv5m
hXvlS+K9ifdYPMdwOBwFioiTiyssTeIaz1Te8tuTM15Sy+/TeS+FddyF+nW1zsad
TqwWX9cD5QtrBQhMFBqDR68sWydYj4bVJ6sfKQnA3doeWQarIJmQd0gem8xt/bWw
/NmGzaMWhJ2D+oNM+tD6Xv6HoknwA3X3MgK23ID4M9HOVKa36jivQxGCV8U3NKqV
RVZnluy2JH3e61kNzrZgf9MHif2C5/DJXYW1IlvFdiDGHD1Vy36ItKOhUlUsXBPj
IDuFEgBfq+vWLBlWESCiMMo4dJ52lO9RReS/Ypfwz+ZK+UUKx/kvykSXimNv/Kj5
4RFz2eUoJRfG5YKpkHpfjWhmdLY5gKqu0z1rVg7icJNsxVktWyDu9ND3814ZxuCq
7I3i8azXE3SvnuGzEptaLe7YxYAtIgE36GO2vKM9ORT2SRtCik4wh/1FdN42J8xF
P8D8Itnxan+z6sg4HYrqdFD4nb/uAEomMekjFkCx32TkCmShdMHq0rt+o5F6L9ye
LGM+BybGOAts1IDN65+afgoDLx3F9k9KUr9UgecDyx0gY1HW2E2wODqjycIoTe5r
7XDBb/qC1kZTkYEA06wHHhbFaISxWMB/ABPtUCGwuAB3pWLymSOuVhC3t8Tl5gtO
txqC+NvKFeDk4c94ijhZL4G8p/sdW0Yij96GfYa6miW9h/w34s3NG3x0T7G+YvzB
x8oThhNyJmxTVU42Rt+e+Mka7zy44k0ciFzw0RsSLZ2JT3X+3FiuS+inRVXksmdS
SIAva7JPKsi5qpo/RsezkqCAW/51CvBxMmgOxANH5fEjd4g25RfWZBWAdfIhmtU5
JGjjPZFSx473a8m0IOAbrrrWDgju3hD2Myyfj8NdVGnM+hKNrvY43CKhBdKJxoNI
W7rnhFo/mRw6cepwhm67brTdGFtaSke/QBEmI9GpMkb2GqcEDmVx/zSCpV99mx98
3Z5B4gRYfsBGgQFzLXCbBqXKALGOxZoGU1HTpY9wPojCCX65JL17TQyigce2axK4
V2wHxC7LCAlf/vE8TsAx/tVbP4PdQItWN7tVGhNyU98w7NMNlxS71Yz9PTfD4JrF
bBe3rlrfutbw/0s05sjNpbX8mKYNrOfXB/b4K1ODbtYoX0817nmXSFkkERfbrcr7
LR161M5KRblkvbReO+eGqpkeq+95rdyx7MKQCZC1la78Kx2iSWjhzQl6mY2UOs6G
qjusbWpACzAbdkdxIFz4JD0s1xIc+TF0iAdgRAbl0jGKELU9PqXpxASCIpexWTHu
/eLtocuNHwx5Q1kn8h8Wp47ek3+UXuXsBNDJkf+YjsHV+mdeedoyIiypmXv2Ztv9
R9L+AkjoMxcildKDdluc9FJhfUg/Rop8DLLMsjzJ04idJTeTc5P/sJOgjbFSIzm/
2TGqt1yO7LnArjb+Fdh0uzTWFqW1ZUmF4h7EFOF0H2DN4TZhMpLsRMqeVCy/rUqs
yqI4rStp7YWlF59XpIukQ6STisTOGxg41/TuKailNUvzBRF7Og1wJn1zK1K/tcdR
gSV44SYfhisN4aVLbVRyMszXCE9irivf4XdxrP6SCVcM2PUzuVRQZCjFV/eqpiNH
6nMTOeHM0yhe4X81BRLKf+IsHmOv1+qVQNxH9rdSiY4RhDZ9dGZX3fVWHqpXvE28
ZlQ0BG8ZWn/IQzwWiqBLZGTllqrNEwvraSkke39v/VP5rdBK7VE2C0gz5nSX4s4E
syZpNUVBBmFGb4HeWHpaC+6VW2UiFhDo0Qbj7rSE1JCL+gR9+ADU5JugEEgpdBzj
VFCpSrHwmXEObqtQs8h8D/mVodhMKKvaLmVfgkEjk9Pnwu8rIEE+XMNggq5z0KnP
Kw0uT+8X+EWuuNTVFviTzVi/uxDeaxOxNso+PlSLvoTmBLuTnI3Kc8wjX5DkbBYj
im/iUPvu2FZQClPy5xO0uaqwDTyl06M1ytVPddSOx4I8coQbY4VrsST/332XPyWc
Tj/vvAlLbgAnGKEoL4tVy6bKh2j4/EeprKTv2mS2rpDNVYBK1oOA8I1DoOO0T8t8
Xtc5IsWP7uTnsShw5NbFFmiOqcfZtkVX4sjLeEmqDr23vAs/pF2T/e8NJ4F6qdfJ
tZw6IAhoBY0gO18FHzX9G8Wh0rnIL/zXeM2B7STbCFxNdi2vDX66B5IC+NSMxPTj
RPEXHsHdcHnKfcZ48Y7kdGsapnfaFEck8mzzrEsB5xwwkcqFqozK/vquS8zFvtUk
yHLxeIrnd5YhVAtQ96z9ahFjav6H3qcxiGSvEadVK5crcrATphuQxXh5Tvm7DLI9
bv4giViF0ceLev8BPm63t+BQ9NVemXDiRDHjt7kQoYTywte+0qcBLdQO3pf0pHP+
U1AhlSaimQIWQ59PaKERFxGYcvcPtQZMg4MMQhhPg57GKsgW0anS/KukDFUux8lE
Nb+ejdQnSHkbGLZ8Jydkx4Ny6CvlVMhPqskJs6VA+yvmDzUl94s/NC/71yjgKiu7
xTgzlmPDnmAXglMFk3tdbUkOJysqjkB50QX6GGwb8j1kylBx1Wv0LAmV/SmYRD/v
T1RlFspOAqSZKD5HYz7JAglobyG3gxdXsmr+Whd4gd6y5YV3hvTea0TiAGI4Ayjb
ZlhMzVFpoKg4eh5Ynwa4htewU4qhRjCsCygsL+pkp97+6r2hYew0Fx+DsaMHHO5Q
rC/dhL2vko7PPAJVjfGGxDNul/V+ZtlkDeZWKnVNLftz0fLvUvsK/fMMTpQqnYBo
uFXLdwkvOw3Aw2FWMl2cWL0wru7kTKgUnRLBeNvgOSnyKpM+U2IrYzswEDK9dAgz
YmZJoWQ6CsD6HWLvoVfrACnoFVM/oKf4M5839LQddRRQPna1VJTqPcComhFSmzA7
C/mDwcw/khLeL8+jZWNPBpz6Wz8E6pL8XufF7HtCp2G3PehJyRPa/aOpPQF+gPiY
qUnJtDj54IOaGJ8S/pKUDKQ4BnZ8jX2ZUYxSjXXqSbDcHZ8ag94bgqRCrrlDnzrO
oKUPLEZQtSZ3DHsLG1cRvPD56YUdESBKVAZq0VmRkh1hAOjqo35UG0nrKH784DMp
tcvRfnOMtgFV6iG5RP8KQ+aRAiNHYXmT821hJ3P9PyHIPUs2/OPpr5Xnq3Kx9R3L
PZJsaRj8W1HjffAG+WMyrolWw50IFCFW5tcHUHbZvWTGa0CIbrUp/OkLOQChJQkm
73E8LGsTzH8deZ1d/SV6XLBIRpfmL+qW7XjVHELBD5MScCdKAHOgcK+iKtWEy0UM
YmtT6SOILecDdYvPX0mU2kcN1UExVccSMWAdOM3hQKa7vdP/g74LggY3NAwcGl0y
yxz9cBbPIKUGjF6RZsWqii11nI84djhHJeDzkde3B4LevXjs2F8vC/5Cz5YZil7q
3SqhsNje8dLKV90N4NeHKCdY63ElZ9OaCkjh/2PJWJM7BZIMlvUqYAPHS5n4G1vm
ocQ3RwUW1g1AMZrq7egaaMX6ArWUfyc19sGbT+x/g4bUzFOmFJCv3kdBOD6nO9MR
k++xj45T8bYxcswGEG7vzaYp1ep3WDzqNC56bMs7HsnE0JR6Jlzg6e7aew9q+vVD
JO5ETZmw7Uaqeb8+mSgDimWdKeunwENLceXHrLOOsZsF4riAThaiMYTZIjRFiNfQ
VUC75gX5XB0WHByc5QIr2QepFqTnMsIEstuDv38WUwmGKusDIpn6Q38p0dXtk1X0
JQAtBcMUgpcP1JZg0K49bVgm57kAZwLv1csCh0KV+gWhz3pIZeUUS9X5sVzPmxyK
6Ls//qtWn5wEWzWImf5AtigPD6L8N9ixZWmQJMRLs0Ui2lkmX3+0XZ2uBabEsjJb
vNxiEVadq5TunxnfNdIiE40d0qIygL28nbFz4dZJQcrb+ny8swkQwBX5cNNnLfj5
kJmpL7xmLATst5Y1E++C3s3KGF39Y3LJD8wV/2EbmdoITe3KX05zpI96kNyW+6U4
im+4+PMkplDXr7rB74Y96rfEkKmY3oOL1FZiI4SmOkz2UPFLU1HyWZYVixSmoWB7
apx1+EheozdkyScbY9EeBCvaoL89sDuoMLET/dsFUFZzm2l2dHV3xfTJUCglnzgW
IQFV51BrTykicGxh64MXMSNZe4voLtmv7hrRxyyu4mGtaJlCW8iJqZxjGdL2OCWK
4yPRLH4m3+txE2ZAVtHeBlmTIIhiPdu8LOntQpMjzvVDEsz0ojWh/pJGw7qDuQO9
vbS1iBEE1Up6qXkvjW9izOmKnKZ+r6M9FYXuGakGtfl2vEhvIhbqtmvmzJq0Ocmj
yNG8g+rGHycRCrB+ROrBYG2zU4QxusIg0ANwZrwcau2tB1MFkPr5JD3Wn5k562n8
ACfqBXS1YNmvNLkL/LgawMetjl/dX1U9Alyuh7U4dc5V2Qtb8+nupxhdBPCvQAnc
DoQGQZPjBA//bGUXJt0BE6V0QtF5hUzvPM/9CDcEb/IQTuvDQVkNbUIyxuXDFxH5
CvaswukX0FbKP3/nNpyCzthJZsxWMayIcqaV9Tyx0fZBwG+MmDicdkO+axBGRLvc
GAACU1YnTLmZUfDsE648eV6DRj0DpjuRUsHgwbiJgwfj4mkIxDOHsKKLiypaMQGL
PgAEQ71tmmq2YzPKQLw4sOI3DbY5KkEYAqGznZV/iVyQgiuHEicK4YZ9Y9l4VcHM
qTQ2TNOGwTEcTD6yxbO+Bx4if4ehkXL+HessqZhRI2kfde1LTYMhfONqZu34c8Fu
hs7Vp/yMFYGd4+F7aREhkNenV8G4RfPIXgnJWFi3a96OzuSHpteb7Kn5GNTHG3Ki
F1gjlwXxphgtNGErz+XXON2Nx4GRkJ8ItJ83KCDB514VhJ0z0JDmvSNSg3rr/ury
c6lR0u5TOlKseLyrMuXPZgQvHSTkVfujXghpqVfqq40a1HhB1s4NVe93XUpkLwCk
M+ndp/eraPNfw6nxAm2ZmNTHF03mCl9ZIaopTlwuH/bH5/r/C2yjk82SFfRbfvCi
fR2cqzrb29ekKpyXItg5l/S6XCS4rZIPrC99PuiapA4iV1GAmbnDnRBRbTt5pv6w
XRUJVLNT0fzgtzHrth92ObvPFpZxxZ6wLScxwM+3ovAyXDbY9KrB+VHHr60FzsDs
rVtyprkGScjiYAioBM4cqK6SVPYpa8kL5s1asJZTekmOwpv3hUOA36QV2fprMIO9
Mb+rwoW+dGnnJ028lNPPA505PqYZKlToqxAU0Hud9X/Sgyp7XA9nCIav28j+z3SF
KO7WnWU3uRUxmhQVvlTqXYrewr7L1X40jzLTTPRnmOJtNSXccA0iuyYZ4SeMn++e
Des7H5GudWpmRhkcyoo30fq5XHSJxyUFE4uV1GOvoU/5ar4/OXfJBGkBTNtsxOKE
4kCkqVw5ifMM+VqsokVQ617Yu8KYAIxj/Sc9rSLRabARLQwTya3ukHFKyafQ+VkZ
d277Qq/JiaZqzOnTFRAkbBxoAh/3VYLwbGu/jc8NM5qBmYlNoKp3gcwS6nzYJ1FH
i8R+uYXXP1brFfZQ3p7QQLM0ffgPyY7XqgvUJRVCKuqj/CbotZfsPt6bHS0VWFWQ
WpJMULATLF8/71ZFj3wxzQLH5Y8QycEo7r71YgRWhKWTH0Av0lw4MI25+wKJlVlU
69DyLPYxmH1BH7zo4JTbzgfUeFjGD6hfNKQtYdl6gpM4V8Ixdj/U50yrpkBIUO4N
tXJDQfw9q/CseullZ92Xzn1I8RH/BtqIN4JIcBoZOJMBr8wZBa+jKikpWyPZ1r8p
WlzfAu/gi2+Uj3efLUWM0cP0CcFinoxsJKykxb3VuPt7kqOq9hJl1St14Jakntpc
52ZsTeZ/w9GF0GbbEQT/Twq4RQ7GtYatvX9JlIlEsE0BlMXXyk3RQ9YLLsKvGKIr
23Oiad5bl1Tgig5g0FvB63z4fhInvoxIc/8vnM5Y3sq3hML1bECxB7eTIorijPru
RHGy93cOBEQc3GtUEkdu5O7Enx2WyL7KJRY0HAeW0oFTbDmWLcKkEwaoCuXqcn3V
WYWc/ptphvyMhyzqLcjuv8+VWghplMIrRGoMleYYUWsmgfB65uieSDWvh7ZMhu9A
vj5N7LqhGuy+Eu3DM25q5668IMYnVXPCpV9b7EfHtyVD5DrEP8X11Bod5IARaNox
bjWxARdZHA0tNO01NQdRvLUeQizxf2KwaD7XHH8sJ33uDcUcqKSP0FtoNZ0F+q8m
cLmeN5FhXatn36XD5izoR5N2BifFQxgvS5ZsyPg8UGLu4+DvUWgxxMAtP+aAhIDq
f5e7tppo6Ba7INCH80SJqb15uvC/uNe55XE+qviduMn/WJM8YfubdZ3ehk0065L8
Cee98T8Qy2kIgtajWyEaLwzqGfLmALfYK2slFinXGsXWeOC+/JvT1GD7wtbGHAG+
FKTxXyuCEQjN0/AiMSc1vClQ93t8nHQDRXLhmNE2FUSOaprxFaNDqiN41R6usxDq
6HxpyfE/4FRVm/n6gO5Wp5qmiLhLcXzNkrftkG7d8CeJIa5EPd+3p6vwacOz/cu9
gB5Zs5n4iPyCJI7j1+hHH0ZnZIdD/rXSGzNxOp/KgT9d0LEzsaMoo0scHFK9St2O
jlWUsK7TkFvD/S5BXYfCbEEkCuiNT5wpX3yien9fs1idBR1CKWKwZBfl5M0BeVdj
gDXymtxykp/CQgQtXKV6BCCy927iMJifLIWwMi/WGgN/rlnY+aoZgm/nlKuxGuVZ
yiliT6D18Cy7ag30plehp2RqWf7I0uJvMBcVqvp+hNG+2XIeKYGy3C4aTu9kEe/a
99A4UERvVpvY2xXNedbDYMXNCohx0tasV/Eph6gxe5XLmC1PYwNUS60brtkL2qT/
WSm0Sdo94Mt5Rra5UtWq+INPHmg4XXnh9fDPOOgxF1XnFAX5iMIwAxWLnjnMf5l8
t8jFqJgx03jFQbhwvHhgZWRc7G+c7BmiJwh6KcWHOAIc1LOUs/U31JpXqb3vyaGG
9C5jpUw75czEJDkWywmGAvKc5gkjCbz7/g9L5987M4LaGRP0j28B06e/TcCElaaH
h0noJQqiPCLjZilJaB9dtX4Z77vDiRUiA7sEmW/MuzG7z+qFRjVVXtuYa0YMbYZA
yUjesqJXB0QCKxjQuHVjJlxJey+iNlvykR2zx1Y95m6DwCRSCUILScUuaXqWV9e8
eJcB7YykwF2OAx5DqyTi/2uWdATrEi4IJ/nZbRvvJFhz2KJo4zEaAfd8tg+pjqnw
uNKnyTuUDAnCIiZumdrcwbBwq8uaksEvHy1iARrI9k1jOOtD6zCg7mQ86RYoq5Ww
pSdpGbGvE+AugOflvIwksYzUTP4mVBOB0AYnGl3Mcny7JHZJ5Twy0LN2xfVmRRoV
qr3xVBYS4/HzOcot1jfgflHuVD9VUwCQJ75bynj1aKPClWfGVlTqvTAv9/4pjQzi
CSRucZBC3ktAJi+I2M3FtvZQ8rkeKmUNRIZKkhEFQtYkI/WX57tBh1MNZJjoCCGg
eSIbKTSf98XlXPsLCZrvo5YmSvxhZAR2e02iDej34p656NPoaHZefgjjF6cMNVpb
xlmuibjvp4v4h3uhYlEV2/kbJiBbgIFvP/d0KaviP5e2NnnuB7SkHQkG/7NX2PkH
JwU7CvyyHlowCHRP1vsQB72JcDJfucrZqKotsZu4X5HAD9SxvpCugU7LjJX7VGEX
oFLYjvtC3gmoclnDzur3yjewcYQpzU0F4ZXxE+oCaCEOa0lcsIL1SnJ6FSxu5AGg
uDbr7wr3MFUcLXg8+gVp6snjSg/dWzMwDKz6GVxFiR0b7vBv08BbKBSaN3OkkgIg
AbmfGN3KlSxyNXmod/7Ky4l/S6svcur7egRA/OQPKQmvvHTqe/aFBom5/cowKnFM
CVlAe6rNzSilTxARqrnAT71oeI0N+UVi33DpcaktGiFnsnCQzRSZZFreCOuXsYo/
Tl1puM2QtclK36FWgF8M0LSjziUSczXtYsZGV1FXQQDIaJ1uWPCALGS5r8IbNdyu
XaVCcyOmdK5kb9CjfCfXxmwOvQqqqEPRR1smOZcbspUJUJMuqrPW/kgENhh23AKU
kWrPP881wLRk4nZ0rr9GjpCgPSyL76QJhavGOPZIG7oSXResTQPohlANbVyAw6rq
pjl67fimzGdKOcOWP1wWeJ2ihhKd6DUiWTaGsz06eYtAdLvAefXJh2rShTZ4wn2r
aWtjMCL6KJ8XxAZH1aJ3zQSsTvbO2WXe8i94CV+VESg/A54Ze+oeavMCDVhuc1TB
Zh/E3fO7ROBr6ZscaKVVQU0+ETD1Z7arQcQJBKNLoTdgrR628gYqw6X/TRrhX5CU
CBJlvsupZXVf8+tIpIbgzL6qS7RQwj6RSpI0YL/TrFQu/Sff8dFwFn3Omm8OJBFq
428z/85wdoMAkU390t4t6B9CzBO4KuPtD52X/zNOWHzPA6qjH7C7WruROQtH1nmz
/pJgBCdWfjEHgETMVKwMzkG7Ung+ikz8ln9zeyBjp7nemrcbuviqWz3+G7n267uF
XrczMNzB+pZBYBTOod9FvzE3Z05JE/LVsCsOE+vydnQotZsFgwN/SZ+nVfDt3vL8
PyNFIFK9VjGZ7AioQI6eLFaPiAUmIGU+dwY38ySmukAMDuN6wjNvU5TZLzpKOY5E
TxFsBB2iW0TQRIcw8+8EmahMBvzyMCQZH07Y9LrMi2qL+T0sj/TxvbVcUSvOD6X6
5fRjhPHR1iextN+Mh5Lv0bGzMUrh3o5HtifpqmMaY81xLMNvkXGgVeioNWNPX3ZN
6dfaao5qadS/lJ+UZcJ62z3bnbKQM1aufTsv1CXKqykRZys7UzoXNK8jonjHWyPU
Cy8gYaQ/vrgEHMeeLTo48p41y6SpQ5XrMWOaeKhifkWMXirUqjcNzQ5pI0O0KHqG
8ELOtwqUdiucvZ5cCtdkkgGafRhp3SI6TQcnymDGWAxdpILuFPMQe7oWnD1tYVSf
yvvB+i2cOODS2s7cABKxIBXDRQIJmLl7Z0fFM5EJpIQzUXXQhGMyyAxoieMjXWMY
4K1BnUpaDJVTJutbB4OBwPynU3u/EUSDt4D7jbCiGmpZAcQcbXB0csgLB0UTrYfs
jH0bU8ApcXtxevpSvOriPeApAj9w+m6kTxt/ESWkskmlv9aLvl7/9D+3ZT3LANJk
9ldSXdLgBrb2PBfWTcumZG6CS4Y9QQAkIDYhB7B8cw6GYc4rqgj9kmgDw6fhdggy
myPz+KBZqRwLHNsXiCTBxBltAjD8HXLuiBVJcAtoWP54DkXSqSuPdO9Z/Ulkq8UJ
TvhU9+NtInKqHEYF8STVZXb6zyO0Gjvc9A6Nw1x6FAmVpmjeGps3wTRvdF6k1aFe
RRlTX3JbmuBX6G5c5nE9y0NzVuXIzEXe4+oLY51qKQf4twEk9VyG58A5zbxZP/sH
PsOR9hl0nrC0wlXZXEhOC0J2+8y15otfH3X5nxSogcJv+bCwmg/v1PJZwBnp7oJ8
FHevDhnYv7HGR37fRZFikuLnwxBcq7f9NIHBkPEFmqrMJz9Dxh+lnIGomqn2bb2L
DE5PVidrmeB01GRr2nX+qaxNyn8M5fXLvjfkxkRwbHfYLNw64l1xwRQ2DywT5UpW
00g6Ei9pYlCJUTNgxDbqqJMSpqylraibHuOx0ivwWApvDchNCGOt22sduYrMfVG7
j0P/enNBD4cUewBB1+0eDLgq/4D5b4+3Od5SGbv9equgiPM4lqopeHvRlxia+bIj
Guj6XNkCEeFQohHrTzvpYabvkZI/H14sN4+R2TnEXTDWHS8OtSCkv7AGmSCO4+Kk
ws572KJubw3Z92Vt5nIJZP1h/PtDgUtj+VK2LAU0Le0bztoz1CfPHGs6TsIVg1Sb
vt0S4PcSNca5wHl3gst519FyiQVKWJAE0+Wow/BLvkG99VUAGLOI27Ut7n3BwsU1
xSPIkZ+XZBPa7OjpjSUbW0+Akan+D0J09CvIdb4NQltKI7gxGvRU/EsrFGFtW6cY
7Jpsc/9qJfoXgnm7bPvC5rEVPByKUuViGkkQImSivTyYtNZg3thY/ej+JpF/sAkz
dn+KhM+ztPtR/S+sSTTJq32GlpJgzPugb2nhbKo0xTfNrmw0JeSf9VSA+mZM8jJ+
x83EfsYG8AxryBaSPD2jh6U1xzAtt6jAfoQlJblh3S6+BFfjzSirSrDvv0khBnZz
8sXP9Q+V5iOgfAUjsCxHkeZdffdKS02+L5wmaNYymRiX3esJP5v/CtBM+xY5KDHs
J3cZYLoSQ4UkLwI6n5EPxXKSdWBWa8ZIjPo8dttf90Y48zf5FXtjqzAHt6//Ciul
C5IczmUR8tZ1j5r0y5q/MzuyW1zub/VMlRPnHTaCFaRJl6byqyjh9NQbshDQUYMO
geIL0at3eIuiclgWrcOeF+1E+0ZvQ7Acq4G3j0lW1DpFBs9ojRFI//CaPxtm4jz4
G9GuDr/rCD9mncC7Ha8UJxA7soSS/UOHqcsEzlWgLhmLUwhmmBArMeHSQ0sYYXSL
Dlf6kQZmVCovn1qxS5DujMbATRh++A9+bKI/D3ClGO+iGm2s+n9e+DFOriUpb/ba
8iIvP+0rnPdfILaEanD4X+qG1rIBmFV9xM4LeAczlsvnVCjPgjyxk3rt03Xb4r6l
/x4svemOGJC+nOLYJpYcx2yrlXOaiXvYwyqvqfvu5tMud67GsnaDytiLSxMAe8m/
C0mvQVDanjg+u0/chZ4bZ4XR/7IelrIzFK5lyJQfMqFv3FQKoAo5v3ih+Nw6waMq
w+0J0lTjQ9KUup8vkxKMEaSLv5OacPJwfO6ibK8q2L3LnnOEDHOhgjCGLxAKGW6M
cwY/KvdS1cex7h9QsU+8KW5IInZ0b45+eL8r+Qxk0K1chH5guxkHSHOB0r1lxmeT
6wt4l0VdszNJc/fdAd9tIWzsnqEXeQezhy6tF2gnj6r9NE3MSS/Y/y9XqPq+rrEW
EZs87Aos8+6x2NSzZo8zA/LjbXUncEQfTHyERZp3RnS/1cyYPwjI4TXW0GtR3gP5
DuaLSkk+QwqdQYgaCVhP9sQK4HgbAwMOHLqmGpi/TD2QQoJajiZ6YtsWwIVKQb/G
C/k8D6aBFyFw8bnk65rVYZe3jdUVFdT66YXNh/irm4BZvD2+PlDeIYEJWPowqXo6
OLXF08zwly98NU/5z2lnuSOi3laQv0a64TDrS56jVP+2n2WScjYb3OQBh51kCVGs
KMmyYsK7sl6VXvh5i3v5ky0azyHeROVylX0R8WunE5mM/dCbXMMcbOLOPx60ee+y
HY/bvAubuVAGqm4FSHAmrV0yBDATGQWTG/YZvGmzEVRtt7W9Absz4384CvCPvt7e
ThofZItP9RqfK2VWV8Q3ZnpxvLO68c47uUdcrLQX+LVeRN0KZKcKLUO/YzYxVtdL
YgY58KtmtvNHTZA26JuvWJmrZUAvITEtpXI+teftofA4+KIui87cYk4XEEEFM1JA
jNHoyPyOxncIvF/HCDTVZ4akLQgXcnScEnqAEq+g++1oXC745fLJBffdw8rM7aHp
osBqGhBTt+8TROH4y8TxRJWxkianRoZwAnk0zG4yMOKEKsPTjg59IvTuKR87OPlx
5qKWifoINhj75Dc2oT5tV0vnyGv3pP/chzmpULSuTVvZ3HQhDVsxuPpIh+AnbTQV
lvMNccOc9PGKdICUKjAeALjwacXjeWLSAmHWujjWboiPz5w0/ZOPj6YaKPKSmJcc
Euh5nta22pjGPhvbffJv2Mxa9R7hsX3b/ae9X+uOY+LGWtaOrTDcclvyVqs0N6TE
xJ7Nen+9EFNzDy5Y3+cNHVA4vPD9V2Ys1NJuWBqLCux7BPGQmSMd4o1Bs2YA5d4G
1O27HphL4d5BvT/XDXOOWOtkT1CRV30SeCJTr7/WqeCEFdZrgMx8aoX3QIfV9KjG
BzuCDxa02qmic7DE/BxPSJNGXE76tkkNWwMcUAcy6+itToWMQN1dESHrvoH8GMx6
q4HTUwTB51ydTdHzat+hTiTqPUEc6aefrVO7/usi1O6iHh8HDht6pn+KTruI61jZ
LJ9jS6RC/jE+8FZiR+pPTH+8k94vkLTKKXS1Md8krXACBkUISydrAWD4f33Tp07h
XZJEenOG01Dsb2qzQWGFUjAepOvJJUHGqlyhMOX6pFyQ7xHql7HGMno/DHkBEyI9
g7W6fhBxuvmpgsTM2Pq67wCQZ2HnxWHqos/IkEmEgx/LwA5fkIu+RYlzT4TBz+sr
ZPfsd+zdH/rRbAkPWV1iNMDW72CKnBiLGh1uSzjUIs5RzXgH376nRz2w+4iZowup
Bx81yBtrIasOqbjLPpRlemxSrNbbhDENO0ae9ITYgrt29OlizsO6uFwk9IX1EST0
UYUmAYlrYqQQM1nMz7p8eW+jF/gkhKHwiRRMm45ugQmAs3U3Rou7tNgc0f/Pjbfm
1I/2TEChDd1/uNW8sr+/4JvsPCLCaxxuLPeRTss+JuRlnFQXIWDg2E0koRbSQlyp
OgM3DqorD8MZ4Q6S+Z1WUC7zcu/gLyO60SyM4kj6BjF5Lvk/spA5kVIaYHCt+JDn
CkRhhh6WKgySCONH/u/IoyDE07DfYWlsMSD8hu9e6axz/DOkga+TuRzizrkjB0XT
p9naCT6T6V5dHE9neZ4YG8oDczv6LjspbILTg83mlU/F/rYSbMF9dSeDP9jL+YAq
6NGIJ4Ivbngmj0et289gWb3M6NzgAmWTIQemDXYAgcyEZnuzUv2obCwUqBn2dahg
RXFNuGGHh58Mjl122dy4KYdbUbEJllTY+wgsLw42MuEglvPt1WiK0uuq4qXP0Xl/
k/qyCzZlocxqF2lzmSy3s+/+PbS2mXI5I7VDZNrNy+G6o9jabEaTzT/QI3xSVB3G
v9dsUhHiZGVtiv5PMibeGjmJNzN33fGgxcQ37os7GBS4apATSl2kzJvyLhRVdf0s
2FE8mpVAvETIps6TqmRTsRoAD5Wj0r1vPNyp5GVoQZq4eiMO4d4II4mKsxJWJL6D
WvintKUj6xekt8cXx+pwIpqYYij/iVf95UnLgZ7aVFrBSXBtuTPMlmqJbxQpQJ05
fMOzNFBrBW8thglnCdbDUxyVF0+2K8J6bjrbStULv3KDwwpO52kX2W6jXNixR1K5
MWhoksTXBApHP9XAKM9xelSPOwR6LKU+4ju7MKzfrvmOMLTv9yY5BVqBBvTnZkcV
tOnWDK1IGrQ58enVlTmvIz4NMHynBkPZgmO2UfyXrZYVHXIOnHVnOkkRwBEu5/Su
6APXmROZSrqiMGzqR1ra39zPDs1EOu4g61qBV2YW+V92i9LBNFS5jxQyxGg7A4Cr
cOuM/Wa7LfYawWkRJ+mCkNx+1Z7QrpBsmxT5s00jhX8wkmISgNQ3nz7TU74I2/fs
XZffwm7aYD5akw/VHHEZ38MPg31gqPHo3P2HS41DEmuMYYwAqEgog4jhPV9rwjHI
TlAKlPJHBE/ZNEJnuTLWTO7A1hAPpOMIq6SbBMnglWV/PBjuYxR55aATmo6g1Iwt
T9qEud8PW1AcYHYb8Lyls5J69FSx5wPrjp53OaPrcLbTBMLEbbwdkpCb4xRI68sw
/FLWddXmEMHpJKyTpOZ+qS60bDGSy+7QOUhZQVpleNBdgwb41TBUE+SackeMtW4c
emF4zvGu2vgOR0XCt0030nzC12rhSVdZmgyOOMrd00F+e+TqKbQ0/vhDctKECLZF
sV0021XgEVkqgkO1OFmLU3+luHPJajABEWvxuMvQbd/f5dzjEkbTfxnM3mtUPQB5
ewmHSS1UCfevhxRnZE236GZVXBaZr/CkT2ufPuaYYhQTEkbYjFHV7ntr9CU5ho8y
4Dz43PTwwxxpAGWUm0GHQCytfXikc3psREcvgwf4wsvDMP3VoWMe4f/82JceYeCo
PizLuyuUio3zdsplLxVkL0mdqoK0qbuqVeL/mAU+qt83GzfJ/iAQgItINQA0E0/7
un1t4tUpk1/VJxjH56imzTxh10rzNadIVbdwsvd+0+3/MK5fH55u1HlXMrml4CqG
PstOFPjdSpCzUL11g7xjPhNUEEWgl0yJu89vLpyiPNlsByeZZEVj6y88J9EEW1lZ
MMHOrCU9JAXdR4dtaZRDaDqHWL/gPe1/+iE+mQEc11iiro4UWZ8GfPUjf9T8Jmhd
aG3O1dmcNn8pDvEsmTdxSjpJX+rtxbsm2b5qd4/PzaH6G1pTYrLobUqzmAvOUjkR
ojIHIh+GJok43yS3HFNDVpmmSOTdgGUYYprE4smqz+v71knui7FQ/AmasJIPntBK
oF9QT+nwaLfQji9JMB6aEoEYPcU99ybFJeUPRtbvHv2XvPXy9+X2LfQn6sEDa8Dk
WIsMlGvbhpVh8vCKi7f0z28tRsKHZ7Mh8HNL6JaCf/T9j8jD48YZEgEqQTpiK5Gt
eteTKbjFW0VzFCRXPD5vpTPq81Aa/tZz18yD3eMEqhCea+kGw8qEhCTeyB2sTzij
JomllSe+n7PoGKGo2RwsD1ue230vV9CVSXAvoJO/wQD4RIqowb1YhkSp6cMzwubN
edbHaeKZ5Y/4fK9At1qRfdGxsEspBlhEBnOUc5dB+KZlajG+k+ENSV/BMJ+QF2pV
tlhxZK5r1nIq8cK4N5gZzqmAUYX2jUSASUv80J8tUBzlUCksuPS0FidxPiLkq90u
8q4WBIGTRSkKRaAYCdzL+2byPvzPvvzjdXUauldI0N4EIvlohlP8/BHTLKXuHLqv
9Wi/jD3OCI3hJJhv8hOWcsggndriYH5hBWda3TrzcckTuWaLzN+kqP2D1MIpAT52
zKAdveKT4DgY6F1fPf9sGXy13M8+oaJUBPqXOLS/hf1dRZpAKmtxFYeS/oHWBwVQ
FnMmItO+a0hIpV0b2WpNhuQ6GFNfDPmx2q3OR3bHkTimhnw5dSYn7a/vnhUamdEX
vnheLiEQVu/wdplI1ipXnIAp9X8DCtOnBTVGK1f+p/SFBcLNGoleaGcGDyHHgibb
Hnc0w5tiUnvfwn5+2FpPthW3vGvNqmlvfu+vMj9mhAsOS2SGCRrVy+226F9M+snl
YhIem1Cp9+BPRSXqSxGYXRMZredkOI1ABaz4kDcNqfAutXx2MVe8oSN/2Uhsmp8f
TM/QMCmvUoxm9Li9IuBYXgnvCdYO0VfJD+jXzn+gimPoW91tb9/eWo3KNMlq7J7A
RolTEfaVViUoXwqFH/kn01+zrC8BqFNeSTOd33s5hAvL3+CFXcLvgoGgsHl7tSLH
KOaOrlO8QIagtXbKIwccaZb5rJYpb1+vvnZOWD9CrKNMnLaf3azvmFqrfJsF8a7Y
uD0a9R9YQS8WbHCIKdtkFZFqK5a1Mr1q7fXU9LNgAMwNwYSjqoSzHpyk8eOyoTaD
mhAwm1lgG7vcjWY3coOoEkNlsLKbR02tMULQ+y0LCXymZzRX5kRuFEL9l1Uc6wQF
cCXytLB6dEu7QHaoY19OLnQnWyFs7vSS+KuW06gKWmswbXBBHwMfLZP6ygjbgl39
+jIDiCYRqNb1o7NiJjFtrEdOhPRCAX8p/QXo5Vz+9DgcVMq4oybIdl3Y/1NGwY3a
Q32aUPooMG5IhwDem3K3+d6WqM1+IdLkZDp1crLLZt3tbzk9Pa+6ixMNMjCKTgpG
sdnyMbtKDQBglCfmGCOINpqHYKM6fRsBFPHNCsCQHs2zsp7hmma3+CQI0g1VgOAB
bMkIWLVOfb6bXc5b4S6GvQDbIZwH9RovAa4smyoujYtnpCrO2TQlt0Adu0F6Z79B
ZXmtLt5j4hPeG1dgi7gmb1qUx7nJnieiTmrb1ooAtXNMq4FK01PZGNjNrmbLdwoi
cTAITLd3zP6qlTRgsJNUgDoXAOg3H/AqqLVwKypZert5jm67z10db2rzEaV4A76M
tWMBEx8x5WxDu2a0c9gfEhPPbm8wBM5R9vlsG8KFDBjWny0/sj7QUgxm7S1wHh9W
P03oihALOOxSXA3wfG20eNQEstApi0eWzCMDNzZ7zdNwJ9h/kr4zmsLTZ7i2EiKX
yD9fBSxTD6I+mRglDNy3ZH4LHmyVOPni9suNWcbhf4Z3u4FYED53lv6HV3upxoD+
I/YESJOz9Dd6b3TGV/wZjSAtB3lconoYpUq2XTA7AjqNpY2uvd20xdR+GgcMymzs
rkUbDqTux9BM/r3Q3MW9hbOEk44bknu1JoP4XtWHNKnet+NLxPwcyZXtDWzu/WYa
GvJgyCmiyT8J5H1zmmo39BTb0jtgqhO2lcV48fcFqMV3Ku4qS6IRFudj98n1jg88
Klm64ja69Y/iW4CQG073Iaa0AF4ePrtOxThymZmyDnkA9bnl0pwejU3nGlvqySBM
HkKYehhUaAPqyZvWffTyL6e9QTiyoXIYC+wDfrPfdTAozTLNgigF/t8ikJaEggJA
hdAijsf06dLo5YU6yuAlyk2vE5W7vc5DaBXPwlNNxZxGqFNVq3ua57sOL83dYH/4
X5O7yeAIEej7D2/0BaJ4+4kx13n7SvRQ5gArvRGeg6Te6VF5L8Q9ZNa2P6nGib0w
Nc4CG5AkFQb2WrIHVSbR4Ny90vA4C0wG/AwJ11qUjllLJH4Sy+qi98MHP4bu2Ffw
UjlvSxsoVdz0ENLtKVUYRKu+KIjZRe2kDAmzAPiFx5QMJcdolcuDx/tnjMAbioy3
lHLypBbiJSq0OEFr0HLFoB9LjQwzLZqpEZNoog85JQOqzbVp42/RL2/qLAkS+BBw
6dKoX+3pDYEnZlgKvRRt7DkJ1P77nVOjrDhsdS6S5lnYtoW275vQHHchqrIz4b4G
YO8QvDTmcvmhsU+goFjfFxOLhkDEEjbOWspW3qoGQP2yEEGkKSRkAdlYlLKrQDew
ZD0I+PMHeG5P305ZYYkCkY6yO1+70jFQYgW7VE1UcB5rW2PMwD5Ehk1F9fgMYqNU
5EXX3eRauH0svyZ1qp8URwj4QlBHp656D4iGjytqXdoR4ED+Tj+1k9zLvoi+7X3u
W40fgzVPbvq2oxHS5edIBKfssH29IK3MPsZ2w2rLda/zk/paatmzWXjZ+3j+CrTO
NmQLD/YeOPVaaAlSm7SU5U9xbmtHqvO8yVH1exuij7DRTHmlrv2amO/RSBJ6i85m
+1PXtI0KhP+0gzZpMZ5x/FsO9oX1sAl41TMQ8cgy/+PSP16MKtLKushdcGCKePml
vPpyOOPaZfjGZEIWTtaRe4GYPQfT0OjKiE3rKddt2trjARk8rfAK30SgkfpI0OqE
3W9uCUx417XKGjIMAv/dtZWrbZF/eKQFakqi4RdXLgmnBe4psFAlRZCPngVoVLeT
N1yjoNeE2guPN3VaXKsVYXL8n1SN7sMVpTFEAQZSAGfOO3AQYIv0KdK005iDXwPj
UFtG5sfFBX+Kqh20yh8eIpj10ZxH7twVjNhvtAlsN4Dv+rYwgIGtExW5WD9rLhQz
CqvQQDwLcAHMQnOgPs4TJfW0b4ZQOufvhzhQ5Rj8FW77sP8FA1FTS1Py2HoQ2/5P
rNRS0O3BcaEUeJ3W0LFMNljNYipOUu9FND4A5rqV+Y2rBt/aSO+c8AT7GIQ/Kqk6
wjDnJ5WK3ZYYzJUvXQfqX/fh1ESbG4EaR8fWOyU7ZDEkaoFv/RARqMYPjsoFOi9a
CCr0whvaAHOBsY+G9KPjAHJQXETd/MFTcNVkJI6Rgk28nZz3lehBMV65wNYDpHBT
mr/vaZ4TFeb9CAxOrPJmmm4xw/eIjfOsEvYP/ZFmTIdLQvODK1R+NEjaM0mfFxbY
T+qZ8O5EZ/QRqA/3zIrPuF2KDyxJh6JKH6JyvRfrSGZPoea7WX9nakBCrKgJfP/r
/QXQfTo6Zd5MsFRSb8tnPfMhUmcVenUnfkaWsYUWwIUfv+mIAgZroEqjvGL39S1X
dtvBLWiKmv0imvsw6Alni2FBn0zw6c9/PoXNSivFltFbCXAw6i1F/CC82ipZblPJ
QtsIXpwQVxT5Zf9IN+RFFwcd1y8ICu43nXalPFdVmxjpVhaHSrq8LNUBqxKPbI/L
yymgrQYEcyQnBg8dTsK2d7NKZhY6GtS8OqiLKcekLDp6jUl9Pyc9TsrVGQpbPZ5j
5/v9qAMmtvpwJ67JTVmRUfzX7dH1QDTiUilBi6YYXsCWNVz+6cPgqhq2Am57E43+
9KRJB0a7Zy0QH3eXEDEU4BMxJz/4j5VgGWDPSIJwn6Nab9s/nieQlOFDFW5Pa2pl
dmV+K+21MS3vT3z3BIQbD+Ei5/+ad9ABp72R/VewWik8kTh08T0T7RbEmozve/om
WtZbn/rRO32ZLiGchwncv4KAZ0m4p8c4Fdi1xR/PJHaGj/eL+4hqhs+PCzeCL3E4
ugj/xdszxpYwwNW32KLmXEmtIIPuAn2+ekr+HVkPp0QCDbYamjo1B42Y0RhX+2k9
i749vYc9dB5o6kwEyYzY2REaC86uVj5p6lZ7ksNFnGtr04/zcyeIJ70iOCNvOqYW
8AFcbQCbd0iEQA6gsuHldWR4aRooXNhQWNU4K/VglyiVeE7mselQvghSTE72qron
tddUl0X7BvNSb9Y6JXdEgSicCkEryYATjbGeNOTgMUD19UVrnNZfsol9KK/pbtWY
+9KKvHrVbbmKuz2GVitLLjLBfjrfQg5eiJdHmi8Nig8BJbzJZVfbS+Pu1CLtBask
xDllzOA7EapYT6xnLSZyXW/JSdQrHjEQ5irQsHlT9WzRmJnhiaWuBiEBrPRwTWaC
rOROoRXl2gzXhR3OysE5nU7DBIRUyLlbAqDS2bPm0vTPatWCJp91cSjF5vpDCaEM
ydAv3uf/EY2CsPaclyfHu2koeUxdynOMEclDcmulQQzmgM66onKNsoLiQcXRVMK3
vxKXOUd1EjH1vHkdpAr58UzF8skiwmDJCg4ItTgjxkBI29kYVryWfs26fJGE3JnI
WhlOCTZlDsyZTFrwO12Y1ZOhy+rGoVRkAm+MAOrkg8B4ypdqDa8cveXcZPcs+I3m
VxPwBZNZ01oXbwby+sPAE/G+ceBYuj9BoYHBKfuUagv2VTSEEOMCNsyVhUBoxXxg
ZuU3kvrGSpq/0xtlwN3G5MGr/cTtGnif8Zaj0az14AMMNWpBuKycR2r/+A3Eoejv
cK9D5+71QImp2WQgQFk7lb15ogCVdeLJdYbeO9m5qApwpMzFSO0elIWFy07Ce/5k
zCl+lJZefaLnbmuzZWdsm3ml0Qun3v5v5lsRH8oNvT+c/EuWUs8mVUvlCe93ABzJ
IPl81on2Bc5Vx7GwPMRcDf6wjH2NqtHcPAqadTH/eL2Y+rwMpcufZ0IvQHgJprdq
7yEckhSO1F3r/qYSS+JST6KV8H88UUs/KlvkpuNDSa0diuqGXAFm6wTQr1oRY+E6
+V6FoXPwP/8NWhUUom6SRd6WL1FIrIHfC0nf/B4LiKiXB1P7QH3KANwnT/ONGqV6
ifXDix5tNC2+zbXOVeKDLvbzN2ADwkpxZxevabpzBaxx8+XQD+xBGZSlDOFbEeTC
bLz/7UxVfjiZY3Z+99+Lxt/ekpDkiXFyzPj7PJf//COrczpcswOorf0vjW1ROf0Z
sCCuxE932VNpXGqwO5RdC9VE0dgqYS8pOBP15NMmZUmFw69d9cHQ9vo7qYQHvcC8
B96K/YOIp2qw949XWb5I1feV2rQPfVl9tgtp566hu2Kkv40GUGMnN/msUmF/t5cC
eqgfr1NujsdXnSMu8ARmQltwIvT7lnput77XgEHOEXAp6zgd9iF3ui3h3xgPWhAy
DkFIss/cr7JxJi0HcX1yEoDe/CTKDYl/fJXEnaKYUv7Kr7FZsO2WIjIJX9uHYH2f
PGdySoOYpL+So0/V8lxBNXGvmUp61FYlbBlmzyFj8tjpRB9IZBZ0za69qLu4ATQR
y44Vn9dkmO4UUkEI2aOzI77XOCEbFIN1skEuPo1FTT/DcFfwPAlqI8tdff/RB7A8
heW7PGbpbyuZbNAqgo30nh2qDAXXL7SLFUMt2rXedNbupM5K6+oYMCKmDVIINnQ5
M6v4YsudvY5QK3uSOuhkDI45FszR6vScTpomcH3B39TL543uEL/Ml2wmBa2khLEo
1BmwhXAz3qReuaiqPz7Kr0Hyx3c7t478zVKjlBYPDSGp+BPUlkPHCKBEikwIiXLs
4vmllKQE5fau94syEGOTvs9gRZBN6CvISYIBfM176nUCFUuyOJbFNmdnIewA3ISP
yLe91XPDuRU9gCJusFf1/BbR8ihEyfLkBUjsrbUwIvNrwC01rakLqf2o1sMaJMMa
kCqGO5kwB3DnacBjX58leIFo2nxfqB5fn4rQ368pdjytNn8IijsH6hiyexHP2FKA
4VmurgCI5if2lPKyLuoYx2J2rl3d0bAlvXlW5v1aDNnVv0Rg1YdWzBz668gV3IkG
lAHvpjnX4ctLEohMMiKKAEExPDL+EEzlEI0iSdrBObA3fHU2lT1NP/4iSWSG+cPZ
IgyFq1w6ttr4eQdpk5nmbZOly1r50V9bzFJmnTouojq8M0l04z7Vdc8cfddw6dxI
6UwjaKEUUt+PyYqQPeKvdg79nuvkVJA/IXogYTD3uzQsf5jJEwQTmXi4+4l/o+3x
Ftaw5CvnCurGpdu9iWx5cH0q5ddxaNoRrX/zwKqMR6wuKE1wjxMYd2rwXe1kw2ZY
+sHIUce+TRiXZNtC42g+uv3AaWPnj2SlBcRiScXnaaFchLfVRHN0j7vFtXmiyHhx
TqB6NpCcM6eaAhCo8uBDwyvZSz+RmqVaZcVhoKPhPBtD8KF5S2tPRtrmWeOnbfPc
NJMfTYVyL9RAdA94JlloXofALUsOuWltUDlIpT2guEHNi5xN9d/vMpaV1Qwe2fT5
9Lx6YxtN4RVrQl8V4JqdldV8YGag7MCWJABYc8soWM9KH0qBjcIAV6RuRF6+TtI7
+bJezSv2uWl3Jd71KzPegwh49Oyu/ey+Op6oMbkYb0e9w59c03Q+kY02rAIgehGG
OKmQkljMvz2yyjPs+oiHwcw5Cg8G5FnQ65R0rcSCUvBFMp9UaMzi+mn8uyjyke8e
Lr5eOp5/16CJYAS7NTL7TF+G9OQAICZ+zB50S1wF2qllyCSuaeZHmnPVWSn85DVF
gkVgdTPBVsmjeL/2mdMIS9g0oxPZNCgYTf1ydxuQ9EjX15lbQXKSlzCs9GCkpoYP
vTftz1oMEvkg/2orM9/hv7gyLEsdm6aLdvCzu6cvkgvwp014z4zIsz8nZk8qmnUi
YuytZuxY1zYbXLFRrwSx2sipo9cwmn3MPVmUD9JfcQZCczpkyylgQ/1p4lIfUr7i
vnEtZqg8pod+xJYo8701FyvAe4gkFWonRImtEFR1njEZxSbC+QFgPm2oXJBRp6z1
byTqtM+gy1baruq0n85YKtomrVhq2b4gh/ejOZcsPiKt7Z30WwdujLaYaILy9x/r
102o0vqfIB5PicNoKQYgmrMVU9sH+xBMbPiXzrcoV3+wjpvtM/o3tNoBTjvtWVGv
xb6P+lHF+C1iAr1KqNLt/JR+nf+S80O3Drx7blgAn3OVN8YTsVxasDwc3z9igUiu
uAcS+Fp3wtUisrUjaLumBN+n6CCVElPuBiNBRSb37IdsWfIzaBQicFiw8dPg3Gat
t1n1rRrKNhNFqtqgAmY7jEBRuSYdHctOGKf68b5V5tUMKky2zYHSjzJo5Rkq4xd9
Si9syzOYVnsFpX9P8NyUMrolGlQfAu8CspZKsE/5eRI7mQVMdu8GDS21TJfRfXjH
JJZlFyKQJtbN/FI1u8Me4N/phLkQ8NH0NnvtisLF2W1TtWznCZSZKcv5A07JTOYy
gDbpvPOjl29g0ic/xqTwa3YmVj/ANU/8F5X+9jdWDdZUx0T883k0hRmD6PC5qdLf
woqXBStbmeh+cWSxf8N2KQW65FMC1bUPOE6Yh+BqEa80KiKVjTDHKX9ilg1Ro1mE
5CvMbeyx0UgBK29T1fElBOv0TTQO37qq89gKXc7yE3SCC2XQ2RlX2nJQw2k42Kce
t8XS1w2o2jaUIT5SI+WVjJ11HY5J9nbO1+reHU8U+55s7wsPK4EIiSk2qEGS/z2N
4ZUki6zUQbLczCL3FgLwwF7qv1Zioh4PsRnqlBPV/z4Hpr/qPYfmQ+ugyCjmVonZ
0J8dFoBnuxydC18HE2VjYv73gyhbfiX6fnJPRnKOhYfP0pYIJk7WIFJJmmJ61/1z
Te5pIwSeQVkxBtx/gs291gKUP5y2fHeN6Yx7T5+/z75SB3cpVsyDp6Fmdz4ZT1to
oTuLSDvyr0b6VlHlR/F2JMA+5F7DAQSce92d0tiPi+v2+9dajts7qJ5ttelRHJ+G
vt9/+DXqYiPJvAySTc3AjqvHtEPAKwlUT1wcviTIPhlxz0y7bV2uTDUW0kQCkopY
zrfNA/Z08mVo38+NU2YdUNlgi/cq8oiODcLnomLNpfOSZ0PgwXXXGcRjCYJjFwWC
wa1cJq8MrPCSQnk4Unr3NgtC9dB01rORnYFYUExRLUzWZAZAVEtR1J5gDWXxZo61
IiSEhSriNTBfCM8HQoR4DSyAAsgrbfcJfviM1IYqaDzHuGX89fMZttET4vyBkFmp
zSbqONdYXoU0OkpkgaH/GkNn1Aiw2kRmaSUK00MK6znHalVf4qohVXO1J+hmays4
1bMyUUhHgeGx7mvpnEQkBaFhiqFfJURUYSGO7JEOEfYsGY4z8k7X2Yx+gkyX/rRY
Wqc2lP2SOr9f14z+yTNM3qnBGRzoyRwy3LjFL5hJOBwa9DeuMlNzbqeEadt9u3ud
nYiwNgb+xB9Pe7jwjV/3bLi1wmIlu90D8kmrm2jTmLB+S1s+VLu5uka6SIXyAOin
LwkBi2FJxKtfSqDKipI2nQv7led+YjO7OWVNVzaHjzkOPlm2WucLlx7z0vvVbXyC
pINaSdzeS50r1iXiPZwvut6wknWvLvBd93j7kXCffpA8C1qtCx+ctigI7vCA87jm
sifmhZjWEk5ygITYJO16nmYdJuoKnTocu3VySpGW09HRu2yj8vpqpu1BMAwzSCgA
IiwiNlHTizGZliurGvpl8DOub/9RFts1g+B7MwmVFv9cJsbi5Tj3UPTsP/9hMspn
eeZ+SyuawK+FO00h09idKz/jt15PYGyhRx8OaSIIHzngJsNZ/TKRUYd0eYKHHAOq
KqejbcmQ1QBrL1PComkq0DqfqiuvcsWC4fJbA62jh8KANEQCu/E3w3s/63OLTri+
KW/IAw8s8KGvfv2kie89+XYpXduiAYWBfqmzkrT872Xnwps+6ne1w0kRfWaV0Jpr
aKu604il9l1ooz0sAXuaXQCUREWpMZgaIH1bpDfqiUeS7YKMFlXdUqKD+srX9x8y
OkLaca1cIZ3GfGvzp7BzUF1tk4ZPh6QOdfJO1IxTiNUmIojydhInGCUnZPZoRMLd
z5IJcWrBLhr89J4rxwH0LRuwjbXkVUhEdE4oTTxJ4YdE1r+yqBnuqsVTkyk3J1zx
xe9ohmw45e3gZIChdIDqmTVQ3sJ9WGqBGkbpAlxIzWZFrvNcZS83UsHagBojHpzL
kjNL7NPxUdAX+VsPptb1osxKSptxN75GOqw1nxTxi55R/hr7sqRJqIcwWYcZyIWM
czDxeHhKjfO8nKBL4K9fe6Sx8bDoK41Bar9+i81uaNlnE0JgLmRrZsEZv3aVXwng
dQit90RjBTCQz4W4b+wQqTGdoguc+bbq12lCqUXww/d1B2hE0N57kAm+J2T6+87g
OAUqBt5jmEjzVorrto3Bjm1CbK6OMrfgylOqKbDo+pYjcH7oIaDsyIszTMtCIRKE
X9AVEKk/oqZfoET8dNi5HEGMfzgdpXBqeSdfC5l52TaqHDi8eO3cffxYtN0oXJ7N
CD1BGz8AiUB+fgLWGa911TTQyikELMq61UIpsbdOcEA2gKfPcUeU4xswfvBIycV2
ct12y8ddOBVWGxWO0o4FeW1z5L7UWmqFa3g86bl5Ad/AuHSOF947SPwsMtQ4ZMDG
OtWKU0JCp2ue2q2/LxniBEs51HQ2YgKV4ZmaK6JB+TudBRi+xE+HWMCGZFueDdEp
aB331Ne8veVYPz4Ty3BtAybQ/7JZFl0OGOpDEE+dQ/B+79SYzJRRPFaJyJyjc6DG
O95Lpy5wivTnKhRcbEl5EEOskFOiXGbdBB+E8ndXI4ujr1DGVNzRDkfINmvOjBIB
TlFWj2YdsDALhH35gzofl5fol27Sb8TBVG3d1MWiJfTCQZHXATeWH02FnN7iEbR3
zGHpj2EIbhZHrOL97IMqqA3EAjb1W6sfdcGufNCYiewndRIEiBJIByGPBNelLVKh
Ec2BfjdEj0+WvVsxv7HNpWhLvqdVcptimOB6xfC5nQsMYDWvHgfRK5f+2cRNTqoj
eiKFwok+OE3YncRlT9HSEseHGRCNvV0Y1Aj3N1lUIAXNOFMTI/gZ/pX9XJFFcUHM
q010qsKijdS6XdEQrO+1C3bieqH5MOBQbncftoBBvyb+Jdmtk9R4Dq+e6HELSwJ0
2sjFSDpBPVeYPhH/+Y1RcqdEiIyjOZJxyGm4ZLZbgySY98L+oJFhA6kPwt1vc23K
e8G+DTwvwObuN8x4/78xGIzA3zAFRBEcVzLbc73HUhTMp9IsSogLntRK8skVsQJv
5oRDLn+gvl2KG30uEZ2j1XtzdMYGYRRvKyK4RNLxsFgnvm4oLLYCEaKuRPnsD9/h
QgtUCgDpuoLtduuqReZ2ZybCFv9JTuD4FBL6+hOAmNhkTFTi/zCcdOplPQtK1lom
5c3PPIInWGX7z6nVga4WwQJ3uoq1NVPwujreeGt/Pwnt/it1EQC23ZmBtadO859Y
jbVu1hseLxjrC1c/yh4dN7bFtuqplj77BbFZlQHWG4rA1uZogovv5F0c6L4jIn3x
p5HVwJGF7HVgi+cJKIUwZvQ122oE/vQIhKJlOh66BT/ySdFazHmsX23dYsusDN7x
LgPjR62xZe47xHexGWEQyzv+3XmpOCbFwfrwqDUA+9CKsYBdU6rry6buGOg/pYlo
oPh2vNqaP6KzIbkYovOOKQy7RZaNfyiPKYpOjhkPfPzbNtJXaF3UgYWvXrGaWklk
aK56h1HrfqDSApPsHwZoAErm0LnZRz7mPX0KL4fnrIy44mWOBz40j10gAKLno2hn
9i6SqIIvnECHsNlz71RAQS9TsHbZVYr/d8gCgFG9VMtFUkxOj3YpmReMUZafZEjL
SmmjwB4NV8HsR5JSqFdnnzfL5VZolO/UEborXVVCmfmmXeJoHJ6WR2n0zzwpocH7
uGFFMhlm3dDB4exgaFpf1hZ8AWc/hON/8i4I+soGMOinXrw8m/9c0nmT7IPG6zTg
ojSgYrCFtWmgQjkX/6m7ERhOBp9IrHjuzSzZSw8fX/avxAul0LH/xJEihlml7IZk
zPu+jPa8IiOAb5yVz4K9Tu9Mp0LtKv2GT945/TrzjFLnPo0L6Yxn+o1b3/R9qX7k
+vjfL9XPAXYug56cAqKGcADdhHZ9SFbNE4DQjjTJfaM852dxIxwuHO45FQgaFnNo
nojtm7DFprtwtMHUzh1LfQ19gofZtoAwhJJj6qfGapL2z31S087JtjK05YEbMzll
bny8Ae+NZ6aluhRrg41sSKZCAMl7F1NwUawchYG0IsFLEl//gw9my+PJrtImE/yC
FZQv1UTRwXdC1+kHNXtGuQlUzF84Cl0Kzd5hgyRqOPHovkVeLpUnwSIkDzLdV+rv
eh2TDyhuL/DufWyH6/2q0q7WXZ/R4kKO8N+UUonoHpSkVkp0OmmWNeeS+tSGy7Rw
IlN0Jk65BAJZCRishEQRSYnqX+FHLYtKNNiUNJRpB+VDVGoTUqvUhWPcc+TpcJJS
37Ih3noFwuJzX8BNxjHfFpqJQZEYW4IbTqaOcduDTaFlfS15cIkM167tnpRcovYV
SYKCdkE7JEUZ8wqHNMUPgTiZBMAYhMAy/IPhPdHzAlkOzrMha8r/D/SscfVjaeC9
XDhgaVWZx2MIy1O6DZVlzSXIOh/y2hiuhlarPYWfdpD/lMPPcAJOEd9/fj+oJaYV
0PF/YNbQZZRSZZXx+0SVv0BN/T8gxZu1xNZVjEUI3CIZl3ymVXyrSw8ZJqA49q18
oA9JHClad0RBfLuSCXIjJNOpCA9b5NkMf+7BHBxFnibpbqiOSOY6rZDrbnspqqzi
/1YFG2E5WdSQXVnRKWivnFeXAKuKHpgnE1nPe4vs1lS6TtJBkYZd4hJpGh/mEk8R
v3Izf3RYudKmeCtW6j/Y3m+tXQCn5GIdPNOiWXWjnfjCezMOAWW1HsB9badZyudK
BOE3iM90J1hXtef0GoQxhpi63yIN8XBeHnZrRDUVlpXnphJ8sTRN39PXOBEOvt5C
8HqN+g+xHzDM6ESiondZfWM8Z7cuY99C8PfAaJfWUv5xae05iWlZMgdhip47pb3T
G8tNCPso1V0Z5gFbPmJHqjdadsxlI2zQyzm8vfdNOm5fbQQDXSOcSyX/PtFhSt9W
kIy5T4bKJJ5rb5UMc9vM+BgnT4TOBnaHvUvFpCtQMTVWW1gLLRtLh5OkUp6nXZUm
HQdRVFfTXlq15jhNXuHssIaGWAfCekj3TsF4ge7fCP7ADrESZP38UqjhQqtAxZ+W
UvUMRUAMfSMFQl4uMzIT6wo6SFjxz8Ym2pqBCdzA3hdl2R9kjVimz92+IMH9Rl+Z
G4wllS4HQauUmRNGMPEOEVUERq2L1033GyaGDLLd/pFhDISzaao/ypig73LPe6yx
vxdCUWGUxQ/m56xJ9GBg5SgydS+FNuDtOeBFrSXe68p7ftEhFeuIm6o6+zIlU9td
LcNX5A3EJx/s/VT289U+JV5FzTybrUPTJZlduWkzpSP9F/oZPRB1oTurNk//Dlj4
Xq9Lt328QkwDlH6SE5YJV1SuUprpWbKaAsHy001nXeFqse6wZPrTBUAQgB8QAEWJ
iYCeLu2eYAFu4DIJ5g2dSZrJkF42mb9QIPx3Er7zz2FvUNbQUBMH78W6NraNX4bG
gLXVj3gjytg+p/f/M1iCUWYwNMP4NF7o7Fq2Xxm/BKnggBgB8cRemZMZHg+STwvu
TEhcBoPB0oGEHbXxRz5wQFNEft6Pu8eji6I0KeSy+cKIBJoQ58yApQyIiskbLUVb
GZLKWQ/Lou6Sxc/DGM8axdv7E7+CuwVCTj/yVMAV34kN7HqCvUokod5/gNrVynes
hbWwQR+JvTp8JsI1nioBwaRfXPfBqe/lm6Y3h6CB40oTaITxDjZwph7Pk11JuPWn
AkX+jviWMk3aQnTH6kYlRyPFFTuF+2+pCc/oDnO3RhmRVAdoPrfyxAkSM9irxVza
UmwJS9KpbOCpbdXxbjlvriU/J+u1SSbmU1hFrENYe8oxK9sRFnyrnxTSBbUBzXjO
Ef9wJ5pmU2YiesDPZ5BeRjAIKBugfDxmUTjnK9V/IGrybkD8KFj3OS7LjjsCmDO5
JNxsvX5gh8USU/wZSJE8NQP5PLAvR8McH+VndkfK7qzsH86sgftoV2HM99C9pA6d
eQ+XG34wLagShN/aAbitC51CxAUzYbkDSanDpUgUA/HqSYkEZB1jj2z/cfdk1v5A
msKCqDnS3eoL5It/kqbiwA2jk6+s6VW445SuHFDv/gXPYkDcwt1zynRCvJROGc2r
K6nmdGga7ZUE1Q1SSlpXh89hH3PeP8IzREE1BlvSZYdE4NgA2+QGpw994/X7lzI1
`pragma protect end_protected
