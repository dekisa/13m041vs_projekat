
module system (
	clk_clk,
	reset_reset_n,
	select_export);	

	input		clk_clk;
	input		reset_reset_n;
	input		select_export;
endmodule
