// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:27 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QqYK2EL03/gio3jduKNi8t8NmwaasO2TiQnja5+vNVLw1amghxMqGCvRZNG82UpX
qU2cwr7aSxO5I5lJ4VvgK1dcSYpWzR3AKB/2BgxPX/MfVcY+DzpGNhGVws5gXBd4
MhX4OCz70ftbn4PgKSQc/puBsz4whpX8C0JlIP84cZY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30528)
lXaaQBVPax/vIK508kMBl/aRDxTcjfGij7PSo5U8lLMjUVs3M4uvQNhRjI3BjMiX
D+1OtHccoFgGUxk7ys/lR4wqp/lsHxR1OBLF3f9xS5oLzcnN8ODtcMCs0JMbx/yu
PZd9pYol9lzjRE9MjGq5ysVJCj913O1WPxPStymrhQEWV9e4FG4QbEC60r+/xSHG
BRP5kMIkKiGAonI/3XMpJYI8drvbx7kSiEA6QhBIteDzcYA8idMoyd7oW57p+Qsz
0x3WFhZrkoOx2UNIPaRo/6a1tvfB1vDd8SPDmG1T6RN6HtQt5ohdMnVSOiY4qulC
L8QPUNn8vkqdVxTy0pEnk9vVUa/zhGhAGZ6eSLGvzAQYBybGaHJMHrufsdqNMpB9
jQw++juOVQmPzymo6Fbg2QOMmupHywhJLWqYWRW6LqBBmiSKsTtgCyLwt/otYJwJ
5fcE+OiI1f9r/888UxsRPykrUmRUxT7O3gp0yFFoIM01QPP5a39L9v7HVAit26ko
32DKcyloMbT5wcQogGtYccCISIo2HOP9kcKLk69at00xquxrC/tIw9dUIbi5L/NI
cjIrtiqvRPKg1eixPLXBkflXy3vA1KVZlR4XzWFxRp5MsvFHmkO80QllFYVfudCr
ya11ESTgR2mMzCLypC7ioc5OShqQ+GTnbDYTh2pRPf6cEaw+ElIToF5Nn3O+MvJp
eo64Tbs2pievTAkH+0EA05CPsZnW/+rvXkf0W3KO13BE0trI2gmuuk3mvkRFJUzr
AiQyF0z4vRaUoW/UI20pStlNZA2QvzGM6sC4AwXi9HGYfUNIcKWlZnUmN45Xgr/E
7mD9mAPfSbZJX7+dKc69MCh73BetYLA65nVsxj1ffhZoNy97xmc9+Zikpjx6DEfl
PqihIJptCp2T1qTZSUDWxR8Sza+O0AKXvva4exDdYbdoALlf+8YRiRQQq1qR2Gtt
3ye9gYzsFeJjQaIkgKlEcLdW6OTHCz/AKKQe0nFU3ywONfdJRWcgH2GzuhrWjQCS
TH9WEgPQJyroZuHYeAnZG2wgI0eCF4brxvL5iI0FsqRqJjs4rJRg0AZWl3ODcJ1t
+19KCPcGOrdZuoOSZ+k+8Tp/7wYDqSwX6w/Z8ugHC+KWhV6uZWZ+Uq3F4yvysiAo
cRH5NrAcwxAP0Kr/FLR/W+bkeXCgxCAoQmjTgImlCVfpgUBcUYFukwGU16jHHNJ+
e/8wgMkaBj+/yd5/tQm7onoqj72VF/S5p2zCEYPR3lI0wXZPp800M+ZhyqigEBvJ
0QgTrvBXx16fAvfoX8CmoKSjH5X6vatvgwnsWoeiOBp/HXNFlyhgCl1RKzlYNvjV
CjMF85bJY7wSPYoYWYKE/WgfU3WT/VpeSL3diF6rdFooi+TQ/6CH+JE7PRoyMuby
cjwZu1cjg8tXeQjfLMoFxESd7mqvdc3avS2ahwlsP8w7cHIsyDaSYrScd+hAZPYZ
s2oI6dZfFXHIr46+VP3k2L9fq+QDhGP8mtsOMSiXvBGVFCgfuc1TxNFLbbowpMMR
4viOMztj6dZZKDV4EKwEgL9TuZ7U+ua1XRx4uvdF1O+PGR82DBDrtsyj+hIDLtDu
pAK/4q69az4S5+WLTHg9MUAXYU3Aw2hoUbcTc4s550MQn67CFkc6eHlSss7Qp3eb
NAVeGlSljmbxy4fT8aBSoq1jqJRfJpqbYRRDXgbuiYZheV6uBYO5qpuDxdiT+bF2
xLnkqsfUwCCJ4EzX86ctk2B5kCZUvxxcU3X+olOBWs/4o5DY0RkF0qnjvnbh2486
saIqaZX3JGCBNi203ZJzvSOC6k3THR80fl4tnOYHFnsk0UsYG/Vj78gcWdYlBj+Y
xAAo3I8VmFGGNZT0Ox6qhOhv04NqhWyY+seO6BGII25opdLf6OphbbhbzE1TFeFv
KhHXcyj/JPPQwxz7MfnXl+yTTRbrj/Jej7Ykh8m+ZOs7PlAOEEryn60LOL22ayeq
FyPqrlbHNS6ukA09IPkKgqHcXByc+mUo5eQ2PC3+QMqPGyc3ZDjd6USqDERqy1JQ
2oHwNiA/BdvPT5Wi9P8o6PnAL9JqinIL9K9BN9cJkKU9r4MBwBDVBuATqhdc7QH3
yT6lCaCrwxICVJ0NKEK8KlyjgtnbqSEkbmsIg3bUg4HiRNC+oMJRIshjoSpUgqMg
r0KuyBROV91vBofTr+0aRQbUe44nG1aIrEcnzY3vawLUOwD3RdcU5wOjKeIg6CI1
wftRJjkL467/NUe7HyD8ZOxzKiwqeogKra04Hyo/mLrCNhKo5JQCv0Zc66P5YLeX
FrDYdGKWhNIEDtmO+P3eG+/bbwe9F70G/FvtSK+EzugfnX4YFsOf8Ervanm9Kxgo
HudTToTMmMge9Cpden5u5Nt9ixNNlp1zN9kdym8XQid9eJDNXFt4Y/20lLUff/Pg
kl2A9exIiM0WQ1I4I4g6CtZ1ikX2El2YzmnCM4oz+wu/SbS8Je35Sw2q0AQ15iWG
/hcpuSNbijbysovxlwkOiCFgbTL4hMUw/F/cu+oFvkwLuldThwJJ2xXRI7+kABFa
n7GNLGHYaOySmB/fTObbyWRsI7t6G4MYFO0HBqJDo8wI7K0vRcdG1mBXueBKakmB
9zO1faIeit/h//Dd6tl0AfuV3040z6cq5n/vtvLQs66YIpfvq72Pg4YgOWWEkyyH
6a0JN21+shjEURUz7CawE0H4wglJRXMbyYTss1YerrBKjCUGfm5dT0l1dxXzgBqu
yMUrAcnXVxxi6fkvcZxYgObs7kq7YnxXAPMVcq9ZLqsxU40naiPuYckqBnv5v3Xy
ZAVA5lzY6c2UNtUvE62InKdJnRjhr3bDSoWhsaP0StxlVjpw2X7Z6+rIag1NXccC
vFQNvhywFGBDJSyWIBKhzgSiawcXFdf8eh1/IXi/8xp3wnPAa7tCYai1DLrBnenG
qGAC6pRehvpo9DwkV2oOlBvHXOl9nosfahgsxX5JcOaJDO7dJP3IDeJeSGvL2jOy
q4SHffyc4tCxUYqJMeqetTnH3wbny6QoexENbyQCUyj1d8lZvXGqLLoVpYF94KMz
QerT7BPHB4+v3HE0Vb4KiV44SRU/4uzxNbNuNcfZvfHQ/iVNeTSaaAIfk0HCH/YE
7Zk8yn1AgftcQ77ejjqsna2NeyCOXJEklPjWyy9je49atLQf4OvICIyMCi7Piv4p
fK76/ns1wFzX4WrQGGfaCeLyzXFIH5Gmm6rBztzY61lKGlSEqoP/hg/D1OyDWJNT
XOqbZPLoz3hDM69eymKZ4QEYT9+BMf8H5TvWAPYfAQIXl4MgYRImk8DD5FRq+sun
VLO38SxGlzuuzXcyE0TBvl7x1LrBewwCKLOGKyvmHMdCzdl90sFXaw5Chy/+arus
Ud+/kDlctdM5w6vWxn6Vr0DsxTofJ0QLwIxpsyZZR113JhAd9BzmBBOv8P/wzCAD
1RCuS0IO/Kvkkm8mldI1JaYYOZepOax9ZDdkPBD8+ZXmKdZD52CRKXsW8XfxZZnj
Hs8n61kUGlDmEQmi54aZ135GNUPCgwyi2/ge7MVn0WeVwnUsDlC+ER0weWrvzMWY
fYgN+OqOkMJzQsxCRQ+/LhISv3NBV+P2nniAkSTbkryCnFCEHFg5I3AbSHzIsbHY
0Q3smwiledwQOTGfaOI3frdo8Ec/y0M3DCexnpSkktjXQ2H56n1LmgN6epGFKSfd
hKn4BeJY9+weDi+W2fE182XWtZPqsj1IxsVtesouYcwExvtmSia3wCpq7A/jizti
yUM2Un4vSxNC+GqaWoERy+XLZgGNVujKMwprdos0lOO1lP4JWQAOUnBOS0AnMtsf
DtEW4AY1nIFr8gskRL2o7gbhHXAVIPY+QupHSyd3OwZiQYPJjqubseMZjFvjBHWK
8qOhDeYc037xBU388tDwH4gEv+/yA33qYONO6h8v1i6LyPHyyW0UTpXN8iqQ246+
6pkbzf3hc+6feOFsbzneVj2gavWnTf7x1chdWYIcKWMFmnCxLQlrsSzAZEB7K9Jt
IC7aKKl/Ckuls0dd3lGmhlrkXbQEvwJlQoLiAe/WLeYOR520CvneEZzhwtTpX1lu
YsMGRROsr4P4OBjt60Onox3WxowQaG4u4kQXprp5rDJs6euOmilVbAxNvovt2JQD
ZxmX1RT4znODHLA09x91hfQf4c+3qtrMe2pUXRJCevv77F1NBh/GoFhk2vSqScVp
9szA7kDllcaJvI4U0rZne4YnCEnkeE8KVZONMaX2GTEpsTTb8rV4twSwe+d51cXe
MW8XkS8BAvnuTK24pJRuV3qC5tEIBzQD1hv1DHiebZBAiTzR/RO/8jXks5NfRAOY
w+MdEp5M9YhtsuMcUAIMgqXEqibGCm/HUfcPiFGze8m//b21Xtd6oGC/3ygTl5oE
wgK9isL5bJ51xSTaVKx/4JhKENMLBNVAPXy/MQv5QhirG9K+pjk3lC8TaBKwhYd6
/SVAdKeU40BH6b0ql6kqakDDdLFF/i/m0/gGX4VFp9otOjWnccu8VSTfxdK317qX
F9J2hcCdhxdohbXPVg9x4yuTT1KpF9ZI1y0RA9asnqjaFkxeRh9cTI+DjdmPxSrf
nrxqFnKuGKhyXTiHSNfNl6hojuuZcm55UvRFrLixVPXkQm4GkntwHLDRgmJz/4V6
ZN52XioDTpUFppN+KwE5ZtIURCWyVu7oB1MVh8XNRN85GmDmB5eRZ1vmMVgXi6e3
tSPn2CUemwvaJvs/JXJetgzSM8fwBB4qsKamsAXXO+PTPXRbQQdcf8aOM20ZdRo8
CeMPQ2SatSVney2UYEKwr8IIDUfWvpgMeYMj/MfMfAb4TAOX6TCFPP6sjpFEshN6
fCyZHJ5byNEK42OBy/o/CeRS3ojOlBcU4A9AbjiancOpTMqTXQX/AVgXX7vXIH0U
vvk6lV231WyidlUuflV97cJrvsHFXnMMTF5fN5R+d3fK4REaurF+hC25IyRnFS1s
Yy/uffNTKJkXMA7BX9hBOyjr/kutBOBA923m4nZXAoi64/XX0pNBtyreCjK6jCBI
M5Pd4TQAthybxiKj+r9j49txf84L6KkCJzyY8Sv8+iIqddFolAN19HBX40/6neNE
6V54XV1pWFhl5IL4ra9P0zLmqe/Ugaij76WAx0jvB/RCn8hrWqWeQ69CcusT1hwB
qSX71VdzvZPZWYHICCle1OBvo61gr3XOCaeEMPfGwg8epz64b/wrZSyL2z1UvpUg
qIUKGq8k1szUznel4OswM9zACAhPwDLvBHT2nUTH4ybUn8bXnfS+qYm1fux/fy3H
LVEylo0DBSuvBu4F6D2yfGBSU39XNIrUyRYwuUZfVTBNd0qeqkqy3htbUd30uUpQ
0T/DobvX0sWWGiA75pR64t8S2AzT/XTUlofTfH+3jYhmLBDKMqisesML+dYzodXQ
gnctviXFhBfweIvfxQg5AHPU1Rncy0SkkuWo7XivTpIsTvF85Ja8gOV4lQ+MBzRh
trq7G2t1oc/9C0q/nTtvUlXV5szgYkj4uH96UTDK175//+f2veszrl8Az9DwYqdF
7ISWJrl1OkPWuQoA8tGOjAfsLfpUfOcJ6vaMcr9AL+rRNwDBhYKkITdplFvg4byG
ClWCnCkbVNeC3aKVOz69G32u2PCb8ydYSEVws/RtAwZADuq+IDvw8YChhlTLzMeT
SkrWgtGaGSgnhskD5fa7oefaTRNLFVMZypsOQZc2rHMKFCgssImNAu0IFJTwArXR
HgmqYROinr4jvGUHI+wpuB/L25KLRFxaxSooiCJIQrENSOEyPeSEOP5HRhabB/AT
OKLkhzUt0OtAIvrlXEAbLf93Tg0bjrYmAXDDgyDUcX+CXnkiaN9VK18n5XJBfFZv
hhFMNCG8mfEcMEeUV6JiYlQkD4gqT4N/rKobE3SgDcyhrSfw1TeoUvhWTOdBJXXW
0Q7MI0s3l9+LQ/vF+6Jo1bKhadA0R5bcNvi91X1RfcpAoAYkKipLlXiWyUrUmdeP
06AtD+SDIeO+jiRkRRmYn4FfY/KApAHetYR35lPXhEaH2eEvdIEo5hUK+4l1JCy7
RqPgKn6MKPEeo9UfeGuitKVKqlVnnbcTXKvYe9m5qZKvNlaryzY902bpwLSn8fwa
JAL3QH8TToODOZ+eOdYcsWtTQvfD2QSO+83b58O/wVzQtzC29auvBWICLisVNHIG
Ed9YknLJ4cvG5nPVTLNA4y0hgCAndxYohWp4rfbLo20q7qtYqozxlt7LdGjKj8nq
u/gMcrFTkJ4HhakLpH7LgjEgPMhHQ88MOId7EHgOR+DWa8RCA5WRlZ7q1MGQEGfV
Vrn3dbkrVk5zyeGUXbOuD60We1hVaW681kQqZ/Mo+bpMxPGfVLll3Z7o0vtBVzVH
rQqz1JPMI9cLwFP9YQQZWQgyiUJ80Ea69bxZiKA4CUNvRSaEhEzk0qH7Sqr9ryad
qpROfcOAIUclTQtd2YreRTjaPqjR98DDx2sc94ZDztO9CLdYlCR32WCktoF9D7sD
UTosRMbFufBLhuToKagF7xvFM0xv2p80+ZRb8WwPDfxtD91kPkO1nSu9bRXPjH+6
N5gw73c8p9cuY7J/W56/dEA4/RUwRCpoNAwoH6RG3ZhFK7g8ImB7zpsv4Sbkkzlu
JD9qpVFH8/cv25gFJDCWFbdr78qYzdylQdNvrn6mp0OGFuWaqUQY1Db5LLGwG1OM
ubp9VuZmSmuOmvEO8TXPE0xQRigH3cjojnkBLpRbKUKJhD+6B0c8gSpbUF8oXEH+
xzm0qz86EpFpF9kqcl8RGvjJEx3f+Tt40wrL54QzrAINJJIP/AfRw/NRBBS2b3Eb
uzlq0cXCLYIVFB6u3fWctgkgXH3BYOp+ySlvG9O/CFYImOdWZNsKWXiztm/whZ67
JvyybSJApBSo7Gz41aaPds07cqSBvuRPpdTu/8ToJM5jeGsqrD5uPdub1nS/ScV3
NbnNWRLaTmpbPrmfLq7JX/1Cz/HPCdEdQeW2WH5MAiMyY5UtwAUEtIQvs0Exzqfl
Z5WK7+9jbvdPbw7PH8fs77aUZTjUrHfxbAxSrcYufmll6c5ewiMgGSLhkwJ2AWwi
PsL5s3XXEf6eSNGRRYVGYXX/U1yVr4p74XyhMTgipUOZPKKotaf9+294VOl3n4S2
82sBeUKZ4+Iu3TUJz92+4jNkwI9qO32pyHsq180yB/L10KFcmsmg/a+LFX0Xb4M3
Yftmuj5p8QSJJv6+hQzLuCQ09JZVMlq59696jiuRukeRu/MORj4YVGvUqy6VdFu1
nhAejwzEK7NV2nsjcAKPUNwVUmvYg2DAy/gr4std/+3bM/H15uZU4ptyL5/C0h5Y
nvS22vGwPOHJw0XU6ajQiyX5KPSVo7oNuX/h35osRLlXIUsZGzOGGb8wT4AYxvRu
tKIH6BVTqMAyEaIIx0wqY+RsT+Jgd4Ti0V8U2E8NHqWqJ9we0KjZ4KQmnuwY3veC
2pUIm5edvikpMaKZbCa2peLj2XxIFWd+ge7q6uIKHXMV7/UbGeH9mKnDM+HnOJiG
jQuucrDeLYi/8PrZD3PrVOQI4ynh68v5h7zgzxd7Dp48PP4eTQGArQR0K1nBPd9i
kjFtcP8Egsk1CAr2IvVNHp/9S/J9LIv7fwFmxEVcXIPxpPw29u1cZZWsxd6N18OI
qHnE9/2CfMIdnC6GdxhGiB7TOpEGOS/EOzc69O6gLRHUL7YwSOdGud2QOsBlCFZW
xLueUKV7aM+saGOn0NH89/Shjr7Wq/sNnRkkHKFsV6I0e/A35P+D+ODtPF2CF9Z4
pR4EfZW2w/ghJndkFstXVvGhWSYlef1OKUWft2/CLdji4S/DmXVgRCTJxI40GlQI
VjcWMyLD9De8HwJJiG5V7e7+FfaF1ikpTQw7sz8XU6NxsmJDdRsWoJhhLipRPYSa
PT7OIuNSXCzk5b0Ngh882PpU5ekhgmhLftZlsThUJ7MvK96PuH3ckivkuW5vkvu7
TgIxEvP//XDd5Mi1xvPScthwyinOjIqAF1DB4zu58D1gI3g1/r4/ckFjKw+2U+5Z
emNVEAox9yXUsfo4U8pY8OCiMne2Cn5EpQ59nmMSvlFbD5rgNWDlQmZ1XUGAF28h
UydFs8DUXX6PFH7vuscbV3OPNyYQzKYJj3WXifJW1rNsfJUHvukie4uImH6adDzl
yZntKvedGYaCJMp43oJbzFyLznQeE88h80TgP8DGs6ZwRcqBixrN4Yg7kg2qM/hc
KRX2kztcLzNgD/Wpc6Axrlb/CC0QcASgNsixGsIckZpVpa8DAf3PkHwQdc5XQXgS
fTOg1qy+6BglZkFWS3dxaH490WWV80YAYXqeuPmPxzFd4vTckpldaJuG60AAZFI+
tEMY0YAPziaayEOxiOw3uJfUAWEL2A0CYiqbETlj89c02j3+nyr4jrg6L/zEudzt
jWZxLjx4kqQKmIfZWbSw51vGH1cg2wwCYTtW2xDvqGXAYXMPcK6F9Atq+sxaaBxn
Ul9DA8KewwNcKvrRYxhfFUN0O9pwns9ZqQ9LJ9PRtdUrAD0Yo6aGc8nk01C0m1tr
H6HvIsirmdMm6FEW2uqtOzInnsiVW94D5Eb5FhhEcvIp4EgoZMPaOPrNAjwyTgUD
LX0HMk0GvqUNvJn9OuRtg95UB5jRv5pIZiLczZvtztjiJNcJO5wgqHIrNJ6N8RYk
By+AHNASOiEpHkuQu/Z2wdVLK27+0wjgiWepQz62zNO7Xk5wxF8gZ1+FXWGlStck
bY7FONU8qtuZAW66lBJ9j3I6WChSt1acGwLKqzRJ3fzsvsv5qLSrwVo1SvGpzpVg
NkcmwtYTV8Z5N5SQ6KFEmNqZpnhs+h1pqycXy6ov0N6KT0Su6mXNzKntcKgjcxGK
rU+3+r01Uy2X28T2qy0t+Fo2esn8ypnyFTt8cXGxITHIyro+PYHMvZ3u9G69q3Ys
YwvLMwrVlNTeL3zcUKJMcJG1YUIdPOAu4FrQXatuHVYdTARPZEoX35g7Wm/nZZIo
JcJx8gksPFHZwpn1f3Tw3l28Zgdqs7ztOxOlS0z8meC7vCJ+ePgwH96BZu5Ox6Td
CbCOGb3ckxGj8l0mLsSJf3sWwq+hOcSBP3npf5gnEfUnwCR99swXyzPi+CkcOBZa
G6+pZE2NRdya9bEk9/fr3Q2l20SuNjr0ZQlLruuKqxutLLxadRtxNMplLn+f3Rb8
prWpOiBsxMVussnVFnyKy5qRx69buobWHyjOT9PON4IQB+M3P4497eofYMoDJBzM
Q6PqjJeMWJiGurhVHF4V45rm6Gq2ATfDB2BPXiU7Fe+PG+EGjr8+eAh5ls7Cmzn6
ZKP8nsvRovTqKDgUfQ5rtAZ+DdPmMuyQTYwOjQ469hj77w+fiUQgg3xdwqD08mde
/mGVyJqj/lkUjYFro3zBg1POF9eyVsJ8nJo56FxwWouyLFDVGKehy2s/UKeHwOOv
vmYm4cvkwgDfZKvHZ/MfAPMH81/vsdPkIncBUJ/JQKW8SGae9hcvVaA7bIK12oIP
0amNO5lDQkZUCnpu2uzCqyoMcjBc1XBqQNAESC4IYfu8E/wySNlsZyV3lOnNCXRV
g8mGidAkgg9WznCI34mBTWRzEfNhIQuk52g7jHh3lr9If1kzUbanQOjndSZow7r8
MpxL4Gc8+lg+sMKslrJ8hsRhOrravNymRAfABxIBzzzVvzgyqwzecjapRjtF+Oo+
ZnybD6BfBH5jkplM6yoSduEegj26Mkbkg62AXO6aeBlGaUWz4R7j9LKNDYrgyZ8k
ySkzQ1YkA6wALYijot5MIuYBZ72Pw0Sz72d0AhOnugnmi4l77gRqLiZVQ9PpNQ3Q
0+ERIPt49L/8JHDruBrclE1ytAEOsTiwx/7Yprubp0T6npBVI+frZhNg4E2pBsoi
e5/R7dmpKUGYfp+l+gTzFV8FDshwj1FTeqOaJ5EjBb1N6sQX2xzbuE+KslnKcUXY
5NxvDHk250e2z5ShewebPTt1OUi6kKZmpv7TcCzUMjjBx2eR/eL2nFIWRDj6HM+j
1DaxyRLSNLIXj2fvJbgRlBAz9NPyARIuVd7HxmYqp0XCDndcU4xX6P570q/RVYzi
EuVbuwJTyZ6RDcV/cqunN0tLyNq/UbzUzDmde1a+QJjcWMCa5R7La8gc7JLVOtIS
5Lr1Z6Bm3+zDdZir7QNQXv6FhWhj3c9Inl/xO93FEK/USew3tLWkm1Do1GHRvgXc
DqoTPd8fKixP3IPgLFurGEyGfSwh/GK3mdBBN+01hnUwKJ75WnomUDfZaBVBvUCD
/JmzpN2PHpXQX2WpexH4GugzZqZ7ldjnQ5lOdjUwBWeBZJjlL6Lb8YpFvS6TR9cK
BgcRZBUWYo/3alO3fhCvXijf8bsKZv68+ik4OcawR6rv2c2qZkQTV06VBdpF1B6D
aQXCoAI5wKTdy0rAMlmNyX+Alim/SeoeR29jD0GjEGnYt6Jc53MvtjSWw28ZLosZ
LhAYhIKdEyamHpLwVLFSTEMiuPv9prdDZguXe6DQHV1n1iqGgP7QwT5qXnbDd0KU
sNo+XHKepIjXbXK5RwwXPDZEQlNGbfbSNz84wE+KdHvY1bJVeJq/Y6t+YbnTbSzq
0zNI3sopPolwxcCm5I5srsj6n5AwDqHSvCMyTaF2bkwziTYBZSxAiLCEaa6sdNYx
9RGMBXHD0Qki8dr8vXX6eM1V+JpGNUQKDvJ35fkQGZzCIy+NE1LQQ7ztTfHfU4y1
vHzUyC+UuUhn5u+k11Xp9rBCRAK/YCxdoXYDt020Qu/80yupWbrjgfXM1KsLhOb6
zAQuo196SnNODnQ6+Ma6WhitnWCC3abw6M0+rm9KPYwAg7zksTyNMVr+VkaNpLi6
bbyRrOp5fwxNevbUuPX0sz32wrBVWAsIgkd8vZeRE81jY8X2Md9KabkE1tgubQkj
1xRkHFjOnAXwj9YDN6T9b1Z3P42CpcLnBFu6vSw+R3L9/QWif3NDSBA9tLU2YGL/
+XOhuDWMhNSD0uQ+O1/WGwRzk+99puRiaN8PgVKr74uoxHC8axCapMsTn95IXbxX
virjbROienBq6N4fuxgZFzL90urOJ5o1WUCGdluGftFm7GaXCv+vMo6GnVmaBWz6
/Y3Id09oYRTB190pBntAeuSiy1gOk5XT+ixXXuQUUNeaf6/0it5VkHpOBZFAntyH
Y1gDPhvn/eW4tfyLcFEcualrOjzdKZRQKzIvtuRuN9LksiHrc0IkkfgQigXJdkfd
aOD6iGQvSe3Z18KSdIgj1T0m3Frwhmt/khhUle1DDkn4jb3nPbeZErZotQPG0tJu
h1Cyym0kEZcHugPPusUT2MP0wccBqquS6gaMcQXcQye50uTCCCOEAUUD3NnyWpSi
ij59/Y/jmCTUhcBeiWjC5PXk4cG5gtMAnoH42T7k1CZrD0c/LI/Si2Vqk6/+FZJd
1ERbxMY0FTlFm0ZIG98fTsyCCsw/iSm05cbBuu4b9TbcUfBvuJLNkngVNYoXmpZs
VetDJpgj65orCqNZ89FP3Rj2pLtQSWH5JKNW2mNlhVxt7+ROvnvega/WfPgtrblM
s8cwGhyBtyw13aQyd92aG5llEQXlo3osZtohv8IojVIDJ21enBWxFwUYeQX3lvXG
SYvWvFRLNyEaBIWlCZUMZM+Jnsv5Dex/szQ6iLhWNc+/3voNnWfUf4VufUw8Cl71
e35qzINdZsuWQF0Iz5FhWdatlCTntz+7nlwLT3+WQQ3R2dEy7wrRyAaMf/Qk5aYz
6Qa1kX9EMxL1n5rFJkI45nXV22x804mI41J6Zpl7FlU2bEUyq80Sf6tQvOu50Qzu
YD4KZBxqgW/2p28PtVZizrXHA13GUZaBZlWsUynucRvst1gyxgS+YvC9QJso4RxF
so+xSNc7o1LXeNFXJMhimYQAOKy57VevKQ8zk5NpLnS2vOMVjKqkhC6fRmM3g2ts
7Bi5ZkBPPNIMCaZV2lslsXwWdN1+HG3F6ad8xInTFB0832A+D1Uwv3zYSCQFjqSc
0mZvy7Koa4qw05OPpkMYMn6dmu8PS3xaOovu0aC0t2h584v5zJ4+rggB1s+xcWKB
uwcC84tQtg/suy9D9llv+CeJXYC5LDQZaOUUK6sFT8/TQ1B8AHixGf00iTNln6C0
2X1QHj+pQyramJKYEZsxO9itYXajhNyhQYqt0QEYCgzmBaabl74NDr6SI8dpezvT
yeXF8T9M4XD+A8hhasQMK2+tDzpXKm1UUjQbtsKw0OCJlaZK598DZy5PZLLsmcv0
AnON9RYeb2RQRcNQTg+/7l/OGRaJ6x0I7ZeLto5aTXJUkRdQIx48A0k06wadPPag
+4KZScRp8yI59EW7V/ZQV+gt5kcEm/PiVMMgcldJ/zO5jiHVpYPjzBX88SWcPHt/
jR4gynMLt1b+pq2RV0wrplxJZiQdS/kawPIy26+TEqbln36HnSNKw6Sl3kjGJBNn
W8dQTZuMo9vsZfTq1XqbVx2XoeO5p5tKBHFQ5vJgKsAI9hueSzb0lrwRp1Xune32
Di/zsMBwYoKMk0AL/eyBAviaCwwU7OqHqVbiEvqsIEduVfYXgTqN20wq1QF02oQv
CPw7HJIgtATfe3NLzQq1JOPz93+QlGnuGOQvMfI2Y2Xe/CUAZyKn491fWxtwBq+/
UBDMGCZ5A3nfy+GJ3LUIxEHaYczBCI0+fcOQnvh6qIBYKTxIPvsJCIggE/Avh1Ox
Gc8GPsE92hCrw4FMM3Bv19JXuJWYRnRzUFGiPIZ4UoevR1nLzSEVB4O2BprX29bp
kCHDm0dtGt2dKHydtxHUMgsQzrMDy1EVVLt4vpPZJLWCMcSf+vU1CT4+D81pkV8P
JzEC7oN5Zx7Wljc2/nlmsV/OEtl4mMAvw4S4ww3VLRzCjcrvdw8ovEE2ptm4RSn2
aEI+QLqWDSTPTv1b5wgu9h9TPdHheh3LW+Hhs8AGPqvYF4M8OJhgxiRjS4L87e0Q
rqlxCixaNCENT1M7b88qPF24PBCZ1QjfcMdFFf1MQz/WTgPKl1Z7ujU9wo72j3Zg
sfKxjU5bbAY86q/tC95+YB3TF8LJlogHvBO+gmhbS3ivAU4rcYy9HrMYRXNav/K0
eSaDOQIJwe+1eJWruFD0+43ECnmrd0eBelXEVgmxss7FBrziMMD5LqJzcX5jQ0p/
Ew8ovhOYCrYM391nkV5M2WOQ3Fn+HEhKn/KVGWtoYZuOhbn1AfH/2sAnzDqt/p+X
ccT55HS1P1ce5BHUVoYOk9pukwXn449VUiaCwysZlUjjJ5h2XZ/Ut6K//JHyedil
5nSqiAO7hvUaaNapBspvL9jmAtpCLlwix0juyTv68OnUbydIh9jyKKwy9qfLU3DP
Ks1xvRFLiVfoM1gQElufb2ec2DkJnXjItQ/gk1aiKHC82U09H0YN7lr7yg3/oVwX
37HszUgHham5E/8r2rzhUkIgm+9NwmNzfstrWAutqhME/l6XplWf/bDTAFmPjJbj
pS8lA+X7TcdssJAvDA/xNlqe2lmDoi7g0wj4bIhWrAmycWAcPuknI+MFRv1gLoAX
g4narP6rUAqwf1znxxgsm5UKIa1WkrBxPpO+a/ms92cGVFKxug3dkZx4hg7jn4oJ
0lLnaVkNYKLO6m+ilANOg8ujK44GVAmTfN69S+v70qIqvXFxQR9V1ue3u0MYo5kR
L5inM4Zi3p91fnZd2/R6drNI1mOjJ2T5iP/jlpfUp5KDSVl6aU9ztNToGA2O1YO5
DN7EF50+tN2MhqIvCSGTomOnUq0m4zjfJRVYfvjd5rKIRChnsIASsbtDfqMga0CD
jO122z6+xSGwupIW5tzzsF0TDpryibzUUthTBLgLmWs8qPWfkwCU6PA8XRmZZWtU
ezFTtdG9QLOMfYXHqr2VXMR6hrHv9LgOqgJHA9AjMxJW24n/YDpobPsF784mxMsY
2VTGgEOkwNbx8vQVDUX0b2jVftfXwFjWTA660ygXNdg2SPi+wzwv0n+38lIBhMp8
ONYGceQX6y3Dr2F/rhdEMH0TUYr7IS2tcFeyPu81kgIuo9dj4c38LBaOIhKBxkPq
xNRhjppPMbzbojYFcOQpyxrOAb6koU2oLtMdyd4NyMMDFf3qGoqvrV7Ph9HgHiAT
Yedj72pEMO9DHPdRY9V2rt4/ibQGdfqApZTaZ3wlq9DBk1ZR3tGB2Y5JpLcvj+KN
OFO7emdsXYXxp180XbFaEjmRH+vWNhOX41SAXmzE2cNqoxm7mdL65zEKOqK42GeG
rTRB89njv4H9Gwzqf+anyJyBgXqFp7jMJYIdUjT0cZAFdBLJ7zqKD/HK1a9bRhvV
EgCpjs+RpZBnJwSKrXlgi3oV9fxydVl7boEh1tutj71k31gtyN6pPXZooH21JXWx
BWZ8PlpHlDMxGxZW7rhc8plAV8rxiRcd7GJvcxG8oiOmcptXW5F3KZx5o+ghwwWK
CStU5JGcZ7BgHVATHlQ5A/s8F/w3SVefEAuGyXVBDbUovzRrUw3WpbdbwOjQEWuo
XwmTE9Rg6wXPe7kh1FHqnGEzJADDTCcWBnvYWZ199CWcIPUIl7SQSwVfQsXwQFyw
k25O0RV20CMLurM6lCWMxRzORRg02BSPVICcGgb/C8vNu3OHEE6dR3wYQrmL1ZIH
ZDEySqgPU3KCsfLkfmFWhxi0LgihAEHns1PDL7861YD+qXqCI95anZriV7Dmc4fg
ZfKiI3+Pe1AzGOib1UDhKhB/u5VqueDCeEOnMp3UAd4PeT9N/4tRqIehKc8+HhM/
aUNmOC01ChUiHSmjy7LSMFMDoa8en7zP79T9K3EhMLjTmp+Cehk0As0V4y3sV8qL
8K4Myh3XG32sIwe0l8/B5fKcoC0BLvgBLZfCOS45a9Z/xydaYkU+dkbOvNVWCFME
arnVsaY8debJMJlzbFnedEyrzSh8C9sQ7pnCexdsL0e9dKeUZRN4rw/qwkLcxY/G
TS3RXhhuvCKjJLdMQkDA3KgJDlSmsGj5LwyWRL2W1p4NDGQjjQk7dBtAOAG6Rn5Y
cYPjQB2jnxnLNfdHvNi7RCl20cXJANrWnOTO7FCLsgFHnSU8Qq7aq8b4tsZqw7xx
iSGuGxtPYM4vtkjPA2R11qJAjfePTYzbpTON4SSGxeuA1Fy1MGVYm8FBsT8dblf7
5UshpgpI5iE/PDxEhGDkkhnIw+jWHe34dV9KirsLP45ywJUzNBXkuOlOzKebg+Jt
Y4n+YWRGBxUIe29UfMLzp3lD+igAuV4cpThoabhszqEKUhGbm5D7OJUTjv/nmagH
+F+YTa6+XmGCi+FZ5yf516tzvdfZObFPW2ILMQlditoUnJph7tDt+555RL8DI+bS
h29tJ3I6DUuBlk6g2fR3XFH26bV/BFI6kWQQlCq9LntkLHAJn46nH2ik4rE/s696
i1Yp8069ivXU6myd/j0KAeMI0809Wg51linY3xJd9JiBSzrVtatFHbod+ydxnLSe
0Hp7QICIReDifMUlONSg3uSHI4g7FCNZ+o4HGu8H3OHUF6Gr3p5fz2b8+muGQ6Mw
EsQpxJJ4jhekoBNHPhY9JqEJ103++FXAYSQRExiTSGE+NUbgWjkHRnKle3cWemoV
zqan5PGEW6y//WnIBoTAHK4xtyTvH8wUhxmUTGlf/LIIzrv2uF0bmBzJiUaZDbun
NXrbOI0RJq3dIDhMiR0hHT7KLUqY8IOiiLmjg3Dl+gW/aUyBUrFj8X+fwkDXjToc
dQLTXXhB6WqRYvjRK0obQR3mvNClO2of8v2YyVQvfXvVDFxHdzo0KL11jr9dDmY3
5UjPvwuVQVHfSd1JWu+nQZyyasAqykzJLqn3tl7EP2zucsZZJPkL68oshx1AeZJr
Gyk1uCNXeZD7ax5aI6dRALh0FIj+SRLjhw9v24AX3MYZ4i3Lzbo1qaFzRfV5xI2I
Ye0y+JGDTnL5zfz1UjbWFsmFbxN5tH1YbpTYn8o0EWN+zy8AMu2gTVdBCx35h8yQ
D/h0DFivMNuGaocAUHl3k3Bvxiq0RzOh5knSx5pg1fWpFqlQUZioWnWFp7i18qJr
KABckuU4p4KC0FEcqtqAaXrmZX43F9X8pN5ni04CSAz6cobGQA7yERu4byOuBPEY
Hm/fbl/TUUcvuz+VedMxgnUfFTmcAXCD/x8yzmvq9HRCW4XfcVYELLjOCqQLq0OY
IZSgfqyH/UjtSC6LZwKnadoh/8IllqW26gsLahBLaf8Cdk5l44Jn9qJmkSuwlFCN
DvwNPUIypIvrvG+JjpmoSDjPz2JXRD8TLmfl4Lt7vuqYPbLD75rc4uDc50edW15N
A8naTK+ZlGZOYTfj3/j7WFGmjxrlsSuG3zDWF4OrK/zOr1IDB9S47qrTTqRl9DTV
XpGQ+DnQtcQHCLzGXT+0PgW9UiQr/mL6FjdF+mp1iQqQJna1BhtcObK+5q/gjxp6
GICNEkbN+rpz8xVHQ76l+CBEntcRrHR1XDFFDK3y/It9JBoM+SN/2YbyORVivqO3
bDUg2TNajKvk5dRlc/DGr3RV0HOgc0Pf4C2JXPppQFgL8B2D7AMMLVmNLRe30909
Pigdq6SL3e5nFMG2T8Fa42vlSJydjU3ffv2Ul81rDVe6NQiSK+1b4a+exWerUKyu
ZBUdu8Ep68eLTHxVl4rSPuUuG7CyxPGsbXss0/buuiiu+onVq3GGmMOUCwOTFeCM
TolnxjdCTSLQg+zYDBfYmL2rU53k87wiUXnYsmFt3SZN0IkEpubrxueaUc72CGXJ
u6d/NOfMOXa0F4TaRMANAOy0wCds28GGGPJBJdkoW0rEC/rDMaOt+V6CSj9y4vpK
aJpVVA2H/OoitPLTGKGb5w35B/NHk+vpMvyUT9mqSmrxm2i0GvTAYTmvyPPdInUZ
lW4OqFmMAPfEECye59SdmXBIPtJLSBc77AD1BLYPbTR3w8vyOoo1v6J+b2tn1Uva
F3Cwusymo30Bxz6V1QZp2Y6rZHIahZUpdqqiVR1O5myF1GxQml6fSs2iyxWVRCEm
YZzoeh1yjTSF5ERke2sfHVZ73dIB+RU31PKPnpqsVdJ0v8+e9Ar3vndibVi2C0An
XG4rdw7tmHNkAtzwKKzD1Iy1H/BDkqe7fkZHkeAdlR7eNg6XZXKgubIrzTioiGRl
tVk9DcDao0690Gs+cVUqzAjRS/I1Qni81pxQz+m1AiURaPNbuSx3xES3OeWPMpRY
kY6E7zs9WhRuW7QniZk1/aLhOvIZdhetql46oh5Whz7MlOzo8jLLYDbWOtRlQb+g
+xR6UJrreWNnHGBFs5AaB/jiQrOphekXqhmQurEbKNG6sBxm5XDNFRgjK+wf6qhz
pGXbskNmxMVBJls1piBJ+kI1+HMCu+oma62Ca6E6yxPGvq86+pqpViIlcT16QfsV
+kD8TvRpWYUC4TAyNDZNi0pQFoIzdQ1z8iRwoJh98rhrlErIdZN81x4NTt7ekGLz
f0x5LFqu8Yw66zsfj8kkH7oZ37BJnKaHlLjIh6fqkwkytW9wqGtmvT5uwstf7ToD
3B5BMEcNFZAEi+DQoTm79gPYH9c5P0N62cW7SJES64r/hrxfJHeIDLjksZxzDKJA
7uV5NCNGOKaep7nF29M8QaESxDcLS7TYP5QpePiQjtJTozg+lgwKrND/SSs2VMtc
WdOPBG+sKgPDTCUVjCOerR7hxo/FtlsXUUBrQs7HdQsbiY9sx9xHPltAEzF4Jgkd
2x7cm4BrQiCwwp2OhAPD8mQfrqXd7tN61ho6C3sHu8EzYEufGzvmTBxdRXIc7Mdo
PHBnHxnLcdvimdEwaXkOXKCgdYJfeBAZmr9xxmJ1wxZhNC8MUs5y6kcFn2dd3dL/
ZzJ2bT5zXrQJ+35uWmgEZDjuGsXzgcsNHdN3rw1sTBxq21ydTND1EJ2mq6vc90yc
ErIETnJpKJkR178wE7RovyW1hSK1gOsQi+3SvAyMvin7QVEIOSxwdYNr+lCHXj1w
PNHsysCIn/tMZhaKBCI/MMax5aiwG1tXbTk56d+0JQzvb1KK+IBO7xxcMpvnQdV7
tu9YkORGlMfLraCF+Fu1sFRp15juekE1CH3Vr5XEBFVcHWaioDZjVp7aYuwIawKM
MyrL9eVrNMmR7R4J0SIa8EP3UfkbE50GGydpVcdnKW0WSJhklWnt/pqGpU5S++Zm
dDENm1Q8MyvsEWnEvN9hf+i3SEieuX0k6HIfB0aMGjQxhxKLSkf5FPUcRS4x16Dg
W3ULDyISwOVP6aC8UKnocejxg3KSNQUy00cmVc3njooCYYYSBVby5SZQq789j8OI
t3IIsbgoCjiA7dTrfGLUL5+zu8XIlJefXpipDaIdGJ1c3krsdsh3jqdU+Yu/eiqS
RA1rmMrsh7algIvW6grnvrnF1xlj9eSg3Hl0BPjZCN14XOdi8wxmNcfOIFIobym+
xx5BoOt9Gi6levXmrIu29BC/GzFhic6zDz5T8NKQ+yUojBO53gk/y3PgQIWRFFXp
cuTVPAOpr1Owyuzzb6Niow7a1htt7L4wDuPIqG1nENle4sSWdPChxqfNB0jM9RsV
qy8JHeoTJC+vvHLh3MRAt29crqAGitLoxnFRpi7xCgYU0HkPMVtAY3ZVgKw19vF2
3DdQ131bonZegKUsApytCk7BBg4hu9j7l1dsxs5Hy7qWlDliJtrZFCX32aUPxDZT
RdCUrUMtm4wUYPqlAxxpCnMQY4dxqsEeC0H5DNj62n340I6ecaiNErrlAOG8kbLB
ptqEs3hFkh/8Pg3dGDUI/KfImc13Up9G2Yx/c/d/7uLPim7fqLYhzDMSAa8CJc3O
k1zowIU8s92K4+DHeeRoFnDoXu6RXvEyctdesVDIVAGX7XXVhD675m82ZA1Elsxy
3uFvGgO2Ukx7msMdp42osKSyky9NEa7FtYOvFJdTdrfeftFP0o1fAmikQyzG6gIF
O+sb5VKkYnROUhKRbhQQGS6uv9yxD2So0Q7mgh/MxeKHGmI6+rhO3Q1Qz54qEDk5
8MvRMdrEFLBT78paAMsHGY4bQETIIhjQUdizmt6xLHcV85Vo0qUivqlUM+ERj1SX
FIp3kztotJExs+0CBKkmAoAXoA2epGlo41WuWpUVb5k9VlmA12ZbiptXuYXwFSGg
ZwgXpWrYll67K+HtbHKYXzvxEDlrASej5tArAUrYGFbhwVpLMEpsreMMvgJ8nAH5
dN3eyxBi354VyRUFPnUBhIZ0pdxTZE46CcEkTTHzgmJpQ8e3u0NdvwTEG7+Zp0hM
etZoyDrDEm1IwIO5gavSN55mJNSeLkfHAkudu/5A8Xp8HuDzOKcpofLNboX7Qa47
Z+iF2PnD3Rwop2TwuW0PyhACctCjkkCCeqWykYYjEu9S7H6pp2ZNn/s6X3syGD9E
YIIMzHl9lQcVWinVvAx8oLf/OrOhWS50swytmgbr5D1rSUYdyeM+bmDootMwAcMP
bjVBAOMqQBovkK0SSLkiSJ9kiqYeSdoi36lBzSUPsxh6qtApFuFs/l83m8X11mce
morNGKyETi30qHhVhh/NiJ2KOhpUaDfi9hisu9x98pwT2ijVIxvMh64dgg0l+Hkq
z94XmKGrbn4R9mh+30HjHR+1LkQdYELvaoUHp+v3A/wiZlBqc0sBx3F3PuHm7R4D
KT9cqk8EUOFaUO+OQ9NuRxzWlK6riS2FKULqlHUDRP8HVYh0vcdOgTNPNIzKrRZO
FUYtAyq7PzhHh/FqyJ/4271r3tpvFcUxcEs7X+Gd14A+4L1xV0JBzy95u3Y8V2IL
msiBH9D3MqdZQX1w/PEkMeB1bXg4MpsO0hYXXz2j2T5MlFkdxvEiM0k2L9kbDpju
7y+4tQcsOUMv8M3VsJyBq0IUf3JBlO7EsPgJKKHcwFf1HNgpU5ojNPUGzF4PXpi7
5HEPjaMEGm87A+7CAAhtoDhkLmeIP3Iqva1DX9sR4gw/mC2lI++UvonN1cjHPNge
3QXt8aRhUQeKexhJE1F0m0Qs5VZTp1u8crj/5QFTfAx+hFwntSY+q6GEblgqK+2i
gt+XHvsRpg9QOy/74y+V3OCh8q7oyDefykKrw5u9SgOfTnfF6QJcvWInVoAiyDBM
VFxfpdL2fHlo6WlTWBsbVXYT8O09tKtC2ZhcFxorHTzng/HKkrYbjgchv/WWOnf6
ihtkBKv8J6/P/qtWBthkg2Vote94/o+ZFdc3kDigc/gyZy1ev74mBLTiUuFwR0rC
hSM6sIc1OaUws4oF1ojvHb1TjRJioUXloVJb3jTPMFSAH1PYoN5k3L8teopwHD5w
ahTZEprnRn4SHPUGSIDEKNd9NK96t3X7ewJBP9YVwovvoxosRPUjLr4hAAdmsbEL
bT0xG4KWuXBFLBHp0bxyfQvrcUWpAt13JHJnXajGilgL/GTAdfaNJZX/2LnPImf9
jHt0R5NqXH3mf+PZcrxl6yTXAdKfGb01gjKWph840C8F3VyGKnCJTeLymVRAxFK4
oWGiQDeaDLFDOHukomkbFmxprdNn5BAV2RVTCJxfkT2+0LPEXYosLG14m1pGRqQH
4D5UjkjjrXmNLLsd3M+CYxaAWQjr4Aoq3eZL0eSbT63/l9kWaH6yRqiylE+fXf/F
K/Mi5HZL1hV1kHYhCtzb3tJB2Iggnf2pfKBhK1Jc4001a0C5E2Bfs8d9s69ZkZI0
3cb0v4BP+qmIz3QCKS0q0AHwg1zK6o1RS5rlTq4gf1Pbs2OTda4x55IJIuyz9c5F
XjDk5JmxhI5tLhhkHzeVsev8nxld3mZE6FgDCtQScqaMnuGCPYkstpYWYIQeFvu1
zN42wSq/UVY/BGiPlnVvZu/tmNdbT3ailP8SoDDr2MgzYqqpTDMzM98rO72hhpff
2ClesbleUnNzVZ3+gZG4W1sg+GRLmQIMvLp0Knnv6svlN6JF6tZYR3dnHqhEC8R1
FMSeVd4FkLTqbiIN+BGJwWOyFl+lObCCsyYg/y3jiYz7P8DWlMXH+2gxeC8OsFy1
w1w50lGNdw6lbIGwqXQBMQI9rkVO0DH0HK0ZolEEXTNAM0oYP/2bp8ZhqOcCliFI
IXPHSJG5jYhvnitWpZdV1t1RFPQ7AOB8qok7xZiusMqVl+sr1TqAmtYwUhoAA/nO
cTeSHffT/ZuNKiw99UOV0mD12iShZqMRh5IOo9dx+G7rEQpS9BnKEiOaaaYLYj8b
7N1p4n0YzYk8abk9mBFv6ilBDxPMhBAOJB8Z/Cv3Q2Fbq3qeaOxV+drDern5bQGT
9eRiYT04mc1wYB1+/de8rYo58iubh8fKa3Z98VKNjgncntipUB3xWxSxN6BIk2Ay
j997kAfcFQcdCa5e4wl0APbbcn5GqEblcJZQHYoV5PxxxNs2fLNU/STQZKuS/ztG
heNTs19wLnbzbM6DLS1Hds/O2+/Dj/BMzU8UBVI+i2F0vmAwJfI3ieir/l3HOX4+
QEhaZJIzIGNYK+iuDvv9r0pZlaT1XJ2uiOsn8xVJTrSxNhrxAvgM79xyaJZRaWCi
8AgbWhJWLAJnHZFBLQOD8Q9Qwvvbxq4JKDUOy+eGlK5OELetTkdKhl/1KS/Oxggb
x47ymI2VV9XctxQrIuhnFWYaJcLTByO/UzNfVAjov43aHxI3tpd3CU5xyf6TwP7U
luxQuh6AGrrmUHBdNMfY8/BBaEpiHfV3DeMzHu+t/iZi/wCAeul1JQ6rzpmLnv6N
wukLWsJ+Lwus8rIP/S4LUTL0AsBTEF3lvxqVNtw6zij9EYw5Xolbf/76exwi0SyH
sICZcnmHgMmYKf2ARed6/vHL4UXPd6M7XdW16Ld6MFilC8V5h2iJtGusNt+lTzRF
k1PVc56mneDhJf3yKiYrK/qw/rPLkNRSohgIz/DmIgv5zHtaL5osuF3+uKzDi9lC
sOXR3kIsoUsTFKIvPDeXoEtwAPatCIUCDaZszKG2pdIdSl32k9rNlkBIVw/YioRl
XVLqU436tpmU0y1z5svXNEZMwhR+CPkiOYCnOv5TSZ4wYo5TiNxINjnl7rH21u0q
S7QSMynzpf4PesoWepfkScFzLKsM+BJtI7xKcXXSnuxX/sCMz29tTlg9nVAIn+Fg
L9nTa6SaGWH2VJz0LWz22x5kdT9vX1ZiCJdfENsHhykBQC9rAEWAambIhL5kY/ia
ynm/LigPQwhFAmeMLMnP9Tq3lKH2//7Nn0OYHWmpfqHepujECxerKhzduYRgPaJF
Q36BlM1WlZ+8+FwrBi/WHRF2sGE+WhihTQSXBFl8w72lcQ18cPCmG90sVS0G3Ldt
Z+Ci2n03zoY1AYefqVwIe6X1+ignvGdkNyuqVueBkWgsfTzwIHH+LLlmTHS/A8B4
Ewll7UmFLIVuNiiADJ9a+YcTNUfVdLqzbQyivt4QICMo4eSHt0tXYWHiPNlAG+aA
Jo83TZl6Hs09qk1Pxabzumca8FxKlDohXwn7PdRXxYsHTkWdzx7wbkpAtgqA0t1X
rhnvvE25Z5QbmMt8RTl3xtUZ7wSG6k7DjOafLXiNdKLITGpfhuxDdqAqb3usDrRK
zzq4FpoWrcTj3FTJOZ1cK1rByY0jC3ba87wEgub7KEfcvl9WHjJFp4iFbTPYI638
SashMOznHSKtwCq0HkAiLtMIuyllCo2CIXnATHTxVCfWCDj3ckmTfRSahzwYglXT
BTOhe5mwmzAfc6JBSAQB4huKojyQu87EbbEHtsnAzmg8nEQfKY6stsKz5rV/gfJ1
i1nPx32Yg5JS1mnsYypEpvOCBQwxNTpUGOlkVk+/hRXnlxeSTFf1z441fjYatsaY
zmbDsNOKPXP4k9TzS6F1s+QY4AmIgD/yMJM20MXoaW003tKSfPT+BxnM3I2mhura
ux62X7c/DtTPNFTl0goqDpxCYSFKhldGAnxjzmnS0GkNGjymtMs0mGNXEAvilXiT
SEQMxgqEUE2R8DNDflhpiAQ6xvAFo4UlvBqzTh8dg8GCZgQoxwYp7gcz9GLETh0M
wDC/exN2Kv2K97FtLZcb1SsiinzaPdVsbXrwE2kQFLHUthopiVTRWuqQfxmjOqPs
Pa25F0d6ofMR4a2t9RixqWC1TswxgNld8BqKWAkPnH2SlA5cyse31LgcQcTmPtW8
TWzmINs60ZWAas4Ewpl/3jf814kE+JlX3qd1Kls9uh6LAu4AgDDiikLqe9dzM93o
MrGGYZW/X/M1cHWkjkp8CQoAqzUDAJd8TuK1G/O0pLnjleIPjhR2p6B8CtWXVWYh
M7qSchAeKkc5rGri9ju6gbrtn1BiB2zau1yObQ9n+sbVewhUuQPI07YwLrkXqN+X
JYkIHJBrdgj9G2FDmzH8dqVERtgutOK8abX2EcPwuvKtEzyMT5ZKhm9c0O8XUMcp
6tTKht+2Dk7Ul6gW9doC7ycRmMVCRefru7/UTLzIl18sGe86QnF0lvCK520mqX8I
xaDyVCw/rX2TJDWHEQ3B9WNWVoDJl/v8D0FaiBlkJmuAbnPSteSjWsyGM9QD/Rnp
eveScxxp1d4q0qHbW37DBzZqGzDlFzFl5h9RNehEhQR/36TD506cKdS2p3NRzyTD
9EJNEsiIXHoX44IMao13P9vnnmpJWA5o0gQRkRDL2M7dHb45P9EMYTPmek8yrP/d
IispITNNhESvAFXcPGUSn7oSTpOQNsT/4UB6WsvtjnQWpqaPMXj1V3q87iq2oJxm
EWqwF69JXH3okaYevF8oH4CzhAtnwHOZHRSsPiWx3M545STaOCo5jegStvIP6ouM
k9RN9ZEJMgYErn7xpbNM4ouUpAI0lEpoeEj43vxJ9t3UiBPlTIH8Tsq9KA3jZqLW
5CyKlCZPDHVwKgLlvSRGom+qnsjezfXXTJr5stefbYmqwb9wD/BEvGHvPEbUD7R4
7u7TK2ox2g28wxbmBQMe+VaDaH73Od56hoj7jCA46TZaqcAI01AImi1sQYowvYaO
is6BZvAg+oKlOl1znTx9+athvS8d3zt5M07/E+CpYDQZ5Q9K6iwcKhn3zZsN78DQ
DsIXPZrs7x1xZDPV6mIQgk8YWfppr4b+evLCREH3uGajSl4MvgPQtxtBdlClnED1
vy6a2kTAd12SSmFiQke/wbndoPZ4PabUy1PvsT9MluorTLfip6fPHU13/XR9j5uJ
gLI44vEF3lXXhpo2lnwQiLksN4kn+WQUBk3B4jcFASaDi+AfvtdbAAQcycbF4aoH
CZQk9jNkiz51ljYkPGTOtn4d+PDek6oDIWDFWKLQ/LuMrkTI1GAc4hYRoaGBOysf
a6qMfWpIYRc96QE8GIQmqKq72MK9IIeZF6uqcAFvKIicewfabL1whhb68SEApptV
IQniE5bYhaD4ZBEtYNY0UQKHK9hGuGwY9AqYRam0Swd46erboMxZKqeOsJJOq9Pt
RmcZBYwzDOebyvLu2xzdDbw+3MClILtho5yBBUMcwJJ85cy8sRiTa8tGdJnF3ZXD
OQ2cCqG0e0zQyl1Hc1B+jtBKJxrHHNUeAcpJ2Gl5AgfLo2WDiAaxy4m4ZdwE+c88
ApiVbaLQaJNGxqZuEJeUrSuZKdxgMF5c5kAnS9R9AWqNtXpPRAG6SxRC8yum/AsP
jLsn0c7jr9xIPMWhggcmCS52zZdPtURjoEvXZRbEkJCZ9wePi5G09peRGbQVTpVe
NZluY4wVrvogmpjz5htcuTjTfrCB+YcrgllGuin/Mvn4a8luZjqigfVvLdHDLalC
yLFUTvui3URV+TxKPwknpi1typRaug5WDVpYzapWV7rdpEoygjvt1SpMKw+9+eOV
MVb5DMAKERE/pthBwzZ1T8M9hFLhk1JgORnsJuC6Ndg7QalhLEbiQOxlbdmNRf+9
l2jbwVht0W/uLV235t+SBI10kR6ohJD/LNse+LumohctYFV9EaKlyhM0VZBuReNH
2kTXHxTSSEKZU72I9uXW0P/XS9zuSVvWvjDIPOGn2Og4i5mGg8J9e0c+3FroMzQA
bxE7kbBIoybENZFPllmnxp+hDagpS91AAYobz8MWM6Gqh5eGj9q2nSGJ6o8TfxSC
unc2bL6LbPerJBhPX6u5DTV3snrTVAF8NQby4+dLKpUvPdXBkpAcXFcyD/jWXJ1L
M74aLUNyqYVijyCmxW+uvtW9a4MrU6xQC+XrQo4aLW5GrtCo0j98NkzLHuQ8uImI
wKPnueUy3KRKQNoUhcDjZCx7EmVE3pkCFbdfC1DpHu5xMVk83LopN28W8oq+xuLP
oNAt5gU2bhasIfI0vsXNSYMCz+FiERA0VKwuE0BiVnUsFZfuatxfeMEyApjA+tpH
TdrRNSZqoWir0XUqe9QU7r/EmeXBkTR3qcZAHDbgruI1z9yrYI/UVFHx11YK/GcO
LROrFG7uuwynXe/nfOG8GNkVIReFJC2jVHupX+FRZwvl4LNfTO0deU+by3c1ne+x
UQODIQZJBKO1PGkbTmcLMJRbhErh5kKyyo37gXE4FFbAZKUOmlQdPuKIECW3SBy2
aO96cRBDS54tItmiOHAmVQ687c3v8JjxSI/qxS2C84QKHLHCxNzf/V41NAv7s3wl
wPiJxPCW+1ChfG3CzR9Sk4S0G3/DctulYZ0dg+PtCnMhd2MVT2EHPz7biXvt3a2y
ZfavvZph9Ofd2FYvE5fhHkewzryD9g/x7KpPEUvkkhGGXuenvgLPQrkCbDLXWqvA
bEXqYHe0KQibYKLL8vGONm1qdnFUrgWYYNBrleqGWaDWIFCg0uchrcSaLAeAjuC2
tihYcAfmkWUQObGnhsdR6NuHs8prjR4WmbVbQmz5TABiQBjLuazc6Wj+MeCfv1wJ
QaHSjundT/aeCEG9/CikQGkxpTBt8dZmm9Vr0sRPOEGQoazkG7YzTZ86hp/TO5oa
RjZ7SENCmIv61J4IPnsbDRHAfQTfab+DACGTtqQ9b+VWOGzYxOQvKcHmKdzMwWNX
bROWiavZNnxZH3re65to9aSBnGXShj0ODgY1pHgXPRxGdsiidRaPi/SALqlBwtXD
Mwx5mbN5xjVibayLvb3CeJ6bjdenAIcGb9sIU79IQ4lVbnPdCumRFHi2zG5/E5RF
WO1rlUgDrCBcwNZAZ4NCn0IDyUrkFMYb16qxe5QiUoInaEdmDh8URiIf6VMtMtoQ
ASs3biO1j/6Tf310lisEV6uVPfkR49RzuEOj6ST8hWKsygwD9hBUfpfgvjMBR4Tn
L1GjGhKsQ7fGR6/gkOTNmN5EF8cn/mkyugmuFQTN3ZL5YHJ1QSopB499wJmQ1IoX
U2FRsLSOBhdzJC5J5OW+8ufhYorVIn5ece8bsPYsE7osM7V4TcahvP/FCglunnes
YaWoGqqn09gx0VVo7rpEBHlMjQNqXnHrwRoT7/XVoMqLWuus003Vs2cI0Dt3nH3q
vfKVMt32REbCfH1zxJOAb/cwZpnZM95I+BhhZC03gIFx4FA74dRAjeDY9XQKwSsv
gEQWfFDOXYwXx64wKKSQUSecbJgDaV9VZty3eTgLvTW/UPzwM19okXm3s0YgF1tO
UHJXu9dT0hZYpluzMhJQXDXhNrJLsiNiEyZpbpHFTTp2hZAWVv98EALEe4Fxj4y7
oVH2YWa3ui2VzqghoeHyhwSb/4ng5UDFf5Ix63ESJlXOsGcbeNY2joomEDOnaTE4
7oSiarcaCdiRcGxe3GMv1EFb02PGUMY1BOKg0REQyE5NkZdg4Sle+Aee0QGyoh9P
WqG/9wVV03MlINjCLozcp5gHznjicyJ0xgBl8Iu9xUfvXp57LZN+YlbnVxxr4r/r
TDrrHHaJB4Z+8HvTZJFfEkqib6Xeo/zDbSbea6WxSKZJL/Jf/Wh+DmcDEvhnNThr
nbklZpJWjaoSUFULSj95ydyqPI/WZkbUPrGMOpDJFjW4jvDnQ2oigciHtSODdZ+s
duWJXQJ1x2MVUwnFbmGH7hGWauhws4YkEJDxBM+BZg0cZgXpxQo5zU06TnkAM0Az
OEUZXm6fudLzS1ccFdgbL1logQSn92B8vdTrFJADS7g4RbDXTxg3yeJUxAWuJNDJ
Usnk1nSaoSzrtPTnU2mvL396spmg8bOXtb6wkFqVGCiMfdY/XsuaxCUpUoKOSwWi
LRE+oCGWwM1T1HbomPGwrhq2gWIuHWxo+RKFT746dm1YnkqoCQMlOfPjKL110twU
ys8gxnxih9q8e4KyjIoH4tqnToSSmHpQ4jaB528nIXwVOfTPqmTFZgTHsmXP+CRG
lrAwELeYEYwUwAatxH6QhBCnnqmTGFEwtXgd9UNPvEdJv+Y0eMluHGWA7+/cr+eb
WUQDjQgYIQ3P3P7AJzpZQY/q8Ou4NeLV1Y0stnI5AjB9pm8hq1MWGX5Dw3O42uqt
f0Gk+kR8HfVjn1df9vjWEvpdsDjwbY+r/mZEOPeCBZTq71Qhacefz/F6zT3mRHlP
JZTheiMtYkpLRWSctMHeISY+olkOuGipVGlaOhP1263Ujp1lTjJOUuhlqgezWfNE
VR36eSmANZsEBvqxFIbCzcXVQe7hk3ufwKsd3VA/TMtC7pyy6ayUvoaz9NxWtGqA
FbihTOmrDcu0dvfrr7h32+MjW6f5QkNas+Fxf8xxs3emPgi//vrECHCOj0g6fJ0Z
c3Cg6c8iAmf00XmVAgtAQvdOyMN2tMYGftVuDkv6VOqy0ccMmZ+UJwbF46imLTgq
uYkYcFtDgOYVROxiDVvlV3IypanCj+JdTFDhnwKzZ9HI/8rvn2vk80lm6BNSmClC
SJgFSceItGGirEw7Pz+AJ25p2+gUZS2ZHPTlCB97sUrGvhTfOmSJuaCgnOCz4YCl
Nnd6gCbk+xUXnxC5f6nDJLSlG81ZAMhCtJIjr3Oe6TYlLBXEvjlC59DuOCjtGoee
EbgURXWaBFxO3jZmYgJXPKNdNxG6MBus5p+QFYhUvNkGB2JOKmNneGNVcf0Np3ws
p6fE3ojAPIgjv/uT16JEp83ScOpM2WM2YGJGovRj6/nmKq5DotXlfEILkEjsLH2K
0OrnlGpdBJEHmg6BxiMRBcZxgNbwPWodQShen/QwZ8+R9IiGHgAdKEs2KXJKgTkA
CalCyWGBn6sWs+ZeLa3nJI5798YI7npHqSCSe/nlR7gwX00yommezRH/bhN69C7v
U31HUsi6PDR9WeKBfsVamw9oTpE1YsWCtQdRNxWPpTpaegk7IeK2fXxD7zpNuxKv
EBy8Kq6F4I7WPz9gIs1ybHrDS64J6ZDeYaPDtawb/qeKkik71Sq1j3n7qP/2EQsi
UdrDQkkcXx52dHDOekozjyMIYyhfahwE3K+SwlxE/RopAp4I/rYqtxKRBjZAVNfb
Wj+SG5m/0ypIT8iarwfuykE/pYmc0evaeN2z29dhwwUTVn3lbZRep+0WLf2Br87u
M2IPVZWmdK2l8nU48342C8LpoWajqa4YAgVl2b0nmXmYIPLoPwjEnBhsR37QVBI8
VD6wpYXCv1OXdcU07yCQgyPe5j4DJCEHXCVuoaeD05Mg/ITnOQSwOYc8njO7f2bp
ARKK7clg7wyABgMWh3/bdheXYdIQFi8jCzLkZ5r7OEzugVyRQtX1DfJFuHdT3mWI
yBZ8P1klysqLlbxFs/LSQ+/SxayC30Nk4+sHGsX0URwxWv0Opx5ot0OoSnKjyGqX
VGzLin1cGmlVz5Vu/N1xUTzzGg3NBTOXkrozCAXVQvjTMpDG48fIKe4/hkZgX6eX
qZr+l+xCrVCgaz2HQG2wMiGf17JScQqqdabPK1iN/qPojNoxDuQFsM14CSUQwXJT
rhR42iwjqux73CL8+lYZBxmIP5VqzZlN6UfGAx07EoYfE2q6RGmRAg/IGJdIpWx4
YEHoh1HHvQJk7BkbPF1PfASiF/3F8gshLygRUisdnxZjVe5Nwt62IxHtjNkNpyLC
yIE5hDMt0sMEIfLHa0pmXj59ByeEmivMTZy7FeOfpWanNmSxl46ASbMiwLOaR3Z6
udrzNMyocBrfHwPwXuBbVe/u2xadFxi+lXtm6gy7/EyJ+noHjNY0VEWdvuLXogKT
1Kce++o5aeENzciHWeg+yYuIiT1s7Z+KslB7Hr9eEqf4DCbVZwjTMBhnBLgjSupO
vujWK90mn76lA/BKLrHTsrTInqcONgJ/xwooH6GTyADg8BoaAQSn6i/LwCzfOg1T
r/MGMjnI19/UkgO8A7cs4ixh3/evFzlD5VU0gXFPJb/wVL0LEu1q9b3zcrdP/GQk
zmjU+n/eGqGAEmn3wZuR4ENqRjNi5qKLS2XjH78EYk9WmpbS8EEvdevPcb7Tlk7Q
sOBj3nhhSpfJ6b6uC34YCFCOXPlT8iB5kcWwtw3SEXGTsDVIe5mWtOHdEHwzMwH8
QZTaYalgznTL1HIBeElBvdQ/J2lCW9Kv0pVls02vrC1hll1/WE+oGkFonEpo95CC
+Wyc4IZpZtzGPu69K2Hb6tD6pyvw7ZRyP1+psNQoWoPvcBneIKL2jBVhZHss6YqS
Efq3qBAsYr3gAuxZ0HlWTjfIdoy+uDJAewA+BwmG1SjYG2xn841mf4oWwZQH9Icu
+yTsvDO0bfVsnN7xr6HYc6i9nzaNgxPxYdusjrmvhpk7eNnkUH96nUZLdGe0ycMN
wwWfeAyrFpzMyzX/jFoj92h2o9oyaYIePlSDiOSCLGFWWgmi3H3NYzJfJ07kEDml
fK0Zega9VWZiLrVUmhMymXgGfJRnyWt0Bhy1aa2xDOSVyg2GB57qbhUcJU+ZvD72
j3sMOEI9bVxDYX+w4pOKNGIPxEA1cOCYI9xtI45lGFmUV8Tb4tUHxHAHQMxJsJlc
m5BSYNzaJYMt64lSEWSafIIolip4DHVQWV8YNl5SRmmNtUGMw1CusGomeRdSBXHe
0upn8oXbLRiJIlYnFPlfoKO4L4QgaHyNCtmIG9NkeqZoNL46pLnLMaIT0wvoHpW8
XSnLE8uoJOTZa8IIHCUB0gUAyqsbrVoRnlC9jXfyqR08mGXvGPUVd10fpqYv5jrp
KirL1I6UTrxVSFIIayxTmc3vocclZj5/z/KwOFJ3i3NF8s5knrpHr57xIA2DCZyt
sMw+l0GOL7zt4eX9zX13spKkitlid36stw9QrUKHV69jYeNReu57I4fUYQ+BYttb
OBscX3WxZtLxmoDEvYal/zzQQXnCm7UKN+dCV1wrVjBOGNoUDpVsqUw9zmUT6LeX
NEc1w7AURGA/wap67vjaerY0qSxrppU/VEh1LS4YC7evOu6SN+Xm9CPW1YSID/TL
CA5JwIOjwRIDu4M+hDeL1fAFZ+93/tlIqEZPqkVAbg48ROX9GtqdAH8ExlNZgHYJ
+H2IYGiy3IDAtcGhG4+aTkdZdfnAsRmuEkXXlZdbNUDXJTLqUnTN8I252c33ua9y
va4yhQ6V5hzppy6hXP21XVMgpC0w3ZU+SKnRfHIBpSBh8WGSLXUrFC9xJswbh0G4
3mFLxDJpmgBS2UdkfHjRmPJEojAwv3w7adGPtFqJqx0gr+dPw7EXVAr/zi2f2HVz
b/x7T2TXFW6xOdj1D+0UI1UmhgOAaZS5//5W9fCBI+u39gUzKbKlnZMy4LW66WiN
w1cAU1sMb4510cvAc56Mk31GEvOqLk2TB67v7O9rHXoFW5jYy9w6kEby7ZvO5VV7
BwNhM1bLHBcUDTQFCL4pTSWOEJuVfLPjO8U7K4zUPwoD6QmMY+ngfVsE1lTaOIUU
jIzBnUjrZURGE96T8P+r+wM8M00UP31CLqS54D1YUoaTKvBFGW45yhjUV1P7MoNM
bfaUUqmrdeKa6nIhvMJZpFHC6UGfD0+CLrwTJJPupuRHxMChUffyHwWt4pDaZksV
3NYoneaTNp8MqSDnDa9UcslAOnE8WFIV2zcww7epy1oOhUYEUHvHAh68C4h0Pihn
jx4k/jbxyoByYprgQXmI04C2a+hLPyPDx9WejbdjUCkA32wGUU32VRuLiU+q6hSf
ytpiokIci8wSg5kVCniJi9Ro44RHpP9DRbrq9BJGu7kjW/a7KL2HaVWDo74iofo5
K5ABaN1fTbkJos5mqAJScCUzduAfivFGhAaQCTnXG86ZbqwwLQPva9HVmXYV7/Sf
F/zl8O00GBrYDlt2hV6jq94i60tvJ77/+fpGckaiBjpmGX7xhCNbUI4lhQ08id2X
PbzljaKbO3InWTeb88di/1vgaajRVMxrzos5PRQ+rleRWrB5wS3Sjah+HbTl0Vq1
C8M1aMUVNP06QVRjY5xhw76RzEnJXG+YUZYJpzKegfHmXnc7jdynTUAXZunnYDdK
EQV7rj+sgxP9sZMc0ImgWwGEgbESStjKHnUYRqOGeSSw/SdH1HoIAf+VMlButAZt
LFT75G3dCi9XfVClsLxqZl5IELQ/BJc9ZpAooZNVUAjc3dP3ViAonKZIvySh3VtL
gOUuYhrdTAw0levhuxaXrypho0HVUBdA6BkRDbIlRF7gALOSWdaAn57XAoNoJfY4
DBIgICUD7oeFXaF1JPXMCMGOLMcmMjn1nrqUE6lImOsWShY8z+sA3CoowRDfv0Ro
72pXWpUxdsx0CBIIQEt3Yx7ZtUZk2qy1qMEr6gj6rvpLyhE8RXyazu6u7BUcxkwF
j27KfV5IM9vNDFRxbyoDU9bjar7wKM9YuZYccFCUO18LZhQv8W3Io8HD3VcqvbYk
xdSr1KSntMtMAIde4Md3efcw2rjHL6sY2qdT1QKEDJYeiGgnGcDN7dL/zYedvQ7F
fp3CcdLN2BJ+MAd11FfQ70vhAPNAZw7q6lJcNhFu7PsOv7Ly0lMAV0Vc/4QYYzxR
KpKKcsLovPv2Zi0CIaW58wtuwqiIrzPKAvFCU4D02NTXOIqqOcdK8gTEOViIsPOL
UJ6TeOZLEKLHLavF0jUS28osm8EfRJmPjGFReJ+9LXoztpNCMgK+kHf6tck+TCpw
duag4n+h9XqeJZf4ZO+9lzqKeY4UrUiHasMf7PYq5kgj72MxAbnz5787zITLJEv+
zkp3YyiHoF2UAwO6pIlr/hWX5nOwt7qgML6Qiz+O00NSsejBheXFCdkK7wP+L/C7
V7qwvn3lXqxGz2diOhshwC9UIbSlEIypuK+7RNFVfLZa5QedFBc7eovoLQJ3nuRK
UVjesSY05SBp0bUzyPU254PHmA3Wb2e+LfJFUTieJJkQelPtalATjFpF3fGlUxc0
SH6/SbcpP4Og8N2gQNV7PTexgUZ9hG0jXRWfcUDQ8UFqjoCEr9NZ6Q8K+LGU/PFd
GLwi8dLFfX6tOjcqP/IIuq/jVlKkK/tpIkriVQWIudCo2/VZvLagRBbgI2trrh+r
xXWM09bvl6h1SwxUzzNkaAj/gujcmk/zeeN3TnmGe5zgxt4VvjJI3JSqDTGD1+c6
S89UPeMayW3+Og7V5XJbPtA5egrsvMRuPGrNXdWdsEviR6TJLqKVHDSHWawdTNe+
65FyHUTJk1Jve2+P5sT+Ff4XRxo4zfOG7D0HaS2NsI+R/42tfMgiN+gU9ws5+/6v
h27g6mGMACGWgDlMtGbgHLz/OBf0BffSVRiR1jgj4QAGHLKGWXhe7IK23cnFiwcl
BmrqP3k3LmlR6TGqmSD068q/EHFCnLWMDTay/Ik91DjHTmWiTH41DK1vbnTqGHpE
tUqONvVFLKPa1ryKQlxsBfSUKdysW6BA09zbMfM9zBC8K3DtimwRNXXfh8Ee183m
XZXMwGtsgvEHmSjQH75I5x7OANBci9SHyztJJrTtjam+I3Eaf0bB2mEgKfuXe1KP
YLGWW2kmV2h0horGKupOGpvBHQMPjdP83S0iQtbworF8yEfTlNzB7L/Ck9ejAWmz
P109t59LoAb7gY751oLA2zXIrl4y9xYL4jOF98mNEz0hIb1SxwtvA9R1HZSCdztQ
zBCnG4PRGJASEFJ17J877Ub82JI9Qwak+ALbHw63SF1hGciAUcD8d2LVjXzqzb47
nIautNW8fLoQIj5rIG3Z1475rT5Kgp8h2FaDR+lALWwukW7CUeUDHvcTciwbP8PR
tV1j4UTASq1jf3EOKX1ppZPV6agjjtNbAx7s6fo7IroX6l90DrLTuLBGHMLh22V+
gjqAy4j62KeWHNWN/VVjfFDjbsbx0h6/ewpXmvZ3ch4NpSZ/9Uq34VKGFQf8/oR6
LC8Uoy+QLCaPje3CeEuNh3pB2FSnDTcuxyL9BRm+p508ttFeUr/Nt/6OngwEZDem
RbzMzV7vs8al1xquM5/sSqzyRcUrrh72prF9LdLoiKkcwE1plwjhUt0MYRF5tKHS
I63yjVkiKj6y4/kSmsce1Sza40ManZdSRHIVJt7nEafP/e2l5hxnfHciUvnTIcYL
PyrzRcRZpeXCLGMFpQllyQKaQ5CqognoCxcHEA8VoeYg09EPoXMGIB9ZoYkZfxSH
1qZTCnLQvnhdxxjH6mmz4wdc+mIhDw45RUnoKR9bbdCptjMV0NPv9aOzkB8DiLnM
Viu41RZm88Jnf8Viz85bASf4WWO4MX7RbY+tBdsxIjNgPsah0Va42Wg6qdtRR/1T
BXsqNVW6qECKgWxkeAfy2vTw0DlMwPPfZe4kzoqclC7Fg3/rLm2U8fU4+/0wXLy1
BAs2tyicntjUgYw78paBScj/f271b+gxOVm8ZtKVVDpoK+d7lcCpg8NhCBUL5xFZ
rLao9pO7mlo3GraO7YwCcMq+rPS6cEK7nwQprkwL0XRs+aSHNlj9HNjXi0+he74l
BRvTR1nDEEmtQTr0BMUJjUZko3hk0kk/gSvcuTHqcDaQY6ONcv0SHXay8Iy6RE8Z
VJac0F/yqiYPLcF87LpyYhxBJvWEpcWMB1hghmHsWyZhSjUw4Ef9T9Fumz9D0rPo
5C0623Z28QBLPuG/KvVab7VRLNRPuB0VTesnaFGmCq2INgbD8l6trJFHYk0TiwSb
yElErjHUgsMq5CgWNDK5oS5bo9Et/6z1c/gXlaQNXMo8u1SbLX8xyYTvs7b1rkXp
oOscRkTMF4mtg1kQ7jL2mmqrZ0JsG1BqjqgsAOjxgFoT6EekmUz2U5z2kimAs3Tt
yVZfZP79126yQqzoOmRYBOxBfSkH5fQQ9PIolaRnLYIduXDDE1o9VbVbnOPxLHM4
xVzmN7Hbi5E/fLy12t9CmeghwjXt6FxOycq+c8bkLCqFzOtiOxisnAxkPBO/8CBd
ELzwMkG77+CuYN4CmpRa2djk46iZ+l8LkhfJ5EivaN+/KKX6sZjOT3aubb4xzeZ5
evFNQLpxr7mzulxf1aX8Ad2gFZgYvys4R7i1BZVVLv7W7yZii05cJwGO4ipjJeXd
7aYfGCW0MS6Upq7vyQYFUg1BMidzMhGLdFfII/mUnjN7G7uftMp0De9BbNHa3Bdh
laROoKsBwAAYoY74MlGz54kpttmBCtuy6LAfl2wgyethPYJmnvzix5yf8YUeL6R+
f91AoSHH55S/pM64m8ekddze1hyLCIfYfN5mKRCzpr77D5vWsWoWf0/CAd7IM1Ye
Fa9LBDkEO/4OtYBGV5CkDrMC2Y1Wf4TFNdTXSPeZiDqa2s2piLgiGdSVUk0jXWtj
rJwH6b/aVwoAYZkSAECn+qVelMzGWtry1ohohX3kH9d2RkiVfOueXD5cfFmuOCTk
3b4FVtwiceHZn5Mm3sP2jarKfMWSviu+9ToHXuGn3VYcdYO9VtttiiGBSGRv1MoE
3E6RQoF6FDEpheFPIesLaMU0ktqjEQGW7V9OY9O2eUDj9mN6hxE4BZYVS9Q7GQ+Y
7dTO6lUG2rtif3Mg752lx+YSlomDg+nXOVYtZ6SHCXDIAiTmegT5lFcxfFfhpYTl
Fg2qKRNfZg/czBr4kfa4Cxc0g8r4EFwjvLUZoWK/VmmVkgZh2X4K/aIF+pyMhYi5
UeEMKKxF5r/rHPHyJqfkGjE4on5xtgDvypkpCiaNM0Axdx0nvE1Ybg3vvA3Izivb
nP7pBIN2OT187ftx9qKKQqaefYqBaMNYTh9S9Tup0z0JtOPucgPZMn4Ah/zI/lxM
rtxbmiQem2gFx8Iubwd7F3yYI6uj/vOV0gv9B+HaMYq1cnZxGiZMwVtGfR/mMOmZ
UpkG46pSL8OImSX8CLWbkB7clrccv+72gwMbGVIomtqFUsHZn4OIwKh6rVTgmT55
umji00Uj1g5mVokz/1/bJ/6L2olpDJB0+X0HT4KblyRhq7cZlOnO3TKF+P/mDiSF
F6rQklvSQN2JjAdFfjOkfIbE1cX9APGdHGnFO6KOy1QF+UKEzgE9UMyl0MpI4fds
DoI/yaCUc8gtOS0mnqHkC86IR71iVFtkwTCCZA7FV1ujcZ0+YYmXz+MlgSU7BPAw
lnAFDSEQZGEK+ceC/hUE6wC1/oapcoKAgmyM/Bp7c4cOdEnpjb+6TEcUwyulKM/f
TlI/WbgQW7Htc/SkVv2eZ9A12wFXUkG6Yi+rFSmR1s7H3oD0KjvQmeavSTmDMO/w
2LxUvaBTNxf9BtFHMnZg9+J8UVafsC7ZfyD6KmdMOcXF8J8a6q16PJYBHNhXQW38
yr5lVQWB45LvipievHK9c72TrxdjPoCTeon1/oqZioLpjMMONnLUin6FB8hvRP3P
oon0/ftZh5n0dRcCfYdiLWXtgauE0dRrQ3FJXbIhanfm8tPWX7B/678MN2TLZYSr
p1/5A4RhfspoQgpjWfNi1+vnLS//LPoqpTJfoJkXyXZRwhpRRVfAqxFDBj6CMXli
nmy1jIppk3Gz1c7TGV0SHO2/qQqrq5PKyCtABNYt0O54dYuk81iyhio+iUQ1Lk1e
ZGByVx2k05W7GDcKvevEYQyNaKSqvibS0MKoRALCRB5G1Ec/DIR3prluPK33bppT
qTYhtjTc2XSojqv+yZEX4dj0gyCul4Yl218g5MFrFmU9B8IlMiaSUxSgr1i0eiT7
NKuC5OWxw67XK+tJZ+tpKvmEbYYHdxtebWo5uVE99hIVPErnClijnprzwAtxKo/+
PKtlQjgg4NMBg8A2BII8HYakpPw7PFvPLLIiTj+eFKVc2nFOr9ADULpE9Erof28F
CUyAjLoOeYDLhrBJkZP11wIr7hOG8t/XQOdzcQmBEcUakHm7eYLMKR9OJDayZGxV
kHb1ZFXo8TOjryqXDj3BMNIJ5A+v/ZlUfBE0Ki3u3WtK+iNJoFPzOUuvAKE6dorK
JuQywubksq9wup0H2WNS8hvChj7S/s7GlCO2hsGHMVNhKMebycc41yOm2uGzPA1k
0A7TFWbEiwgyAchDOpXq95QGSBGoxTBq6L1vfDkVWpYbaVSMZXNXB3DOhk1bvxiW
78+acZADvr6iwLs61hiFRg3Kl365fqvYPWOzRwyJ4lmU6OsOxPfxLTF1KXqLQ632
yFh3wLpNC4zg9IDDAzRw8lKC2Z1skjZ6d6FQLlwLiQDNxqf24wXUbHGCqao7yMzD
wcguO4tBBS+Hd3uJD3Co75b6EHMp3dddCkXdQTEDaR70F+ZXL6IE4xDfwFT/rea2
u4zk8jW4am4F9/8ovU6b7mK4KIETpORYyv7au3QCyngCki38l6F0cbIBD26d49cG
+SJf5efo8CwIlUgvl2DzFVqSg6A/fd1gQzV8PSGuGPREn790r5OBPcQFNvGFt9zO
uM7jINFi1z9eyNulrEYqqcTjNMjdBknfkNX1Rjg2zaZFjN7R6DPUsUcqqH+QdAcF
8VnS16zIPg8AATuUXJ0RvCgjx0lPzeaPfVA4OqZK2LvLkcoZY3YRKftyT5F/ljn+
TE+8nPC6AHHrj9/pO2c7/S9rP9qoek+9FEuHpRnzr72N+tfAt5kzxxccCafi+tUe
gQw5mekDD3cTXD/fRmhciNVkR1/oGl8mk1MSociaNaHy+CZRATBBF+8X/5FzmEnL
e2KanVPxoduXJBeQzCgyG4fB3Ij7zorEh5daLfhZj/7G+sAEmlKNUcSNr+fNDI2c
UEe0IxWhtqHQPw394CUGRcR520rvSYcBR4tsAgGINHowGoArSl3+/QkpE6b9RXwU
iDxsNJqESmFF8fEItpplTy3YP7noNYxDiiGUJAjRm9i7qTgoRFeZ0qdPHtp1wtTa
SOiDH3vbz8bLpgXZQi3KVTlWjw8eEfbI2EGEsPD8z/+kr9RzTwAsdf2acEwzMkOI
NDYPWUoX6rY5AdSen9jSFFbCJUslqOUictJh9ojl3pWHQgJEylh2cWrJP5lcWbTS
DryQiBw0RD+IT/0kIswcua37xcQ7e+kLghYHy3KXCz/CQkiKlhkWuzEZmheYgFk9
WAxVCIbsZxbnTZiZLc7+/EFj3s3YmVvGNjosAUtb+gB9Fn7KIkMRueh8lvQ+s9li
LJmFDxzkWQWmglsQiD+oVTbiBGEQPqAYOZrwmF5NY08g+f+P1BE8pEMWGWVx2AGq
f+cFGRSIH4bvQZYqqURaBFH+wT6pxLozCOJe4re+EESoRZAh9Wji8dKGej9FNK76
JymSH1YBl5fqFfMhmkGdFjBMyfSBK5rNDK2WlVOaUEua3GUgJJlR8l59xNp/BxJM
7Wm6rBxgqTXGM8H4VjWO5D9YNmoNrnB53BQfQOza9HR/X2npIKk09xPeN8rH2gdD
ig/HotUVSws4l9S/+BdqP+VHenLIq1xJTzhzgr+GdwZJl8+0Xea0o4J4NPUpBwOV
f/oeswm55daTx1sjci5yeojOQXo7o1gmF/KfXBZRwcza2U+U/n3L+fUpK9Afn2ac
uLuTWhzaTQK2NsXl1YySIn3AWvjMwv5yf5WVbQJ5Ej9/KjDBQhv0BFK5b5RzttLl
5koz2T3RJIyy9cIIkey1BuOyP3j3+vphTUJGU5LTqeezxYSjhVm6OEwMYECrg1Sm
HZX/HS5YyviDS4n0oCOPkJIfOSV+L70RHhT6XqRSAK5eHbouUS0Deop41ZTWpGrV
V9KhupmkHo3GSMWgZt7cWPGCBRO4ZdRipbmglJbjTc/KOpiikBlDA9g3WZT25eo1
Ct1D627a5JRkgkLtyIBmo+YMGKKQv533s9oatxyMHmeS94H690YTY3KJCRQKA7nS
pD+howcwjuP7gSJ6j1I3U2el/3uMTscQkExYLLLYjR1ICsYpFwbi9saiXZWgihnk
hrlTS1/pFUPWQ3AsLOIJB2lbB6CD63y6yc+vcEu1Fg7qC7epnVO1G1PRmzU4wkTt
Aw8D/J1nz2VnsJ3wxNM9NU2jK246koPQ1L/lI5URS+Tc302L0uA4OKlcPdwKkX2d
KZHF++8u++FmDC9xfrFF7PBFAuqLHVNoOnRLm79orf+7McrjtOJwqBkul7scOViU
b+wCABzqq1ux1kx84bJg9AmHc3U15fflogKkw64nu4NpzPm9lpgwcC7i/at3HqVh
5Aki+CUJmiC7Q/fhRztxVg4jdeZuYpCpQCRNZXrH2FnU47J2p4umtghmkDogwhvF
sSgbtxATToqXrR6tjzA/Qj1JWzWLWKiyO0JdRoXpcRMLtRjoYIzhUvJLFdFcnwmK
M+TcKDHr/jNyWbL2X9f0gSefC+Imm6l4burU1RFDTy8K/8SfP0V2jUs4wH5NZ1Xt
gkLlQO8cqdJP70HFk04hpEYeg8y3l1yRXCZpgDuLH+Dt/mxFV0sEJPgSz8Pmv4WK
geMp4zWSl9ZZ/UNt4SjNNUHRV2f75/y1+CbKnPn+vweWctEfXinXs5HWjhZEwbJx
O5YVcS6aj+t1V71cPH4Q1B640FXwRTwuSACv3v83+K1waJ3L3vgihDp9GT5TAoWF
Pc0Lmbn5O8cgwrRWSoiCOzGwzwPqKB6dAUQk2wao59nJpMTsrxra9rCkkhS/EjJn
xDci97YEi1XNwyNmmFr13PoQFAI1nN7dMfPuKRI0Wk2SZOF+9IdLCmwT87Rk1lyJ
lsNQfr8bfO7NiK677hynV/yiTznRYJ30tbxoRGFOhRV7md91RHiyWV82iGyo8nHy
ToC2MWg3HJdNxRIhximTm6H0ooEr87bI+i7uD3YB3gkYTNxsFmqnBZ0U877ibw3t
+szlDa1cZU+zki/eM3uh6UezViriDrOREaIdM+00h7B9gVKsBIBrQxtd5DdIyj1C
ZjiSc5ouPxy+4mJcmZqT/VxRi++IxLwQ2W02UJnJyp0KzFMTIxR6+AZ6whmvYU1E
uIR1pygFtfnghRSGsLYIo9CE6Mm2GSi0FApUH589HA0FE4eEZFakNR5wKZ3K7TR5
DJQi+O+0qBLhukPhv4fJQPyf7wWs+Jkq+XtKx2luSl9+tIy7XkViouY6zvPAAL3H
nBXTiRTEJMx9nZQgL67BZSgxfm+4NiUOrlKU3/eGhhp+c1bWDXwqS8bg4QlSb2ea
KCQI2agQ9yBklHNB1FmLbrpSVcLhVoMy0ZmYc2qmNc7cbig8NnsFboa41UUit3DH
ZRZeL0iYhXDHF4OnFHlcIo12FpdpS+vBIK0OQDqwGPB0QKUGiIacdCQaRA1CsAOu
LkVl3YXaH7SmHzHcerZajc4KpB26CQngOemDwvlNuGFCLjMkuKjWamh28w/T3qS3
8Nzw/wK8xl93hbkO+5FjRRn4hJgFGWMSY7nGQNRP37WtmVmOhy7BXlzdTgi9sxkn
hZURO48qTQWAwcGJh2W389lEHmeYeTBzkQYVCSNm83KQsfMuAvxiUxg/kDYqn89R
pQBhRhzpZib3+oSsW6IraeqnyPZ4Xv6QmoBpjgpDE+N6fG8dXVO9zzLOyGXvQOWH
+E2zaHjjU5qD/bhv5md1T77Zq5DTYMZh8SFmj93UUy/Cwy8xEyI2xDSUCl6TYqPc
1J+AAjiCY9mRe81Z5q4wY6BrNFcYMl0X0ynTdqme0SS1j8EUXldzoYZ4AMNt0Cq/
xrbkTFnc6gW6g9/+YRNowY21/d4lUbltYiegazio42D/VE33pzFKV15r5Igz6EAp
UNoD/RbXNcxpAz1BKok5CYE8R8D+z4MYQ0Q1SPZmJwQgr5uFjnGTOjC+bzZ4aMyD
Ef4RNKTiV2vAP8o4Jvjt4suup0L8zKXGSthrY21RJEIdwwGf38bf0KMq3oltnaZT
KHphwg5vG8LtW/JWK3kyUfBdNVlqdljWwkkq3g7UAih3+qvej1NaD64CrIwzh2si
bezYqXO3xlz+SlrdxMa8BU1YNr2aR4jNoLtNxgxRBf8mor4ayKTAylNOD0yTalLF
eh/yab6NC6WeE/qLsSsIA0FoJLwTO3XSIJLH9AgKbXqohGWt84BTNzSpwH2dqH/S
swIwFbLP4t8LNzLPXaUfX5XRxdcY5/RFoIW0Fd7dLuU88HN1Hf7IbspcZpUOGsr1
FbxZBaJRn6xW4bg9Ame8xgu0lseyCLG15nOm+Q6Lmi4g/0Nu2luUyGY0I387UNXy
DHMtrl4v+c4UKPKpXzlIHmisJsm0svNxkhMq07LBqfapYO1iOImxMReFJcVaGbcG
fGyUmNtJ2NCvEhNl4Hb/1G37k6/1Fwt7EJO3RU2yN1I2uDliTFMbOTIdH/y7s1fo
K3ZC0BTzFAUR86H6sh7ZZtSSnFZb0s1N3m8pPUAoVaNMYERfR3qG2gDV+4wVaiWG
NCx69i/56ohWpOx6RdGd+aGR3WKeup7DCMBsfuou2QkHxQYHPa3pnF+Fdnu0Rn4M
UH3ekAJyFF4npi7MqZx0qg9OWiUCp388G7sCYSVHXafXbQNHvOEHvVBNJF00UB91
Vh3CbKEBLMJv0XUeiIICoEGAvu/TZPBc4Sn56oCAd+l5YqlaL+gY+h3Vw6fQkw44
/onnfYQrt/v/PD9Ljz+iHj1tulV5elsG7hLRtMaZu09tuBIHK0M9TcPRKSt9bG48
`pragma protect end_protected
