// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
nTmIN4ZVa8N2A+VDVKAiKS6+4EFgqd0Q6mGPE5raAGsqpmD6+0pQwEwb3b17i/XLG4k+5WUN016U
canV3pqX7dgJegyxzYoH0XupaE4lsz52ou4pjz1WAzi9NLd2Kdvss+yGSfx+qBw/50XYnqS35ogP
rq9Lr/scPeKFGFQtkge8MoKgzJwy8z8wGAvBP432PqG9RGoWPWY214Vkq0PpvZ7bFGKl0xQMXp+F
ppFqerUhEkcuPkstZJ6drhnKqEZ8oeRceT3nXE1dXbuAGNXFOB+45DQcmqoZNtxy2KF5dTKLkoVk
W5KBMvzWHzQq9InbJwwuvicpKcF6JUlM5iGszg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9712)
qwEfONf/iOmNj9CD5Tfuoo+yh9wJUvJ6psbpLNyqSA+rRBwRFMVRbRTLxnLhfgFysEpQi8Bnqq75
Ri/RbBVPWsUQQuxqgEuWlOlB4VCkgTQIkdR7OTd3hWkRBQQ+P53KXDROfgKtREMdy7fz3lqF7yS8
8HLzV71aVptAzhJCkP9lMKXsefwEwaSkzV7CqZV+RRKAThxAbQ4oeo2lr1FwprPNlYx8vNRqb8Qr
EDUrtdgetJPIYLd+KbTw70OSb1ZdJQkm4rSkPqtFepjG1edw4G3SXOChbsHqcje88PDa6uDlHDBp
wr3RB+5FRja3vFCLx18F7iaXIpjM/B6ChafhfeNM6HbIHVXi1eGZGadVepj9Q0yJ7mnSAzMDfhg/
fy8IuRjFDbZIwyFuG7GStPPdhCunEvRcccPVqsatFUgWeVAh/lqosdqoUTTIFgKlykGg2XTeZroi
m2ve+bpCD6tWragXWCGjN/BjOGJmaq2eboE+ZYTVjnggCF+NVYhaJQfvkxFxAHXsv3+Z2HcahsZO
ttUrtWIdnxaEpBMNhX0OAVLsMJCHjZ+cbHFtyMbCGlIEdkvvzcb4PNSg8/AiXeJZnQi1W9s5UtLX
4gmQ6UDchBS1RzrjLFXmMYePZvwvke+ZURRe+edfRGbIm860XPpAlc2b7zwdvF1XC5KffvPd5442
UMc6xr+6xEtVn865B5KzdmIuQejlX7Y/Fv+WVwv+3ZfmceU/zPDv1Vajo03Frjth8hFDCQXVZg/2
8PfY0XsjOWqeLnYh8hGotiAinh21LyNVzxIpNOo2oAAmRC/pC4OXrw9M1vEQRKeyJweiuiJs3u9m
UOrY8uTNPt4ZonFe05RNyANqSWAoAKxM7FFN89kDr++lpWWNnKyIJBwzgkqwSd0/mD8wfe98++6q
YLKXJAl2xGXvd7/lSwnvz7a3wgX3CF5zQj2nNM2Z6lctG+FYRHKENGP8q9EJO+nyirRj56aWS/C/
yWe2EJSSNRLe00P/iaeQpiJ/VBeqrCRVfg2XjwPiivcvH5JOlVfH7D9so278NvLMOEnkLleg/iZp
VOq3RY5SvI0ix8n2fpX+5+6cJjpmNIq1xCpklIuUtAtJJ9AQ2OB8cRD85nNNOcQnP8uJdD3tzccr
YOHcBro75wK2RzmbMr6kH4JSBgb3i/+z4LxdroK322fHf6OmJn+22cKZUtx+cbUcMN5gcuQJPPcr
KfsssHZEE4DOUEAZrM2Il9CTJeFBqOqDrt5nPDdBtCmVopem2+GX0+Ze/s9LGypZFVLq+KEh3hNl
En8axb1BazX39HUbLYvEdy7hY1k+m/Vmdpz5CN4/2jBOQ2Ix2N8pUo5mGVnAwE5PLIcgrRiui55X
qnUc7WMKvlXrBlR4vkF+e28vywIW2zNNjhxs9M54vwHu+6wUIzRyibOi9wRgyOfZqDfRqqDneFWu
0jGPvL5TR8kI1GxpEjIYo8C6KN+wT12W/6mmnvKxY/wLqrAeDd78pYUtVnWJmmbuTJINU6ntwJ/5
1F3/5ccKvC1hOxZRKv+1kbzCsDUeU5aqcQ6q4V1+bFfIDG2sbJm7hr+WbrlJvGwSLoysVmed9GnY
wgWrhq9cYHSBPjKqg/F+dD1D6nsu9HRuaMBw5cszw0XisOxkX8YqzYrz0oQCpXb27bUaf59XNcla
oIQk7FZ8WzsIvplBrXccqEhHDw0Vys2nNFe/CdBo3EBVqeDzjNdaCeI+8nWRirFkCP8Y6TG9HLxT
BYRdNCSjkiyHeocQLPUcDTCTfKJCR9jf1dJu607zHo2wOIcHOf5zOQ/1vUphoCe2/F+3fN5lAHiv
xCLdpHimHDwZjlZmAfR/pnaFQJOjbRTCZnq63/gDMhh6ZMIpkNGNc9/1UejNr4wL+RuahnZ7gYrT
BgeHvkGrcteb9Ak+KH0K2xqty7vyHaKtWqaX+iegpWBtUUcjk6ZCLrwK98nNvyARVCv0ptdVPEcp
qap/5ehklnaZp4IPHXj6GOoMhGsEM8SbxRzYNqt6JEjQ1j5nqdzEil0H25CmGr/R1XaycLfH12bc
K08caBfdLMmnlGAPABvOotWtwd9qcX0Ia5hqrKE0GGJDweM+fnzPiE4P31ESip/+1RifQaB0AXH9
utz0r1Nl43Kgk52aAuVW4NFK3AW3Ww2jdzQS8vWPdvy+9as+1wuR/0DM+VP60CpM1tEgVrEfDGSd
bXOdWpgUpWiz0LnrEOOH0R6Xk6Y7YZhXWQx7ImXSC75lUI1T1fVLnFgLLZ2LXye7gWQRGGLWawKG
AFUlQICa1er/lpQn6IzJjN9kzcK1yAKscxChCq/vD+v/MXccRHYI7b6zcOQmXYyU9ZygGr8v1Q+P
uezRxDFAh5Aqhqotob3aF/9AMbZxy9hies6SrVtccjl4LJ9NG6mYhlazq+5qetqUkX6VDJynH+Kk
L0OGxIVT1DcNeO824KsnzL7QdQeQ3W0eElD3tCJYadY6v7mltZ5C+L5/lSSZFx3G9W13bdpC0LtO
EffDwt4/G68iZ1HX+hToSXE6Isv7DI2VMrM0ftZ/Ug8Cg556LVg/CvQ5lMpQcz224l7Wfwl+KN0v
3jn0z/efyWqimj+dSSlT3NLcFqTBL0VtEYaG7eg3tuUskBYNPEQ4SRuR11A87fN2pL4gAbAn4+La
BB0+/dq7FNY0ttbLLwB7i5YpyIPmVQhRyAC7WwggI3TptHzLJ6GHJY5UAw34NhjoDB/Za6hPtjxl
zX5jOoy7fb+Prbd1smAVO9A5Z9UP9eiPXLa0HSWt0KfaZTCfrP4jPkbWCLKzI1aHCH3x8EuUACks
lLOvJjvDZUF4LGuWVJjOWH6CuJAnQ//K0Tl7zRKdSkHWVixUXO/IZNt+BPlvPHv0wG9Mw5YL//vD
GpBjS40eHbLY/NDwzvvA6AC99h+qEs+J4xsoMX44D8VEx9reUw0AIk6jDbzHahqs0o6JMp0DCSTO
iQQ3Cw8Td+kkKj3BOETSuIkAv1nAdI2l4gHhVtHRfHTdMDWqo+Ic7M5LgVr7Y0pVE/sWJqmyhNEn
vENLVGoozndy9Jh/rZRNVI2FtbeIWrorYLvtACXlgRNhlmbeMu4+7hQsPU58tqiW1pBdg101QhW/
LrqD8fw8EuvrAfVTCCk/aaBmsp6Ubf1BzV94IlZjveKfAZ1Pd4yHjrVKKJyiUFQJWTVrwUcW6ve/
3/ATEiEGn3E77stVWkl4ybINYLt4pRdHijlu/ynvuFlWXMrnEbDwNxAFrklVY8I4Cgb2elIQuLjg
V4T94LU7OaeQwrx1gyMVySneoh/vL94zjztv6Db8xS6UToFMNRDjX4tXvLVOI1JO2YMAZW6N8WDw
YwGjG24FI4zux5dx0KM1tn+rrVKwWxJxMg9enuLH48/zBQWRsJIX4mWdr7Qspzgv7xhR5+aDdCgi
xogYbagQthFFNfelHFyCA2hn5W6nwRRBzICIvwpaQS5KitNi+Ao4M1d+jqL7yxBJP/QoPN+Km1A5
r7mLvdQJUHEmd2XlI9n9wE6IDILc81jW509j833/1uCl/cHE88abXShL0yu47Eh1gb3SsY4Ir6/g
oTbbkdu3JnW+UM1UM9cZcukgfMXPCya9Azf576UVKxv/W/eQRPh8b6vkychMrNv4UjsMa7GUgepO
v2iumk48lBs4EVkcmosbnda8tBT++jHeIfTZa1rcOQgBbLgIERj7iBL1C5gtMg5gpvK9/p6JUCRA
wkEs8DD+9hR0EjE39OFDmUW730K2T68VGdf49WH2OUQ8ZouGSIQ+of3Qky4T+RJcGZzdvFJSC/T/
M4chVCMjP8l8prxVCSHA9NW/Q7DgVyQi8iO2akT9prXlyyviLs4OIIvUI3AO1rafxxMyvmTdDp9d
STWXxnjeo2RL4Fl9EfpMrV9sCbotjU4vrXnh5hdiat7Osk4leDauNYQNyiPno8VxoqQiKcCsR0El
c1Afk3+8y2ZZnJXSN5YLf+6vh1Hu4fHYW93gCdflm1AVMZ8EqyNI+enYM3lgJfnp+bBCn4Z9NkdH
NREZh+jEO2v02MsiX07ApQFo3cOhxx45aFKxd8kN51is6Gg2ZUxnKDKiED6sBJO3Cu+SxhP7+xvc
5MyKkL5UJHKXxHhR+sxyXYe11Dxv9pZcWJ+gRDg0QSHGlEa1hlnyNidZV1Mzh6Sb5KQx5CmvD/8F
AKdKXYycTdlJrd6gE38qu0XkC+LFG44XHGhj1Oz4qgosSFhzqbQslwS6hg+RlTxKYqXC+odapICu
zaQXouiFIIYuKzJ/H60/gUprK/FECCn+fUPra/QcP3jAFY6U2iaRoU0A4XdeEpEBMW1SZVoKy+GU
v1Nce4yfKJK/eT2KtB59udKGBE0f5aTaF2VFlLLRVxtQjN1euZ5W321O5gleP/uH9u/JU5iMq8Sn
Xfxgp1NUaYZhLpZMeWzIv+nwtw9AtFUHrIDxLEEyYis6MOnBFRSMHoWbmAJaH2ppXoQ7NeoluSZv
TkdXw/2Oxmpi/w07sHMpgsW3ogMLTZH4q4aXmRLABoSFD2tCQrUrU0Xc2w9sbstljyuRI5q+ubo7
x9niDU2uimttC7dY1r8suBEgMpP9Raz+af+cYlGGpRFZHXxyt8+TljBE3G7sgp59EAgdy/bju5oS
hXjon6cXT2oRXMJnPVmpfREIw8B0ilqxPzXRYLnLS+gibF8BbBdPjKu7Qu78YEbTPDUYe2+92mxp
L782pwZIghNLQyfbB9FtoKp7CrVV7KsRRhLDMrOtD4Pp+q3F/ewWFRnbO8LB8o31Wgad9y3qjI94
naQi9txgyRuyNxReGHhgzsa5ld27uiN1059faddetH4eeMqM7QJE3y6eRRyPxdg6fSKt14qc/IU3
Ie3QybfgFGS/qcc1gyr/yrsOuiNgwAXiTeWLVPEwo4ZgoWqvHGfjItniyQ4Xu49r4LwxnPP0hNYi
zK36bNJbU7eKrJQm64Y0xDI7o1IWstzewwigbidzOegHLYWQBbAmjpX94bj5VK9HRcrsGTTBSP1n
7cVG26RXJ2WjKMtfEvg/jvT6i5PJr6fTYe6w08aFPQ+5sKQIoH6evcRn1MVl/63IqqFEZevLMwCr
LQhidOA1BNP9YpvrssM6et+0dWRm2Gim/cd1mgC0oE3N5xO5ufCghjQB6YWmbX1O4rFYxUipjCbp
+8Ces1MkntbEZ1CuuJdFxYmYd26jopC3PjP+A8nreS8w+W0biEP4bvS1iFs2K3xZvr7GtRxuw74Y
9o/g5u95k5FnfHb6WhpBqzlv+R3W7WF8dKR0vpt8uBYjekpx+s6D3aLKumwk1N6ASkBzgnZ0phqQ
27aGjBCQ0dnlCmvhDCNhYAAv33kk4nyCA5KInt0aWvOZlRq2OmrJ6udqyMhv6dTiQXmLnGmXek6w
HnwQgjbzlyR3iP/ewNlDsbfOH2IM1iFn5qe5SI+u4bgS/XYePVOBLtFP03Ejh2YCM3JelZBElON7
Z+87itUHQnvuW/fFhMQoiwfE3SY1SscmA+JfaPIK1nsmt6e2DK2eURVzUYH59K0JfjIA2Ksp0MBJ
fGbFqUZDxx8FnLFuyhx7d2LIJCag/FR2z9fptqfxmvtR8I6702aW8c0159FHZEggYKgcJgtj2iP6
ADUC+/XHTx5qUhI7pna1+MOwwz5Re7cVKLVdu+2+5sqo9Qc7MBxzEjifSFB7Pbcgk8qb0Z7y4R76
S14GUi76+ReW17jso8ljr+ocmeafREVzhxhtiuB3jYEOWpu7LIOTeqt00T1tYFdUOQA2HEGPI5c9
W7RJpF0UJAkg4IUeCRG8cEu3N/SzNPt837T4+qSPCJKVJee+y+0jq9R3hiA1SORgdVO0FQDIHCWG
jGgDOvBfOq17IomE7epJtSjch69CXrqSQwrJKnKk6CYotHRVDGEmmoJGc2ymQWi+T1ftmO/47YCa
mvHVLE61FF77p77Pi2vgdLel/lSH/jsE6bBK7IQEy6oFVyj1VZ1dbS070fFnLSpv38C3Ofn3dxGr
O1vJKZK32p2X+g6IurcB6Ntk9X/BMzjxf9s/Dq0A9LeWpxuuf4r6GFSLGlIfbfmVxX7uaS3RxnWP
NvZFAJsCZUcB5b6N6YEmtBpJ3FvvoCyZ5StPXF+oDkLBVy/lc1GefodQdPUXbWjeC+asPCD89dT8
vbn+NK+dNWWzB59TDwhc7oUKEPp9Q/WusXx9MVKXe3ljXt7SrGKRvwtDZ5eMfdzAj/XPaAQtp2Pa
yaCRdgu++sZlPZgkPHjUyw2ZS/dyiDc6mONjdjxFgYuF768l1bYpgxF2YZgYFAEopyteLGLBcQCJ
3uDHa9dvW9992KNdt/LF2sDsBnq6nuNoyieNZVghT/09hFubWfVDxHe4xynJmp/PNPuzTjk+bk3t
4TYhu12naXDF2gjFMtSQhORDdDLNMUNFweU0RvpcQzHA1vre+PFlFIw0GF/3yfFN8dTnzLqggQ2I
pu0UjjJcQ5Q78UJKtEW1NnsoE2npzGn53tNkzMHL9Ox51l0fYxg13zApqOnxYqwc5eAPC5YZdU96
sIrUGSxshShrsOLKOgExXgIn8bRJiZYeTzj6jSh+t7B27LiTUCvJUuxylHIGRNh/bld7e8hoVMBN
5CFJxPnmx1k+qkti4JiYLy0PUsPwuR2uAXKI1j47s/qjYNVJiPtw59NYCN2d1nkAXyVCZJsm/kWn
zD+AcWN4DoHuh5BVQivLtsBSaXNO8HL4yIUWr6l4RPfSpFAs29xvC0MyQJ5kAl80PNeqW07zr/KM
4EXxKVJtj0UUYdN14PBAa/M0r+DQtC9a2upRzVNY/MuCsnZl/4zzu1xSBzlOOYpytBq0Ao4HFobt
HcJSviiEKv+22BjT/ii0IJDbAQXKfZZsndCk/igKlvYoKabqg1s4WWFe+7ErlWaVc/vy0GM+kB8u
0ZGYes6RIOds0jkoHztvRhHM69l6JKTYeUCbCms+YPZpyaSzRan5h00Ps2hTKGp+yv3RLm5EUNKa
BIkwbAw2+H+c/mSMyRqiDPH3MH/CSwJsSBuOREbV2elM1nnSagLTJqKlFnJpKikAU8BtIGGqWyrs
UHDWKRxmfhhpVfmCpWub/KknImKryAXbJeWXP/MguYIgwy9nvNwbgyFZEyzbqmX2cFOMLtadavvG
5dqO75yTH0XN9yFbSntpTrI7c3zKYmSk6/DUih6MH0yS02EB690ecU1buaj48QwpgQCcsuiFy09X
M4dIPawEirXaDI9QDYlq8zBICZ2yCgXxwplLD1nV3k6N6aiU5ecNA9mTPI/Qpgu9WUkocqTG7qjV
RK7oqOiZu2T2PdVZCsMezA2c0LikPq+TAhnLeNBeMGg7OU7fwZUosCviU1CUjHpzMcN/9vNIIuXQ
OGx7KcLzmmA3jAqCxCEYMj3d2hBxzv8hC1BVDsLXd0QL/G8sNMLAW3bzTwB47FdV+iFNhYdLXi9D
R3oAq746qg9rlKBgfJqZebkM6K9gy2CF/2zo06kwbQvxY8eAFy/pQevo07mF/9uVP5khKR1pXip/
IcsMcyjwfrzlMWnYZnUwYZwwOD9jafZa3ToGvaV4lOXhyH1a4LSeCFT0IV8Ea4Q0e70UOWKSKcD/
gEVHZcxt5tGa0Qoxa91MRkCB6NvYhGFIpc1WeMxpo8NSqBl16ea4qMvNwl3Dow9HfRYEBOjsDJwx
lQNXbEurRmmZv/6RV1ao1Rfe8IsbxoWCpHLNCcvFU/zCP/fxF3pi6gqIlvMJO8xwXL/50Qnggyv0
brsHgd8jt7RJrIg88tDv9Ai9KCVP01HHMTrMVHYGkt2TfMs1XEmQibKRiCNV7x4kw5cqahBYWMx4
IHrYmJCnUM/AjVzbQIX7IlZUAFvlbIIWkBhM3lPlYe2ohk6C2On6HSxE3OaQjcOHqYuutdUAARdT
ABlTTAOI3j40vROy5dHMwxn8VduLY7Gywm2bUdgWmazJXl2O5dZXs/Sg+Qc2RYAu5MML3bXjFFnI
5hOGlwynHTRIIuYEyklOmfK4+jUNFuvbkoIpZbvMk1DZ2UNOEtPzvP6/tkQDaa3tkYGf4TrP8eU2
N6Ob+j2MGFHTc2z91Ujh4pGbzHwWtBfQJ3uN/C9GmQfikzkWBDax9HR2ctBnfU8moVVXTx1pXTsJ
g+Qi/WB5StQdKvpVBSTYxYHdngDIqrcvRlD07Nb61f3Q/h4W7v+a+/Qhk+8aUmfThEqCFnlErbJF
bpr+1TEgqJItVOG0LlMb6C5FxfKjggAOrL3KB1hPhOz3oyznzQ7JQG1dzmUJB8HMwSDx6qEti5LR
6HovSipX8Z1FVxJSkqrCf0f6luvcnZ0LCVHLKnddzlMtPQrdmtJk8fMwwLoTMnFsNrDPXpMNFzEo
perSOFcsmylENIzgIqVucNLdK/U6TNo8SFedZ4RsiAQaDqkaLH370pEdX+stO9oDoy7saFhya1zQ
sEUwTHGwv7AAKYhV9TJO3kTbNLA97kTzxUwAVhz9NOj81CdISfoBa4w/craMfPKzh0HwBvBLKgHU
xgaHr06qwEzap438LGkYMKK1oywaJ9vZshfEq/ts1qNKhUU1mXpKk7Z0fRckV+Oda8h6IzUZBZ2w
mix7p9GUitylnKk17DlaBhkux4dF7UaSTMKVwk461vMIc8eTpgacmhO1CKue5XhJ1FlqphnaqBVJ
FtDVyc8bwSsSjqUElhhq0TVjk5oyAzrSwxaz9LCexnV575ySg7fjirB+Od/5kBXWrJugmPAeXTbb
oAKN4vjXQSyO1qnjav2/VIl82bjkmpHAxzxULpJ7gE3F0tsAK6XOh40SkCnTtck7dPnxQiff/Zun
faNCSbJ1OCSTUf+6/VxhmOcr0a/7J7I7HpmvNFS/cwHvaihsj77/YloC5jjEX0QvJGDLv4a2tB2b
K0va8pZvP+Ihwt9AxcV2JUYuL3M81IrVYCrDfQAVW+ze03m2AqUYp/FquBeuia2bMVPQdKcn6MsW
2TLwjwVTewrwzgxQiRuJh2D2aSI6Ja9nxTtw7h7ZzycVUJfHnm20BztYsmB5wlVr3X9DL8JBW6Z5
I8NYrCwFPGEiLMzpqRh0AttUXPf3KdWOscVsIqMTB+UaJPrYQzfTAmaKUz+gRlCS8HPNRoDzg4uh
0niwmMfpTx2o0jpmmVhQB/jlPFKC88vQlrQuG22n4TcDkUP50SKx8a6qLHBcTIoLZiLaOEGrYIWm
wEg8AvgyNm78i4PXeLwnVFWW8pJwlMQUKObs3nqZmy8L2vDW5G49MYilVNRDlRWMAspjjgkXbsV6
uiNUCxB5JKg2lWrwV06bjG2RzE9YJ0XF1UMhISiSkklrO94rlPmj/+mmVx8M24SntKQZez1inqkC
W00IlBqyfe3a4HwnYUahArhudIalgnsopTQp96OXcyQ8DZqDReCeXSlKUro12pZdOa6Ht52JYBJ1
EoxqKrd9mEFopdnpqqkExpodvi6SoQ+5ZOuR37liqtPmxfcpEkj4CoJyR8BICTPquHD5iP3jzcjM
DjLJQ9u3+iLuLfManY/vBV1wZqIs9IopB7ncddQZvcN3Ji5M2cM/Kjt8yQI0i7Yv2g25/DZgpTtl
f6FWOjdB+nSLhEiUNkgQ6qrdQhA1NdwcuSUhRjg39P5ZLwpLF1cry8pu+CvrixZhMDZfKx5pr8KZ
u7ewW8jy5FKH/TcuWZySLVXLF+uQgbAmgMpdIVB0FZTs3SLNVfpojRBESerqj0WCtxs3qJIZngJs
mSugtbtKl2ZDhdl0VcHUyHb05JrGmuSKpbBK+o9jlLw7jyOCRVckW+k6YQn2ikuuWa4pDBDoOkkr
XbUxKx+JBAX1TWZwhJBB3bDYaFW8kMyElMth5ioTyHDAZSQv16c4CBxZ7aKcBpmYr2BCkYgmh9hY
VwZPXHzZbJpMbwiYHKNzm1lKdwEqC8H3Y2JQblvxPjZ8mQWxjvSAbmdUXROEv7KMz/kUxDdxgdKK
RQ7rumBY7icSNVJF3+QQQkl5+Iae/Nw5gKUYEvw7Xo5rm1CGYaIVbqJ27aPT1g7gTJ54mYwN4nr/
R12p2BLqk0ujbiyjNlm3K+ARvYrMF9shBQNec5AvfpBI5XtwWPBgHfKqVTE12SSlaYPGsmB034V6
zadnbSUMtEZc2O878BzoHjAjsNX+ljP2yXMz32DEiwrdQt+7CC8j0/jfwfIfulIJhM16icI0RAdm
jTWcKk8hgU3KiMtvNEqMyixrFS3DI85b8xjb82qVMNiBxrkr2EX9Kw7DefGHcaQWd1RFe0GUnMjy
MVamnCKIpTymQb/hDBIhEHzVC/zCgFb/fokQMqSsueK9SgEyONze89DlsauUEKJBA1BncH4U9ahI
nYDz94TakKjyLGZC/0+iPdf3/oUTLVMG/FvX10vxbYdmillXn9oT51oXI1dsX4F/yGSHWSa6EpQd
iO3PJAxDPfkw9ZE+lSacNBbxjBQ/5/Bqsw3AB3HEE9SLqaIj7IfK9loFKNcdA2uk8G4aL1e1x9bT
Y478kgBKYzq7YfPaXN/K37Dyd09GvQg9xXA1kn40ZFVBYSrbDERZx2XR2hopN7Q6t2YC7n9acVlh
VXp5fajycXiWz2So7ZlZNn7UzIrYhcVEqKrLqzoDGPw0yDhi3gRHJaVFXyIAiaYOZxZ7/qkU9D8d
pFUlOdCvzrNUGx/YxTj79Iuksz7h/uLO6xAi39BURD+O7quiEeSinEoyIIuCRumXzBoulr2rvpbU
3c3941gYrV0HMblYkRzWjR0Ux1Jz4qV2SlOSDUkiBEpkHZobDgU6yZIGiTn5DH4Qi0QcdPIJlmzw
8YOXXtG3gG6srXxNXMcK9N8JFXkQqzStsnY87VSqiBSoKR13HQMjGMhrLhoCmWwbhCa79hBMv2Fp
ZQbWmHAPZSYGgronemY1QIjCl+EoBBiMqiWnIpb4UllX/HC2OfiJaKriJHgGgOxcUpztGO7L+jYX
nzYlAujsJHnjkZhyk+/9f54XB9MM9qFqbpa9Biu79WU5vU+7slZ3LWBf1j+hMWaDCyRCjVlMLevE
hhRUrh1KuQheqGXa9Ip/Ve0YH71j2Twk4Mfy37LdLp+aNMuSeAStKk/FZ6NW1n4IYyhTXmkt3nTb
0a068KtvcQMTlxN+/IDAGy8RPOAh7JnMz2tExA8t1hlZgTKk1Czj7k+k5T9kh5nwBHJfydJmJrxw
y1NLSye/7iY/UqzVhDvYRXnQTLiR7zWXBspeCKIcfwWxZH1U0RghdzN149EYLi/ixu2eYFYWpom/
PurCQe3OnH1np6LKmoKGcbds2S+dqRx9REUnehe9ugQs2rO/JSG7jh/D2Yn/OTRIWbWt5mAL8gzD
i/Eifq0sAYWRciNRfDLk6ZVYr1aw/gb/C4x1iUNlql6TWg+cddyqc3BPQhWDDbie8O89VM2C2b8b
5z3f+0gjzjr24Cdq8a1aKCFm1NMMqn9MCrs6TcLn1TBIs2OpqGr5ghcqqCiTiUV0zXrLvDTwuhI2
SeDfNcc3FDpaMHxmfVDPVRcy4nBDvgVK2zD8Tmc1n3Iv/SikunAxYKFEshEJwyfwy+zxp8tDJe3U
lSK6lyo+UYF7I5uAlg6IUBEWzSb6Uqhnbo7fLAYWkcdNwOTlc4QA1xKUMxGI2go93gfsasMocSFg
bSUm0FpuCmtCEdW15DCdg+HRPoKd7LFHIlPCGQjlla0nr9ebWKIaLQ/7Z3LKtRA0wvalQM4SZSlY
J5hnZcG+h/F5AJVdIukhFn4M/woaVqLAsMuXEKZISjoKImADAodWA3yAZuKvAkJxOnlFiOiOYvmr
VyEGWgg5gXj5vx/WESI0qhlZz72O1iPmId+EoDk50S0cfBu2yzpNb6TnPEPUfzpcXnxiVBY9BEv6
hxHhc0nLbwjkE6o10TQUWqO+Ju5pDczxvt0WS6aJ4B79AEAeKEZVFi+SV9YCc6xAwD4/atvgosvF
jM14TFvb+T1GwS9HEc4sfolH/bw2I2gwyGdhZr9fdY52VjP5gwGgA6N8D/qWQuwewWgMcgZyGpxl
jnbAAUhvv9oeC1iI8cGaeMsmFo/EVouwqWobXFOgkIFhZkoiLE3lee2xJicionBtwAqKePfj6EbM
xSV4cKzNKvLGidxd66L+QtLazbwIfg7OfnqW/dJJUPgZ+DNXP5DSIEu6fVuY5AuX7ceaMW6K6e8u
NPdmEG5nKH9M27Q+06FhWuH9XTerluijrxmnpkEUOmHXE6omRd7TNsuriyQ1+/T5madsttTzbT8l
FJF66tXcnfsESX7YbJ/tg3FuccWlQHzYvXaA6Chjur/fnZYXrvzlfGr0zSB1RLfkiVQOMpfuT9h9
soQas/3ebk1Pr8fXvt7PTSHyFHUnCGmh04G1DPRnWGzSHQ+7njSGSqlTFJDxJiyVDvNv9CsKvx5p
93yYSnwVBmS4/50WNl8NTlVzlRDO2AXXnGdeqBaAdEgJb2UVOflQoV8JcKIoHkRgi5ewD5kALz+v
AGPxsmXyX2mPecGhZ+m1Aa07+Pmt5wLbLBh8xVYSdcESah0UwGi6Qrss7n4tpCQdyX0BlKxV6dWP
zlnyw1t19XVef784tC+0UHbLCLsIppCPXg8YTbbh8JtZoKDhx6tg6zd0XhkJ/Q9YZgnu85ey7oTi
Ysog+hKm0VhiMp2eTWyjVxE7X3TCy8jyTZIbvT0V/sj1dCh0sapL8YKYRavVoJygzgBDsdz2KDgv
LZlrU1UZN/48NdXeicn0sOwZWYjSQiI4MmMvEeqVbs+M7hvoJXk+k9Wv1P29sZ5IB12ZJ5Yf+Knu
6pIeiLtJuaVGNZYD3Vp7PAkx+Y2IoWYrFzNZ10KALPu0m7X3K3PAvsodcS+BZOBOzIgy8DuY5wWm
TaeZnDukW+3CbxU4dkV9Eze/G3IEgQp28Sog54d4LC2vqQvJSr2oMhtv5s83/gBUofD5NE1NtJvB
fnQjD3PnlY4LE+Vf99O78ODCLmhawg==
`pragma protect end_protected
