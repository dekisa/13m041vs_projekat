// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:59 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UupaXmb11B6mDVcGspks6OmPu5w1Hx6PLrz5AyUAow9/3H5AvCVijcdjgyO/cBZr
yZVBULC75Ytxs0VvOR1GXc01FXLhvaO/xRnJgiSDG2hcO7T7yqPzDVn8TlH7I9ht
rUq/2noCmkmfacCzjj0ILYdakmN/o1w3CLp4zYyaTbY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42544)
i9B4zYdxPwlZstKWBNqo8xZAm1bEj4NBpD0vm0xsJxWhQx1Oyx5i+xS9Ve2sFLM+
+53V//e35QyLfRQjsPWbdr+BTHxusyUmygBSWIBLlVUuWW0ar5tVMCICKMBMJ/sr
IcVPruhGD9FV/OE8nOwNu0E6IaXoBskVLPZXal+YVuGfbFejdCE57Eo4ze/gc4QH
95WttefVf06krhHTEeguCdIJQTIJXL7plN3AEaJHaVq9r8XFit4zYoJOq1huhDi1
A1ctgPEz1DVWsfm/zqeJsE472rQUXrRt6GvjgsKaCJLmJzE8wMLdrO0kF9oQZnFm
Hi4H+4z0g7+cA7IYWMWb8VjmrWm+nqp5kMX3huoO/8sHPv05qjmo52U5uRKYtKOW
5CmZrhIky2xjSryveJrKT6RJvTiw3gVgqFlwv8mEK3od0e7N4GodweE2TXSvMwNq
5Idlo1vzxJfX0ZuSOgHO/SNVlRqcUyi5+AXtO2Qi0xJH7xmT0PZcNtFwED7RqfAl
MSHDVMpY2Zn63vAjNlLz6HhfNSF1VNX6AHNPosnsb3zRkjlzlCmJ5JMs6p9hWBdo
GK6OvTWtfs4zueC5v1u1KltAbtxY51SmUPx8NeLBL+ambO0EUf550OgLk7CN9DD/
NmrlBRNYVOXl9gAE5Wec4ofcHQJFgLBQ/xsf5bnrS/6SnayRV/gs4QjL8sWIAkJy
4xi/NmWrHmY5wa5PTTRrdiwecZVLHGcBlfuiodFdAgHRblD3QzeE0R6u/Q5RO9Y6
K67WfZHE8ekExmXKwIWAUOnMNC/ZOhiFlFseFASlRTrtv06XKX+UhIAKgNWO43fO
QyDr7OjirxmDQCL2tHD/pVDLc9ynrAVYQf3lzXyUZggwh8k+U3Po83D2pJdEmPmI
W6JX4T8liCNVqdT1H1jsj1y/qqmyEdl11qPG4JrL7/iMi/G7+b5O3vreAIxH3g3y
dg1F6n3RJWVtb3CG2RtKzHp1HciyKYijLZTBsiHtwW15t2x+phE0CnR72PERK3yy
iyJJ1x02gfkMHdJerfrxRUBIZ9Xz4kDf1fApE0RrWOAZNMPRZrdatljUl45492tb
i0rk7fVv/Y3BnWvqgzIN9NdsX8bLDkdzGYFHRv3e0ZVuO56Tw4Q/4mFYQwvC6fKm
PwowfDXS/ESMhJZNdmzF5AslWJi6hOi8q1Lvp48D8SwKIH3OH9//D4gR4rQXjUjO
hOtYp7rjrS6nIxNnr4iZ8C1rhngWr8gE65kQ4DqhZLzCN+e/6mQVabIAgk6jVh5X
HUjgbe1tPg71Wdds2MzLTeWqGG9iXBp1hetz2iSx/r1w+U+ptvnj5+KtUtixqU6K
YDYH1tNADp8ohia+BaKgNwxhM0QgnyMcWNlBD5BCHV/4cV8TGDiRO5i7Vc/mJxCl
ltJqXTH5tB+mIjAF4NQtWHBcO2QlMwzKvJp9ob/sK6VSYklEZwU3jX2UnHxJ/rL/
9wErqpDS6CNH4UKrqUn5++Y/WwRCHp7td6XiSRZycd+mjTVZS7dL6o60YADOJ9kz
fzGsWdLnexTxkv2XxFYFwY/AH2lBhTFkG/eRgRrHwjFeA+Lp5bhvo14PrHgPYVSg
PhVzG+uzIZSZAy31LDiAgyBXSEax14dnIY1061SKfx6Mpj3cBY89wvqac/z19iHw
ls5gshbBgxkDmh3bZVHCxdtkwkfUvFdFkNGyfiq3VmRNyEwoYWi7EiBSssppUixi
XuAmFpUtilUESzZEreb4+BY/WYiKa00Y8SwLvPSFiQ9pdp3cEpjsVS4meQwrHwOn
5pi/RpldQeZvamhLYfSkFAA1FIh715dPEbuFGZa0lfKBB1Z/gXJWcFevAQVJupE6
1McE8pUS04mo0XAn+TmxzSWejnMcoDEpUy4sJpl5AL+HFlBJmFPhEDipi+qH6XKI
S3T893ZzmQOm0Tqhgl1fxeaENgQg0J2iW5u7cOr2KhBsDSpcymICvTnq6e7CqTh1
m2fK9nDxK/9jwGwhRcvELwDOec273FNYNB6/ATTMaROBACLUxMLU2R/vMiR82m6W
xOr+laQG4sv/KHfgkOwTB1g3bY/uw7TJsERuThwUOp+jiJdXYQZ/gxFYrUTJ53Bu
72A7G2g8gb9fcgPZcTEjkiZvonKFQCdwrKTVO8fWKanw0jgcQ57eXzzPktHS9k6f
tG5LeYzHOEwIyhQagtmP05c3SKwLJ7xtsnsj7I5b1uahslAOFYUM+qDXviOCM9NN
8qho317UlwIbjwMPnY6DPRJ6RMd1JE8i6Y5m7tXTT/7gU75CHqfxEf7Gv+IA7CHA
aJHiFft3UJ0QqU6tLqGk+1QyIBwRI8g54rm1v8yrsV2zEo8D4lZwEPuoRtYaziQy
zAfe2u1pxhrK+FfOQqVaeXxhLrVdiTypBqTB9iajLBgPwxJYNwiVopwdY3s/lSCq
WMWeLMkDJBdcqvQdj09mTNuNiVUuITzLmMh1hff+i3Ri+r58QPvye0Nqh+tHgSoX
B9OJC0sFT+GXMlTjr0czs/yhfEZjvsCiRM+sWTAkZhfMU+RPB41VrHwIs47MmCI4
2AYQRhIhXbEgpR5tuxakSV8+3m1o6HzbmxYb9VhvBTrcDyieTvnAgUTAQiDPpSoF
bHL76sFuf63A9n64AJEYbmmP9ClDfx9vQT6W7hc1epmns/gN1W5XV0UuaqQuaptd
y/DdwpcT1SVVPVxlsouinZKTVoIvlkURHPb6UN+AYnrx7i/7EzbYpbDxNKL2da6E
VN1zGqYdPDrIwKvJan2UshjaUi/FF4qpZ+o9tlGFELSP2T/bdCbiBkWg8rb5l5PZ
I6wvaMnQ2mIzzH3xgVLnZ+6+UvWEc1gKtlJbTnxTRE/b4ch3gJlt2bZVLpEH2L5u
DaHptXvoqf8X6qqw2QfhCel4bLJpdBFLu11PkYaMMRWfoBN/vkqcYZQp1v+f0NTp
heX+6LVwijVd2B4Ji+0pXgmLdjrKUvMDimg6T5mDMzPMHq9bL6pInjtaDNo1rD3d
Wy/7cFo6kdX6DLQrJC2fnd6wOywYPhyInNunQCPpXUW09Qa/neb8IBkCUlhEdZAY
4LkcrrLuslGdKIz329ARm+pCnJOpNcs/zRUEJMpjLnCY6q0qGUOELcQ1uvIZkXsg
7icolgyWzftlwNnd56MtvP0t+vWYmJmLZdB3EyhuG91c7gnYXZhQ46jTjZmvy15+
c9PheHM4Z7dzwoG6oVmBp8Mymknc9l3caAXQwIHK3tviv1qcNoAlFNjTvf1BVzQh
CunNc+84PL0LivsDH6JE5t8MaqbE9igZAKN6zfuorgINDO5rP09PmXhxazgB+WWU
5bW7dLl6KZ6E6Y6ZR4n7ZTwuBskA6VKhFvoA665TblANDCQpChsVhpXUl8nIzId2
PPl5h0BTU5PVf68A0Xx8nBr4PdiUuL9c/eBqthT7Tsrq9BuIiACC6jDwm0R0+dKl
bIGb6vXUktPgayiRsczAZRK6qy4HDKz8zhxdTxuAgOAhtiOgnANSUm10tsAlCM84
YDCDt5TOGHyvK/uqfAQxcr+N9ZKutCh4QJvHbcr3yS/6EjKE1QpPtng4Q07QjnyD
khq9EX0enrYf6Ylg29hivVu3iS1TTckK6KMRgtNikStgBag6jxxTxakPdAYGzGeA
sXr2I6Plvyafw5krkdmu5MNYzChoSYGnRlH+T3EmYKvSpO9MAPqc02LDLxmxpza7
XnwfYhJKAqvDQG4k52jMqX7D4yZPHMO0O7Gbu02WzorKqHC83oPZfmjyzdW+T7Zr
YUxLAKd+ks9BygKrxd5I1OO5YasS8tWbcRqYSdeT1TJylhLRwK4La8Fm8RiKpmkW
oRtzDZYmbKGIKTh1f9w0sTouL0SjTECATtl2HIfcn+XNS3PEDqAIYnUSlS84BKYR
ttf5jajTz3U62+rUrzdBbHltjw0+Lr+F52DaJxTiLBYgG2T+PEdR46U/Qg/Ch8Iw
vGUEfAeGkrkYH2qUZ5+uciNPkVOBT1lsmN/YOifcYu6GuEMYZMG+akAbq3ZKhBoM
ZOj8ZgT5ko7YWTS83hDwgFVSyGLtV5uJOZ8dmEi/aGt1DPXd1k0sK1MTvxY8S8dy
RsB5Bj1OTfJSjK+ZmVJl8VuP/SSj8T+zY0iB+2zf+GqycdvgQ9gGb/GR6N+OpJJs
8eEDeT/Ygp4ZwgQt0LFdV3UUZbYXPoFuAPtexlPOseV7r3ofH8fa7kQlsF/XJWfL
z594eM3I9bCKwoHs/AJgZygp6eoL5xmbprIq9uBGINAyM5vfH+qvqC5mndNgfWiN
zzQ19Zpirbnk1PIw5BD1FrP1xLXd9TeC4Xyh2XgmRvDS9d3p0RV5tW3QuVvr9DAF
Ajehf8COxEG58mxYxXm8WbDZ0MjxX8KjHFc4NsUd06hTaC5Eu123eLGTOZAqBxMq
ueEwtRsn8Z5RI9++LkaCigELtAVTsXSHqMOg2WjL+uSdU+zo/E4GfJsU8O7cOeyY
K2OCIvxbpe0vrP020JMH0Ry4NIdILkC1PviikcP0DEurhaUjuwjRcUWXVTROp7oV
0b1FvDDkF8uBvHy+EFyKMgxi85iiajxMLA5Z88EASciD/YfksS7dar9qvMbDk4ro
IumisXMpuaBvuMfva83sb+CT9cQ4ZEjIMW1bPi+z0mIJewnjXnlSYZoCRH4/wIVQ
FmAPDNxVF8VIlAXzRQz1JHAu2LrPWwmEvhWQXCVaZjemNWFtBsDGKP/q+1jTzQnn
AJd71cbQEjo239pqTBk3OCSy53iLYbszIiN7rlfGHDN8RdgPlcX67754C08yMY+C
woXf480oERCnWPBr3STg05Df5TNUQH5gRTy6y8TsAzW8oKsXv8BFqaH/h5ih5O60
OGutTI8qjwWWkcnGgWvOvnoBj3GHi/c+sFdZulIe2BsdepN2i0vxFAxgcn/DcPFi
6Zms928ps44+kyqgk4cDRv1kOZJSBAzZZzZ8TUzAv0EJccI+T6Gom+9Yda8Thmvs
kPjCjsyW5BWcpWBSSr+xnHGJd9s0X98L9vWrl2lLL88FBlGyQYwkn5ogeJGIsrOP
gZHaon7DGlLyUukFijkmnLpG3Mna0Vb09c9iuOPboQ/u0nEc7OFn0f/j1sQdQJUs
RDn+feW90tn/v9KocOULydl/Z0WLvp+76NBrGinwc0Pi+lX2Nn+ADoEGlyJP3C0w
7zkk/Yhu+MSMkPwFbo2CIm/nGdJCwOwpc8uuS8AsFK79/Xa/A4TtcUTpdIH19i7M
2SoDG6ct9yX5A9530INCheqqdHIr7bf9cDa7jyBi9Yh0/N+jFD6Si4qGURwt2wV5
iVbo85fIR/d5L2StNo55FZHH9iQaVX18W6OqLOL33+Nqm7o3lSfVNRjbbhpfVuwk
daltz2qr8V0eGroFN9UhW1kqSJa6xhExU+pnVbTRnbeclNeTTLoOEr0WD1yVojMz
wD4CZHqu8EbrI4eIdM39dt53YHZwEpcGvrxFzIx9TPgG3dthjvfydeD7D/AfcM1E
8v5gDVYTXzKBrtyOX5uSVlcT3GuSpcCwioxEHxPAdHzMxHIbaWxSoGc6nlIGgO1U
nDACoal/q9j5LGy4N557Bbgxbg7oNvAo1E3kJfaQLXvD404QSp5ADKE0glx5RYKd
1MGV2nfLdPG1H0hnx/SGhY7HR/NnFbdqVUAGYpzwiusD8rSp8+2ahSfB7ib7Ws6N
+xkO3flv2BrKM8ysz9OxIvD63kbr3BYwQ8TUgAdLHkSTe/oVDFZvq8ttqHkGi5X6
Mov45vRZNXCKsbKEkKf7xFRm1x49p7auTx/2yFpt2+/ehGqbruHHr4oqMgprh+Co
ptOtYoAwSTRAuTOQG2JaFAlfH79u7GL9mhGTfMIr4tqwgwzWdpJTfcwcEW1IkjTD
r6a9vmPU7yBLA0n5Gf7Rmh/kmnMhtXFJiG0dYp48IrcihJmduMIV926kFwLXeKFT
/PyV4i4DKBK4DxwyCT3w7wqd28ImnpjNgPAdpin1nnvEF4TjC/S8c+k7Ezw/ayPF
WE3jMEhR99+K1QbAOE1UB2yzZlAJ/sdspMUzlQXAFhD8sTkUZ9HpAJWY1ikKI2xG
YZyi03eGTcJtZ7/hbT2XbyCsiaacYBpMOxAAe1Pw6rqNA4aYF7H8Sl7rMz87n4o/
UVZ6nYDjWipEQaGIwxGtQvbqIRFZykFkDKlUepcwIF7eKKAzF80Ns+xQTtSTleu2
+kkn/D8rTGggTECkGpB0v1+/lTQVbyEjZI6LnbiGaCQNfYTSy31GiBT22MWjcDoo
JasJ2ec5T79esutWhOGreCS9wuobWZ75IirrRmPKTDy+AoIhnQN6cOFtDAuq/RKa
2lX48+VbE2LDDqTPx69eX8z2ZcDF73ouXbAjHtwBG+SuoPqHoJOsSxrvkZPlcSNP
MDhG/c+zdlPgIcGw5eY/xmsvqGiW8IHSyzJtbUl8INzPT1edpH+XfzDqjdqAwQfv
gQxmd/GJ0C74wmUQA/3uDW8eUT165Q3XVqAAdKOM0V7W5Pyl3it3VcF1etWY6BGN
nt/w+kY42Vjgwuf3KJAJ+kDWx/gbUllQKIQ2mg9ZSR7Lf230o9jSLPassiHWZaJ5
vRZGjSQ2WTVAVHsDcj4lkTkvVEtEZTaXtTHfCNnSu600ckkgYpBUI8vOuGwkCI4p
60EpTogb8kgKR/N+H/RLNc//N00Crd3E7WMXfqwuLBLvAhudPYeF0wx/9HLbm/yn
+teLT+eTs00z16F0Y1vfG+8oQhIDu+CG6y5FGPrFUR8l0Fsho3dZkERUbVsmoLth
tNGhxVsb9sL7atwuNROGhDKlvQkQSg6MihBDCKgqPTzSwsQDX/mNUfvM3NGFj1d4
9Yn4yvvOuuFmUIhiH98fQCo9PksDTDCrp1/R4uAnqZN/cbIXsTZUuEcUg9+Y6akq
0gTAlClAbeqVVem26WY1OejfNBWXnBcKHlbFcYv78V2HyPwZuM0Iva8Eri+t29tM
3WqPA0TQbtuEHtSn+f55RnQJ/Jb3EW5d7jRZUPjykJkp+kBSOUaqm1ML40ZXrE0h
NdDPLfDTGO5Znjuj3ij/A4yAEsMgoWvbJERq2rNg+P5RJrSj2p4Jz95JSrJbdaB5
UMxexKXLNww0h/aJENLWvO/3iwaQoAsD3NlGyPK7Ei06LeZ1Eroe2MGBbWvqP7dr
29GoLSFgrPDMLVK5t4YA8osr7tXbn0ZD+H2WBwZiocKgEkYKov/ZfBcKhdVne1Gg
BX5AKZ+dUYm7nlUq5hMyMiFOVIEgLzP13JrS427LaN4/NRA8aNjQbQB8Zve9lc5A
uFbUQAWXoHqMbszYd5+VVFgy8vEi5dU6y6scSBDKsS+Pb+kxlUDiYHOPvTPfe6AQ
zC8GUZR7gLGArFc3VU/n4mGoDR2ZLSXCkfgi6jRrkUdHy5h6oIUmawLCvkqGJXeS
8KJNfYUtPD7lkf52xYZxPZXWwyDvJyuG2KXJdHyvuk9QoszP5LjK5YA7/taP4dak
lCU92/lqygvaTArR85bJs+/sZgeF8uDjuDFPGv5uPJM6+meh+MI7+xjw2EwbcCrI
zdOW+DDKa1bEzBTUWqwuJmlD0vT9lRrK7trssQy0hhbisbS/UQwkub4r/ah91gda
QO9hgSjk4JcWnqGibZ5YrR5D92xOIL/RFmiaGIwF3FUl7IDRg3BvCX4UzTcHp8pp
/jqPhHZS9kmAAMF3SYt++KHxDc5p8lJXOF/dLsSfwSefasXoxXxayp9INph9QmfL
UCcXELACz4KXzQcwtGJp6BvDoUsBNR802MVOhSTN43uDd5sNyXFtojOo0mekbDLH
CAHHcqNYcA+T+GJpcjSJsa+un/7qTpxdtTW4psVI/6Y7L5bmDqNlWnr7J3bdzXnP
9oqQqI9CmfM/Ku4vMXWG4WhOnlMna/MoGZwFGZFJmBmWT9G0/xPV6cJJ1vRybBtW
Ttr+iMojcyDWBSufz7P+I2v9c4so9K2xZHiX2j0GG4G4lCMt/8ZMzgvJ+i0GyOeR
IwPQetM5jSmod/OrqmTxxwtgzQVFgkgcjLoS04oCfgHo2t5BT8cQWSMGs1Z/Kleg
BNo1YrjXM8hKVcFGWl1BCcqyIpyZCUfdqguoA3H9n+LifIXBjeBsD7mEjyHi5XGQ
jIY8CFruX7ZKNudEIElXVKpKExo+K+3ZCKScSVPfGP1Br5j09tYwnOA8HvGvyL4b
3Qkvrza7xbA6BZxi/6JLd4o54VV7xpTEM4UkdNtgvDZMRkivch5QmfHh/EMI967E
tS+4xFqetQd7kRXoxD9MGkBSBJSsRMRmWHJ+vkvPXE+stOBi/NHp3Nv+4rtv33vZ
q9fdtiiZXHyiu740paHPH1t58AyYPJfRLJuUV9Tx2EO30tmS+hVzVdcrLgQ9KIjS
GRNRURfM0gwbb6b42l/Spm+usQp3r2rn3xpVB+WtnBb+lUYJh3ccIP5wR9bGG2dJ
OUIJRzuLmzy1gr8cdVxxRZM5tZeNom5qbMTvIgE1fNQs6vvBfv7rIz+klJk7Lvuz
iWnngHMVJPPvCk8bj6rUoMTH3e95l1WuoUUhVw8hQnd3LpWYq+OhVa4vEwcHPhUi
dJMkpHzECSqp0HB5TWTp45cfcH7GqifOdElPMMDbPd6gLuDGEtBbXXU2WjVZd9kH
K0WRJ+JGyBv7uL2H+DofZiHlVSruVRW0DOhEjLCFyYM6rHRmju7B++/MwVzMbnP+
KRFifIuEDtX7gXJE1tXkQQhJKp/eFW+pJQ4rTZjpydftB0FnAZ4in6ZoMyX0qoCo
pb4F5eHotcki85+thW1gF4oEga/ap96qNmfOXypC5zgObzdQIfBVeaWH0RKCt8VU
VpCOLHl/UdDicQIJgZcid7C+BDVCdXxCt47VQnVNzeBInx7MuBi3jk0V2/VNnmYh
TJwGApKGLNubpNt7T3DPRINuJ02J7SIOhv2CEwe4HP+LwtZoF9b2UFUtmE5BtGlM
d7KLKil6re2dlscJ8oK7DKqZlG7ntKhe5iWKTln3jCKL/pIGMF764OkMnqGDGDrP
rkPiX6o/xBjO0qehrqkpRH6m4WWprhm9LOXoHUBIWpbIV0gJxeXQDvbmJ7yue/NP
eTTBsxwbFmCi8rc9WGzPaLTLs2yffMq+7xtpIA7QH62QnygOLnxsdpu+Ww+zdIQ3
SX1uX7wvVCCa4SuU9/ux67PHUJqZW40fEODEroIPRlQY6ETLsuGsDLS071aopxF6
gRULVP7WSfkTrbw7W3lp7Zxhvv7SzFSuF3YsV+s0n6FNQmjYlnRqJ6rylc9ic+Sb
LT9YbUarSizZhuO1wg53RUM5Jf4XJsrRCWQ42iJLVbUDObDMpf48BV2JeWuFR8C4
2L6HF6mV0T4pQuGlsvXbyRlrV4zZJ6pO1yTgZz8F1kHtYn8QaGfRyb8GDth+RoWk
8Gah6CCVm6bqUdmJ5Wl2Qx1PgNIuNnq4BGpJWQKWLls7/NOJpZWaAigm2KlCEwLr
zb19LMIPG/SNp5zm2Ezfj+jKTJ3qXyfdxqz2A/zBRVqf6S8O2RoszjDktcfUR+Zb
cfuH+PowPCUi5z97wcj2V+Ikd5WRskNriEwELMk6BV+aMDTENr46v0dd9ywVWekn
EKlVPqoEDTz7qyCa3s4Dc8kyzERO0fH3xKoLVxiUB7EBXV76Gv6/aRZo8A+CtMTN
903F+suDhvZ9xGIjrkTAcHSIy4XXJo72NUO9/rjyb2ZO52pyyqFv3AYCU0dBOKFJ
B9oR6iR0Es2lJ+mGoDrM/lNrk1vG+t14b2ozQGjKsk944kx/8TsAp5KW7WZ4Av0V
bD1XDMLe2TCUjNXw8gexE0sf51pvRLpqczkJHg3IKm9p1j9tO7Kaymv4wH486XpS
n4uZitJD+i6VqjRwcGqSFEjWbthf3PQwxZzpxsq+5t4cGIeNKdjUbQcPlmc7ZImZ
QRVQyOXNdTOz9gblPTtBAHWqON0cwlouA1aJ6odxpnHAqeh0Sy6Faa3+54tNYM40
ihEB+KsGYRH8fyRVcdZVFZMPxuO3lLzLzNvuHkCs8+ccT+SCNpEwWY0cUHA56Eji
ZWxZ+o0EL/1WGpnS6uidAxhq66lMz0HVzcgiQzK4ZbPC1pygEHuAIh4pIvaIquTK
7XoyLqH963h71ChBNyGvEFhzAxUPrxMYJAY/u0Xry1ag5PaudupLnPPw9qCA+aQG
SpR1vJWK2qDQ7dqpzCS0gQ/MJADQDWNHatXUrELeAggoa+mo8aAz0xPkMTi2qkRX
zq98eswYo5mRGm0tQFJYqNREa3P9MFu/CaOniKf3jmq1c7HpSJ8/97WD67CotfYh
+n0WNq5Rc293uiwN1ODfH4xIaw9E2AyRwOgcXxnxfAnzGsmPWkHpFr6etAYp/TK0
fka8lEZa9GQldLPyCD8vRgQmRZ2KRIOBEYK+7PsEeQc1PlgPJ2SYl2tquqsPFO+M
L5JweKKNx1sl5u1Jp9LYnHBK+Yz0VdATgQyQ6bREacWfxdOBNWXdflKIR8CY8yt7
l7jRQiEiuJJvo5uqW6Bn4xPWdpgLGBJUXkoPgdzeCWXTmQJZB11cn7GrGdbIWfJx
ezosGy0UvuJKll0VgZWNgqfA3qWsP8DFCSDJjkOLDGsdYfM3wcU6Km/Th5zg60wi
CKqIWi1L3A6ZOUShyUYzh8ulfNMLCq69LIyJSJyZwDhmUGwyarsdFLk6XmhF5UJU
aLsNKzRTkENDTTC0ON9i5yPoBZkqWi55+Fs2p3HGXbSuya42XsbOKCrNir1f0oXz
ncnu5n+h2bcLHFQ2RBFlxlNVeUx4WyXuUKZZvjUJgLNgNo7UPhxVyDCprNFz9LDF
w4SuCVA3Po56am2xMfMgrSjmL8aEYHWhd6mLmVz2Th+ZhXMeSkP6n2BNxwdvywFC
wBKvtoKBCb6yVtfxyDFftAnEHRAGb+kMewGBmXF0fcRTTdfgmt4UkVJUez4JkP5V
3t1qATdGkj/Dv+cnSq+mJudbouUlsUfFiZ3hIHrA49CmJB4gk+qb5raQKqjy7Isl
Ptz13bowlGGYkY69qKOSpHbxtQUDu6jfpgF9E1J1uwG+7ReFfVlFPAfI1gT9Kw+t
WIDaOLXDEQaXFZXSWEfRgovhevW0APzJP0vIiZi6xVB3FLIGopHOH7UQzsGiLLVl
vznHekG87nsp73RAIzNM1SGeOtQ4flhVc8UMc94U2Gtgtxwge2VOzvHNlVpS7SWZ
I/iywlVRos4N2jmvE8FqEYchANjCVqhikAR1qekWYhTwAPNenlHFT1HO6E4r/7cM
ma6hqNRFrLWm7DDbz1ZCl0hp1jJbZwhr+bwZRE6UB8Ri37veErWBfMya659J9ZpW
AqmowXG2PZ9oiNZnEJcRIeC+0aGiMmeiqNhomMIDDKCwE1ys4+HAEMoiDhJGQDLL
VkGN0qNOA19CnDf0sq3WiypuLCJEgxr7AeN8cm//ArG1x3fKzc+N0pz+XCtITDaN
WQgqBPQaBei02mk9PE9JTxtPGYX7k5CNCejhPcRU2iUiYsVfx1v9d7ldRj1B0bZW
y/RUkA/pFpUY3kNnwJYTES5X6m7Iuh+0ra+d0IIOvwbTWbVhPvhJ+W/0512Hccpy
yD9F50RLOcoMYSCUqc52B+vt3QMnQxgqArH2NtCHgvKphy+e6e90kP1Egaj4/Bj8
+X/fkwYbiyVJWHz4NGQfS9K2h+sExSJIubIfOVuADF3oXJZMJbgp5nP48YaNm04z
MnhcT/BZMyP64oieTvouYwHdjfHex9GtspzSQ1A6rEhiZD0awBhllGVRgnpCsAom
DroJrsPARvLgXNefZZKrVyiGdAjK1hkJ+MypZJvuMcraOK76U2OAxiiCcVy1vGZF
KxCdCqs4WVuBqH00GrjjtsxFzHkg+rUEbOZvMT7cvCRIA4udg3bAHJPdplkwyv7a
6CK0vuw5VE2YWJ3R+Iegk6bAhmEvsscJL03aHgTpzEDDo6wQ0YoUbER628/9VOX6
fLr56wwlZjEsRi9B7PmZHUVJlkW00SyhXAOOf/4BzrlE4hHsvRClQOsFe9tAF8fG
pmnHY2tqgpHFNUEgu8gboOLpUyvfgv8OkuUfIduXd9lwFvkV2Pj2cPWxSQxmbtJR
ov5I3QMpJVV2C79/f/6F4vFdT0FYT1XcNqHJPzrxXQEtQsygWoiIGLGHzinYgR4T
+0L2N0As3fmDCkeYn/Pq9skt5b8nlLuf0wNu9EfoRrPoClXnJdQ/Bub9XoTsWeZl
6D3r8MgbintVwSEwhEup6FE6QLyczGb93Z8dlrGKf1nKTaId+TS7gL7Vt9OGjAqR
zqB7Ll5cJoGNjsWscmkJcBvm3SeErXQb7wjc1LBtK7x6GArgFC4V5bzRSEQas4xu
m0c1umvNCWcWl8EP1jR6pl2uGvAcD5BpevdGE4yV6RzjG84f2IAgv9Y3gspK4JvH
dWCbPc0vuQIq4idSahHiBZSbgpafyicMHYHJpoivzy1RrxH0x7p7xTQP69xWaIPr
IfVFpTMiWqTPq5+Qr1RE06Qd+2OYYnZfOc/uEr54xb1DT3yfGhyieLQB4mVkJ9RW
b7E7nhFL/SpqnhIgqkNWFHLtBDwPNxG6Iyf+WsWIkrKGi14buUBWKdF/d/2pH8g2
vo0hPNQ8ZVyUJJOaNGY8jr/Rlzqxpd5Viq4feYnhhsd68ZANgVheIyijKAg0gDhg
q6FSII7fYezFxberwNtAJKEwqf6bbijAaQ/LhJf+YAii6bO9E/Ox0TNiu40l3sFJ
SONsTiLN3JHg/LxY7HIFFQzAvxIUSYwK/BLrlHZoX06Ey4s2zwbRZyVOLeTZbhue
BfqZTufdmF7dh/jcW3WBJxXXYGCQednxvI9rZnK0rA5G++BzCTDsAcVhdBSAWrdV
HJtxAZ6q2tkyOCWJDaDYADFfmtCtw7JQrfAl+E7/IO96WQEt2hUasTQ6MZOMAXj3
q9bhkMn3gu9A7qID30tFIrMn1E+pwKTJCk3NNYbAdFZZr98edd/imKRUmNV6V90e
ciMb28fyVX1z5Dye+wOMrRFgqz4eMgRfO4gMW692NTsNukEJlrWjsCITAW9ypl7a
+1IvUVMWReVh+aw4vWSM2D7MPRqecO8nuMs1wOl1WxRMmjPpDQuR29SOLFoIJqv4
yArsIyJ20AEga2YGUDd4K8nCpH5YIGKaPT9hdjqaI72T0Phli70RaXTBkLZUwxCi
9p0R+jibGFTdGsePkMBon33oP5G21vHprZWrnFNsgdssYDc5wxxRV8R54UTCSUB0
pUB+V+2PXEJ0zvtDzPT3sFmzS/DK6upqba90Wcntuom9/qcZpP3VepDVLadIC10z
8I9yRSYGZoWnV4kHXzgb3gd0G1uH10djqXqugb88lM4QpAuzGUZBJ1bdnp0MspwB
5eIieyMsXtRRJd04Y5vkvkZ/Va2sb1aQGEmQTu+UBPr1jMfrKbV49PdqcgyMR3oM
N+l4w7DHsDENOdtmmIKcBqaAbA5f1bGiMMtZUQdMT8StXSrnvAYH8K4Rha/f13nF
Ktrfk4lcN0bU52nIbAKtKQoNPA5CIJYq5MbbqRWyhStatuukW9BsG4H3e7TaZhZ1
vMUuLe0IJZMwBQT53+7aybklvU1mNt9udqX4VYm0NEHgJKEwZugy0X4NRto+MKkf
8aS9zQyJ6sMhXEN9yaTv72jFoht7uitPxALkoL3g3EuWnPB/q2PcHlvqAZgFHyW8
si7xATbbcoUhIBZL1XbDHiGdS9USJqQ8Bs4qntiVZFznlG50fYuOhZK+Z+Pvk4NE
ObswhpWID0+/7Bu2Q6jg4IFM8VgaFIQOieuKKrRNvA7p8VWGj+y4TOEu4yHw65nA
60WDX/aeM685In/Y27enph/N2KykpixE4l+8RgNjFRGzOw55BiY3SrH2gamNjRBr
AhorMzK/QYfyskgLJSqw4lSsWvlzzK9dQA8PDWlPEWgiTEmFDwbq/46csx/z4kmy
V/IKdK6z8rbyzUWBfyplfrpGs5lZlVcW0jkfpnRo5FKKPrl5RUAGlAZj/VgSKWcZ
19/5GfwNKB/FQXDrJ7QWnZiXW+iCIPttyc5uVCS4MA2v3znFMdPMTpFGbEQCySrw
4omyc0xGv5ttpdVxkxNiOhgyELjb0OE46VpSiCobbtIfkvjeLiVziEc6pchABb+I
6g86mQ1Yj3n/hFWhG9A6nPDUa987fZYNrqJxCvT8M6JNWUhjT11ogiYXKPy2WjHk
G7PgRbTs9phi4a9ibtJdhOpOwjJj0DXDztvRF86rcvMz5Mf354koTALKoM4ApAIU
KswnROFI4Ht19ub91UUA8wFTG+w99dfUoOMBIHde6hFpPmmo8teQUsO//1e/jaRE
Po8hIFdvjOUmK1PztzUj5R8LL7/zib8rWA7ug6eg0IjcAsBnDgL4fgZHDg5wjA4S
ic48uw2dTacpxk3an3ri/au9AT+Mk6H1yOv1jCZNvjgvCn3GJfsAsCPdeQfUYeE+
EjgsxRqIBJ+q2R9lqjVsZuNp0LXewmXo7fXZMSoaqAFNauCXMUvLIsC2di8ELRZG
jQlrA/4CAUnpq4O41N/vrIXtABU2Zp14iyZFCVlOK26ytMb0D83rC5oaoDdWUU89
+swyEf9MUEYfigg2Qt3nd+EKP5ki5Cu8HV7sykUvoLJA/qvHRWdbLEJaDfYIiSzc
Xfb1cMVF+mgfXe3K/+1xa5BE3sj9NXcNuO8ki6dKKRsHctQifoCvMqUBaW/vnKrU
ayvswMPROMSgTXAvedhGfZd2kD+R+5KUjYfyll0fJBdpdMTvHwgogZxaPqSTGL6O
dFbPbZLUDPXInIreOQquwiBu5qfxQAUlLcQkvNcMRWRu25Z3+vUFPPnGklHdwXs8
hr/RdG3/mW/FrE1dTI1RCfcHyJj0JfHkqzKghqZLR+xEJZggmGXTWGL9wW6cX2Nn
ttOB3MuDhC7l+6QMzcDmEq2TSuljFNMQOoelIhhV5pMJv+6CQSPYQNLXy6W/yx/V
nqZHgm+jFWgUU/gBLtE3MUAQkQP9K48IzFl+mfPNkiC+NpExBv1wIEp/4hwvwPmR
elKcMf9IT+DOej6pAoYODos5uVNV2Q9w1BYAvAynsmLtuNmBF/AKI6O4T7in0EbU
5qAiLxaezm+aO31zilOGfE7bC35IYARPn6iCYhAEu8q1pacP7nUwQfSvGsZvV0CG
9TGcJnItLDQHLBW27zxEal9CjYGkZ3jEUPiup9hN3XIaUmdm7UljO/ofD6MIrbG3
NjRDcYP4TrPV0yy2QLbD6Zh8N2Obpy5uc7/4P5To9uEvEzsvvIBTauSf4ZpfOF77
drOGB3DcmvEKZDhG6q7Rhc8/Cse1UUwmLx+5k8S9cNIFzeaJdJay6Vm3Ay4HdFkY
0JzHxdTb5pJq/mTmk7WI3UfHAx+fXryFHuQOo9LXPc4qQrRmEna0glw9WGzIdR3V
IpY1KG04fFQGDNIC9mMUgVtFhdOpH3HQPvOgSp2i/u7KSw1Qa9A7FXgo0EIYQR5m
HqIy+4lwCsD0YLZhkWXp2eAH8wXexi+itBE0DExG/NzVa7e3ec5+uss519Atjxj1
A1K96pnc64DIhlWtTl/wtHBeuq1DGCLmaWAf85HSAmiDLJ73Fu+1WB8fSmUgutpE
F32amDl0617orenuLouSGQJ1KWRU8km4Noidn4NsD11cFMfAm4HjO6dwM3dZAdO4
TKjlmeGYx7RJV0v2nNMraet+stRTPVqO8VRsIaxiuXZHakvu3f8HyXXibRkHvr9r
4DU51ptsIXk065hSkBgQOoLpQ+/ipWe0QbnDdZe8lYaD6yknoRnKE9pzjrvqkpSw
W4JSsiA0VADQ5/tlQLScDVgpUrahgi2PRWVRE1IK2LmtJr8sv1RaHVrDMqV9W/v9
TUWU8LK51mxRUL3czKKjYY3Dy6NsRbvjby2CfbLJyv377/Oedlej47y4MK+5VX3A
L3bTh8cVjjCZiJ1RDEDbnREuQMdwqyP1ITpicn4HqW6mKhP/DiTHLLq2wpZ59w4i
79zwABnvEeYZfJfCda97lmf4rzYL+rSHl4Z0KQD6XmTaEp6sf/uniYqqhTy8m90Z
TFusNf6dp717/R6QaPfP60Sf3zhgpyBhgKQbEjyxFxV6YEc43cFGkIE/oUybCcUW
nY5wgCe2JJ9iSpa63DKnMdePPajv8xH+J1oZA5Y1PyGDhp+jbDaHn46vUflNs2ma
C09AGWtG6+FXua+Ha6LSuq6gbILYbiTddsLTDS3ffAREVjHPG1SI/Bc54flhN4YG
uoDnEJQxHC0cM7ITN966nTWLyz+Fk/XPaNSR6gAns/J+BwtS1y0Z+Ijw/Uow/218
nMuSo+CK/GL/lsjXm2GOmtMtS+msF5fHqnpoiM3jlk67hR62A0V1TKp5OZ3WgKVc
VPGRjp2WmnRrlC2SPm8lnTQ88JnlnuqR7q6zl2Y1g6OeXyyHeYxHRyYJ4kUiA/og
XEURN+uxczaLCl6wchWFnpJ4E63PAkqIUT8U8rOLRANPs2Qx32xgYGxEXOrki/TR
HCLfQexq8KRV1O3ZXQ0w2Rgvel4FYwLSLGXE+cf4wEhxubl8DpsqbLL58JuxnZIL
C+ZvmnTSvOHWZW7tKtCrVVM9tmRK5OpmvhW43XXeYHIyHdlpDCXDa+NxMhBj9TPp
I3WzKJVVMqCc9zEvX4npzd070RmozO5YwlZoloP78l/V0/8HrUt0hlrifXWnha1b
do23ZhBVTGQ+3l5VrUx4rSGV1ldY/NPbP13SAQL42xLqpGaO/RZz1gsPkVkZVKsn
GiSWOiyKtn8SBL7FoX+mNG404M1A8bsE6nHzIKpS0ZFh/PFWnncK+3ocrjtQGg4x
AEoJ9AtmcTvuc5hgKQrkpJU/2GeQ5dq94TtiDhBepKTerr3zG0F3ihRwZhy6EhKi
no7TWKPAixxZ2r9W3j6OxkHYZqaBiKjWUbTRGAgdH16ApUcXjAEFbGiFJ2FVZhP7
i/L9v5stdoOS3+s8DE0AcUOhgHFHG2/yBQCnEH3qxlG5X4uoEOXZxlnZisgujj4P
HMzNL1bdXAIUqK3GEP/J+QG1LYdGGtyaXzbP2Eozm8oeHhTzmH4pTzNBnOPHETRf
8iFlwjJLLy+oYmxg5pV/nNIzCoIdoqkKsvM45wgMtJn658/n+tEiuQL8hR3+3NVk
xkfhJXtjXrtCbIqCL33CoRz/KL7UFjmds/Hdh1lp3BEqI4GJRsvfL7uLVx4AJ37q
hJWk+OyVEg5FPwMv5trtWTx2jmyev2GYeE+kIVkpvtefJ6T5bios4j7i+r+gX1+Y
iM3P6gN/gJE7a1zSmVTCFDKIcb+MChOgV08NfSWDi7CuVUVmFaTjm5t4vv3OOgkJ
pWuDWSwIX4btpD4z8WWCecuNjgOeqES6RXJ7M/uFfI8/pHuLVp0BzX6VJFpi1iRY
GjVgxtNS2TD0ptSY/GKVdIPY9quStvOzWXQsVazGpPsJtovNLLSe/GAo4LrC5HCA
v5MeVVmo8zP7T1TajLIobUMMX8MzWgocug7FZ+DpZnqIfygxUtOIF9KMg8CbGm9C
kdklGXGjFcJst90p+scmEtzRV66kyRCKzzqwC5tuJmTmXCliA8Yh653V049n+ONs
JKu0UDYQaIjGs7qx8YM6BAy/P2PTBA1eRABvvunm9aAcvJD68khYp5u4zHb0Ukxc
PxUCAMjOhPUx7gHrLzd+XRAJ2OA/0Fm77g5Uv5aJvUqeNumzFQ+mj/TL0q3RBV3j
ri3ScbEFOp2PBl3gaEmZgUF4hHjpWSg/nsIgxePc0bi/IkXRPwTOpxsJCt/RR2Pc
0VoQiu6ywK/RmCU1mfSSivcnqGPYgZ76XV9Pr7/m0O7uEN5R0kLJske7Tiyr9MK1
lDXgSMqM/Hsm4+qRehB3p/PRiWRT6SfCQ84nA+nt7NKTUUBQo4n/zYTiHTKpRkS3
xJw9cU/W8VW1iOPm0Y55JQL9XmT0Jomk/ga1dg+wIZ0NZMGYxcuUpjwyUofT2wh9
Xut9SkhuyrrIjfIoNL6XGH+IUyV+DXsLYCaTRDQXEJtsFsaRvmiZQnQcMrSKw9iz
GWlVK8uNedtMy015T4ycedfGwBukv5a5pWLElmovqEoeWCBjdsrI+daOhJcjsHWj
TYlTABrJbSCBiH2clBCalGF8WUpHm88jGTa+k1xT/4PXzdn94LNnUHWnWOG41Pjb
yEHmYMaqvwSNDkbmaI8KwHApgX1HEn8HNntEKtG0gVnSMm/ua0BYuL5kfVw0Svyr
k2tEB1n6BcMbLHAc7b6BcrUZZz8P8RJl0WviXFwCxgGFllG4PbhqMctlSgH9sr7I
eKuokVE9mC25PfK2Z1QY9aNTKHpAb9ZhXw31kmkjz6phOOIb4WbDiUYGqBfxQz/f
OSGS6gJWDE56QJpNNNrm85cX0A0UxZ5yzUHtO5S/ST3MZXJzYavVGmVK9YjiVW41
/9NwqpEdJ+aoeZSwMWf9/lUfWRCXZ0bwnGHvH+iYEk1V+d1iEqW0T+VJ3BlpBQTa
I9fuwFzlEfxTOT7MQyT0yojYe9LDKbL9UlNhNPNrV0z/aNHrv7tCOeE3n8v/c1lk
OQGGkmKVv5TG+gj8org+Ox0V2GgDbreUJSdf/OCzeKqC7yhwrkTzGGL1l48IavYd
7W5EECFyFCgc5+/kdaOjPEfTtALYJm4SIpQNME1MflawEotOz0yJHfoEwi8yakCD
Fma89mjijLJ1esLlW3CXxaHIszgvoj68Z+BU4jDJTMlFHl4nr3tadbNbP++KczLP
9ydAuPO1dpdBc5S9ZapKWJbpl0+Me1OREmtpSuk0K//3LVk3sg6K4V5AtPcfm1AL
/zE8wTod7OHAwLnFLcI+QrVDIgCQoUIYo326KluFsiEN+7TmqCB3lsK+MRLbRVVL
gBEnQKL1eu0k1j98Ui/zUEy0bXiWSlRkvMUYFoNwdF4TGJQX1W6fZhUqh38JRf3r
0dnoZsNnrJFrT9EVZstZS8W78ps4gN/y0gOOyxMQDzFvlesIypk+iaRx+E7UBYJE
vnpIjFwkqir2NpuYp2lELQwpgEGCuNZXcl9ZLf10wsGWQ8i+WHw5gv5/Rj4BGldv
KhbGFG01A80TkLZL6YF407oyZPS5GKINK68JTkpE8gAod/yVMSlDHZnNbYSqpGdX
i+2UUVOO7vmzGVsb4EG5hRyLU5gPvtXwqFsx8/ddAY9lrUQz2wJtYDdJG24z0PXd
fLFhcF7335NSrvWFxJVqoLra4KYm5TFoOUsTwKTk9TUlq1qi7QtkB5M1eT7hfdGS
MWtm185vuPxnTT2B8ABtLgYaHlG6YtkJUjWPbquRCT10MYBeuqUXpB0/MqkCF8iI
TMAuI6hcYdA3xe7OxhU6/HyvkoOwvRw2FNmxoPugsHwL4Ge9oty9lnSvcdVQHLKT
oiNVGjAQIvT0GTgQ2xMXwsUZ+cVMHASbdwCiig9G/xz+nyHOHrQDNGaH1CohH1Us
PJsxBNnvS0p12E0m3J6W4iywR1dYphbePzODukuZ8EOgsZRd/IY7oo1JdB3sBYuG
TsxuHQPin7R9C60nGG20pxR/O95FjkVsLn4ztMKQRyqLocauo1eyeHfWlzklABTg
tKsPsBUlhfzVws+oVRUUZ+DlDCAQIweDRDDFSTqR1+2SXwM1hfX2lATvus1dXybA
rfY78VF6J/+Il7CMSCykn9loj5Bf6B6fSuTebA4XnPre9kFphHeTJ7yrFQeIAowq
fDnl43IiudqlMXLkKQA1JDIxn2pgq8QAc/VY+3uRS931mDYxwlwzpZza09vXwQNa
2er+qXaCxlkF5HXRTPnb83HW8anIB0VoM72uAxL+sOIS1xqAwWXxIt/zQ7TkUL5N
4PN/oXjrxWjPNGZZI1b6IagXbpD7VK07Qq6K53ttTjk37v3FcgqIxzwqpqNibCbq
DVrnHg4rIuVAZlF6YDqeaHf/TzVTfQdjbjQQNJjUDYz4LT/F8IyMec1OZNGWfXWQ
bFZRCV24qj1Ht/kfCG3SFkIsh+/z0zFRiclzR0VLVqjaaElp4qMv2lM/x7/avHbY
SN9qq2KJP7H4Gmb4+b6Y3Ezta5sZWIZtbLLaFEzLzY2iShF4BtH0hUrrIksKcwL1
5yB6QWbCQaDEN/yPEkkQJmQXD48p8Fi75Bc0LM90JNJDYTiTJD3DH66JlHRGFoeY
u8TVj+o0I3aWY3hrWwZOnSP+PP4UPcvpJMznyt1fNHBXpHgayo9xtwu/WrdHAqOu
4JAv0N7Cq/TvpH2cp2Om4CUD+uHSKnAhsGp1BNPqgJ0lr35zqfHkNnB95Zl91AQ6
vL7g+GJlQtARWiQFH9Ug1Sm6r7dvvXpGLaL3mdyeh2ywVsZBWbA/N/t5TH5DS8RC
qBTbwc0WVOKGR0yolEsa7c8vt8jTXBeFiQMq2zQVxiYYPcIgX54hz0sxrMr5KZOi
4+auqQKJZ4nB5hwrmEHpTOpoyF1+wRENvtZVIzMA8svLHi8hYtjNGwGRWj/kgUQe
egSKHbNgSi8u5l4QROLl+5HHNVXFe7HrqBTkXXi0S3g6MFPD4ZltL72RvobZAdxq
aL10W2bxjz6HTGghWCvP6ELspc/dzCc1sSwbnra00q+tQPiCo4Kx03aY/0n8+Mfr
f3ZY/8ABnTcpQ54l8+H5fF/7I6mXysqr8P6kLL7GFqs2HLdT7VioxruEpkysksMQ
jJcvt23apVS+wsD2/TsTEH7nOsMJ/HM/xFkzEU6IxpxITKzd0SQosrRTwU0n79IW
mHIcw+hfqgLcazV3jptH5gmRNSvGAU2Hl89JwY4o5mIgfW2z8y4+SiUmSFCDHukh
B+YLuYSH+xcxD5zTVk6syym3gXGLD4UH67twf6U89Kq98Dx/8GwDVhT0nrTDjuxO
4yWSkiZs0zCShJPDw/JgzlbvFVkiWiEMFTyzJy9b1ozv3egxPSdWQR0CaPJCspXT
DSRcNIrYQ8dn9dVvNXSHPYc5oLcI8XujMeQjofbhALUZgHpbxeesntuoOmdTjcKJ
jCPaccpVoYVMiKyqVVbptcVl4RnR94wFOsGI8znigTNTdXsT/S+XlcEPMJFgmlPZ
XMuNbLP+1FIODVQvrP04/oP/DSwfIhcSKwZaLCMMJb+ifztsfeouhbSgOyZ/LOCN
Gmh4aMuUR3PDE3ImZrLNXKXqqS28nAGiIcGuqX2aXwyeamYbfrN1/8Bcw9XynBaQ
4kTO+uGw5PCflfptUuA+pjSo//43zhKtEEUBmwZIAA3JGvpeioONllln+iFh5Mcm
hujjts+A93kOignAkEZ5PyzOIcs8SqMbu8taxKf3Fty0iXTLlYltv4eTF3KnL4/P
glaeYJhxDUWIA2+BUCAeJAhbs3c/gN6D8r4OYEXnnCMY5D+bXQfdIbdfuemNt0Ko
FJVSVhU0KHzycV4GeSIwwYFnRTwRStv49wNzTVCPd3Yq1PDMDzjez3RX0YNlXvMf
VnqQP+Q3M+XA2ChdH3UXSnXQO7Vzb759QwziDl4Si20+YBQQoXBK3kofXMEQITND
vBPu0LkbdBfQGC2BWQz5hY4yVf5znzhkMw4aIEVZT5Iw055VnsdvISO3u0/XAMDh
btzpYL8h17EU9fLePzgiwJc8XVVvzLOF1Y8mUOKdaTnt+Hy7I2rg5kcnkR1NMOPA
2XvrWRjqyP1sh3zZ+aFH1yZnvHt4dkVvGKYwmkzB4jJDOOs3SCX00srvBGcF1oWD
cnI41EOG5bmkgRnhLGlCSo7OdO204RjRBUOkY7slMkkA5kuoRKTjLqHYnAFejCiG
klaC6ui2sq97W7Y7+v++lgJxnISQdjojASgUI08LQANwV9zgl2Ik3wIiDG3MOnzc
0pLYKceH5GJOisBzCWPztbEw02sVo7GFXqQ/AD3gaTlvdSww7Rv4lOMjQV6xD2Vp
K9PDNsOXpZSkhhRE1IWt15AIWNm8dm84RisMuRQ1Zu0YvIGgAjOb+Cztot1LMU6k
s4fPDdwECrgZXozimEwNO1jp7Y/wD+Bt9mkuMG1x6I/UHAxOg5INTnyj9n1W3JXG
6KYeMxMLYElREf/X1WFqHBxPs28EBSxElbX1xTAyM1b/qR4yNloHUDiIJFo+RvVO
cZI/THTwQbzcBlUpJTTsnUmI4Sxkce5QMqGwDyf2TzpNMovDRiD8qGFWqEOItE7M
ZsLNxAQ8+cZnT5uBHJ9IKC7OLkvflTEZfnx8oKfv7GWIqVgyNaVfnEibEV2d107X
l6hNjrro5tfYJhI8KiaqEKK232+EXkIp1okSpAVK1fQmwgUxT4kw+GWdPObTYTf0
q4c0zUNEDYUmEmG19RcMxQzSBDN0JkC61WM9WAWZnnisQWSwqrlbZ6lm5aoUUNL7
ev51yVnS0G1LUswfv6bsUyHnm7ggdutQrw6dkognqWMddXCkaYxB9z25lvCcWswq
rRdHZ3N4hyj+5Gdk/hcEUAleUUF9raf/cIqZQuNOVD/y5SnbadfEhFh65IvdTFs9
FVmxM6hyb1vvHh2miya6uKPXjHcdIKGzV1amrmziyVzwDBLyrBAUz2BBdqrvc2Ju
yYV06YLDIXZIViXuUS5bSF8CciQ7VIr7hA/vQoOXB7QQfe2MvyZOqKlzIApoysvl
6PC0QHpBDUPfZKMU2YW1fjUGtkajxADQDQEdDySz27nbP2FMKMppxpti/F2L2jzW
U/qSSc38WZlSpm0zhSUg5DJ8V547I8xKyWCumI76IdJyLVnUAyGDMA+XSay1RscJ
IYcNVTC+2LxRSqJy79eAO3Ii/kZgTnnfwP3lRpPrDVd/zoLXMKWWkr6gOTFrqxl+
HTrnryEv+yNyhn3tXVxo8eAvCp7HFGdmEtJKlUoOkAPNtHURR4wASthdUKCZfrHt
BBHaYwfH/jQaIifEdXHra2Z6l1moP2nxM+rRnisSiAqDibzHHydjZtJqJtbToM8O
9HZ1uwSA8uxFdruR5tuzbgjjpOr3Hq/a0//BlnwwAly8ZMpFIAifa1y6bB5KorVN
28jUAVJrXK5HbURhZ0PtQ02nCbsSX19FSeOuIso0HU0sEB1R7v9wb9Cka6TSlrbq
tAYpRYR80g3bN7CgNkNtQ9EgLzYnCdGFWp+01WPZl8Gv6Y/ycXIWU9Ry1lL0L9Wu
b4Xm039uySkRPExz+pQYbLEGMYM9LW81bzqqMKugFjk9FjUwicAQsDXDfHvwGDKR
4A9yQZKI1QOv4dRrVHgAjFvIVqmaiGBS87yl7nIQapbJ6eBilOHwiL0GY7txVc6c
EBi/s2+IOhPRXingOe2iqNhFLODIZK6HxdfFS4E2MBiXCKtH6/0uBvCoDuvatvt5
fZdrvVKXbQO1qk12wGf1t1FDPSQEYytGnZmHf8wSL6mS0qWvHJGS+k8o4UbpV9X1
BVV1dBwrWYCXONKmtTShtbhb6gzB6mxJayTTzxJyoEWDpaJRPnZ2us5V4lNr7OnN
rx75rWw3ljFr9MqaYEl0xawlT7ZvCdeFwiNcldqtgnl4h/9vlwryfKlTNEdGlIWv
RgAN0s02lehvUKZUkw2B3r2jtDOudbHF5ha1kFD+ELRL6BmzzzBHK2xpNzAvvh3M
AiT3KY1H28SHfYE6dRowIHNRlB7NMbWWOUKNukjXSV8WmaY60UOOzftUOmeC/wOb
9nw7ZKztSGDUJ2LoOcv8IzWU7pPls2pUOzGc96/NcKIPBF3vIwCqFFDF3oect7da
OznH54Ulop1zvZAKVJauktStAALfH2ObsD0rUDIIzgVgmG1mdmXI/xOoph/TPAw/
HnA40Veg9cMXXKOheZwVyk/Q4TL3kTkI8do+NSO4DWCdQD0POezYZB7wAJCD4Bwn
hRO5z7FOFCjpbQSCndkWH13fxEiL2sImWPF1gvexff4ZsgDjV5uH/XHlVtP4m15g
BplVkUu0mhvHLguj7WOuzi/xb7rcsOTJNVQWlzPZTCMQZtFVNdQUnm6v37db9tmE
vTsTG45KFZrr8yuNyn22uyy300dl0QRIPA/auu/+ZnuQMbEqROpQgYEb+g/GQKNh
VGyduiJmdLfpFhhCEkz0DPYXAjBYdMQKuJYvNaJD5Jsr+x4eHvXoVLCeqaBvNEjf
C84aC/+hVC7XAazgbKaZPfg2WSsO12kBTLQ2KxxUyvn65D41NZRwYG6dpTSyVh6H
Uhb9dSxtJfSWQIhHUoEBFjjEoJU8XmzAcm0xPS7SHCt0XVWHiqIA2mfq9g2WALP1
7iOLuLgvwP2xErmDxIqUqbYnNG/h7hZwdS8s6o1h1QZ6KUGHyG/kI3nCqKIj4Q4+
R+IYMKiwL3cvgTZ0WUIVIyPXAiHI67cWxqzZkvF/r249vg7f++X1N8JP+GqiXHUq
1Ku5ZiKEMdN47oMJYhXWQo/cinzkMw6/jOjTpkKhO8jqHooRl08Q7IRtfGErICm9
5ag2dafIyNHaeeC97g5JcxvK9Wz/lcTnfe7cPNzxTt/86snMPiBZnbn5L3o2y7Bc
V6gTvz3ox6SrACZ0Ta7qP96xFeVRujPRnlFxgXTQhAZsvEybTYKYFtJzN82Sd+3e
z5+gUbpPXh96BE3ajo4Xcit3WMPe25oDBGh7TPtGWYo2XHY73nNMmcB8cROdkDli
bGJJG2NCE7yoA2y5QXUnbsRPddht+2iBI43kTW19ieTBC11b6jVg1g3/rlbo9jlj
KB9fPW+OE7tZDjyQRqGrULCBCj6EoTgyDHXZqT/ImQGPTD1kbQ7RSAA3jK1gax0v
PR1XKEZfCDLtUeNQxo5LQomuxr87ygM6oRpr+Yv2aIVOxdmgu8h+SNswSLioEakB
k6iAkisd5kfAJ7VcPg8l7XxcEGu56flgsg9grXp/vwYb59KD/N3ZYLi5rMO8i8/N
nQ5tfFuGClyb6JiwpBbDMal8LAE2C3YEAN1v6jTHJNCAYB2wKVqUSAtDY0wMeZI0
4V2Y2rjs+/ogMihkk9EFaTBGcz9DBBGK7rXXfIFCsvBEvUT0M6Wb34jxAFe61A0x
j8CLyahZkm4cYzEgYKhUmXwylpSkBxHHQUGrXBM+JOBXkLTMETjUD8yqQE4jb8bX
WSl8IdgHM3dQKhuRiYPwJU9vk+QDMEX4CasfsR0UHzBhvUNW5IldU2KKTenAigio
rTGHBjndnzsx6D4NjXGhtMKwnTY+EQKIMmlyrZ81Lh7B9qjztlf5V7xSjWIMf7Wy
Rc5eMl8nZQ5yPIrqG50ASlAQGvHZMQGT59pzJ9kKqdhV1Z2+5MhmKt1/6NoXwGgG
wUwinJtLqWq/lchVLwcuKAaKvoNXjxrc6A66xcOMBP9voS6y0lcA/5HCUqk8X/fk
6lM5JFUbK8HuqSy85gJT/MC9YQOFM9TPoQP7XOeKiUUkgpddDxijv7rQC1gXKbIK
sPulFkBd1McR8Yt2p5UAA3CKi/y0T8gS3Z9ZWSQkuNc8UsCnRmfVvLLyObRj9/LU
j7cmIbnKzFOnBgN1IytdVBarEvvUF2g+sst44/b2Gfe48JO64ep9czDZDt1sdlYp
dOR47FtR7Uxyi3P2EIThtqNIJl9K6pgzRNOPSkFi0Hc7WmlZeiaNhaRsJQD0gSLQ
AVEDbsv22f04XU74yy5VkCY7K9VxVaIpBA7etic6eAy8b3+g96iAIy1Hs7TzE3uy
OfAvumvlRk8tmToQdaP5bSenVybcab4M2b/JsXI91rn3mexRsU6rb0xz7ErA6YRh
LD4iHTKTf+M2ZxE1xpDj5+ICfCKB4wIvfjSwUDP8YzCaJ2nc0MzgIr569OWEVV4q
N9G7TFnFKtCoTiowHZhVnm3N3t8D0In6GQSorwdtT/Tkl3ZYMMP2lajYJLjKsaTf
nSDWMSlFgHxtuyJ//KLC6rkpc/kS41enUpCeha1S2hgFTWoOZHX5FWUIC7/SGWkH
aYbzEossaYcZ952fgwXNI90lsiJOcAIcRDsmet0M0mCK6svWmR/ekPaM5rhMMsZD
giZXdfmyoXfx0RobRVR3HRLXW/xGqXbW5YWo46tbCtX5Ie3V9n5jV1AXH0Gp3Czj
JRPmK301qzYJ3f7zGTpvgP2PQx2YN6Rn9xsO8vSTGDHuSM7y2K7XjnaAQDjka8SA
RCGwt/bvXsOgilXSkn7PNe7f+M3VmiLyDz9FZaJnOd/ppD108cgwd4cPzVIu4r6w
FgwNrucYzZqmCqaTmf2lN6iqY08mZ92l7cCMeB/dUsprHzT9lwNgPiN/ktSHWXlP
FIEbsntx1Fs3uElf112YXxs5iOiOzfFJXl7jPxunVgLJ9IkN0rxTPR/TW84FxEaR
GCJoE3NVsTHAaboPpMFrh5cXJtWpCMdBcNlC0ylkMR5rKCGIlWutCjo8hTPqo2d3
SIWATOL1E1s6QJP6Psz/yRfPZvo5jzxn/BlVNrC82Fsxcktktoai3XZi0gnHm2WJ
1TfTBAK6n7ByAE6uXxdhMthEtq+BiY5ef9PW9KbtIGMvda3OgwGLVNodWEdNyYqA
VXgYRFE9bBuSlCpbK7JtsalAmeK6fxh/A1bGAP2kKS1bc5DtMj4DfjnfeLF5oeOq
whx6v41VUJGEjCzsL3G6k3GR6F61FOZkRo1Ard3rgUInM7UwDbc3qwXXl67WY2K9
qT0xgUdcinHTXsHPtJyQ1+BiuDZyMP1kYTsQW+n3g7Du262Wc+9utDseKhNLfG5Z
XD5vWaoxcCx3JI/laPSkZNh1MZWG+jRmWiCBkA175OemdnosIo+CF6eyzltRM9Ar
AqlJDyrI0MwZgkM4501TBXaKZUdioITBep8s41MH34MlO3H3Ui0HAQMHCmhalJkr
0yJSM3hyN52Plxc7s0jl00w/q6u7X/gxO78zp04nihbG7IJYJpiRyhdQKVjOImMc
FTxa7xjzQsj1UA7WWCADMqk7Qi1Y3memTYJHnFLG5eVan3xV9rl5kk2LgLAPnwvQ
KrmmNDKYuD9Ip/Jv/3WxGzjwlNWFu2brDmmvhOVvU7YbpvOyEKK5ItpNqbqGS4hN
+9FZcLHyp82VLW04QftYsVaUzkS9S4lQRE1pINswb1AhYLNqGhXZ5Ciaxd0KTxUu
ZUhR2G9XidA1+GmzCKuKHRP+sb1yxKchY7g5ew6UnDvd9bo0ZicDQpfrCoUCSFv8
0jbP94PKO1Bw/JHPaYDax9trsP8m85o6ZY4bKAGhfaHmBrBy18FCUCJ1nlxV+Dy2
s6uu38g7l5qjLL/1h3naK8tUu/oKu9bBQsNAG7lxOZU4ZtiA4V42iN2MlX9kP4Km
gC/3vpCL9izzm8RupoV3Gs9w5q81RGFQtcEve8ZpiFwF+hH3DT7tQWuvRmRYJVXO
c92w9xr8sg+JihSh2OV9OSD2OHEOLLslbk4G6GPGJwFeeCQA3wFyypMUt7scnA2l
hFFP/6+UmNH/Z9cpZWBafCSDwtTPVwNofXF0NLtZRqh2ClOf2vGie8gduMy8r4eu
bIlQjG3joVXiVPYfRKrsyHBiUAnp9Pva05SnsPHC0l21flYN5UeSELHkiYqfXEzE
NalRdJLt1ZyBgOPZZLbF99DtS8vpYtxlEOFSQxBJZY1narjBrmhRJscYd38BouZA
LV9x2dqjdf7kyvk7BGbCWWgPRuSGcsM4vHCsR5XHWztgCsyAgRDH4Zi3o/Hz3A0f
ehvMbOSTwikry+yBdwmX8VrG4QfdxC/L5JdKVB6GPrq2QTZNx4E4jyrnPX5MBXla
gUSNMssajLS09nw4v+8vCrr6wuZE5r/X4d2VCuhr4lcqXGJbb7kvho2d/lh9GUdT
wb4y1oWC/nia9DdRBROHpZIwhJldeH+SeMxoF/a8ARfYkpUnrkTYLvJeDutGkLDm
Skhse7r5Tb/MAC3/tdN1gt0qWIOXeRtJXy6ee+2TQ4qOTg9og3hVYcvT6JMu0AM+
fAI5hQehhXbZ6fFwe6U1qKRkdqAV0i67pDZKMYFiJ0vEyjME+pw5+Y0h3ClA2tLv
uYwCuxVKfj2riyib8HL4beh3jfxFVB8URq0OyA6h+4QN1erg9hWsMaDmvkTtl4KF
bXwXZa8bN8vbh1OiaRbb92pE2WGpVQp5KojE+CLFEpzJX2fS+lZVaRAy1hJKDYxr
hqvJSkqSSsbeQglV7J3++IjdVeyyiBPRbH2zhQXGKDnHFiXTyPXkKhQrSHH+fu3C
iFcGDi+iiuJSX9Nd7vJPkyHHnGP0lfel9fmw3439TL3NWuTmWZz1x7Dd1yn9AYoD
YvNk3nY1VBvVILb7/hPXa2BjZp4mopCR64gDgDDingq9RRh/6yX3e4LqHOTD7JNP
l/01UBdJvKTki28xNjmjTzRLOsHT1yXKO0xx+vhK0jmHc9+4P5Q00oYybHKn9hN7
9dVA12MRsTJ8APmOV1PjrbC7xiG9envSHlbSRX3Hm4q/aCz85HOjZhDtKwtHAmK1
KQOZcX+TuDFJb7ogvQOYcerWfou35tud9V5+qi3pVKBZbdVvWvC+gVMA8OVNf5Sd
mHeWzS6RWaM1kkx6/LKn0T1uCDiwcp6psDLl1QvusyDnyznJYoZPWsJ5Tdbyg24p
RiUSCgUdGw1CWClMDsOiEqCyQCun+voN/qy8c9zDJgbYY9Awm7HsqRVWiZG7D0yQ
934VXupUztGbdRmdogmntPT/xnHz3lF7rT+O/37tVY/J0pv0AtrPXi3yVz34E+uD
mTpGrQm00alRHU1ZaiQ7FFKr6XH7ZqjRy/LCJfizDXtxxNKLeCwA14+vprY1tARV
gc80gOx6MvHYv6sfZ2amPTDZhqOPnDRMn4IrYVZ2hnxDwtdx0lRAaEq+dyXdHzXS
vMRGCggPpcPGJDtmTKWHOD35GGqPBXKkyZbOE/ODHYskGNqe+XKgP5tBoALHSrwU
+ySD73N/Q3v5VbS9rvmDh0OZZaPdJ84vKigkYQpD6ldJZNlq2sVBX08q4qkFbiWp
OnW3luMW7PQHXqxGP6FBsA+GcmaAwRGf/+cTR7fAESq1s0gB+L1jr6TCLpaCqita
EmQhqsmnzYe2NlhJT4h9Mj2/GKx7p4K7jz8Slwtd3EybpEyQ0V5W+A1rIR5nWqdM
y5aHITLegsNAAS7+6zSugM5k6t9ATsoICDb/zO25qNiQj43Fbyavq6GpYBtSdQAz
WGNhmurFFCCkItZ2gQd3AIK5mv0cyoE67llH0/R1ocWJcTNsOXF8yTahLMw31x4k
mdH/k8zYC7TPQGoNsCJBY/ywoi+XVYoP2YKHq7M0Qb5Y3n9NS74DVGXWkAc8TFZ8
TXJ86NQgbvFoXobCc7wQLQC3dWNOf9j3P4PYml5A9REOhHNBv0LrBq9ddUv9Fe+f
uCUBopBMAx0RhNlA/QApUKAjTZRAUlaXGJjHJP47ddmWNUTESohuFV/0Yafwt6AI
dvQsuaKr9OdjLapHzXPzMab7zsprRA7fG0lJQTVwI6vyJLYgUvbGiE6QzGEsb3rm
iCunfnRzrxtaZDDQEMm04OL5ZyyQUUGPkuU394Kg9aJ7Fd6B4pYTD5s2urzzSnJy
2uHaDywr7GlLfnWMjDLWrLQiWKLgC4ip0boPu+l5E94M88wtS7jutkOcVIkvPkvc
SUtuN9Ps4NG6VRhA/tevU6SZDTj6k5XEt+rJ9Xj3RJbWMU1i12D6I5hX2jCznvUt
IXHvsvn4LZs/fX0FnhuGuQeA27NQhQxxGQqbNJC5rEllzg/+v7XfHyyYnWVaI6r3
HMqb9Qlk+yvS6Kh4W9p4lDyCNAKb5dwoEnWwhwtLGd+DT5xJUwAtCqQZd7JVmsxV
jAjbCEJSe0KzZwIwtrMsUyZXtrBLmTDdaIgJB7RPBL3hOFYRj0wv060+wR8cCGYI
vMAgY8bzmxYlvt4m9nd7/YBvHlQ/IP9jGrH4Bokn3q7l1Wg8XPzypQRzuBKvBHv3
Oy+oSD+nPYH3MzMr2BV8V8H/fOpt0PlOlhrsCcgSOWK+GdPBhIysljAuVVTqIcDt
wSID/byBpHJ06jZa018j3YGGDiK1G6XroIZ2UfHWOJoLh71YhWKr3kTzizJO30wh
EZFV4lMy50ZpS3OnOq6MTK5lOrNGkb2Phn93YNHbEhTnXcSNWmjq/D4TEl6a7rx1
rGaruRbvgL/NIWpp53le0cndhQ3XLc+N40c+snldrVn8b69P+OAsEOg786xgG4zx
HAJk7DxLMsjV0BP6wTJe6RvcVEz5Clzd3Q+mjh/YfYyG6WExq20UBxVZjYDvbJl9
bPbBbcvcKiLWXirBUmfMjibb3T4rW1+PyFoXuVSvIOAYS8X0y4JhA8Vg66u/7Zd3
nNlnmkc+VEax2t08nDzMrfPfjEVSN87XH8p18RSA3oOVn53jdSFVvBmrGZ2D1Wot
Jv1ZEHvNjaQKtnYpr5wRUb0siELx8SVz199L5JElJtCgcpp92BWLM2LYhRZFLXfm
79/ilmp1++K/qMQJP1gd+Fx9DkSfxJDd4r8yJ1bmXA1qpsxkmNXo3wcbv/2TSuQu
GHsBXvz0zRZX5DYrlTKp9qwS1D2g1Xnr9JXZ7kL+yGrPTfx9Dv7iT+WTSRIKdPUN
vyFZ+wspewyx6180uPAKdeovqnxL+3qZYNH0XRoiGrkOhwA52GTfG7Qr6TkxN7vJ
xtlGcC4KHbuDqEHfoDxdN+oOrvJQIBU1WHSsB0DxmDH7wHx81eeUwhfAmOEo/OQw
W9a9D0Rtnb22Ud7HxpH04Ehx/PkGb/O+Md+rmyKy6iWVz3pd7Q+a86r+e1d463x+
dcdKOM4XsftLh+aWhKV3dCMjd9AmxZuvGsqNrKQOwKgiXRmeoF3GJiySOwSuL1Uw
5l3Z6uY8dqFe5UYKQldM3yKovu3XRmaiJ/esWs31erPB6jRsTeYzYptFnQXoftcS
T3qLDc716FR6e+khM3HFyZXmbOCQBG7WAu93Ck/XytMbjOxnZkWP2jCjv7sjRAp9
tzxEtJHneQvPxd7nHJtprb6CWWs4BTPb0hrVoEGISz1KVXYhP/errFZz+fAtqXcY
cqnPzYsI24tVkd4ZdaB23E5656pcE555MgW8u13PGn1/p/G15G8ZUA4nzo26cYEO
uxazWDtII40NzK5itsjuVuuv7cnshV7nwn8hSgE5U7SwauwwiLnk5SGdgpiYzUyU
LP1WYO8uzHes1eM2mp+r2VH5WqvO9P8VIAlorekSAcrfakUJXbAeIYWgX7+4xj6Y
zGcaLbUiusqrm84TCfTWUvWe8bFLhBXTn6uCFiO429DBuTsGNvLMTICW1LlXHLFo
r/SK43HY1uM08QEp2CMmpusWaN2KLpgwip+rdDoKIguhmKmUBqSG1OV17tWCbbQ6
pxzCSQFiniKnYczox3bZcrTbUVyBttgw9u5O+wquGPaArrp3b6kQSCStaidJQi7I
RQ8TMLUahkX5nguD5kOIBBvDi9/KRlvPpJrb1iFcNF0py6sW3iy90m5YJostK4rJ
lYeeJuwPsvvxyomEr7hSOfFA248V/oegR1YKoCHnpROpvyg/kWXZJtCow1bRqoQ9
r/S9aBKiSnqeS1I0GBx2JvYM2tvlj5sYDEX3yIOWjnk2Kvg8Bf260NqN28qoVRBm
8iIc9wjxy7IWfSkNh0hTAkpnIvx0OzILfQCwvIqGMjgtIdgf9vvSNsd9mwE++KEo
+RMicn6KLwDalz2edRgDMPZitjMjJnTHtwbGpR5o4nEGgn3GmL2rRbLKSThkjCa/
Jz3QXAWrzuYVAGVjRNyZO1U/r0TfcEpe9ZzCXSDQ4noYPeS6DRq5OAnsPBKRH5Fy
njMIn3ukyNjb+y/6oXjUrJbPFwFzHC9wr09PCMK4NGmxGrx8suHV5Ef3AWWdCa9r
u2NjboalCPSF2wHHS4J91879UZBkPc4bRdpttpRmC0UNjz7Jlrkvdr7RinNtAIM3
fP7OgoOfTBz6v7H3K6bABR7fwqu5S/ORhIEYQp6UTRqdVHpr46qa7t67iv2zLF4u
drYQAS7LwrKCu2OpQuf/8vIPsTbDrkIxvFNL4cdh+yYF/QBk6R3nEEus8oBn3MU7
P3qLvlXRwfKQOnd5QkXhqH0Crxj8xYFZ1l0OdoUbDiquwWsL40TLJyQgzNNPbF4d
oAj/6QGa34FwE6KoW0hBUmbcAgRtdEv39QO+YbahFi3r1cs8HvvEQbMCfxMWd5vZ
Teco7hrrpQbSiJHz8Gf066T42yxmALSLItaOqxzegIuS5/O3JfXPjCwVwj6b1pRv
29S/RKbDqtKwN8PALZYpszNcYLNAMMrC8bmMbYZa6LnQgbC/wrtPOU8fqLPOdlEe
eZFBWIZuxP0U3r1KM8Wri8YctHSS91fgeRq97oqGypWV9lq1bBxAJauc7f2ivt7G
3zDUawDjGbFm1swciNKWyaSQ7ASNFjqDKLbKCobqEC2zKMz//mGB1/htv8ezvnZW
fkou2ekzHGimcCOO9t8cvqM/lIDQRQ4zYZX9eZbXyjTTut7j9JLZVJFTdIyMtlWE
Qpis2+7arUKKU7VUuTutI5P6Gb4f7MSIoYU0b+c3hjtr9M5NpHf7i8PYoj9p3xnA
qpGf+M4CyRGCRHOPD6ReSYuB+IsXWQTlGDLRgU3zEEWWjpOAFFfxeCcCAjGaGPcy
PS9fgXjzIS1CVK0UzDbgR7wWDZCyZO4r9Gw8xwdVM3XnmIl4YLMbVEPjnrbY8w+Y
NQAVu39064HA0pSesMQHqx+fannkQ3uduhB7yJqWgFY0S4E/9Krm2cdCZVMQyl0E
9ZEc1MOZ/TO9Ey9kzdDLWjbn/XNOSkI5xKE4QKunUvvOwgJU19PlQKuvU4BoKgqv
BuvnOvcBCqutQNjGTI+TUPb+ytvrttautdO6xmfw9hGiLkvHYYRPpWnfaXg96CHv
s9KupMlP2KSxmX3HFeOMWLhIUVokcISaF7aaAK4h+a0R/EBo/tVjxnsmLjPko+Zh
dUgxm8WmExDKJ+dKMEavwGBnT27zps2/keRqcjTOrmzXROhIbFkVPyx2CcXw0ILi
n5MsVt45p2DIWAhXSJ9PtR84X43KeW9xaMcJq68Z2ZX2qtMvY+QjQ3E+ACPRHkAz
FBCWGUiiSGmmrKDuWBJZOm1PbXdZojDaFhpF/FJ14YxrP0dCiVf6Lr02hiyJ4ypv
scQSqiN1Idd3gTEkcaiC5PGAuF8otMlttdNAbgueJnVEuOmTbRY8UJzpNzQPkfxG
Ie3FdF/Lep/muFIXy5gwtPzdDLVhFr5wh90sHN9BZh8geHbH1oXGHl4Cp8NctW3h
vN3XmIYknEfaQbengJ/k5YyOROORorfVmhcUOifEz3DQF/Eze8j+G6iFOL5TtXTJ
TDF03uyqXG6W9H/263KNjVt6Y1KxmhaQ5t7cLIv0Octe7WUO3H0bmVI30QwzSb3W
r1cmUwOwgT7ioD2UTlUKck/92tnEW+QwUU/MP5xXggLfD1XXdXCmPXZ7Q1BEBBPq
wLyOCBC6iZcqJ2w7RH+Z0HlTOut7HnQxyQN7IHQbciKRrnnnhnJFMckkGOBh0viI
ZmCUWmRA+5N3CGPVhoH9rI2tI50/dg6AtAJhfgFZN6HF2dLaQzfDG5kZ7fhwIpPR
Qowm5NJsIsIIMbCEjnhU5mC8fCMtWq8Dh4/dKCAFUxs+ZABEli5CHkk0OitnUXeF
dQtq4svqKl5cWMTM4iKflHKO6xWH08jKHD3zB6+cJriCQehjmBNgFVMcV9w+rAcI
uNi5LoTs/6fK4tn3900r0Wfs3/JBBGouJk1A6AwFoEgoh5WqjP0YsOridze9Mp3G
6Ie4v4UBrrxmy2lExi3fYLYhtBHRdNRpi0/gkhAUgloMN3jUbdG+5nmF+DjT/8Fj
bJByqW6yYebyglwOHoa4oMzjMR76UDLH+DMYmHyRjbul92dNS/O1j4RukJBE6lpC
uqAtecs0+zxbkqtoGKZrJnJQv9UMmnPmgc++GqVMEvt+GFMR9Fh2Vkdul/SQu+kW
r70lFK8jp2zXNFy9Int9dw6yTt9ZgH9qKBKl+7VYt1kBuAhI/+Kif4szAiPBfZCj
S2OyejKXCmIlKfnCog0hQNise6yFbywFXQHF13GvaEo9X9kOdesisvsaXYLMDUgu
iV7aqlz8tzLrT7CuuRzmWuvToO8RecIMkD2+glRgAkZavfmNx9eNquGYLZWqypzb
814XQ29/E4R9ovcM0ol0VNPu5eArHhA0GHSZj/Fcf5JDE8Vq7I9OtGO2SEvfeMBN
F3azNfbpDNFru3V+EAo3KVUsAEn2cXqoe7J172bBuheCMA0ywF3cksZK3AShY7Dp
h4UWrNbugKPE1W9bBrdQLSZ8mh66tqjJoHE3cYRLLKdBffkWrZwLycZGCh2Z91s3
6twFPL4JcXpchAmiaFI2gkHaIZJU1MqFyOKSAGWPwgkTfViPqQvMd4WzIAM2FWWW
lKksZ0iRJBYQqO4Ku+LK/35YScAJN/wEnpmYAZTjzrHikYY+Ilxtt+IP0F2M4o2b
MWcrsA3Qo1b/nGQDDRkbnoBT12HygQtm7ljRUmO67fvf8OCbjdalmw5MXNddm8Ug
n15M49g0fHn5GM8zWAI9PGr0cUSugJHIuOTKmEdlu9YowJ3zHI0Ob16zDfnrEIg2
V1/ji+UOJWHYNb43EBD7EWYvsTTQfkHmd5H3XKmxEgoCz1xfrzH+EZZ9WSypSiu8
NC/RE+lrRiLeLkMS6+BaLUdTNzkNGp+lL4sziC96RoJ6UEXp9Pn7lsEzLVnbq1IE
q2hGI3HPvqxFGGV0opNXp///2LcLpdm4wEnWLuL8hpMsfvSzyeOj9Nrccmy2/0WG
9KIZ3fbqpmBLiCLl6bablhYJrxt/O22rlg4QvyMu5E5P1DIxLPYb8VK7TENDswto
nJSVmRLSBNitYkkfaJ14XF/Vr8S/fDr8E7e+Oa/MP7+ifLun218Vlns/Boo3F6eM
qutAJIqozkg8AdCAVipa4WP4r84uLtgvrAcOhaBtzy1MKUmwxgMxythgNjMf3r4h
+MLmHgi4SvLXPgMsJaHidjhZLiKrFZzzqL6DHi3edDnq2Ff3DMaXFakEi/jM4qQw
2lT4mhaVzJzJMtBQ+jxGJvsP3X0ePhbahCsuOj/JW8PhGioyHLxLMUK9dy4Fv8tG
1dHQO9LgjrEHSTIz8DWDfYXpr0WALScSUl4NweMAHU6GEyfQbFpXWHRwYegTb1ju
kIU/m35HUz6rVQ+MW1NIwNfjS1kyjo1sw4gfvNysd73X9fLvO/ppt2LjBcpbpkcq
IcR+6kmfUHvpCvPcaKkv2VKyteW/IROBv3wx0xgHzNDDb3uaymlV9dWLManSHshX
FyY33otZPm4YGiAjjAf9md2aZ1o2eaz4uImkKja1hdQ4IJzVsZuiBt9Zrk63f2iK
uRHujtkrAJwyaqapXa7z1tx/pwxoeVTe7l07mlPgw0nMTH93l+fwunAY4DyMSzld
Dk+R2JMh5r4fpjxCm8cyhaqkOar8j1TUTrmVfhqJPkfFEv4eCrB5bcdihpEfslED
MJfzQ2SCUiZK81U/Y98yCm7NWKFSaAOjM2WqUdHX5rFD2uBSNZnWp9ukOEA9DCW7
HKuGwgXAYyVIwIrBYOpPNKeDOnAQdads6oBi36xAb24AR2b6TWKefTp1WmvgAg5k
dvtefx04TyY2Sh7vs4AHqT9nMtZ2AVEPFvNXE2hOo3ltw4LGj6Zrwg8wImiPIqbT
jiu2PaEmcaqUlr9bLToOrHfFjTsOUyxtqrIq+yRsXF8sFx3w6OCf+dJdDs59/+Q9
c4R5LLI77KkvnFKwc2h8ZOgW0qtgytoDFd9claYsAw+v6mVl0UYXFp72ibFAtnpA
rx+gbDPuTgQlFFHoRzMm2XrbUW/w3uShVfxXRY4G9r1Nl05Sj5bmg435VINaXHZX
7TY+VPVCmaYIG1iiY1spWJI01CgoeOLbkqb/9VPXpaU7zrec+UME7CcffnYKze4S
L8ll0dJOjsE8YVBOURLmSDdgg24hSnFwk+3Aqb7QOT4+jeFp7sHks0xZXIwgkaQr
3NQVy73uHusOaGoCTUAV2vWDNxgH2yd4nXToRnZINKpGvVhiC4/PNQFhJyIbEA1w
POBW3FQ4dU0k/01DFIKJjO1+kY3RMmv6SFvNemTbmr7T1TGbqp6HBl9ibUokzpt2
7Oe8+QKZYc17MSXYDuV9HKqg6O9KWvyCKOg55rdXRdWMP5IEpqtOBIY2HJxizdw/
tMl4fzw1nDNKtayL1brtLgEhqr2wLia6axR9Y8iA0THbL0Wl3O3MvncMFFHa+lSr
mt3I+HhgQd3zFvx91B344tST97C39uk3wlEgO4sg1NY3TX5nJ5pzZmy6GpOAerAC
WGJDcKDXL6GUrgGUTuMOoEOrod5zOCL9K4Z1DxspJLzCs5Qhl+efH4q2GcKeUZIF
vf4CO1nVkFrx7vE32ohbdE1qvzvPrRVqHKtdcz+NEVTgusNZNSygmXwpsjnFrmCO
8h06DTyczkySCSuzrdg2gPxk9WIHfX2ZS5t7m8NCMfVXLFH7y9p9PKQk0aAeCg7z
1SH1MM/rMaPx4hfH92jZ5T3hX/lxnzeIIhPKdDUhOR06a+7lV9OterEcTizygV1X
rVu3oSvf7szeDkxKBzbGBn7dMcX+pLD/cOE6iSOY86WlGAAZPQtNnudJktVged9c
dDo577J6/cadnaK2d4aAwZM7ieZGZRGc2ONmYKtyLlc+HW8zw/m0WJLil1GMH6oM
utYFoekE/Wfu75tZsTAkC9DdQaQQsK7RKpkw4CzSSmZ5HrGZ5/YjQeLKQ3YRtPpw
cmDudfJgJCTyKpuqxusoXq6MeG2cZf9sKkKhj4p7Teca2+IyKhiU20fhNZEpUv8z
pc0O2Na6UH7Eu+dZGL7y5JfgeTSUMvC+eNjOmuROmAen6pAKw8MjTapjC3QPOdlq
ac9xPoE0/3RXLlgxZfdnNRPZ+Kkn4eg5vqRyrF/G7K1qFCjwD8BpV1sR0Mu/stZC
9FaDAu0+AC4xQp9O5ZQpwSlw77D63PqrXBaHPdriCgeDiwgbTCmcxk7UnyCwbGbz
vQ2H328An6MjHkRqDanYx9mKDxF7TARmWHHjy3aWnERodFGXz77RQJrOVdXZ5Wt7
/D0mfMwXR/I+BptSlbccbUyHqZt6J8mBPoMKpDpk+ZFfhzOHIi+kLxrNy0weI3qc
oz8OBpLzuMOFgFMqbnPoH1HaV9DJYIyFi5c1HNq5gobtSJgfWjdTbNjmlVJUA0QY
lVtRg/BBOMqpI13TkWfJ0uaa2cEWEC8JoGOoY9JfAQo8IN7zazQ71OFzymDkdrdu
kvH3ZFTKYIwknXCH+hu2J9Nn2yxHMfNN/3LqDEZdAJuVothQrO2A8LVRoMOxe2YH
QCuU4lk1jfgtKgF5V1wCj7DrVp2lAvVogM1Udyu9ZDusENOU/DXJ5fP5s7IMDcEU
rnFAX0AEYYuO4mvmJ8xSY5ztApscW+jJzgNioIeizpZaKIW6CmdZnQnjSe6ZORmv
o0FhV6FxLZuyrSM5lmA7pLmJedH7ulBDD4yFTGR+9+oO2vNrUZCz60TTnLQX2PSP
NjfjEP+adJBD3rZjBV5TiYpMg7eVRi0aQGo1TFvBMuUzEi7K6a7wJRKlPkQiawSL
uQNzWEQE7c1M3oVvCTfG+5N4FytItvxt+ky5nPze0s18W0jxfeNVIiCiCDQ2zKil
So8eKiQK1HuDt6lFehVwQHCwB/Nq3Ka0FAmNT7gRVPlCiGdJIR2HAqUAh/Spn9/O
0U+k2tL0goT7qOYOLSlOo+0+ZM2K9hXjvKBDSastvR3X5k2g29jBLwAdYzAj/DM+
zlQ1Tb3MFl6v7fD+Noh6mzRlX0fWHTz8ehGsTkJbT6RTJnRVOuVXC5xvq+Fga/kt
kqKD3VpsQSrpAP7VmyPkuJYild2yXTA3A7WWfin9mIZWGVzvmeNBgBEI3qOfyKoc
TasXmRoJu5NjtuuuyOVZlk5TGOghL4PIKAkU+Yg6Gj2kBgJGStba7kHPM+FH9Ck7
AcRMwtk1hdpNDg2rovLTQYXjGFNcPJxj9n6UWE5lyv6EwaCe6ucGvqSfgDtPG2xJ
H6JTmd8+/XDIM//4s2agWllK/K+tMKLWGHR/plPLt2s2maRaE4B+6aU350mXH6JN
wLJNIeLlwV5uVWuySEpVfhGOOoHSwnd5AjDStyYuT1LEViXEcWGrbvc8Z8tr88k9
Y4BkoZxJAAtmZWmj9xEiHdeLreX12xAzsj/+I1oemAX4Rv5sOm1yP2yd98dtM9QX
DmsGeAafDEErUycXHR9rhtRmm3Gmh60yh28PiVyhACbGgTz5uX8t54eagLuRKHVt
rFfM4CVOAsGUpfN5uoHUyaYhi66nrWAjV21W/uBqTL9ItPUE5C0DIlsvzXc4gMz1
NnXJNWWnH34ppnC0JV4KJ2qiKOAVOH3ebSruAMPHB+pYvNtKM2Ic6PYbszE3jRyg
ZdDdUn9skKm6vwlDhBtruP6QV94ONa5cevZo8xXemUttfUCcvDpsPtEResx21Vms
gKZ0KgHTjldztkafQmby1blHnWjilaCsK183C1UFKANp8QLJeRMDkvnx9QuosCdl
4EwNDeHzU9i4yBZGOCEAGq9qcxXQ+sFvN0uirDKJ+27qTfn5QESXOFhEImBoXVea
0IOjwYat0zvseFSYXyleAsB2zF5mZ/6IR9NlB1O/rJnWlSmeRC+CrO4cRNj6uoMw
2JmQNDhgjFiX1xWbv+r0iAifYgzjQyPIyAs0DIhxi+yOUOh2a6QiYdusNrfenjpb
dzpzv1294qGUmHCFV5K78OCBekIHDpj4DRZcb0U7ixFqdYShC4tc7b/E5dIFSani
bc2VznNnPLxSLzPMnzOPVmgm3EpNwqtutJu+uxrebN0JB7QR66NXCmWLKOqTTJMP
R0p6NgPmrgPntzpkZzXOW48+RS9KDBhRpBMJU45yG5LouDIJ4imK2f2OOQA4/yyv
3mXH0jodjU2SCxibI0y7V0ZW6Q3GZs7eP6/nIASU512yKQA84bOFHwyKiF4a2pBg
O3HVc1b0ehdbNE7Qtpe7ou9vk835jRMaCJZrWcb+8+Uc2npD/akLumbS+eAjNYnn
I5CrBfUqcIUScFxEGhi04jH8DVZBSF95AIwBTKR5xkRI/r7tEPRkaDzLYWK5n5Se
p1lcrgN53oVOlLVav5aQNSwfoR35JlEApzoMxLXPbwkGsnoh0N0u8q+10/ve8slp
WKmJlEp+TWxKbK0UqO+NZDQ5XSkx4GN64oybjwX5DhWjnGS/OLDZ04u2BnmmWDAA
XYegh298N7VTW7dsGPjMV+kXCu0mImGR8kv3XKeiaT//8pCljuXe89J5Rzzy9QgL
bws7aXBQ8gHls2h6Fa4uXjXJ5FRg01pRT9X0IuOInL/f7IeIhmAgRK7+yc3nDQ8K
y2WbDgZZHC1xtZ5YkUOqhFYqFn4fzdjP3KXYk4Zo3j0qcjHbkKuJ4T0QvnLzOazg
O/CAO4R22YXIhbEe6Mq7eLCCDIvReW/XIxW4N2LQfJPYWFrMtzw6dfdC496GGVPE
IA/8NxLhwRkz4GuY3/aSvpQ50gj29nt9TnXq8TGBT5w7auo/7ezPHrlvpzJ/UZ9L
RpbB7H65usBThK0nQf0HoNpdvM+S74EJswmBqD1+bQpoC5R8iGuHU0Rs0au/iLpD
ty9B0pm4u70kTg+zRor9sNxuw6mt+8OJTkn4s9TMBRbT79n1pUA2Asmr5e3loq/z
hRn/j0j3J6MDJyMzKgAwXTKCnRea/aOto0nn0odwOuMH6OyXjZExyiuDHRXhhR6o
BgFNf6hWxPrRuD3z5tVqCbEmad2+8j374Ofv994y9qGxw3sjJiIm/ooIapg5WCtz
VUFeGE02WcAQqJ1lj6LIHoP15MhBqCWiemfhBS9kYCpEd0Fsi1wMDtIPmQbPm42V
y7n9kVt1nwqWWv7KEKkYOBiaccKi1GZ4KIsMiDDzu5nUVW01Tlk4gT9PQLIuCbmB
LAiKdkcBB+1pBF6wt6sWmR2RJ1aha6FAlq8Jw6h0G0v8ZOaAKMuJKMlhYdK5tHfU
m+xTJNcngTgo/qnctgU80nrpTSHq86RtluKfOtatJITU4KzjFakJpVko8qVsLGSr
U8FHnt343IV0e7AsUGk4dBMFq5NZAH51qNtsY9PFwO8uH37DomVUm1/hvd37LF9Q
a0EP8HWrxPsaTKgs1w8rrVKwkdhGBKXKpdwjYg9knhyfygUo76P1HZactPdLlsYz
iOPsf+j4cLF/vjkRXe6P+RrZbbL+8lo2MGKz45oi6ArS2s0BEpyf35NvZK88jEhp
zXahm6/xh+umoI3g6Yurs/u2WgVOJ+wQTy7/NosGLaeh6zwv4IP1foK4CXFrtMwo
fuBajhkKMZLlkNuA7fOUMNQEhJRrgCmOcK2Z4cHpFGO6qBzZPlUN9OurG8AQaBLV
jaxPVcfCGmRSLqrQgA2Xg+wA4DEzz7xj5QVShqYNguB4d7pYNGtO5PWSFZHzTpJ1
zsHDsh2cKY28zms93ABjm2Oj8gClYaDsDP0PGeyrP4AkXF+O3pdaGvoa0grWBi6B
Z7a9sjytBLv3GV+3Rt5yv+i0MXSjhGrLaNYnY5v36uA6oQTMUvDt3TnoY1vvjG5R
Doyrby/dAmVkRzL2Ter+NpPVK6FSb/cTFWNlHRGj1WH2ltoQyeEYuT20bQwE1GBR
f5tPJzHD+E00dmWaSHCaN99NaXedUkkItRYgBMWa1kGAqFN5GzT9qonsM9VDCodL
DSo2xxKkoZ3DW2y4ZIZcZVgqlJ9XUPun9bVnsC7q/6Cf5P9y56E/LbSSj9CZsOH1
l2x5khwmJWghHW+/L5RsWzCUXHn/3TUc5EyL2mnRDLbjOcN6wfVG1be/djWZdbZn
sq02bXIQSiJ9McZEmsQ2zx05lieVI7uFNPb4MgOue5vVYr1Y7WWLERItvVISeNRj
DKavcNM1AaOazZWX3ewJuiORqLSqOukAihASSUNa6tEOtHTav6iSM997cf96k4Tu
SGAHmnfJc6q17SQNmLNg/nnCQZk186bW2HJmQ5WqU7CbcPwvDdAhxQbvY8shhtqL
+0uh4wHDvkURwdN/g+jzS6wBUZLHH/5azsB4B/ASL5Y5TXGsSD/vvby2SVlTGphh
vmOXWbhaf2F2ulNQ4zkhlDUjrH3cAjMlJrX0MCG71sgMFOJeg+7SRBDzE8WUr5lu
mWcmeY3Os8J7ZQVjGxcyIVheHO1u0ZPIQQRLrvqCK9xcgylKTJ2qeinil8orQox3
kTV3maneSYqvzbIClIAblLE9kf/Ii6jlYBX33vs0B2B4Z2dlmdm2yfY9uFro5LwD
Z6FhUxEpamVBFQCK2KmWtvF1JGbMQDXC8SjhKOCzH28Z3hH+xnb+4sAu+Z1O7RWk
qhKIEPMguiNb2ZRXpa6w7MTARoBmD5LkbRm6uyUfbvC0finCXm3tw9ZOIJaMB6n4
kDeBiB/MsbJXTyuhyEwNfykIjRtbjp1smb6CbWkdUR0+Hrw/8dK95p1dry6WULPB
2j5KWjii/xzzdzwr/zNjBgRZm3rFZptTI+zzwanxVPBqfVuDJxjQ4hHLM0sTtn3N
SLI3rxVFuqpPkLQQ6obeLnf8GnVssZFGYQVhKLEBNY10KYjRXxEo79uoyXbpxsuR
jsG70w3iuMXGeRw6lppPOY08b37082KzVN5yYRDMyfizkrEEq+68fSKDuq+dacuc
PobGTDxSbCFa1RItzbbLgv9OPUDj9OYaW0YzRwyzicKYHGlOBIr5MgKh1iqUFftT
KLQHMYnSUw45kXBJlIaW+ca1KbAyiP75eER97N9LjWjd+86XZtz74KOJROhcz+CF
65e2nBhKOobdiehGEjQduaxV3FfVDQU70SWmGm+pTkQs58SyDCLvPguhQBsFQ2o6
al1FiNX1QuGhzVwlQtl2BUc9DElS0kttJM8G+lWBdSd4+abmIM7mSs1cU03dYHV3
5iJeyBkIF5JTqy44FFRRQuGIZL6gDKGyUjr9kY0iEVrgVc8zgYy+cxeLouLsC9OJ
Dk4iIp/eU1PZQh6n+AzfEzBbjGrbOZM6tPSj6/uj5ZXxKRNKyz9wM+E4ZbVt5QE9
IznkF3j/wBgJikhaLKraZHI2B7vuq0a5XoeMYYrJOUD4NG1Dr+s+Pauqcuo4hCcY
DdvN15+Kkkv8IMZSNr17BQcKTeVam/nkv8dfMAVNnKLzLuqerIImpcAXK40Fp3VO
5OXw5sJ+lTfKM6+UovS6iSFlpC2pwaaCihH8gZjcEKk872wZCMSjdlRSy2VqSQGw
d2e1jLuPr+zf4mw0Ae98aBFamZrxHbSBvAbbpCt/t0oUeR1KlC22HZ5b/6/ykxA1
TtYGQh8W4TkctCe8SNmkj7zCGWLkZYkcyQUY2jROeTpFLmRcNhZLIHeOKZUpvQIo
JyYR48FqO85XqM8SaGywM2h/EJKBwgGRM5BPOAf1zaphzU4ZL1KLqP8JkzpB+tdi
vClKV9+gMhUgvi/DPOKxc4j7+JYW/W3ST475PdSBVfcXTJBwbYjaMkG1w88JV9rq
7V9qGnUlrxo0iY+YtPY4dIH5Z02b5yKVtRtSuBge7/rTAuM/BM980YnDiZFZ8nKC
LRIiGGQfAPerWQN79gyefFZzGgWmbB8IAm+x+ytJrnb68FCcj2e6xoBpxfMB4HTh
ol2L8S8KxoqQqj49On45zB792gEWstOKLsj0pjC1/hZc+odL+6sSfb5BZUqpRRdR
x7gLQZwOEnTvWrW4Np+TfHh8N4HY9vz4VSZih1dF1CWw4V73V6BPqmQdAZX3F9NB
fBInAOTNimH/AG/yrd6+RzIDjijjrMPlbifqLJF5aNyc+kBlAAlxRPbSmhUEnFw6
8GWmtKNWIz+y5lyKff+mcFXrzu2XLoSRm+/pHzBC7wb9Enx8J/vZaHUbjTlyQSPD
dJP3j9k5vZFkJlyylzVMPelg0B32aX+ZYFi+aXP9Ym0Y4wUBK/d5Jb+x4ZFiCTWO
SgS06nZmDWCGU11UtAOT9S2rMHIQ7XOD79XsF21YIT9Lt1cKq6nmcG8OeH8gF9kq
w2JlqIkbQypbhcxq6gVFWWYoSe5Tx8xMyMoGQNY6G3Kccyv0MQcyxMC3jQNgGxka
TBwws8xayMKvhPBRFnopMxsZ3C79286kHl93TBcW4fyKKN95Jx2kyV0MEa6k52nE
rE2OhIdGbeojVjPAQnbjifG0zp2opR7Ax8GIOR17kf7SVYWzwPcVhKJm3bUle5J4
NW1IEQDtOO/Q73WSMkdbZTBkpnLArRFAU0PZJ1Lh3enLDMake6hOAKRpfCxZ2c5k
yvvIIXzemwpKAS8dosX2vzXuAesfMX6uwPolpQ3yxQEZaQW1+24Sz54Ztju8TPm+
6sTf+zUOqH27PVTa+3uOyqwhDFfElc5kyXP1Al4qmjXvegGA3Go+34Akn73PBlxJ
fBOYxbi58B4mBFf6ipwEI8mR15Z7os10d9wMvfWxvzyS1OkyBbjccqfbmPNw2Hll
BlfNyPG8tkTB94RIcPfld0OS/+2AtdOFfPwA37xKnF/2YVACa4qA4NPUPaNguO0H
Rq9CuBV4vCGf3oq3CbK/msQcY43JdWUjRei4GGCNa1jNVDDB/l2BNpjDKly5C9Zy
xmuVFMrLNDY1u/OlTX6kOSWZvK3BQikmn6v5fUHTQIZ9KDzuG0/U0HhjzU4vF8X2
YXsBa70ZtJt6MOig8u5PZMZxOxNZAHMKGDJe3/gNkmHjUxiaWezdUrgfQ59fLktV
9rbawbGFGH7X3OFLElDSO7M3KB5AVBSQE/PKj7O5sTMZwmjqDsaoFT3F3tL9Ul0L
tDew3wZHTZy0hgtnXyzfoLCk5jqGI6bHp/DGyiS738fpJg5+m5rnPNyn+42qxhan
KVOpiVLyGknl6KwFDB+xcqg5VjT7Csln2fjCPGL140CbhOLLYjFVe6z0o1rxiXow
r+kB8W9TZvj4hfAeBwpt22XWKzPSMfQ+SyvZDedR7r37/gkAFp6e1Y6YyjbrrxHc
9KolRVjUwuj8d+k80296vYcgokJ4JScChy0GFIIv5yo7DGZ0oN9pNbolVhjuJspM
D8vj9H3hUZ4NLAU8XnDg4OsIAsgPRJhdNX2fpfTr3DF/JQajEMgfuaiGsKkDnzri
Wl6ieNmIk8pNqlYEiriqBaA/g9OIN8wxBCSXiJ96VqXWQr6y4y7El9SrW/UBvWwL
itYnnOb/0uK0Z2gQUzshLt9bLs9ZgA3PhNQ1sWJoVsuAuqTtPxaOJxtnQRbEnHQ2
AwrPi0EEz207r11LODRUubptvblQtImvi0LGBz8vq5LqdZsYl3SEto6JTsME7o5G
klkJOTpxCgy3afekWIsT/ZlxK4dLnWWIDuvsj1XgR/icQFRQls8E9sIWN4wEi+gi
2Oqjxd6SpFoGluMvP4O+y+9HT/PNSAXM91JeoStxynnpN+LmOt7+7E8zjwvWeHDQ
bJN3KdavuivTWxTj7OR9VVWoDbZcg2SgT3ovl8Ea+SZUbeHNG2UUSHGu+Hdw2ggo
OYCGNuT02eXeXsqFQ0OKERe3mNckKkS+hJXO9OirD2a1lQzzq1SwCQHYEMYOVz1o
6bdsLB1RVAJTo+rNMIN+tbpJXjNqvGHsLh+L36Vtun7Itlnbw/t74X7Y2Lf8m7P3
LSoMAP6gOydvT8byU0OkScCyjefb/1qGPh3Vro+7rlOhniFv02NvqHwVmfPcmH5W
Q3SBSqUDK2SFFmavkYATdLIf9os37x8wDF++yg/zDtTiTJhTY2enwzxxjThVPcnI
RRGzAlY9v/jdUi4PddTpruE79IkrGVlwLbp+8gYJfRzT+wfOTZ6EmQ7t3B8gb923
4EtaKKqRw/yq+2G1jfws045xL0E4pT6sIbmwieHjgEMmNZeh/dAXQaVJBSFH0uAg
0j88U70Ha7e8XSyn7shh1eaiY30ny8NeHhHe7kUEHEjwAKR97ijhe1IuLtkrxnGo
1Ktco+XPLwYyXPS1zXrMaPiqctsjJilIEgqozeQkMBeTodjDG3EEBvmISwi6t69O
LDbSZzFM3Se5agIhmGvf3JyQtvGoll+u8M6mATfvJzhpxlXC1rnEmUpXNO0hxIf7
tLGr7oGfgsoNjdNfSQWPY7i2GaQuNQiSixhl75txGBOWjQL1LVaLcbN43o1Gur5+
gGcPgZXoPELM3S19VZj/KldDFpT+kxKK7fzgsW3eBLTuPs6+fYz0hBpzEu91375r
ZU3NK38gwZtWc99SNt70r0lC6SKQz2hgC9H0F/LiOHX1t3YjqmXXMnim5aP2VDkC
ksMU5ch+UtKUVHOFbmle7HTyE4fLFkKmME8NSpMrZESx/eEEjYb7UuNEHySkDJ0W
hHIHTJRRWtMMwUuB7m4+KuDggKko+gcZiT9yuotOLZfm1QfkASnoBK9JPeK2pr+0
UAc7tQ0gnr6/VwmljJB2VGcv/3Ill3+kiCkqpeilvELnjY559YZ9bUxh1AxiL+mD
lga5C2qwo6Z0yvNk31MLvHbj4R3pWb+lUc3rOGDfmRZQ3yRFHBlO2bSkSvjyXZK7
oj7m6HTZCZflY9/zuUu9jgZN2TqAYovrB7TQ/1/NL/+/mlyvc+liJu20jkLjCEmx
ayZDG4hNJKL1Dwc/wscP4ujEKPQXW5StD3VO+VT3Spq19zCKiHiucLlns7xnwgNw
FScwWGCPbjw7vF3QoSDQ+PUwGYVdfspKomx7eOGP4r+ITP/BTbVQo2gRqDa9wtE4
b4IySNsekwT6EpwXAF5rVE0kuBN9764PGrgk33qA7eR7wtk3KJga8tLGWMwyirhk
BC6aFzD/sZ6VhcFKuFauioVocEkL9+G4iFpg/r0D5OmsPvjttcZHHarmj8FMWydS
+vFO7TmObK6EqJ5hcT7kDQqVQniHFmyFwETKfKjzz1Zla2By73peiEP/18le7d18
U3+vnoQvnfrmEIoZJ5uaKnrgx6yWLiA8qW8vJjmGad05bHth9LEXN3QTvBLGK8KQ
6jB9t3hfjQvCk+QYxeplZQGqd4gnL41w7rZss+45VpxXmSUn2OFB1SBFmJ9iANSc
2jU07k8les//CSpvWyhGa8oNwyOGjYsoUTzkiEl2dTbCV+g9gpy5lENwcEsC4Wiv
PCIGMtwFlpDPBLNIdOH01yeogRVDkWZ9BNZEXevbesJA4OpjCzGL0uihCgBBUFdS
pEFpfrE4bwe0Jalm3VmxJOzTqS/RaxSuUu8kfnP62i5CtWk/W8Kugxjttb9eTDhc
7M1cp1B4agiEHq+nAQB+aZW+ae0XTLn8PaM6I6EqpSCLDfoSxcDIeLss0IZAkWap
ksyKrEXq8vcQPNb7PeKaI48WdciIb7yPdRq9u3QlHhGLxEIKtsLt8fqSACoZ3Gz7
K154GngLHic5CSP+sk7PiDWe1WtEExvagOZC5kX4i17Mxe3+VLalyuYANpWbmsCW
GWLLem/z4/hWrl0bm/IeWXhlr/bQBH8rXzOB3nRQk48DWHmg/khRiyInFHx0dkH0
0TW0l0aYEMtpUsh4gCy1LUTyhU7GmjahQ6SDusFxkFn6kJJg8xoHApraC09LCSWr
yFI5UQGsvtj4a7eKdIKCIOAU7XX8woLqDVhg1wWedgx/cnKmYXNo7PlHaI/pb0s2
Tv3YDPFsaS30P3D5oz3IrIeFwV6M6hxAXvNxBx+zeKUgP245IWWpdu4Vis/3USCe
grp5YTBY2Dk1qznIDsutBPSFkAmgik9kHE+FOuBKHPCcbUNfbctRacH4Hr/izJgA
OxzFU90whvTcPWc1OCpFZI3Da8r4cPilhSjAcIfSSkjZgORA/Yu2tVjs+tbse3at
2iPmghuIKWRTvwCnqIDD8HglpJerCj5MJdgudFvoe4qcD4LFnrU3al2rUXZPFNMZ
qJ09urGRE+tTrV/SXhydK94M5wQfk2aLtexuZcU5WPsb2U278Xb/TgUvPPJXSYWk
Uj7Ezm1T6Rty/CiyPQ1humztQE91Rb8ryjU5OUJkbrtgaZPXfEPGIAvZezdpOXUd
gmuMiLm6ghktaLGrnwtmDw16+K1aDPJ/Is+nz2Xh6i7rCsKwIHW3SiPhEUnun5CR
CEbF0BT5ZQ19+sNNwQV7mEdGLcfDHiIOHYhyBz1F+qqowkR0CQ/O++bhtdk8LzL3
MCAIwmRygu0Q5R5Dk1JvLsrXqAdN1x4DrXzyOk4r2o5JTzdro0kpC40934DInG14
eVVkw75emBpbio3RcFG5XJH8s0ByOMY7lfiZNOaTEdFR1sggxF6CjlLklqyNwJmW
AZ/ShJKJSpxYzJR2QrgSo0Jh4AHYn2W7cwSIPVQCALUrk2stMQpaazQKgqarLFHd
C5mr+qKGbZGc7+tQoQ15chtFc2d5wygkxK4Jv4LTdqQz9ZhIciHRGNXZsK2YiRg+
UYNgcey2idz/FVHpg/2cL7Koo0UP5JP1yVGgA+jGPLkKyL3ubdfTd0Az8y5hho1N
HTOIqc1rh7AZzct5pK406XPOvSVcnnahzrcdv894q+N751zGwvARSCbRMgpAFNqz
C25yUtcIk027pRRvVYQn1cAjphgagJ+Z3A0lMiphe8p/+KQ/qPHV6+LiX1qrqxV0
6LZ0wD9LPnVYNlOXPR56nbAvuszteJVJ8ikXVPR4Z/7kov1+wutczvezuOUI5cOa
8lHS2MmniMHb8iAIG/wFBLPOiW0tuOQNHlnXWaeC7JUUIM1HlDYI1lGmE9xmADND
Clz5RUpE5t41uzlRuOas9d3Zlqpz4HIZHeCtSl9+prifqhq6xK0IPM+jRr+xCsJz
/AnHVHw6WaqaMviTjq/gEiNfuYqmghCzKCt6FWvWCN6qeHYGLXMnpeOSLuy96VDn
mZfBI2ZltxGGmcv+LB8vquKSCunWOf9revf0NENOq5xBEVW+sP3R5pfV6a6bDn9a
GWAX1cmZhEWG+YNwKTFFXAmZ86n3BnTxhvJoH9bKSWaxHLfm/mraDNgganc3Tj7i
8oFjJYQ+/OBHdGbqY4HZd1UpYPNEIK+S97PCoH4VsDLAfiGunZ9kVTylvz5XGWNx
Ax6pdSxVoRMr72rmcaHAa1AqERCdVgKjE8wpz7EaKdHLGLdmWhB68Q4krk2C9gG6
uK/NuXDIhPAPO5g+tb54s9P0buGhRL6FuPb01MPQLuVfcgnXEyqFRA4Bx5Y0C5zU
OdwBm6rYY/BBPnPH81AUezpmFChseOcCNR5LtnBqPVQnLGMDpthF1/2bHVdXJtr+
z2CFPsoQOiAIPSNCsDqju23fkDaCLLKisz/E3ccq4zy2PtbUBaUThGqAp5Q9Xxsy
iq/0JDMew9LkBWGUKT1FggjR6g+YfUn1JWeMEHPwQi02PMvEso9h2kDWomJquwHV
uYU+/dB0cdUVsFzNZkEvU1czCVNypyBPh6oTVmKqJP4wpZPSxxislWrN57zLsh81
q52M/blvsOjaSCy67UhkuZw2uhkO47lFF1aGgccRi1ai8cm9hBnj+7Glm8NfRkW0
oe4L22V2GPYhg31IoL7iLuI+ImD+546JLwSOR7WfKECQy8SkUgTdGagL6X68pAbx
KOQCZYrnQysrJAHufk/2iVSiqJW5fuNa2OK9Ky0Xu7I2D0rsE2KofZ3+G31BHH2R
NwPJOLDpbrXOhNr5aF+pV5ilUsi9RN3GpM+aYgPgFOZQ4p2LWiU161h1oIXiP4y+
ghxQPYXjv0O0YCxxaSG/cLBw9C5+HU9PF1mcE65a/kOmlzZyDVKX48+vMHQtT0UF
dqx3s2tSk5Q2YHSyUis9Wk0QOeOPeO79Izu42tJGpyMD2E6w2Pr5FsfQRJO/Qs5r
zZHVZhvmPl/FOv4RacNX/giAF/WMrs50muMMr+THeNt0fIMhZt7TIxL4x+woUaz7
lWW1OFZRS8BgOXhOVWEumvVXNRtbk5FFrZcCIJdAysOaRvNdEpt4lmPmX27Ll5Fy
gCwV3YFWGbl+p4089JnRIpzJnk9RsdXpgjTPynTQczfkQU17aDk7YSz4gZ3sD5sl
5RORriMhvZV3fnMI2uwKqdEfnYW7HNxT4N4NjJ29YFRJMV3bEaC2hlUYsxSYuJnS
sYz6cJSia4C7U2FBM2K+8ulmm/vrOXnt71BKhsh1VyDzWUBoWe/hxh0fHwcdtFjo
W5V8zKJBkPaKbN8zFcnds//kRJMpOaV0GnINKVm4Lt46rWkaQbzI0otDcmAUCYY9
4CgcB6UcGcYI/wJfSsxsEEOBjKXWcqtcXsvND0noaRIRERo130ZyJJjLKJVQZM+t
sTXPBfCtHS/cpD4J6YeVLm8/sKkXFyxg2q0CjHBFBKE/Pj7l4DCYGPnkv53J+KL2
Ktvzd3JonP4t/UOJSVR9eA7XtWW6QNbs1GQ9fwBrVc/ciIX4waFiF3l0rV56QFhm
mmsz6ew6pSHGyb3vWDkM8zcIQyxQzFcnKXOSAHnvUqGvuCJuMNRQ5r+stRO+uVeh
Ui04n6LWiLd9fwo+1mmqQ0QNwsXcmejH0U5ayFKGqpT7vnlIFqA3FnEP9tg2U3bk
+4IxxsmnZ2rGDyRkbuCkRMmBajcHM417wVYc0r7v4GY2ESkGpsyBX7qVnWHOmBwG
puO2WZvKGR0eOHJCZZ4xPV4JPeIDU+nMz0+KdJnK7jpyfvIOWoC65yo/35Kv0o2s
BGn5JWDG602ee2ZfUxN6ueVs8XSZbsoAYF0cBiezIy6x4oyYcBL2epCKY3WbQ8Vd
Fn7fWCPV/4gqB84Qyih+fbbkCf6BrPT8BzIHT1rwxaEfjUkJW867Ckr0630vx7mc
F6gY4C3709lwKhaO8BlARQtpruiTotP8MZ+16Y1YB7Kcol94RngD0Ak8vzZM+/+H
zm2Y6cF3EAmfQDLiRT/dM4VYnFC8BA/5vOxMf5VI5cnb4nK01QyiN/jeZJHVqV5o
QNnW9V3JPRYWjYCSwIMzTWKd5UYuFn26AARjbMYdYtKzj5OmXOTCO2EKHUWI7zAZ
KKkdrRcy7cJTzSiN3TNkP7Kthq7RqahoqPJPPZ9XyC8cHNjjd+mbHYYY42+oJX3S
Gi472f45jNFKWYj6L0PCBIF8TLaxpqRM+bzJ2gRTGAzOorVU+XvM/OtS8CgE0WAt
DNdFnM76tFdMSg0cCVZSqmNiSG7OdtXu+3X1Z8N738XpCkT3rfGEYlhQA6/ynoqv
XdiXQ03L4L5vHHMwolSJZzDO+Gh4e8EWDACtwqlXEeKsQumx36SQetyqp6Eq/CA2
iQaoHveLSB3s4kOJLcwGBAVFTSnRwEem5CMoYneOGnLHmMhz6SC91K1CVFBo2td/
SQ2ebM1+x3jh57E5nPit3uYCU9qHOG1C6pxQF9GodokVFHw/+YL/IJ99VyagHhzH
vBUDJX/VyeDaM5jOdRj88jMI0ECK+Q/QCqa1Jr1DkTJAK27oCCBBpdh0+nr+fMUp
YE+Mr2yKsJHSwQS6DwiPr8y/Y5D8B66CvJzaMM51TB9PUEXUIO7vAe7qhYQE7kCa
rGVeYMGfND3pApwiSROGKAPbOktyeNgL/SnOOQ/0GL5nFkbu1SjiSVpUiOY/FisJ
y98aNPybp2s0lUfFkg3XXgHjOarUHi6vXgKwekc2pKz1xvzYF08f4LrhqAZ/C6U7
d9pMkgs7RTGjnGHG14C0RW/cg7TfydoABLbkcbx7LeYeQDKMJpJt6s9/i6a7QPJC
mJsh972whaSXRxSSpFLnXHi6HQdBNaU0t6gqZAO/29TO3LA6WADllbLcHRvJEdce
J6QEA4lw/AofXcN3AOP1ytQE0aEr3mR6jpSvBGpMaQHVmJEBXHPbw+xxf8QB72kA
Hpe2qz2ZLRcYmwdFBjLnCbe8Sv2lc1Fn8KYqF6Fzz/f4lbosM830pfMU1By/8eCd
BCUp34bnOB9y9Rw9LRb8PWFXVYIIGKgjTvdaSeLAOjegifXOKMClrbeH5uUZMJDk
6FHMrgvAt7vXWXOUMelRj2hUf/qHERflMSC+OXioWtBCu9F5BBNPKBZM8xxH59hD
RExcM8Ohgu5P18kWeU/8wfp2nnFQKcvhlrBzaQZ6PR7oPgylMPE3zD8yYLTEua0v
uQPNiuuU5P3j8KFtjVDMluW3z68ZqvZPRUzHxAZaAK1ZWtxMW8TLVThvndHa7dfO
TFZLVnRlLtmi45rBYM44c1HN6Y5MALagJRaMCItsZNod3/4KJbCayQP3O93ErciV
nCe87muuokIphoj4XOejxkTTynCeop+aH5br5b/ZLs/vEimTDbwy7ajYli4IgH27
bCGryyRmBDC2BN4dhGyB6gnsVNRKLHBUtx2SW6jXevsqF6xnbfSPYVnKaXImeV0i
fYg8y2TPS9nYfIrf5sipsA55JSxJuTSEMMOWNDGdmN3plaO98/Ze5V0ZYq87F97l
unHyy47mN+JGMQxiJsbdecMSET4Hs0FQs2cjDMWkcyMWMdIldN9qR32HEaAv3OCF
GlxLMQRsFbtaSlGZKOyQRzV2TXOt259wAT3G5Eg0rOdCnpRyk3zKl/99u3Z8rd5U
HfrhSaElu1kkcTrN7IY973gM8zm7oH4HbOI24O1+Kdg1OEDbgr5wBA/0zjZSjJiD
rvD6eNu/NEr6xnIZoiDdz1VrKJKcaJWw36ryUgs21GuGZ34C3gTTuyRcvTQfBFh7
4tEwW09AiQUBuQKbQOiKWpu7sxhBNIiPbUWzcdXJnsVfN6F/NVxktpsFIuv7qIz/
S8xVWH5Cv+4IEMzdCU7UDyzieGlln9ZaiKfrn7a1qDo3l8/2lLOuudZFozVasx/Z
YVK86PTSQcWRrbpArHkEcZRwunFRW74s8cH36pQ5/NH1FyfClFebCCTbVK1Qg5sd
06NaapRAP6s7lxgmxtY9Lyo8KOw6ftO6qmYjVXablYFTDRg2iha4k6Wyuz9k9LWE
lr0l3spSq29xxcZEnRws0BZMNUVkneCeh5SjZblOul7a9TCNgeaFcaPMDNanOJ7P
APk3aAN3GTpL2VFNnlmm7P2nkqY8Btyau3BWOD3fHpmwX4tJ5+k5BlHJ57ndEvh5
5C034zzM4klpTDYuU8XE5HKG3g3RN5jZf1+5V5m2vdDJ+FvRBUxi5Ysu3tZhcykl
VJLJjttWmftIYjXXq+7tQ44HQxBaHfSfQdcILHP0WamkfdDOaNNbW6pCm6+34RxS
ZtDtlmZRwDwW2a81M4c0bOap5Twl1eDHcuBg7vlLm53k04NT/x3EixXuL3BfcFW0
Mzoix+/X5BQgdXklpSi367C9bd6uo/r41dTvfB5p7ofuXukA5cAXqgE5Rl0/GNGJ
ZmSH2PUuab81tHChU/V/BHYRO4AV49oHaSNjWPCMUmsk+aENY2V0W2nvIHgWMRha
bCAuQeYd8T0+7nHwE6mL/k1fBDseJ7uqP0WaNZxOObEdTfZVF3Vod1Ni3XnNteFK
UvMHWZ8LiyXNkinFnPoHLbcAWtLm4oK0ygk7TWlAJrcaZdTf7mTZNU32524b0POs
FRguZLlO0/SIkblrGwaMOp9L+qNj21gtPD7BfnAQOZI9lcf7Wx3ZpPpslPal518n
skjn22kHkUPATj18rtVtxNjLQ7luhbQiguBwfVDswh7VXv94SD8ewXQdVXDcUGcV
N9848F475MhWhvwxHiWW8Z9D/yKKiujK8ueJkwFrb+b7TQUrgaMi3bugYxzM2Hvd
Vpr5YHPTp3e14hLVq6r0Nvn0s16R+izM7md0VF7iUrqNjetNSwyIAOireBUQuyAF
NPf14CL4ZAONWLlMh++COuphU+yxapYvD7JbQltiruio7jKmycyYi/Q2kn4/TKc0
Bb189XP8yKWVmoFh1TMGEWFWPWIigigRBVZfsm+sm3WDOQO+zPCQ7C+WozYo5oL3
ZP+CAf0fWAJMlvhqNHUAisPCHEGzLTOs0Zhz4EQGCgWhQEOITMtsGVJdGO+pPcoU
D8Skmpa4uZ7YU+3YsDZ3fPQ99cDWNAMlJkZfIjsMRypCg8XX4mSb+RxqXq1FADAA
BvwofNSq2xZ/Rlf3TkK9NnOQoYQtKgoLPzgilTo4jVw4Uu+PmR3LCaowNYwyAASB
zgHxOpsiKE19YynNikeU9bsIBIxy+sah83N5fqtB90+2hgoYEE1udbBDlWmEXapF
HEWlvemGb7YPrYR4HPlqrn0heLGqe//XPwhtXxX4CVdTJ1h0cWkM5oXf+5E1XHr/
O5P8Z4cAmYN/uWcLwSKKxyGzaikYSj/lv2Gw5LQyR458FQlnyE5r3OwicgvIH/+0
93J1idbzyPZhNKdIjT4lrLrq/qTD4591tyhmCcgJIovAYFzn3d9mDHc4xmqED8RE
Be1ETR4C52NUyiK7PRDJ3zh9pXYR5S9APJV4OEdmqkH2CBgZDc2dg7ImsYOBcNZu
iS5I7LHRPYSZLa3kUZYNUOXv1FjA+YLUOXLoOFR46Lj03kwh+V82lsJZCdK7T/1+
lAxr/CQggwPooEmMiqz4eOWAfbZ3nq+QH2m07os53gDqBsx8mgVeLar2bh50IQUT
4WjefYnr86Jweg1OCyFSFvNynMwhHNvRa22QJsKMdrpT5cd8ULRRaPyqKVe/TK9z
EgsPU5fpUGlYAKkfTbbNR96K+mPmhmdrdjXXMChBnS7g4muZ/XFN6BxxY4KJWb2e
uzTU1ikVDtLAd/m/X9lwAnnyzSEweBO2rINCCRdenrjQlNtRJPZkfwZ0gHrM8N8W
EuS4SjISYMYpqE7BMkB1uabzT6Hf+6yAVlt7CLC6XgCCr5NSYqIsdpukVklcGCHo
K6ZasOjvh53tbYZuhKMk4a8yOHI+SP2zpZwx/tlDM+1MMYKjFNgVmmlkAdYZidVR
+jeIWMGXoKF66NrIUiVWs7DJMZK5i4kzDwQfWaNSnyiCwXZ/pYv1x54XVnA3G+xI
XsaP1DjQAmtoe6Yzrrwl2TqJrvrdXA/1nlp91MrKdqG9L4prLn/N1vGHi9n0SEFp
hFkKcwE0NOo8ZUJiWsNeqvF5h/i/eBNtxV+3LlDKxHCBFL+XTfkBeseFwrRyUpi/
DjoUtJIN00ddEmBJRvDaXMuF/+Pa9GWprtA2DHmdEku8hlJ5Hk3SAaaU0KFDAbbC
M5bSnwjNYok0bGWXQUPowlPxHtgRwRfEbAeQgfi2FntU7Vet/wqu/arJiMgqo9DY
ONETyrhwvjCibojOU977M1A0PoqX6q+k9zUrV9NRlrKckfuJwGlI1TFM1mh2agtI
Y0mBf/VXWpY/JJXBBnKbgbm5pZ0+KlxgqL89CFHQTgEEEt4cinShL7XjMCb9kxOX
Di8i0YBqbch7jgnBPGlxkLJ8lJsjMDf4ys3ZvPkyHrJVDgN+QVfDC1dkdWeVAeb8
bEt1zRSb/McY9RGn9DyDEc/EjMBrg21dUq/932dd8uLsGkn8tOanRV8Z3T9kvsZ2
ZbjaWvztgnYHucCyuqikX3WM3RuS9Uc/K9tFjm1olt7C8WpNgTiF0vyRsMFI+dXo
JhiDJLf2kaRyBOI7t3QQbHToFHTznJJzNWB60pKxEqAIebhE1GS+ZQNgazcq/+DP
hzrdp++0anvioilZr4de4VFi8tvkVnvwXuVITiP1FTe9VBjdT/NnXKb8SH2MRDws
r81mHBZcXxjaP/tCfAYAQvX4uEhcTwqh7jsbmrY/iyWWfgRp9fqyx8tCwAZkC8B2
Jjl9/YMkxQ84KntWcIrlqg0Vnk9KGXkbANUwDjU8eYdT7cGMhDUfrigpBAKNyEo2
uf/tnPSHv6Il1DXBQkb7rICe7gKuS4lT52QO12h8dfPgoHYr/vm162ZbO4vUzFXx
IybrkftSS8Vt4BnuDk8RBlkk5tcslvw3m1/edYfXvu313MJ5mjgZ5oD+LJypCFFq
kaylwm4V2zedDx6nYOy+Q7teGqQJprH0cmsexBo4N697T2RBCfqnRvRkSpScrtff
slIf03jUrJyFmbrT72UNcbM87P9/EvIpTXw/X+fBxrR80UJUgWKXDHJNavO5sa1s
VUpTDXydDwJ2EhecET8uAZ7Qd+LZfnNs2qqWqf6zYuVT75OZGW0eE9rKMolridcU
LOXpGAEuTpJbbnltUR1UM16urjz7FQTx/kp9k6gb4siB7tydkZiWqfXPJCtbZRWz
bwrRhA8NZpQnB58hRwv4ikeRUmDy4sEC1aoZpwCOKTO3FIunV7zjj9ousgegrTRg
vB6Jo+Sy7VYAgItSFD5Ykkecq9iZYKrg7TxyP1lfDY83RSWNj8/UXvTmBGKXYL5S
EP6Pgl1UF/e3qkbGkHymK3n2eCMkirEqEWHUOMefu2rRVvPuMK43fyxRbH4nbdRl
LNgCp5ZrE2WFc2XaEOOhM5fTXNVhK3knZ11p2fIJ5b/vfL2xIOotIJOAq9a2K+f6
NoYLdFnoAGMUPvzj8VeuHD7kMXcHZVlvKWmq7mgQaFlEff2boC4UE5fusfYQw3L6
6so6HQwWy+5wCWnuKr8GP4sf+jOgFRKgLCN5OsHjnr353VF04tnnlP1lKUI4Knxn
uCuBQBmwLmivgI15mu0NRBPnjRc0ZUqbyFIGB0XzdhvDbFvvHXTpQhqQ3iGJWU/l
YCw5mdTqFhAnzBD1j4dhJP/TvPerFcuZaI+Y6UbJ53wZ9Op4sChQJqTMoFbHjnEy
Ul5wT5K9BaciKeIntBlJAHodjK/9Cf/l8aOH3aYSxAegCjsajTWTMkzNoc83vKmQ
DD+CP2UJSl1GH7uKy+oEjYsr66LoXVDyJzysgkkSRT6DDF1MppeuL5bDAkHpK/IG
tozYUSvBkYEkR+NaMLY1HS2huY65C1LFuKnYWRrHne3O+8kX8//3KzWqdFB9NO3y
a+s3ZUUhV2/TjF3o1pyMv4EaICPVwg+ODFqflB+QM15caSoN6aR/v0NF7ZXWZvp/
1wpYynD6OkRX+bSnk3ElLUEN6inE+IkdPKeK+Iu7fDdtGe8GFXMFy4PU3celTfxE
7LE0Suq7ixSjJAIqeenO+lJTGe6t0Q+GOEjw1Le0MFGVgm9My7oZzezD6DTQGdRS
b7+1eRX/VyfD4VtVO6ZCuB+wc3AUfRjBi7aYtML/5MRkSyCWqaS2LUQWOrn4XWz5
aC7CFOYzBW3Eh5VJmo/CpeXhC93a3TJmNe/rcU4XIEa/Y3G1n2G8iul/5HxBUCpK
hOc9M+NGJYtIKC0SPIov0rDmlBnww1WX4NiTQNP+W+EtHJUj57KdDK+/9lA0nwb4
08v3HVx1aVkJKSwAwjttiiVYYp4LFQqmkMlqBRSBqffDWRIR3qxd4rT3yrJs38Rh
qAIvcBew3BEcs8PQm7ECWK3WbHlvc5xFvtJ7NcDO7OmaWRl7E9dsRZhR/4LMkaQl
DrKjKERAImcy/EJUrRaqKxRDCw4FecPfuRWyfQ8EUTlQZDm4MIDDFj97vuDaWrpt
XzOTqb9yvNKR51RLFttc56cCXyOgkUJioVmEXNhHzc1kjKsBuef/LgE6Ui73HVEk
FOHAxf85hI/aD6Rx7qrwnMffb6t8c49wEEPXBDuOfQPsemKzyASlNuczYgEfTw13
jSirdaoeCzIudMJYHqAAWfCAiutNHc1XiqKtMQ1btArwWbtT4QbZidf4QMvOj535
ifI69ndccgtAEXo53FLO648i7cI69+Cem6+7HDL1mBEKH/bkHjOZaN7ImKg5Xh0v
1dg8kIXrqXV7XDoPj95mBpAmYd2jjN1iWHJQqnA8Iql/PHFIMjwimGUidj/2JYmB
b9+keDiO3BEMerip/oJh4UNjUBD8BRHO44prEXYt1lhhkxrzYDvpjVv1yNSoX0y9
byLru6PlXLACCiUnF35XWyPJWnc4fkmo+3lfYl31cFNrot6SNDDXw4XM0aW1+Hgi
+spPQP/jdzuQTi06u/mFIg==
`pragma protect end_protected
