// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vbGGRBLBg3+qyzpD3S+mDLsLmL4CGsj0X++/HTXSElMpexNed8tiCR5MOioRICyRoMcl6LMyIoMC
u69setU1aGhnb8V1gTm5JgGVLfeiNjuNIRTBf+sJzDnSBCPLTPs7HcXkvJp7ntvEKl/2T8SSkQ4d
fgxfq9aw6oHNRBzgA3d24TppP0NmIHjGH5Ah3FgNs7PmA+7uQ400izXUsyrHz/N8/4Z0F95lyxkz
7j9JWiA64C38BzdNB6wGBxuvp7/ZtD8E2a3xA37FXdb+EjTawX6ROx1KM4UnUMKJwP4nQIYADXjR
4OOhfk5mEOMrWUCnTOJMCWpD2fxKhbp7IlHAoA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 27136)
GGzfdx2BQQq7qiQC78HdZVRX5NI8BFZzbvAIO50ODgoQUti1vQVRHh4fwlX+hd6Q/KANRd02qpgl
S7w6IXPsPhT3VWskQJ6TTagHXxa7nG/KAmiUyc0xbGgCRHh5///usVgsYFYksM68O+Az+OCl9N7g
h81gdbHAyZu9TN+h1bh0r4FGhwchYdlE+sR9Svd8S38W9moJXNDTZ6vvuI3zrpT6xLkcfgqsvhWY
PxwXKyyVUxV9cj1g87iUjLq2kRi/EBSJi4TJhbwK3zY9JfD2YW6VvtO9WrK6izQuvR7eNGFaHaEO
76y3sdDDnjJ07pDrQseQeRx1ydJMzucVrTpe+VZiKXoxvaqz6BYLtIP1YthgK5y8uH97v6qtl6R/
LbMd90MKasikSBsDgpqNNiH5mFtT2J8b2Y2gRj1bq1DUaOloPAQz5pb+3O5TEr20UjOsm/KZFFyL
qf5Rn+W6mE21fzM/4kq3TkcqtOlCKOvwS9PAQjyBwV+3TDvDNYGB8XkW5BGCKP0JgMbMjzn8IGUL
735XigZ2xSRiPTllUXed/SwPBA0JreRJSfq36lLd5qtCAPQURgG/xZT3chaYmwvWUYpni6Chj/7R
a+iPbc32+EPPGge1+YPMR/KUU6tAbupjlwB8F79S4hDjq/NzfcrPromUPoD9zrLaHWOoASCjbfdA
YsY13/s0dbgN4P8QLk/bzikULOV7MDaQliZYB2TYC9AMbpH2cQgQ/auIQdZGDgZOsOOs3iKot1yG
1dodDGC2RkqSTOS/q4gYILig2nv9qYqnkxO/vMoQWZtp5IxM9cdJCbuX9uIiFn82aod1kFLS8NfJ
W4jAMUvqfEzxc27LrYNRRBxvGtPifJBwiTVU6idPEcqUmuJmakNFwrk3XdSMqs5+/FCJk0rzEwAf
oRFwBEERUlSnJcj1+Uo5kJb1O5PVSuh82fKNhCNvQnN5z0Jyk4rfXAK4ZZd6U43I6VChXJD0e83T
JGfC+/jSUVGDj6K6wOJTqomB+T+e1pkIVAXPu/I4FpgYbrlKvqRNoa0Mt4/8nfzQE0L8TwjISHo1
ddU58ojEXCtg91HHDB4r/KfDtimN577dZnHkNybbugyaLBqyQMchawAbk6l4RV7QL9FvrP6gE1+W
vRIfbKJr6X14dgypgMHuiwXjFwTlzPoC25JpGuTBF7KfBIRHHVRHQ/AlQndwj9WnqVqNxBNW0wPk
LCiVJ9JzemcQDaIgtfS4diDbAlzb4hd9Gi47cKtE6v9O0C/d00RUp6hXBBm0XQ/dCsv1oonJKb8u
8h28xsWyrnda0DaxLKaRVNFQrjtT0dUARSPW0Jwc4ss5Fy9I6AKqLoeNs6oqutbxUe/yvmfDuC0B
3DGYJQaQPBXGBb/i4zbU/+OUkHT2eqdR4hR58gMLxtyfSTPgjc2MV2corsfx+/RkCrOTov/6IZh9
Uxrdli63SfiVjZUyy5ggqpgAEz79mRYQqHQJuIf9N4zA/FLKKJPC3TRUC03zNMmMw6iJ7uoZCLf4
IgaJoYjQhgAzHnrAUTop2+Bx2Q1NFxjIyVYjoIEjRR/AwRXGKBxaMRrrHqLHAgWSJAGZWQERX3FQ
ub9B5mCsotO0+p0QP+bmwX5jbwTkIx/42yl+U9hd8eRot/zeJ/l+/nGnXt7IEkI02FdnoREUmufE
0BJGckfl0oiCQJPyX89wRPXwJ7AD+J5i7cHW4fjjbK8vi1022r/wJ9Ds5AfudMMM/M/fA9dqe3Cu
zy/Gz2Q+l6CAGQGuKhVI3JiO0nOsM/gVf1+UNAh7PldTzDSLkr3Da0rMaxiVO4w0sIi/7Ry2Yte/
UbmMiepuUwgOC+OCzIcxHpBWZXkBgz4a5AY9F+EDTJw4AMumb+FdtWepwaVbU8HH467vDMVnJwql
CuRZYLzunOpnrXB05XnIxVyYq+Bxir1mP2i4YAyLmBJe/dYC5nEZa8+xTNrADDM8zm+6/QT/yWY0
9xuU2ys6fOdIk/j6A3h+ZD5i1lBxj1FVtbvoe0Xg/4ZC3cVEV7dXOKptvUmq+o0sqW0RYwnRdS4q
1aptkOlHXeJOxNFGZBAuE36AwTQ48a7ASLaRxlQjuHIH2CJsjVVJ6QmTavzkRAPynXNae50OOr27
Qdqe2CBIM4igaUJ+L97Al5/Me+qVWSdJ5k+VY1NQ5WbPaKOOLSaXwakcw4ilP3MlX4qeINAdOqFL
4i7c6GAjUFQ2jmoxUzKAeZfGBXSknyhDfXiK0x/BdkJkaX+As8yIKt0co5/DMXxCOUi+yRXVO3Sb
g4a/Dum1/GnPaaB6+tpEiBqkMZCJ5qNqL4xykYDYFoFZ6r/kgVmlHe/GjFJoqiMejERpxpbQW9ON
W+EhifTDjMDaYAg0x0RiHTxON6bqX4JKvVEy8Yjpim7NRJ7Jjz+rywPTTnYDf1m5xALzpN+waTHx
N1IznWKnXXjd4D+QaWr3omjvgE6xrxNJ2ChxqfIerNHn09zIWpv+ShnrYhsVECIcrvfM4TmCRCu6
cqAZhfMD8sm5nVKPF3fIySn7zOQxQ/1L5/QPdhlia9RBWvdg04tk8g2YmV9MpHQRQUoOJQCNXKsj
m0HvllGhhHR5rFXbuA1hCWYM6Ff6pda2GsH5yLFcFs/sZiVgdzcyOTc3p2dPcf1Cgmy1XkCsCj2Y
CO3WYvFeuprWzbZrLfHYKDNGPyPRo7WMdYK2RsrmTZe09cj9N1Mu1+zm4pBE5E7mbWbxxD456BVm
2cK4ezzujefcYZegberFowGU6Gg1SUXXGrpdywx6veH+wanCYD3KP1sBla4c1HR2G+75BsgQrTCP
f4VLxNUuerQFT4uVr+Ot1ojxHuczBrROQwd365+3rwBqRu4WA/TABgRzNmo/Jld511qcWBC8yVGz
DkJg8h0UINCSYY2aDLom0E2in659A6iiGc+JlFXlU1oGcvvKel4OcNbeAodiTbgc1VftG5VcAqAn
Qnvu5CptJ+q44trkXq35pxQrQClxY+8l+i21JKMPnXkV4oh5iLlNksnvj/agwuUQjCJniGCWSgp5
Xi0QTg5SvMXLPx+ehbb/IJIH2udn10/hAwA6pp7B+P0ZfO5+7PHdfwnhFh5nTU3H4LSxCuX7/UBf
eYT5zNEvlS8SHb2n70cV2gkakSS4Hf+XwryI3kG7pHzcX5j0fn36LRgMAE3AeFkWS+MUwpeEak9R
h9Q4p+x0qSPc4WND7JC/SolEad4fevZ4QDI5CSQ05kPz0t9s4Fwq78jycl2vOXuSsQ0+ExVHjCKa
ChdgQbj4vAGx/HfR0jfkFEA9nN8V0HlvIqZZxNhRMCe5A71SudtXAxb/oznPlLzt9PswWMZk++oy
bKihy4nF8Eyzx0hy0YVzHxZQStulFsw2SHgBfrBHlRH33PesMZYUV3tj3pTsWxxy6Mket0A+N2Lz
gvnUL2Wlzhce9x8h00jDkJ09rZ4dtStGgJRP0DClSPJ2ECdcV6JTEPO+54xruaXWk00zOj8qO74o
4Qzx7RcNAxzZQYQhq6uJORoq07NubIXAWH12lAcvTcVuDhGrvLeeAzMpsRm66Fvz9Cq4aI67AK0y
oi4z0MoJJRg9Hr2mR7u1JqI+PD05VjiwG6U32zKHZSaDftqqW/ZMqR/BxI4y5gJifIFZ0C2gXJFJ
ozz79D7RZzZ56HxX/qpnQlLLZIBLCFf71ousXNv1DJBuTW0a8xOMMLWDDVjH+sijsjYH3+x5h/Mq
RYdI91IJLSs30AK4l47c1wMhfAi7aKa2fkD650jMuVWVnm20PWpHQYek82NNppS9j0tvRZc4A9kp
kuA8i4shhtkb/19deaHgOeKUE/0oOSCmtIPk0zU4ZDNljiBV/wuCdepa0EWF5IwGo3rBeOMDg0RR
d0aL9+gsVOBP0wdTk6+G2LXnTYHNd2yQFMfNiSdDbL4ZG+QG9omYT1+xLLBX5qgC9Wu226bD1HlR
LSZKDuKU8dEjMTol4usEPNocI8Iemgsvvj/fVcIOZuMOTH+PRSTpENW051Op6TelWOPTkQmj9N9d
SySTIS00B7E6ox0Mep+RrNvzIG+HfDuc2rl+YhfipxsoNNLFIMTMR128nNbhZzTQFs1bYvvuJ0x6
GPw/P2XlZJx0tEYnEAQaQ6K4M6RDqtQ6PZRyc+oS6RQNjxHRiVAh5u34nnPTdLW2v00WWV/5VoTV
Jg5EHDjnk+ldAPaSVG+gIvLzo4F6poidnwjuuTDCuXkN9XmsuNzGtFJwqPOdoUnibv+UKZVBthCc
s7XUieW3bI+JbjVCsBQA0i8AWkGAQizVRqmx/Mo3dPraGRR/MtEgzC46beRpenYPQD7XFtfgsqT6
bzrhOwvnbqSGBwVo0DHxL8lvv9TetVyvJfjutpY6T6SPCBaN9p4RLhCSYO0h6tSo8JsZ1ykB9Gbh
5UKWqdr4ylP2oHa9APFYP8piDgZUA2diFhsgjpGIDU+p+JdkxpNDGFoXMeqHcmWiZ3U+/KHp0VOH
ZslY8Eh1aTFsOIFBvxEWrDnVy5cKnWQmt0t90X5RrPFVSdPUF/z4p/eY/6C4nMZZQEi2431p3AAm
kuO6AAdLxWyXAz55yxM4vekW1hqtivmIZa0j6PnUiK2olgMBM5EzwW/f2P0Ow7/aDPO3/EmwjSO6
9D2+uAdA7xQnppt4pYBJnnE2zFGQ1JRS32qniictsFXug4+ex2axV4RIyXPWn523x1Ra5Ox0xjuE
tNMOAyBJhyYEWfkWiaiXNdtKJOybQFl84xOKDFKSKZXTGHoHvSrhrgEPbUIbQPMdbrvPhvONWrg2
0KR5W3a5y6vC5YQcQUbVwsW7GVyq9LRvn7CjdJcIxJkKTz5e8gkYCNzfUwNjQXkD0oE8UWbhJMLU
8eSfQ9a6a4DEwogBwfbLA2gFno70eFx56B2Tm7GOybAFZf4ANh11qCw/XZaZds0NbT/exlGpBhl0
sr/QKfDzalYnXu1AalNjxmnPUA9q9xpkhloqsL9neZL7ZV74BqVSWxHJjvwObmWa27qYTHESa5vP
rcScdra/kJEfYA+Kn19rF+EaNoxpaaMEOwLLup4CAeejrOhf7MaN6PSQiuyunGp49sbqhxExVzCM
H/3h75iaOcUFvVnQ2TXwHzxhLSN+/yiwf9P85F4oov79e2XAaWpDZagqhqaHaNliLMKyZgQqn+oN
8UQdIzU9pmoWlTn06ROfwdu/WjCF8EYAfUcJuGgfy3xtGzrvislMih9JjqX2Kql9p7dvlxxH3Mdn
ctxBQw+098hVJe9MEcoQ8W4TLf5qNSDUMFR/FxD1wXFIC6xs1kWx6lPHK9A99zPtGTs11/hbxkV1
QGhMdVkQ2HeVfBGTttCHBympC1WN+fZgTu2QrYUFjdsf1AGOWD6ELXBMaJCmySRXbOB4P+avaZf6
fET6cVtNCJ7yc4LErjjJEaImW9qADGJqXaPDeaToOXB6qrqJZhSiWEAGMZJBB1v+vsmzixNDnSPl
fTLJDL3h6ekD66Ceg5E58hcTZY4DTIWlNCePp7o9i5EJoBWEqTu59KkcIe1z8+7DWM3jIOJhdoY0
6ixxSrnwwKr96UZhLpAMpH/BPce8xejlDSYMGUbpl58shk8ZIpGLENpmR7f/icNhIdQE00Q6vQlJ
CLI0wkud7CJjqSSaVW7kLDw7dxL0kc75FU+e6nmB7FwsKIVSdJkxpYk4KHPhY1goT7y/ZW34T/eb
8lxE2jSpms9ZEhjv/WZDKOzFAeWlSiAsGN08ye3B1WE5SwBOV2z6Odc2wtp8ShTYx88DWrjZWfma
bpdAGlhRlW6siMsl4y41pVpSinI00f0MphLjZd4MowIcJgDrwpINN0S9JHFTxB9H35Clvsml5nyb
wBmpYsLRf17GPmY8uNR/OgpjwFh2rubpIhznj1uSWnQK90Dj50naD4vmML2ZL9+6v65gOYEhpRDw
tIA9lmY9P/jkmDxyNtOFWkLOjen0QpqmVJtdIPA6SclUL00tsYA+k2pLYcp0trTrNaQpVLjJ0iz7
EeFV7w4977WtyBpJMfgwE4Xo33RbpyKe01cxGczPAhgMKfkSQyyUUIU4p+KM1+ZWVaGbAsWkxKAm
w+FCcJ6ccAOcfTk4pXXYet7UUVOsLtIxOUtgKmHjDWVHh2Wvornt9gvGxF0WtyDycPUdK8SFORVK
UPPYUgmokY56IU71l20zEmok2vvWYZoH1jLx/yEJoi1HkApQ0j1W7d9phOPeOBMjUjcX0GKc0Xuf
4+tgUJEski7cQaYJfmCgW8zdoD1V6HJ0AI3AFv18iGSeEndJ3IXrqGIdEkptaJN+z84MIv2CKY/+
6LYJEgR6VfeHUVLW3x345ICi9JGDHoea59iHGf/Ub9mYJmMRXnuPx7AIusSgfvCDmtNxa/ahSRQu
LXq0W7sg2Cl/UKPrsanUT9tHPEhJxiG/ZaYC/un1BJk1X89pOZgw7w1tPxSh2F8JKAnsNaB20EyJ
kDsvIvhakLxZjY4nyLCqCuFGLZcJCCarf5126I7IqQdDwQ1Ybg48kHAxugQTJOl/YN6Qdzh4VA+r
07YSYuWEO4Ot9YR/7SiAsdJk2JOFMef+dc55qqsiW7IrJJz+ytkONYPhXAJNjWwFhMkoprHpVqbf
iPX+vw8YqQwS9CkiuAVEcTB5tXwPlR+gvEV5v8DYlgxHzEa6TsXMEknaxBKgMNbDpVPFJ8NRnU4W
JHYMog8jsdLVWVBCnCdSCo+nZwD2ToC/R1L5UNnf624aeLPE394eR9NjXhQfcG+vbT+0qg58jyqA
BeVJdPSEARU2YWC8EjG5x1L+UIKGtWDrXUZD4wQFlsWtC/Si2ZWx05bqibjeWRHR/3ytgrd3Q3P0
cNlLYcq0YF5RrAthEtNxF5Dsnws4X1Vl7FziyPJbMjAQbtNtkUTsVqIL+ADqiku314hx8PeBFCfz
NN56yo4ibVqqEP+pt52DSZC4r9aoE0Z6htScFRdjN2IaLgKzkbmuQBqFPIQL6e511O7HhsiNEAtF
eU427Ra0yHARp9qM/MyNp1aECfo63wl7cADF+oPobfGwKF/4LqNZpmZbhE5JLrmjNuKxonwf50Wj
lCzp3Yqo+9I3RlDBfMgtqD6Q0UkZxkv5VeGjHDa2J5f8uxe7y3Gc6g7drrqn8kZ8KclvukD3yfBg
xv3QGOI33xEZ1uMahC7CQ5gqCfRdD+cPuQbyvcw2E0PHUwqHDhROLKo717yi4vuVL6VupzeBumuv
qyc5tngz+3NU1rrBeHTArxNjIt2JfIuZ3nw7gfCNBzQBNb8SfXWA9plMmaQbRaQfP/guLmQoJ2dw
rVTCyp7G1e22cLdVZoUWqwk0ZhPjgTEv8iwH7u5U1uUFA/UTp+LlXRwacU+2XRFTYyGhiznmsj73
AzhgAmEBtu+r5UIRm8GUgYEqBqbvP/ZJOe136w+TWNt9/mdfhi4cTHq/8nLXWTw23DDif73eU+g5
EgHkSXCbHfzaxL2ScifMtvMG6dJzTDVGGL3l0ICWFVcuAmU762DrDnviZJLibZlYJcgdQODBpdnc
yLZ7a/MfaI613g+7njEnPrxCTAKIegwcL59Wv1guFx1UO526Mp6aDT6bOFQzsbCYP0SCabdnsSAn
KWoVHep/HvBZPibiV1VAthtEeSqd7T8WFfAL02xZDomYqL9jahTPvBYR568yYa//UBNcikz2kDxu
LjQF09cSFklKuP2g1tpzXBjfzaUvV2MFkhxkEf9inDqqGgDlA5mFLQgkF6HQdz9sD5z4ZPU9Jk7E
0Hc63QWtIacarfenxzh/r63zZOixmYF1nAHTtKdVRR7hfCfRYNLw+s1NglCTXMbc5a0d6OIe3AdK
o+NYbYeBMKxHsUFL51S5fUh7vIIpp/2jQykQeaPt42js44k14hHwK5SAN5znxMITWFoL7qDCKuiM
rJsnDT5QmIBzqKvV+krQbShTsE3et8GC0KSiHs/2mQfprJwveq9fXUzOOG6YVeGmmRI3J69A9y22
2KaLOSsvuY/yrts2cjm+SEwmDfEmAoIZE034soiERGmmhBhTJ4C1Kx4nUk9M+D6YOmYxKghVLu5d
Z492sk1yLd6c6L8evRgM31tDvf2FmiUQGZOBA/eaqLVT77FVNJB2NjtKFO+dtKqKYHpdsLz9C4jI
0Czxq9sfklN9rsw27NF+9YOLG91TUSQtxDTlzhu62RGjVfPVXHz+tVjvDpVBCPOAl1U7+UUEDbs7
Oje0rnyp607FEWJ1+imZyyZq+OJ/irrNJaBIjFm8srfanbspKRqdPMl8xrAiU3l/PtWjh86MxdRp
6/gopU1wHoJkqfljjknXhRD/lq4neZUxTuNDjqJz793YxqSi0UmauPiT53SgpYjaSnQxDwJlcwc2
mHW+xd3YIwG2JWm1et926OPsaVp4ta/KHaGFNpRKV5rXTgy+YgWv3Pk9v+ozDCgUPE859tNYG8gQ
IySfPzUDlUe3bVRCSZYHiaPUsisJalHoNcQDgjS1/AupECCIsUNn69LVWj7OVRuTslAVe0m7rNia
nTwGX8zNfM1sirEssXE2LRs5RGjB2LX+/54oh3YBkRMrh60VcD+QL+5SPdmGmJgL935Ri+TGCN5y
Hs7cZBwV31chluMvg6gTQQAO4afrID2C/ULLvwjI/lqcOfz9Ezk9yHhQ3xi7ZauwMrJpM16j1Umz
s3irPMQ6mqTehzaJEG8gjJoarXaHjB4NSEmf6tjyRm7G+fjfwZ0FMPMGWuCzCadqAwovKMXSiHtb
JeIQgCw+sZYPEZj9I5xcKV3F157U4BlGHZH+k7ww8qlWSyiLvcBxj0ABfFkVCgOZ/oe+cYsd7x9s
pClZGOOrEM7Eww2LUjdK6C488wnbWnSdPOp3dsZD4FnQwlbaSXrpYD7obo7kILh/xkUFidpInHLC
J4E0KwgWAAFVTieYssWEq7YYGpA+60lmtU3dYtBT1Ltc1y8y5/hXG5eAoIO1ZCTcBx2+ll5ClnLn
NCnFT3KpAOEGI1qAhuGo08NCFJeK5DaodPVbQu+dmdsM9pBTiE0L7TDTX8QvJ96EPEEz/wZBv/g5
G8zFGntavawD8ScVUnkefn+bsAZ4Z9HWO1of5nZFih+chvNRwpAzO/hkugm7ad22kfXNubBqV+Hb
87a2cIu3oIDNl2u06ucULrcnMkO/7XDcMj+qqJT/bK7hWXiXvfOEuDwsXXHDHVR7AAkeqqxxN3cD
UduV34JCz69RyaFac8BcSHNtQlK4nr4ZiBdkzN7USYIxrAnH/l4sgnPR2QmQAJk2cix09KhSAFtv
IgOhS/zFQGOfpA+o7jkgEkzf+bHfyKs2atM49CrtsM0HMy1yQmevXukSe/KsQ7RwZEKZ4iFf+mCH
/xMEe2RiJWXuBtgFEgGEwoMrraIJHczrkWSBgX7bmrzlKHKKtLZC/kgoohA29of6zljetD3TrOcn
yOWmZc/8VQqI8bUYh2xnSxMtCO+3yEYrTyfscHqpxyR4nbPOp2NbbiNoKHOz0CYAnUnVqVC9ZdBG
5wHR/R57XSdDYOujs822oIwUWBDxadNpsaGs99mjR4MS0rAMFSSjF+entK4/z1P8NynSEn2Bof4U
9g3Hs6aXwA5xAa8L9B15M795X5RLvOmdpqT7AG5a4fOsUtEg/2MCKBcRKCGM08S5mAosAnpXh3SQ
iT32Eaxhb8DKH6DsaODUKUQXfjNqDVFkuHWNhfFN42wxsrRmMWsRRKs2wsWwFrqI+AzHjMFBgsdi
ypcs1fTRI9WGv2m0j4OhH+M3+u30vGvSVCbySf/UaiWNsptVtbfxRCaXrInBdLhvv4SlpJdaW97r
KGvuNuGDFDPAjbEvKsZvq4/98rq42iuRxZQEVYylwk8KakLt3AMv5GQg3gC32T4YqNCH3gYo/oeb
mpMZ/VkDEjnkZN6ue77TWsIHjmQ695nP9J87UrsSyXyF5dWucGlABySjSGqukiJ0ndByby6ZDX/j
Ghj/QuJhU9jZStTic7eXoNAk4FrUEzdfwN/gp5xdfA7ni1tfsCPUme8kugXNXc81jF8c+v1kcs0s
SGXJkveLOcHvIRe1byJpvA9cXQdY6+DpyfC32ob0csl/RH6a6Dju/j/qqBafxMJYVTlwDRpR9aK4
loSJcAZPpvOFns0I6zLnFq/GyYDz6UxhJgcq6fI9ksVjBlDLs655CI4MPvMroWfHLDL+peKroprw
n3ZMCIPM1ZSG4BH1fVHxU7sGY0yNHRpH+TZ1n/5DsDQBnSwWdn+HFdaVM1Tq7dJCeyw9fMwasTrv
5jXajU6ecCXVrmvtIwlroGTgQrXl8AIETbsjCHPX5nYvORZ3quVb29trogAKGc8cIoUA43A1CLOr
81AFxe0gJvQ8YgPP4AnNYKPcmsfA5bpzf2EAfDHjVqIKIMQX9a2ur/csXwx5t0+tJC9e0muVAhP0
aMuZZgNE/C6IxXHDFvVN5PvO34BmkhrjnMwq+AFUAHMdgI1+37xQvPGPxDrWbsLwX6WqfQZ1hx1a
GaYzJTW0ATEL5HdkpKrMpXl4MMSjSI37dCVV+mzQ8IaXvtW9XAsO/4ztioVESZ8R39uefoj8Gfaq
K3ijoqEtnh2HVGYZWqwsfOTf41lTnUTtRdsk1HpU+/EG9Qw6FaXOkvvG5ZTlwav2cTGlMd5bC96Y
vB7SLv9CVQJ2dXONk4YhvOwotkmv0ynIDc4OUQ+n3dflOWJsauDmdeIEiQKqWEw6tMdNTbeDSzXj
y29UjNPbxxQ/gEFxusI8Fl9edYt5qkqoGTUnfG119UEQDdgxjmpP62geEG8YhX/GCUZSkWi5cWhV
FdCOTfkExrZaZsZaBTpCtVU77VwUmqosKB37C9YVPdrh0jh3YRCSe/AxN/rR0GjZHT/eESRdQUo+
N88q3vdlWMOAIhpV0XSzuSMDlhj9k3wN1hKxuxsd9uteZYIq+bcEzVhMloSeIcljvxeP2VTVMwyh
QLgwyLdqVMHx7i0ML3lCLmAmW5/bu290SkROlDW/yNJJbL8yKuZ+P/kdYT3G4oo0IAh/nyaZu8o0
Fdk0Cl9i2sgwOAW0cn8xIoBfbYy4hael6/njteSEBt0y24+XfnL527PDjWiAC/GsHzQyFvRADon6
WgPoaBiQrX0bQOaJkIYMArIVA2IQg2WwxPvC/o2M7/jiJwhOlvMFV0ZsTBa78hkKjYz34zxMaA+X
zsipReRiLBnvUh44YiDfciH/pom1itlX8JuN/f6PsPAShb6le57DCrl/pOSopphsUWeWihElYn4O
wKlyz+9nZIQbd0g1HQ9w5vIWcPtOvpyjZ3jNm4Z2Cn45QHY5vc5IGQ8MFsrWrlrkwMii6PPfzhGW
TM4BGSsjqI7yHL7FaeZCIk9a/atftK3o9TIgwAudr/tgLEQOsbpVWIGIkn2sNojLSN3X0Pa3qY6D
KkD5KXWNBMAH1owh/fMHH0ybe/sby97tkwFGvkMYL6TGIz5XAT1QH3bJpQkpa9bpGqaCMXkAy9pF
92aEpGo56KkdQkA0hlCdHyHU/ZI+5/5jSi5o1vJXEEXnQu033TIEKX40+QQeKzFddomyyaO2sERN
gMCuEyD6ocu9dUzwzrZgJLv/qk78i2wUu3kJd1f8fYM42B9a6RFAxFHa2iJsPsnTVJHhQnl743G8
QT61rNUGwnHax1CJB9jmNVsacryaCZW0O7h4dv/TBLZPArs/NZqEe1sMt64AjjATBYQSqy2ybobJ
oUIFkRp9DNbfa9JQRNETPdhMPeEZLbIhz6DtRGtD0gN58aTrUgdlhaNjoHd+0WqxyXpYPpFEjs1l
InZz1hS0PcUO0SdZS94hrPpbERbKYeIe3Ksb18Jl3/+jE7BCwKhqCfumByHPZx2vbChuD/MHXqUH
AayJk7CYyWc3lXP7PXe6nVnUzosFg4i6H2y78SXhiQkzvWcEzrDZXob8P6YUPBm2HQGrzTJHdn4k
BFIeP8UcYASmAFw6Nn1GCrhjPDSOaAEfN6ICbV9pInTDx5mNKl4t6t+jRPIDhevxO7onAyFTHJZe
nt4Bt+vQoVrDUK2YG4FS1etj9ur29gteZqZiJgJmjNKINoPOBnmoAUUqDTg1Wg8vGy3FoULs4K5G
vIpD7291wBIaxOpC9c9sv8L2HtG/x9a0E8jgG6Zm4ME1Y9mAiwORTpUTqBCydqfjCuV4tY+BFE3w
ZFDVB38RrcGTnvJ9X6Fkxoqn2kKmGmnkAWkqjEcyS3i/dnkGESSploEhdh7WglWh48kgrEU/ub8h
gnsLQUepKjHkHsunSIvADyRX1NbfzCAAQ0g7X2cwoP34lTCaYiPAiKLOOLf5COmt3mgDBPpeTq7n
FzjK9xj7RIkggl8GkNftxOX9ZUuXnx9igcuXfVO5euNV9yrBe2KepP/vL/vcDxfop3k/Abkwhfg6
TjQCevV2dXn1Naon214Z0HrR0K6SjoUW7zJJdc6dVTatd+bb4UjVLKgD45mYSsPwE+4GzXmqgcEg
VWhWVqYBbpLwrb1EyEw/O9D99NBLUWpxyCry/ABsHXre5vfYbFLb584bwimIxQ4HfM952sXjScgZ
qCRjKc+HA4aP6MJjy0oDGLqtlI7SpgxuUrXHGDWUgOZptuTYZgyznqhR/N0VHM13XuSoJrBsdt7B
oyv3lbFqslyJPeZAtLQI1/loWDDOqQzRzBVERdfGo5AHCGJgkZ1Bu+eSkI8zp78SL8EyR8kBkWrl
te8IOvJVtjIPurAE82Vap/eMwYOuvMrW+hPoGZ3Q8lEw7ntFNLLtXocsYW4dv50043JWEa+h9HW2
XhhgpulMMnxSwGUO20YTfb/4vRdxTZYoMVQzbFpKILKBeTFgIWZj+AUPeWvbg03zCp+ceE8F3WvH
48nYj/S4SxMhGlPYRXZPwe9jkqg/VVdOZesoc+RFA7ojzKXaz50iQcs6Rmr04xRoHW5ByHL1bKeg
Yf8MJH6ZKN6wU2309m8407RGfAaFvFtk/K2OpvDvPDxw/9akqoHgNWxDSiR8P51yXFNWFiEgbHXQ
B+rYRcFVKXwUaZJaN0pYu2XQv1EBcWarh+dB0OI87Nejbm6kU21GwLW/w6ieLQxwsH/dHaIN6PNe
hc26Jne3OazNGQwSDD15yyUk25OAmfvMmTHUO0Wg5gYseyLP+HDGK8G3WNNDZVupa9eetpDAhx9G
1nNvrN2j24tG2M8kwUAzIUxXZqZmYWV7k0AbcmaHGFzbD/9wtw9xHdGwGwatpR3TdORPeRDQeXhp
ap+EBQBcuZ47t2Z6qUgpEjPWeKN+WzhHkbvCr9xy2k+jYJpML+ngIKfcX5J+aYL1NagUVPiToV90
uvFAmVno2l3JJF+ADTMhdaYEiLUk0neiaMpbEZ8k5tJpwijKQ78Y1QEDdOFZs8BHZQ0QEDzdenCE
NIKSHYVy5rV4cW2v+oZxk5sryZX3LmSBpEL8HPQbDp/E/kUrxW+x23SCw/vJn9zenQQm0921gg7+
PIOkg67HQqgmzDmfd8NxP6KGp/L7+KPWr2qaMAVjQ1fcXRfHYSuIajnPSfewBntppDkx4lD2wG/G
lBVXGXFrq1nddSMVwnWYy+E5LKWOCHfZTW6vsC4R/KUUBjP4JHplOFYCdhm7yonS5dpUKAM4RSLV
17NlOG1lVpRw59ibjW5Tlmqn6E/FFtnpQWcfNjn6/nHik06TZETz6K7oLW3KbMcjVCpqEFs2RVJR
IWnSWE4JjJdCrbH0UkVwlu8p31NZTBV/0W6JmaScRdcn2mPowEQiKNsomHqezwQjZyxOo+x3CSKI
P+qXm76c7dQj8LQB7N7WA8BWY3E+Sg/efkLCmXfKRmMC03TqmWg2H/ztBYoMNX+RwECCCfThcE1z
YWGHmtv6Y8KYaT/iLnA/1FsTI7AzN7cp7GYDMdiqkIEPMPHWi2pCYsg9wl79GgVTUAcIykFyKh+v
d6rJev8SPjwNoGMTVkhIWTXb+QwLk9Rp5n/SX3qKBjDUZSbI5AaBQFfiv6KkqX47hr9bSqWVhPtf
0unCwdR4QRjKn6i4DcHejCj63qpLwyCJ79gEgOQpTv5wVz9h3EbQ9N++lgVPhnW1ZsQTK1ABJ55V
sFL+rafsq+uxWfD1te0WpH8QLSmbBjSydJVNR2hHelxZD9oyu2Tuyp8KOEt28LY20/ANHf/W2yxg
RIXn/oif48bekMorOnDmGbdQb4YbkzzutP6+bpOdmx7/gWcI76iDGngx723to7nQX2OzOu9czcMp
qwGeipnfgEa+PDQCJoPHm9sBUSy82P1C35/Lg7TcEi6GVCYbAkrOeRHFRWGZRsaMq2aCdARe/mcP
qxux6l9rc3kPfckcZm1gj0hu6ibxbHoHvx0gQSQ/sl9CAV0zwn9w0PWCl70JR++q3bSxEXhCXz0b
/f01EE2KhNl+swfTNQefQPkH7UYShJcsHmtF1vf1pLWLFqADHSPvlmwiv/3ZRmDAGX4e5Vi+mpF+
ouJ9WHH+jUvkXXCbIX7P2/+f5/o7KEImc3kI0miwILUJrA8eQO0dUd35chSBVg9/yyPvChoM0fd0
77MxpaqsNZ6AxCQ8Zczg877Tn9xQpIv7X55clJJUxZ/IzqqVmM1pDczbU8wFx8IqQ5CwJR/uEd1B
zCD8FsYPmPi4TgehwecMnpthIAGCWG7ci/8xFn9UbjZBcZul61nK/zrUOhw32W09HTPOmqa3uaAe
dcNvllBsU3NFm5IcV4o2wBS5Ng060/K9j3OVCMJIod9G/wwKioyxirL1cTFKYeOt2RdG8migcbu6
O9aBUsaffshvkz9fgwucpXnJQb/T2g/ZRbuj9N4kZFesvK+GBBvTnoxvTyUQMxa1Hqq7dVr6gBrp
wSw0+OQIYGe1NBW3iIwM3CrBj87l7P67ds/cc8NZlNBsawxrxvzK4jO7UaOoRmQ7Dj3BFUGMuPYH
Y0nIeHPaAktjLoeIQuSWbtybYnU45eOmFFTBh3vGNdbYPE0rGFPvKLxHKQIWV78o4wBkyTa4YwKN
FnTfjPV4DLX2y9C+H6lp1YId0Q9XlSHr4U97tWuR1hh7rKfrL6mFZAFLhZpvPhGzoCo4CpFUZugQ
UwISPJL8nUl+oMeUIRv1sqTNC/RGQjViHddw3rXz9Gy3ncTFnI4EfyWeyTgtyBm4dyVBBRXg8ZD7
RJ/LaPN5OgAKGBQTsdoK2Ha+GU87XMtFnLBptfvesYErOi0KBxr3xN2zeqgZQYUR1huIGc/LdYto
ZNW2exDSUhZ9//vaXk87ixAUcBeN267EVsbipSV8uzQpt1dWyXvor/GJjilzHQhiR46Lg/z46c2m
DW26IR9GNUBBbFL9dLPzGRvM4IC9USPjIvCo+FbHzfIRJZ/zkfzz9F9wI4xBL9whHLL0CTZhRqji
3dEDd6FcOEUiygsoCIufZAfj+EV+dtOecn5MqnFqSUKIuwD3s6vSj+K3cTq262PCdmYW60QdXTk3
53hg+5QZQztyDBJbaIp16gEddPOh5qe5egXoRISXKDjWaSQfXTXJIogectG3PQf6eHlEJWhgU+r1
K8rVefqoUo1BFzQAUyedkk50EAH4R0WWOz3l1wIaYViBaNcLOlRTnp5VMyOEnFbmvVdS87iFagEl
GB0VcxCwJY4MiyrSukV84ETu7mgsFTFKrJZhBf6CGP/21w1MKgQHg3BPnAkCj8N2JYJfCt2sveRW
y2/o1EJ8tEYzkEi9Jj1r9oD2EVw/fde/kniu8GRr0a1UT/467g6DTsISZBfIo4CB4JEHi+4nspxE
/I0HJDzTTLzIbj9q5gNu9FOdQi9dsjUpZXsUH6tDgTlXfF3vr4DyJg/c2Y4WIUBd0yU9GO/lB+3T
UTjTeCUNI7mh6ztBLDFU68dgzJsJaEC6MhDSOazJCDsykjls+agNJ5KDr/brGLbtdIQmpStENkKS
ZRB4boDVbwftzrVfqwo/DvuBoJZ4NdOQcxE9O9mhiW5CoBbfBrlTkSeg4wblGPlc5RYS//S4rHHP
FHPP5EpbU2NrcHrVIKZeRsmIxjSa06HPpXltYbgXFCikDJO4pH/qXt2fpksD3hvXaPqqqI/qvuAP
tcSq4VLWzaRl3De8lQx1VWcxHbNfFFvcJWeT3KfzacAyRZxyoFbcj1XVtr/dFcX81Tgev2VzZw+A
bs2D7WdVtukFb4YMKqK22/kToYz98sydbMjpBRSM4rKtR6fCYuoOEugSSsdGRzKX6Eb8oNzgVSAi
qEglZSPbAe+4FNikuSHFdY5M6LQvJg0J8p4eDoijMNUxsL58zk10S+eRk1RQwuaKqQH+V4Pn0+VZ
Zn/qMbmqmwPhJZ9r0zOQ7aC0tMzAfsJgCnYtmJf/NResV2DJpIgLOhgBtjg1hZFdO2+MYieVwRyH
jj0o1wwG2OE2QILr7mZs6N0e6+JsswupjDsGwTbxdewsDHgGknAVCZkBa+zIzwKbIydv8wzC+D9C
6yiD0yD/WoVkh36zkBgginnJgDCI+zKlFk0ed79HyunjETd6EL2BSGkq3K8PjQTQX51yEE2M6wcs
xNodktxTMQ8qjSdXdlZg5/WhR0F9E2VS8mxR6STNZfy4C0EujLirlkUW3ayXNyzVfOkBpYYsFhyJ
b02VYmCB4u8kY4LJx95s5EtTbsr5YU35E40pfuqJDMvJtnIvLKyya/LGXm4j03FLpJFu2W9F1tlo
6iLdAJPqkweq4bV2nVfgP2aFFnxGqD8RMBkW/H1hdewcMyqT4Rb8hN7yRvpbIy6uxNvlkJiQUKAm
E++Seg18U/kerazxLuYYPuuWZrLnyNcH9c7vtKRauUv1qo1LKbDZAXMivCoV3muqIUvqHW4K5KL7
8Dg2x2r/2RyomoIDcrUD/A7YiWHFt/zRa1jnJfPj1gbEn7GDncOhB6hyutN0Cs3baL2ThtXGHxVf
Ie0r/SmcE8m26DtdHIMrcLYWuBB7V8wJkVE8EwHOUM73OFkO0wpE+gU/YYxDTby2fsgOSLWwolDN
s5RtvOWzy3IdFHJo8Nf8nz7mkDYETvgKIu+g3D4SzoV4pAePqlrGQgi2CMpE2DOgkuzIbVJ26gIR
nBvY/XSK6Bn8O8ctKPZZ6729cG58y/LU9D4F704zXpr0u8XJBUQ+fcNWcCzuyTBeDd8g42DcRxU3
U9pUd00Dhk1hIajdGsO5HuyQk0b8+uBN/DivR43MW+fZSwnbuUdGim+eoGMYFGlYQmnczWCWTCOz
0AVlkqtisQ/XdwjfcgzpmuppKt+3nzRHJBv3N7H7zmCXqsJTRuVt7e4AinWSPGCKs5ohVTn2Xgn0
AI/+xOA5nUONHOTAO/JtQY2dS+D52P25nOvfJWJPRZAyJ/oR0V9IrzTaT3usTqHOyGk72yz8a8O2
sVKdQOIqwL03SG5BP8DwnhzOYrUoSiAw6+M8WeBMperTEi/BFq+q+5b9jM2ey4d+/CHGDrlw+sM/
feklizbOsVhRleGrZrAIUYLQhOt7zz/PBwhqsAejq2BBVpHRHHb6lhAwrHuLzzgZMGkn/4k9ATx/
iy3DkuDmP1jdYzoB8rcFZs0IEaSjXI7ygxU54/gNzacw4pD33T+joPQOGDg73yFDpZEY0fJwRXI0
bkctnfr8SAFF+sdsP2c71O811P4kzXcbol7+KpYmSrg9zaxMIOD1qLmAxZ+cFLPOlWOU1FFp6ufZ
ASXVRl5tPGYdvnhCMwwwbB8Fjw45N/e1Pi+KWakx4iazLAlZ7RQeR1GaXTObS9IIjBxCGU4WK5Nn
L56KkeJVpDrRdklaniGuOs2vuF2HPmUN0vrM/1gbLyMVCNFhjjKzWiIYFblz1KXa9AK5LNaxEum5
fQEvwYQx2dhdKHdOXm+o//xvW/Rsjfs8rLbF64ltfMayJIsUBjf3TLPz1LVtfAYv2ybm7cHTHml8
BrmvT5G4vMST3b3uR5yNhWOyel+zX0evj0pbsjo6zB8Yg+v3OK+TSdatgSybJA9JXuDjD04Sp1I7
siiEK2lZ3/aE0qrE5VDm/5Vi6TrbLCy/tgD5vbu4cdUV2JWMb1Rk31tDwZEx179MwGSjSs0jV8wt
LdqDQgfCuZrgyuUP4k0PfWbS5L8cz3XTzq4zz1wgb6PqDp8t51Pr5vOwLb4U1JXNbSq1dm1T7Hz/
Y959HcAa0d0uu8tw81ATnai+3O6b3YwBss7di0P72eMdiVQIJQta6UAhthQHMRjJMpg956wR7muN
UlV0w9b2RW8dhUk+//3RehdGSf4HImOiq9M1xLDP7+ohrBlWLUtuIyyub2boubEnVgqGRkYo3Q4g
FZJc6T4pb1m46cG9KvE5ghYfRC7jFD5mJxoYx8H/Qhu2Q2HsJ/ietGRUbAZHpstYXx6+tHN4gWTb
TIKKvdzAnSZx/ktSeLhbhDE8h62VxxL05Mud1pgQP+x2u07r3xLmIeCzNP8lZ2AjEHd/GpYqwXTQ
QzW9CEYwazwO93VBr3UIURcF9ahjeDfpVNPA+QqbFbIEs5TlFtcSTecql/lSCoCpynBOPEB0+g0E
d7qpB+vBXOT08W++v9xSFKZHue8DbCanE0Rbbr1vV7PbCPERUGQb+I/Ej1xi1GN1UJs2prbMLRbU
mKPt7GjdtB0vOmxJLvO20SaqCpn9qaw9ivFedHrY4maLm6g3cE66qIdtq+Gi7+tyaLa91REAbKyw
7xqxrEsKe9tm6oS44Htq1+2kXnTJCVaY+28uN0EQZrQ8OdL+2i4FxTYbYdrs072eZBe2XutARuar
L8EvF4/8lcnqohLMO5dGZOfR4aQQRyK9F1qvcFoth7JDtecXfftWSmZYdZoMwJNpfAaD9Ai0myo5
DnPR0ampjAcpFfKVqlLX5h4HMkK5YEeOZct2udjV8Ql/yH5buq9f9Mwbrsv9FG1erVLW4Qc6to2q
ffsZ/WGMNvNJKIARHVph1y3Br896IE7NxB+8VN9VRS655KitutUvXGTaQh4VKpTB+o+WIzMIe5do
XlCCEz7qbd2uGhojh3eVyioazfQ4xGnM88HWqOMsFp9kajwveeE+RA+BP7nIWchIMKEyyBVSQlLI
R++nr7xMFzZFBduePSVf3b8xTn4Z9dpZ3s8ZyugumNhryjZy3Fp0KoHzI7xagMQmEXwLYpyH0atZ
j/ompHx/RPi77+ZmNsuliVKQBaOJLm217/8J5bDHVc3jny+rArNqIOsH91Os3gZDnsrLo3GwqmIP
iP33H+IPc4Eag8mhiC273d0LLX4hWKV7SBTjO4HUvElipXxLot7T2k1rLC8AwMeVbQP0QWbupkha
5o+hJSzBMVeIQ7/UQII8xpOQAVVSGX1ssgogDf3F67X21qheZfXxKpqVrYnPXFGwluhQSncme25S
fmjma0moWMjSy9XQ0/qCqz0gvLeDm9PJXOL5D7y+sltp6ncVVg8vRZDVqPzOPakUdZk5FjNbqd0+
OMVSec6QMJ3sIXI+fqLJgrBZOo31VqyarOT+wzEUYFgSkx+Yo7zGpsE1GHy+HZn+eTzafhAIVtLD
V1FOd9Zjy3xNDkTpvc77xqHwOUkr5MoHYZayiv2B0K1p/fVg5vywMj7zxjY6D6vqF5TVXX0I1BbS
53m8PEtHfOAg/H4Y1S4BuRxS3i5cvQy8lCDWMC79EMubgzz7v+WkfsdmyW+1FDtfDEoq8e8dhvm1
IurtU+WVW24lqyNyakk6UhmY2yk12PORU1PkPQGf//N6lLMp9ojRgVYgCfijiqgiDyZGvY0P/5vu
3KxBQfRu2L63Mo5lLiEhuXJaiFZOrg0KoYVjDh7KFCxmsffaOnDsWKUb5T2rpqlmnhQaS8MHi8V9
iPgfV00ILzeRAapg4cMoVGR925kFUPc7X+NdJZTNoYhy4J6CIQ9qdJAK/uVx31/CshusXqSpgZCH
IN4FGyqJQuPDTgH2xaxNw+3fMceM7moY5z8UoucLg7XHYDQtmW1um7tBrjNt+TIzUkdU1NW2utye
m7/O7yBx3uvjbL1hEDZq6uh2mBu4DSwkuVf1XuYu7xSgsfcJyukUq6JaeAy9uVTWJmfdh2FL33wH
/0pjLe54+7aeQzEv9AyvYa7GVZvr3BgjEhr/8PANVhOStTMr+e7CkHi9aPWcw8nFe/V642jZIqyn
o5AqG+zjEjsHFSyNbkZuWPTWOjNFfZh+mILXmZyhKNC8HrGA25sRxBeyfGtnILIabVxrt1Z6j0Sx
VlzBr+umL4foQlbmNAK8FBah2XCHsutpzJ66ohbjk3Q8ajabjyipuhiwsTE6X9Q2kY41/fy/TX01
Ltk6DAdulEN1Q535tnfOLqTQ/Bj65jHMWZjAY0CgTCcWJW2DhB71rOqIWDx5qZPenEIc8GW/c5VP
9ts8pVrUVyY+OJAYwa+sAoPTQr3oUe/6QQf4n/9c6k4kT8a6qXx4ky5bFyKB1q1GgchU2jyl2Jgd
6zg9doJu+ujrncNsXw772zmUSHUtxcqT2D+2p8ruceJBgAojsmeG/trPYtOmN8kpaq8ilixBJsYI
ynYej2+A45H2vW0pmiURuEtfQ9J2YSKeoqzNs3KSCJhykF9g5UNwFrgezzU7XFvp4XTJSE8h2zdQ
UqXZ2vGLYsVvRm4kPNS32a0sXecVr0i0j2YsZ2dwHcJrqUXb698/UX4NdEA2Z60v926nXBcX805k
/XVlkJ2RKSY0pbrnS/sKnqOhu0o5GjQBL656tWFAozVNA/uxl3chXLPXPc5oMnCKaeBi/73lh4Nw
KtYPR86EEqbWGN/Rsbw9B9K/zccmyotf85xzNYy/0sfENAJUvG3fR4CnYNXMEvHFPvJSJg3A0YNB
Zo9U4bZmJY6260VTwAGdYLwC0m3xT2d88L1RZauoUauofX+WcqL4IZG5iz49GGu8AjUBR1lWBTtJ
BbeZQTImwrCb1fZh+/sWZcTCqA4wQT6kl73KqThoqBrOFcFyEckmGDX1SpQnGYfIO5Xap4IWA7a5
VonwiOCuzJUoPKj4cnDZCUMWGc//vn7hVxYprhfH/npy1Z3bn7e6ExZyk0g5GI2wV77I5K5FhyX3
KwAGO8Sem/akff1vx1RjE80ay0PW25cU+CWIfuGCbPl3C9XsWdexdcTFtI+vKDaMY+Mu8CiZ2B6G
VwtTgkLHb6koMFROgogVIBXlRWowUZMLvmqgsEGg24coQ1W9H8P3bCIW6S+Up30KOdtAdiKjJPPK
SUnmuK0FI0fZwH9Lg2kxVr3uBw5qj26BWXLVGKl7xp8xEWyR5s0r8wqznPjRNKmUc/CS2we3un5S
IRYU8n6xEUUjA8lJJn4b1pnqn9IDg+QjOPzwnQ8xdSd8fV8lm0cdX4aHANNTsOgMmDg8IlQeGalb
/gHvYo/4dP+oEiQwYhEUGqSYTqIU4jVomp342iOoLyl01fJGeherjzBzctu0Jpterai907bTSuk9
4rRFhVY+5xvhjw+ljAkqhNBDws0v6SXUqNa512F0cKmo9i2H+Imvt8q5w3gF27mlYbZVpf3G+Myt
VwKIrMsmpYBm/6vF6u5vC2V0+CzeJNMtAzq8DHfuZ3bhb3CidtxH32569NiRi0Wzq2+qFVdho2WU
3zZaw4Imf9sp3+DdqgRX0xBR7k9Q7jdF/TZzcP7eBsudgSTJ45/Oxi2+hE8e7f0ZAySt8863a3xY
lHOLexSm26XwokhNALMmTQxSI2cr9gbskkew3BshrhfI8fTupRE/2Jef6Fy91AsJMo9X3TDnKucC
XgY93U/g3wQ0GPrdQmLbX1YJZK3A/w94v+hHA2Rugeg/Sm1kGbmCJkqKa2kjxq5mDelY8OZ58qes
17QrcL8e4EqbW/PU2P9Cd29ABLM5+qeiwVEgi0ngIMd/jNwya0is7RhMVpewPPCtN3uZbM8GkMKg
JXFUaSrH3VcJ3u7+tT/OmFsrP8GwUthHFaglFb4bXNtK0f1KmnJzrCIw1e9UOo5iSh2AfABXsOD8
NjN4a12GIqQptI9X0LgIucCJqYFMLz1mOwlF9zjWzMiG/UHB/UBxlwxzfAjlDOpJLYNgGFJIFocl
MX9tBPKdcM7rRCXkDdtjBa0LPHcMdh9n5+x4fVfCPuvPAQ3r91O9KiuUHsOUImLkcnu5dwKCmNHm
psO7X+vooNVBy+53JhIdzm6jyOBM0WyQsprEO7UH9tL/E7LBkUTefZ0oz3OQTiU0cYt7hvIAloOH
BCcinIINKitSIABkVp5VnklQWfXgXDHi52O+/0EKFVH9qaIkt7nHHWhFU/C1FeBKQ5nbUKJajPbr
R8XaVVHOzSIqHjFC6gGcGRMA2a3ejTsprWAbnR2feXBMOPmrBz80ECrRX2jKGKx/1auvusC4kEEc
Mfzx7Vxd9xaA08NRtOjk7Ozq6xvLvdk7Y3jDVmQvyK0G5Pq4q3NZK4ptr5YbQbfb6ZiHi9Y2qRDb
QZUBimGs/xQ2sWZO21ZWCgnLFwwYXt9IgaZVMwL2wyxm17dNY188/dy8WAu+HFrE3nhH2iDu05KZ
lNNmyvdJkZerUnJvzj36TswZDCT3mi0cG9gvBjnBlU+9iaYNNAdAAfspqrSQvFZny3J1ICr7NYU3
5Q5Jk7Ssr82Ul9O9zqz4oaZFfv8olCDOYKR07pJQDFN6yE5CkaY92CWhkLcuw/STBVe8vi2fSjfI
2k8wLQdHtD+Ws3z+qsyOthVPxYjxVRjq5s1eRrq4E7Xp22pGjQ0vxKjRz9/vN6mlRZBGVfU0bCpf
8mNH34Ew4dBETJYx3DcveFLVAeIRZqmZkf0c3UyywCVWPDtXOn305EWDez3m0a7DNXPtWWOeCsWj
fBweW6uVhpinAEtmCc3kih00mny1XjZVBDuKPw7epKbg/80mGfTsVh/KJfgpJcA8zuNdn0QN/9hh
74W6rvP+YJTmqFZ3vcNQ3gHrpDB/HlSMDPNnVQNFwTJN8yrIC3ge/i6Hl+jAXKBeg5aSG26xRMK8
3k4bkPFE0WJDjDOfgwOQnBZFDDphS7CmAY7Kjnccpv+As4RH4c7K2Ud0FEcJX27SswNRByUKCU9D
qw9T4gfFK3NdvX4ddQQ/jjeNYn5V7TEEZQKxsY3AwpvjVr5Q3SmOduLcW56AWfCdxMhL6GkU95WM
F5eb+1sneh8B+qTbVjKtz6Hud5cyxzKdLnxGJouNyoVZKJJWu3T4VOqZt+OuUTfbm4tiBnqApgzh
oB0WN7t/YxX4Nrt4faDMWYROySzT5oAmXl4Rn/5tP3IDvut/qoxMdReXZB0aRiB/V98fRMF/g35z
j6S4uIuDPNGLMzxo614E+TzaNC8I3Cdhvwfw2o35jF4AdyPhQIo7RjdWYKwndpVXf70Q3E2N3Uj2
bUby8HGPSnXp7r7fH5sFlD0PkDnLob2HxA5qZHhJ3t7cnZ8cdsxC0/ZuCrlNcj2l3pZ1fZpgWGh9
gaXA3Ek/tIkxh03vua+pxG6h8CgsK/R3EJ//WD88nOCjTiyKU+nYfJmsqhxqGC2oN9P+AW+Qzcpg
zECnNBOsE8JohE/J9+4STK1q2YM2A1MTwPn6gdq9lIqzeHFQrFpeUGnLg7IrDPd66l1nGYHdhfVx
bglybF5s6KgBlPMOMCPN4/fdmzw+N+tkvpWyJj8QYmh1au/vvxG0gH2AVxbKhLfp6nhy1Qqw5mBW
dgk/XsAVC0QmcRcTuRhxOlyVBEuCIazPUMnKXcmFRmbZXAI+0ObNdgCgRqwOlNyYyTPLMh9Yp6V9
EM5QbSlwIwopyVFrhCSwm90pt6LAu1GyFTJ0ZchBZD5Jgu5cMu5MoD50611eTahwhHTaMF1E3L+v
kYghtvIZxLByiiGQA6wd/2H0tiT8ysGe2Ax/lYa4MQUIF3zDyvCM+kuCDEMKI4+JfDYWp3ewSF8q
EVEZnWXtwtLH9154jnNAWruUTsq0TEy4FNpbFpf93BGRGl4fLbiQju8HkUs33iFMRJGMHifJwV7O
KfXyQMiaxzTQ7AtGB6l0riZ/0ws98Jkqy+5OnP3cW1pHEX+E+F1qYPiSXD62k0rs5cUZHSZzlMqn
Z+OXWYwDvj/8cBbczqeYOoqwZMHU+YQ4qyZU4mzR0C+vZXADqOs2h48nSviODWjGQ/xYXkJI3rEb
Ih274NxEsMSELoStDoDfSDR5Xp37OuxQJpEig5MpmaPVR7eb5VZ7t+hccBepvzWanBIXt4N9d2Et
YlR/E9cIMkwu/xfyZBx6FYdaGCEWgRjK182oW0X9wG8OlRntulAKAvApMenmcF+Pf8XI5EKskaV6
/Xf7kAuZIAMmZjOVSNT41mGCC8MwIr/kSlwqKDFE6n9gsX6zVlLPOMUte5z2s3mcq5Kg86MVQrE8
yYidkGPh/vVLGZFtvdW0LTCh4htnlsO8GWLHVoeiFzbTB8Ykc2Y+MIRmEF44R6KleifCz98XFYZH
Gah7gVE9QZ9yPioSdnOJbLuc20Q9IHsY7Bv+OEPqT4hn3l6IU+OruYP2RROBodVleNzuETEasgjm
5d2yj3j7MhXf8Elobl/dahhGHBd3wGTyyZIoCsmAvEVXYALbYvaP73Ed4gkPnbfno6UTw9pMnt3D
NwaLSDWCotjkwfzPJimqcnBaQDNZVWYZiG4OkO9kutYwT4DvzSZ4olqadRP/KgLoMwklIav5j6/R
hCUycMUWe6IkvfYNiZh54iwyjS+2X09CPQxI7QjDdkRuSh15pJtot9OmPDTseyd1xDW0r8J6TwKK
dNh3cbLheVrEZ6MCci6uynyr49cNPbPu44swn2XtyKPJFegsf8PH43DwpIN0ck1MlYbVXMHeqaef
jSm+9ku+9OjTHR34ARp6QaRAU3OZV41hnQemcB6IfXIqjrH+9wq3HG4aTIQ45HdbISLR3+aqlnZ+
hOqZykabzpDIcVsrb1Y/kVwTzJMI6lqmaFtf3Qqzw6ovxuDdgSmYfguwyDGErXutaC6h4E2QYoxQ
kefwEhRLdIO4MX81MYyqOC2Sp6a0GluTwhUfLoKQas2Bsi18RNbf1bnJJipK/TiZhTAP6x8Rd29U
FiNyrZovxKjcn4SAd7fiSFO0mYLXYhEHOL+u1xapSXrTRh3ksxPZ1rForKOhcReA2MR8ovsA6IHk
SFwBDNDizhj1wg99vaVAio/+PIUKCRX3hFfjaltvHtYH4i8LfVM99HUw1k/uhWlVrfJzowqC3sKE
rNg5BOrZx7WcLHXPF2W7Hu1qD1rgYCMqjrxJ4WiGqCJnVKIZ3cBncUujXdsDaQrfrAHrYboFCT7M
/h0xAZ62n7Scmwin37/ewFo+caeK8/AXnuBsSAO1lk9gjg/4v9t2dvIcA59sXsghUDSLYqXoc7DY
zz83HRBPR4yLYgRkvzCdOSE9Mmdu8Bug60z5dpvH4T/ApS5wAfzrcHJtRq+Ay/nUV9kE8B+EKKoZ
7ZqWE7XTaSe6kFss17sJoN6QHpFOq7bJpXyiDgL3oCkSMhdmDv2zV0XARWd2Rz+gRSpOiSs62cHT
16XQugTmhYz0IBwSbb6yPNcrATq/U+zDosSFQR/TmReItd4I8xcU5N6CiXhZR817PiWsVWfJR1As
Ju53x3jM9PCF39IGlkkRFbG3VAHBHsGPzgWaPEGkHanvD9K1ZfLRi8flUu1SAgdI+zxzw+JQ8PPA
Lh0X+f+NVFskEkLvh7lWdOJ9SQdAfssIQ6YvlcbqGiuzIPYEur/mao6foY0Wcytq3dsYE3DmecPN
RlrxbZyt+oMvwpMwZJ5qPAUg2diCy5fCfNHE7q/8XtdMLNZM/ePHDgWOz2hzgIEaj4cCwnoknte8
On8be/QpTLWGAv7Ws7+2lDhIeCnNoXZ9BVRbqcb18q2wjOijSasbRMJ0w6w8l2+K3xDHHgE+ChSw
MkwYPFoBL4uxtTX2NFdbqZCCUcIU6klILzdCJdR/VeZX1uaTFeKL2Ua+mWVTESHiudg8Ajz8lHGw
YxTUNll1YCAhVnTLfcT+LLVXip4cIyDF7WS8uq8fD6o/XUsQfbLiKtVGQPE2MW5OG2bNmKvcCEVA
S96XjGrM7jc35ZZCfhm/jmuXJuZmcwj967IiTVsycg1sN2yzhs/K/6hRCwD3WeDySkHyFyfbu0GH
IS9v1sJNV7bC8GfyDxy2n/y/O8eNibHQbJOG2cyPi+BzTqvOd81oAwxb75+7h0LueU0I3Ni6VF3T
lptFHPATv6R1FlgQyrmUrBic8Kp3xoo6sKW78Ehs004nia8mXUkqHjMHYu9+4F5lrG/7guGJFwgo
5UikroSvWaN2F3TFT5k6my27YgKSBnz4k1WLVNsJJMwI8pUHErQdXRvoCWtPfvMqre8ehKqRHzgU
KdxYnhw9676lR0Cl1C2MNjYUn4MB84g6zSlAkWl6P+wt6z90WhxeCddYW2L0QgL75F6uBooUC9ZW
HsuR/ivmb19q1OL34YHPi6IQwNfsmPu/AxMK58qzELtCatll50vPPP55OgTa5SJLJ6Eye7MeNOKe
nxqBGrH5Jv6bBMLwLxuGg8dlaG4gKZmdFMw1WmaBiyjURxrr/atqRxip7hL7d1HuUhXD+xORF/U2
EgBNZPYMlhX6cgvP3wHJ7exeUQPom/HL+H1KPu8ZTGyeF8QMRyoN8Ft+hd9KVx9BGg5bjdhPzUkT
Y/Vx0VkCt+xceAEvu5TKnyE6EvWFz1ba5rfWKTOI0GNneVjUhcjm+JVp/E0U0D6+Nt+QfaqYV3FH
v8Jlke3ERf2zi08VRE7j24K0dghW/5ja0PgH6qVagLjHx41+TD2l4i3erKFgVOkj/XCUgHWy1JoR
hYJKSUuGG4tlNEvs7PpiZI0Nha3TLjOKOPMpBvmpws2NxIc9X6N3Q/MSORpvFH79hfMQAuFNevCS
zdcnQYPocHm7qkKu2PYHfai3rTqyJHEXDm52D+xemCFDp46Eg9P4Gca+TjzU9WZEBGc1beqX2fEk
qoYEZCGJsihXwgO5rFcogAz1NsvlXVWXmZFh38D8AxSeuNCFr5opDv2Y2FoS11ssnY8D9Z3EpJ92
ZON23QqUrMC62gKi10nrrYHit2W+wMPa5tR/5o4k2RJAZzFxUofxwCR/Dpkz+A+mXL5ZoNgpEHd2
NeeWrRNzApLdANxjjrPS3nzN3A+X4Fmd5I2T3ycjeOifePBSUabsADes6STyzwZbTRIMVAiaUdtP
R5+Q0wnlBtC+wp+ipCyFFGkhN0l8rU8oIJr0aMdpdplTynvvbelTAuor3w8Su47zZIc3UipQ2TjH
YCmHdZhZRvStNHP/gGF49xm2nGqbgErXcqKToXQCrRzyOEIuAknGRWWeK0LXtGFvcl3gCTIbE898
FrmGLVe4qcu7nUZSehYDL0mRXs4WLosZuMvXuR8W4jtlIULfv4xs4v12XJPx37GwblfGW2c+bnmF
v+YOI8cViF72ykIl2AWQRGk1+SuDKWQjoIxMNDKaTn3/SNj4/LVLptSm7kuVUR8T9+/xaMYBK5vi
ZDKmp1Fh9TK23dFToSH2b3e3V0zQ3Jnn4JE0SFxn5AoHS6EjhSqSbnQe199ogyWwLYnA4imI4+Br
7yy6QsOA1YOPBytRUziD4mjE5gsgsqWHoz6gWzO/5VLnKB3CbwJcrVjRWBEmnRj7zrmQCpJwgm6N
54YjY8AONBeQ3NS8/aWeZYQQaZJxreycUerLYsDZ571b7ZrOwSmTbEow4ekDczmfjO8cEP0Otd7i
e7ZHKqALsVJRGA4XUTTBk26XNl2YLr5kfimLkGq+hhcFwBEdC4ptrlG+LuzSQRJzhUA7uKtnd0vr
k5KsH399VNP6DU71a/g1RbgUFD5e0v3xCITr4ZsTvccFycR5DzFVodbzLetDuJnAwxAdVkWce+Lf
QVrEJAxCK6Fh1ym81sMv1QTVMRh7KgPzYEX4jXRAC2I0PxHScBPMWhE/nEueAYk4YtDruf2UkvIl
B/jRt2mOJ5IxZzXevv/o8RzCOg+hDOytbJtSJUPFfZfRXyoTN0HL5+KHV5lIT5usrYqZpLD3ae/p
rC+xKUfmMXSqQudz8RBQvJez69JXxm5IKpv3efP8d0KMe4IPr+FxL/ulHHfB3HM8JJSbcE4eZ2bn
qkMVN5R0TbJCK2XYk1TlsU9BBSCnzYAb9HGNzbVs9I9xwm6gkNnsvjjM1WAQdpxAECW10QiqxOBe
x7U821P3I05z9UiG3qoeptC8CXZmPCVINIJ9FEq3qgyNnIL6naf6sJbplsRo63Dq161gTkzpdBe8
8JKc77lViCYXSqCnQznIbobICrmCUbERtBBZhWv4+Df6x4G/3+3WJ/VHagth6rHTE8SD9/h7wEKc
p7XW2GD8dgEFUYodgi1U8wo0ZyyCbmkJjHAGTFlmhndBPNZnJHxcRkO7EnvcRjGc05kW+3IMxiok
vIdHG+z540oeiMFHM+3Yv8jS8HDMRmpL90vY7VdGmi6zKvjESef70ed9Vh7mKwakyHLexVXM63sh
5dxltFP8HeAPqrn7uDDrNzOb4VlloMFamzi0y2CVytoTKUwHOdQa/9gLdio8f8DKTRBFl3qF0cR3
Dz5AE1IoUKA8r5X0tBBXqu3J0DEvwf4jzoz0c6OembGJE3rnfsCar3VxmRAX/Z1s8EnalaEUXRDd
O8YM7cy2MTjfl3okQEaGX29XKYFe0D/SbAOQbnNs8rkhhyo5NAGoyA/Yf9vmRujms0JHqK2cIrHt
mgxoucKY0zDWelOEdl4BeMDc7Yf5l/riTqbul36nJVNxwWu6EBcBQs8KSjaMBjNKwNWQcHJ8NhkT
/cRi41557xOOjH3O8BBPfRk6bbLpz+2c1dsn1ZqaURpTovqiJTN2tY6wbaI+F+hmEe5bPvDXN3D0
Bbk/lvUQGuCyU6d8xPmJDTsT3u1ESzyBbQEqFlrcFQNSZ+0Tp2Osp5ty7N2vKwr6uCrjGlhxAM4F
wI8hdMWvByqqh+9dPPhvqA/260aMIXnsoMc4H+vfNT3kPcebQy1B40FPhd7m6IFzX8AWl1gh4mWr
olCVcj2aObWM2lQH66YiWDnrvwoDxPjqX6gq3rRTE7Bs93LYVmBlnDGkDc7tRYbOzOEMnspdZLfQ
yZap8apZxrKJQL07v3kU0H2r51edbX7KGn4um58iQroba+UPyrfUIh5ofFZ+bKQ/7aZeB8Lf6Qjg
Kq2Xtu5AMnIt7jZcX2LPd6bneZjpa4cLjRAtFb+7u4DJl3P0GyX7j9XOHnqMb/xfFCLV+4D/dM+T
do8TZ8jxwAJgczkYTDG5G+vA3vCl9DXNy/Lcv/sZ7ypGXNz/Ql1jtJuBihW/qicK/y+TyypQBQYy
AjWKtqa3c5Am8zSpXIttzxdifiKXsPiEM3BMKHFDoT95yM1+Ovm1m2w9DxFxkvT/IUX7LgXgJ/Bq
kE87IBRbAPeHONEfekJQiZJx4O0/1+NBlpM/d9GLfy1W2PSVbJttmKs0KAOzn1Sr03XncQPU/d3v
OgMHjH+PdAK46NOPSHnHubgQ19QkKoiQm24pCC3r6iqoAGZHtGkiVEWqQXW4qlwJ6i0AeZQaVJR7
01oLGNVN0Qj7kkN93NgWoJUaGzjpzj70X1q9egcFxkm3tK3Db1tp6Nl+kHoFzYq81A/jsqVaranV
13eJRonQ0kME11omGXFgMMsxhzJoaj1Gh0mtUJT9+fZwSxiN+YPOJWpWiP489HEdL4/K7pv9H0aX
WS2idHYjfawe4o40MuJVsSn+HBSXMuJjcStCbFzJ1VP7WX3fHv0GNqLZsSRMjIpbR7fOkuiVFVuk
/bXA+1V1rcR5Ohby17a9zg3UkwalAXOCI3VkYEZFYr02dAS+fGygHukxC+u1HPcHe7FcHP01/jHx
LG3dj7GeWt2cjAZIfn4Ku3OxXM1tiIzLwaO5JnK/98yoXXSx22/GJxqt/e/9g0J5+x22PVsSsnCq
xYWFPNFob07KTnnTSR0zGUbamu8BNDc6JKYuNAoVGQjomMm04mK7j2PaV3hx9dSt8ysDaIk0IlxQ
BFtfICO3PJ50IOUmHG7SNO2J42af+dIB2+BvcH2FPHXCB4Rk4XrpUJ+81PH3671cs+9CGfaYSMb+
OU+q+bsiQG7ZCLWH1hoTYd1o3hHZ53x8xMNh7Ix9zP7XmJ7NY45B5E41X9j5VS+ix/wRTUpk7Whi
QBayz5CaeAu5txDkMzFNyXqi5iGmK6RS4rxwHzPJE3mrrm8L91qrNupTlbNBvQq+LEOilQofaAPZ
loIwNlWGnBjmtdjtqwjNj4DFgpgFvnCDaIp3iVaOxz/Dj5ZEBz7c7yCm7+sDx0n44ns60wXIVAYM
KY49fR0vDaNUcooSVddLWsN0EdNxpKMHWGzn6nLkh5S4CQbWKLQAPzGlqwGWwIopokaSDG9CRlQz
lwQi/OEMgxkryhzbWS0Pvx3FBZk8nj64fvhum20+ARE72NSvX3XbCIGdA5xdkNwz73LNdpGrFrEM
m6xuEzDM4DsBOC9n0MCQTKF9W6yulB5U3rOuPK7h8GCVjWNJTfHDuFApdFQQYobz2kwubK9flVov
cxRxw6YLw/wbQPRQeyvoj12Fr1Eo3N0K9bJdBYtdEgtHB8MVb7AxTTW+MuCMCtyhljLPpDrGB9vr
U6jJMWYD2xekrG0yI2KPCFi/nBwicktp96gyP4WmW74RnR7IDxBCV09Ze//vPZFwYW2Ksu7jVO9C
n0u4BeTav30TS89KMH0VcE4f54nPnBFsxk/QG2UYQwa2ojoJshOn3JtYUqzdm+4xtmgmnepttekl
ril7MrV8oiTm+k+BdB1ySBHHHuyL4Cr7inYwxWaZjDL4gh9XFGhpiw4HAwy8weBjbphWuxwplpZH
6I5XRmXQzvhcciml5fw1hDWIVfjFPG13d4ux0tBSXy6HHtUtjKDAFx/UfU6FdY8uJmCgKFVsVFzS
RbgydBIGJgcPmD/0B+CDbrpOafNb31UZ9Jb6vZkCajXqJplTfzL2LSocVCvCfobYm7hB6cs8TFco
0nKF1BUnYQN/0K1gib/Hc0DCwk6LqZr814nSbLBkAaoNDeRAoybdXk1Mbk/gdu5TR+ObrP7nBQBX
0O9e5TRvAe7HvXXtRzbU6yGz18+DTmeR3lr4yfMhytJUChAWTpV4agTVskB7/1cRCiAgy4oGYA2q
Qpt/AEa2PrfuZDZSK7DmyOXA+Rjqt/t8SKxdZq4bYXiNVCinLR/v2xedfz4BKUTa1wcYB/ZLmMo5
fHqwIXdENHAdHwequwFBs/B96GycfjHPeocX5aKsH245TcbM0CuJzMRo8jBOKXOFQtTOb5uxtBFW
gighflH4bYVKsCZiRNLCiMn8r757Uq1yMa5U/7ZCzzAeYyUKc2vjb8NwB3VmjQ+MabADK41myNoc
JaCpkg/IvCpVj5ZQCJ+GZ8M00FZyehkr5cOBSeOdw6t1UBmaXLL70aMVTMRGY2ifFOctpZ0Zg/R1
qe5GxvEuHORdpLZQgMzi8Dx4bSLISNlThLTQeFBYCZunZIEOq9LOhpyPcBbhBDxNNucy0xcSidX+
ArDzlQpkDJS63yQhBaWTQh/hSfUljZeJKFHoX7VA5VhXrYXOYiTs4Vj6EMWe7nGNlktX5pzYhODe
XQ///kP14m3Am6zCRZ9AVzW79k4kbV4IZMC7byxSN8kpqTYrCoBJX+17NuAclklw5K/1s1GalLdd
xAAL8pnJWupQ6G7h8ZLX8x1MSIpBehbTZrb/vOxTlwVMSyi3mon8rpRAjzmaFJemFo05nM50ieel
hVDGrfz/ssEmJc5fC0HyPeI6SVgj2l0tFoOO22hfloGOqXuCF3vH2yscpbMyvU3UGpzvHgisqwgw
HBw173UGASoF9mwi/KerCY5yC9zbk4cny5cGFYGEcDDqA8MI2q03fd9jcIYauZ86lxUSZTPTxN5v
JzDWrj0QyTN6iK2yOHvWVXFK3vFlQpYv8963aV50AxvkciB/6YUhpsaJGWDHPA0aOb1vFScYrEwm
9njv5MxR9u5NomWuWfXMsLg/EuvAaT0pq43LE2a0I2+NyU89zpFNg3s38u+wq4qTwfhVwGMDuA5/
Y5X2Ra67Q3emIYj2mvJMFJOM/MQXGVtplojxUtVrD9UFFNAM1/NBIv2h2ptUZRiP66PJLKza+S9W
6OcRPM8UbCdXiMygGPUGN7lQqeUqKKuZ8Ta8kO2isZLCJbg1QoDBPVgBgcHHiIZ7UZwEnGb1BJY9
Vxi+rYDCv83uePlVD3/I/WOK51s+12TQXTaLvQNB8jI9+p9RvbHgsfo3iU1/oXaQ+QZKHoHCeKjS
6FeoXtKHd55Hr98LBUmM6WWCZS8aVL8Hx7XESwm9FBhxWGyHfF5C+RziqhO7am9BmRQZKzUrXY16
hqriTjZ4cXqkReVZjvxqGzS51dWAVc4f+BkqzD9fCmO4GxhIvGMnuBpCIQmNtryvzgeQKIjRUF7O
3DynBoVVAERhF/3s/ft1k71Ku2GtB1zlFTblwJw2NSA8XHmZcBvOB39Fu9CG9jl3RvFZddc529i7
4uzdwnVN+e48SCeRGqBszqurtmXoVVJ7OuPLaVpmV8jKmaN8fFu67mtRxLFbmq4+ffhshLTApgza
sTRKl8lwb7on2rvTIAFPMjO1O3HngW606Ap+qsCCLbq0+HYFqOMe5eVtcEvwoEJdzJbIlsxe+nyy
buPTtk02yTeh1Yzp8HIVWEI5Hck0BlxHf+fOHmbQ6MVAwVWsILf+94a1S0i6FL4e2Ne5DuoD6XTB
peSNxiARxUipVHhdb4JlemUl9v0grL0bT/qmZg6bsmWECn9czQ23usgKhvd0iB1YhF9c8LVnt15S
Lxqk5JOuiWfm0An/RTrZUbPraI43+B+3FFA+NYAXZMgGa8BxPyLIW0H119PaHJUCkD5gixBzDrbS
u7abki3OQyeQXgEeS5JG1LfzvPCZ2nwzbBqAr07QckuQXVOIraUMyxZUHunfH8UxOTewnFJMU3gW
VFoiJRvILWyguRCOTEHPZuu63uJz/h0++zTaTbm7sJTe3ydkAj20mhzf/rjZE0hylW76oESUov1T
jBMNqesjGaARRAkFLDQbiZFMuvRHZjr75reVkeq9auFcZID7uqwr+lSMXKAVPJVLQhQkMNP2X26o
wbn5hMu5goQsNELfvkdvbU1yw5NkK0cE1/tgdDbc2BbqlTkix35NY8H45JXYVzO0yg/tQ/tO60mO
1MFAKSr4QqNnLKXNhqT5xq4471OQiZiWaxd9/Yv/WNbVAINB6EcVkSQ62v/2QsFErbWhgZAkX2FA
tLDlJq2a3V0Hs74ZiCx2V3ejcZDWCU8/6Dzd+d9C6i7CD+tvTr4UaOkgaMsl62wO0oi3XRwzJ4Hr
DiQQz6w/1L4nlKnugQZwCSsZ5KGC9tFZbMcwvNNfpdop3GZSKBJECouN3FmOQkcdHhnYq6q2BAeV
05D85Akjqd6SC9EPDeEKmLYEQcWelnnNoaC99W3P9TpC0jQcva7ECzD0Ysnoe7WoV2xfD6CqA66d
T2dIS0TbaB6NIf4vQogKYcV7mBbfV0ZR/VOcSUbAHckMQQlp1ucM044YGcmO4UlyM8YRnxHKnYui
yBB9D6DLdqEe/YR0tiXn1Akoj98lKER7YY/wO+RxJwEjq4K4PLzwCcKn8AJsSefpN5oVokk0b+ZQ
BB2DKzQZBBquwEjZjLHSb/4HeKJUlXWiFXE1e1Gp/TINF/bdz9KguRhzuktUB0CvPGQYrR0bQSqC
+OWker3gpioB2pn5lmHXfqSw2b7TkxUz7LWlHJSXglGJxQd+CGxgWMzcQ3dOrSFmhAc2/76V5Foa
NhRVu8HVuBhIPI6gdGCuZE/OB2VO7pK08ZskBxZaLW2mETnilmiOYFFoL6eh+imgOSI08E/fYGuf
MOV2n17dhtIBdLtDN987D2TRNwMjfP2eh1CNm3BQXjB7xaPnfr3e8vDGOlhQQlBiT+S/awV0XYDB
xinmD86YD/tK83JeS1m6m2BTILqjcS5ZSsBEF2ymvaQQe71NViMrwXhABT+GYvAnpkz+XHsf8TjW
eQ/T6jGe6Ez4O/oGWJfpxNlbjJpHztGFJy4iSecFCi50tsCoB4DrI/SY3X/3Kxf1gdvfHJ4gQ3kC
YITp8R8lmyDbihE30QzKDqZ5u2fd/C2jAHbmpHoolU1Epn9QoKcz0h2gKMJwPdbIqFswRm6Caw0n
3Mjpz8hve+EzCAvrHLECLDwmAbNXTvZIRc6JXtLKzO58mvPIvSZzw56VsNxPm/pyxKVeg7sR7WWh
3rVU/SUMSyWQqrcwISJVqSru3kbR6SIlplMuPnqSD3hlMoZtKjF7yN4JaEWq63gydGpvxwZ12cHo
CCkih5anD8CbFQhtoh+2VjkAhaPYV0n2q1qjpvL9T5HUR86lEMU2/iyHj4flvwQPNiq1uX7VPk6K
0zedKRY+VOw2c+PFGV+OVPp8LWLUC74ovybh6sjR0KWDHO5M/Qx+C5g/X3EHOWOuDzZwx+DWTiab
e1BzusqLHVCOgtlJlYl5e6OJXroBEWy7p5Spw/tvjeAa9AhXX+MPg5OSHc8cAxobFIG5fG+sSX0E
il6aQnM+opLZqN5PB7dT7tAVtH33WT5UuNCfWglKRX0e1PQYxNHXoGqOqVhY8khT8KWo0UJ+RByP
5ieGE5bKzJK2OqNJb1cHmT2Jy+RmsL+yYpD79Upu9AsDeoT4i1LmFJApyIU1wnDlzZS1xln0BI2H
QOPLR4MbsVaOdjsI8d52JCg8jrCEcFwzcnhzcwqM0YPlmPwQd8OzZA1kWis29nh3o8K3ex+sGggP
PuOCMk+HInQ98QRHg+/8w1isP9yMjs816stWKkwdHyeFOlzSwv6XyJ0a9wr+Seg30w1DSsYXrIi+
9lOtU+kIdBhiP5aa7hYMmqMWznI0x5Iz+oU320HK/i5CzOOBVKEcUnZyDiXhluxs1yGn4i3chTQq
+IcCBQ+l3S1JxBdfDra+u+JFS0FMy8iio7YUXwjuroDLq0vM3WzMNZom7f88xKnrgJe0Vwhu+S3Z
P/kEgj4BUwooDfB35WuTuYyvtsbE25ic951MpRlzNZwHExVf9Dn0D4o5rYtixjjawnQ1SnkKSDhi
2CfD2xK++vJoJ/mxEXlI8PuqznMDxsgx6XrT007tAH6EjKtjhDUqLzUtSF93dz4LSXy+XrLZOoL5
/sXcBtPnfitj+KKRH1QeNcElKK4e/xIVT6i5vdwjKxkzJCkYDvoMHRldLUOcswo2UwYlW1hyX91U
14LUICt/+CvAZTQJQJ+8CgsOIrWrlN9LZTp6p+VEYFiH1WT0meSd9ds1Y38P5Zhcoq8O+cTmVAGC
aG15San2rFeB+mIBwqVodyR9bkputrbbLm9tzFbp4aDQ1wNVKXsR7Der6R6/BbPvDIJWV+LuEBAG
MTXdC50N2pEg7aeB31xBCwunoqA++j6d5wpEUKcMF0ljheRWkPQTOinuDRPp/FZTiJ5CYlNiR9uh
TAcxYHM3P2Ok8nAre1T8PgyFYMFt828JQn3+ZDSDq0PXrvXOWQrU9LyFyTHLwfpl3rYb4eyiDcWI
IAn45vWBtqByBRadeRF3dZuL+sCPi9OLLZRb0DQIPdBFZqCoJk4D/kC4FMuPJSM4DJllXCIMb09i
sYGrgtSV8QO8FLjJkxAHyiBJCM8osT5ZYX8nwFfwbUx00q3Lr/FeThHVVndjbFZNndDibYfBSiXi
qkLKl/9cm4MJszYGm5hwSvspJ2Wo5XMp3xagKy0OYjlXrlQojlCky2voD2GUAKWNpTrpu7QV13bj
YCivuK/FS/NAonv3cYceN3u5aors2SpBLayXyA0/vj0nPET5iSU8fIPaBdnwkwh45jXFw82ldBni
GwQuyeBXGHdRyUe1+WyG64L2x24d3iSkJ4Z6A9w7YTwnS3l9NlnM3iBbOn9XEbRMFlnas3lYTTda
EaArhOgLKf7QD4VkPtJwgh7IN6zo/kXZ/uLmQVPZEdnY93BeDQ06JUpTEyUMZA3s6qAT76+ovdd1
MA3BqMekPUdRJtme2lC8xqIVlQVhd0z7dl4tR0/qWkpl6n/Soaqo+ulI+jl16K2hm7esfRZmtKb8
TFIacY3jr0Edo3quSVbQqii4ycGCmoJNcLycvwXKBrCv9miRXgOQEB4GTnEtdbFfLmnpv7h6FGHS
crZmhgHMO6aIiRn9W5R0Q9UX4P6MET3D7UkjtFpogiWbE6ehl4CuErWCDX+82ShzvxKj2l0VKP20
O/+A4f210swKS/IIN5d3JyZGOp9Lz8xQLNz62vnaFDtImhZ8S2f2OXm+GuJWp6U9TuJtwUf/j3kM
5Moezg==
`pragma protect end_protected
