// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:57 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A27/K3IdH9eP4f0ky1Mw2DLk4QffCa8kVQObnLEP9cAufv5N5/w+/z8pr/b4CNZu
8dnvunpoQcX8Gjxb43xC1VOth7/zlw4CtcK6lyNKD9CpANQQgly43CWbkVz8yMy5
8q3fmk65vq2xSdmniMzY/yWRSpFqrokRw5v66bqaKs8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9792)
UZJ7x/1taDqsT5gx9UooZgyMt0bqzBqrmp5BWTQT/LoHOKhpkSDDaCxd/W3H6m0L
Nj7XNAfxEIUGnvtoqt4ETBZ0A8c4F2uR8sWyvc1odGd/JBy0S39bSOz7rj473c8P
3LZxNab54SfKobuNF0XtdgLwxTba6A24Meux0ZlasvvcUyu8Ck54DM7dPE5bsana
IsgjWX7cN6QjIgeqLikul/yin3mHkES2A6/bZr55eJNz7SfyXbTG2DgQ3mg8aloZ
gF9BXsRxbbDMou87GBZrye3BgpssUNLnM+GNFHevOzvYpIrKw/g0PVhiAVFHV79M
0VxeOGa9Wo3UiiBYix2f2kmmyNNdQ2G2Nch/ShU6ldAcYDqzsEmsbJm8EcBe5a6j
trr/trSknv5AYpNEu+IkLU6PYQKMAfOVANlRCqmtt9IB3W1ihtA0E32Bs0Y6UmUw
9pklTuTFX7X52lx0WlZZgCR5/hGz2uPVEdjvjjwtZDGj1NHK/3VxY57rrPHmAbHn
c+ccl81otrYj+euY4Z8KoN6Y+ol+D2qOpSTyJz3Ggk5Er2AL8qjStI8L9uwrCcuU
FgQ6pQ5m2W5EQeKlktfwZ8j5d2Tn6vkPGOG3/DH7IzFpLHQ/AvoZ9n3fiXfetwmp
1NO2OVrR4FqpgRhwDU4oHVJaqyvQqXJgW4sbaWP/U6VapqYiMzBpMGX5Sgw+gSFZ
PaaeZi6vmZIZPFq4f6bqtYRK4jK/z7TBQByeQ+ZqWOks3GJty+g2cqRASXueFve/
s5dDs2tlJdJF+AnKzqOzhKjFwM8ePM5CGVXlakxd6cbR0HS5nYCfm4tqWA8LZzZo
dySM+EieFGGAnv8PWm+motr1dZ4gO5DVI2WmKZacJte/mxgXo8oc6B6LS3nLtu/m
MjeHS2qFeVnme9gvf/iwtvi/AGirqB/1rBcbnk1zQ0iS/z/oivl6ewrPPttD+X0z
e4TbKlhmxfyoasI7yLP8cfC2zMGghg+44JSRroUwib1kp7QS13h9HLeDcbbrXFn0
S2UIIK91slZGcdjunHFzHUZfzi8m6WHDqkogpx9M/q6rvTsoxJzdZ9f9hknWt5CB
Rtb1RNbwzizg2nLz4o/vHKgQa3icAeMY+7gzHnzKS6LDbOl9rHSyxjRAxWeNV5ph
Wu1VDWQIFzItsojMnCBh2AkrHQgjP5qH/nFg4W88iyJZf5kLjzP3H43A9uj2Ltlg
X40uPBtAfkntoWsf96V9l1uG2m3Tl0Kp99I/GnM+UPZvZbwre55EszycXHl1cwl+
23u1TO90sjWvGbF86UQMqF2sNgZnyd/DcBBIHiSjGdMKVS0Hiz/gnAMGtJFUWSPR
y+athrpYOfaYoWZTO/AixrCo/Y12QTBYG8bgCBcbMhRq/Ia9KaCKQQHNd6F2oTaa
z/TvPg9DTfyBvK1870VjUzCEmqmWgToqLctYNw9xccfCjbodSJCmIxHS75oHIodO
B3fEf+rHj7yEHMgptlzZS7RnNJpWRN6FEBB0DcuzfIpbuxu7rxeXCyXW6+VJj7a0
j8jEcCJJB5Mgs/B52/IMllIQjojp684+hDQ4MOx3ZTzynPMF/NKvJCWV1rFMInes
fFMrXbgVGzTKY5j5O17mmby8gktmBTedSO3RVqRPJbS1Gv5XhB7z6yIZAaP77jBl
cQq7xdInltJSsqFi6Fhp0ducMJI0cNAl/CxVc/DyjnGzCC0sNpQFmL0OEQvnyjog
q0eWgsl6h8JblZR8ewqD2dhEkjysEkgOBC88c6ySD0pryKw/tSqKTCoDFQahcvwF
XWmclsMbxlekqCF59tztmS7zGLHLoCSiPwtqJyNXT+39/ymhLsavCY6KNxNPQVuL
5UeUiXUm8i8nmuwJy2Of+GHxZrfbwDp8ea8Z33/90kJZSpIZ20iRAbhh8Khrec4i
SlyGf4VDLYEfgVGDt+KNe8139YO6uzdSV+fuQEIIRIPhKdjtY4Bd+1AlsQFBjBpz
xuBy2Wor8Z/H46jz7cjQBFNnKJ3kqjV9OoTbNbF0VJpx6gFHHIh1ioBULNhYne7A
TArVOt2iHoK1WvT5gaicKYwbKePZP3isq4vs8Sb0efnyQg+RVufgmD9JeGm+l7oa
knglDEtoga2UyBZaT8fZfeCg/WMDNdrAqt4KGXDru6ZlY4FZNTXczcWUz+Kl6PFk
3U3TCW5U1+kaHav5xk7dcfBP57U+NgTQxNFtbxz2sHnKPMC6c496zgXHyAYRJKhX
vfZIPv4ZunF9SwyZ7OlrMCnfq2ENuJopMcLXLTZ98DB4TyexIzzEWI/Fg2yePWGB
eHL2fecYzV6C4VQrQTmDH1DSgsTI/em7oG7oafLUvfUUxd1a63TuFodq8SiBJjZ2
/7TLdo3E4UCopz1xuEoCefhYkbSnwgZxx1WXJp07isJgqUCtHF+fXV5l3StCtGRs
n7YhVThrDGYk67wXMPckJYlNFYaIoRK0E1BelwPK46E7uq5qqPxfPbbiYEdI4RYB
Ni3T/rMe9R7Bnp62NJLLqPkKgIxUYbYxpnOaLf/dQWXlzhTgz+AxjZYCSnoI3Ky+
X/faUHGw3yM9kz5FC2mHjj2OAuFEx0+rix/x9eG4nmTeD2a/RYiiLzrze5nqbsKu
EAE+vNbOC+lEUWF2Cxu9DxXaBAtuSCW+KNgrWosoWZLh7+/rCuTF2GiP0hf+674a
Q6Y9k3KN5YzCe1WbK2AS68Hq84O1dghopHJd0VyVXHeUxZqELa0W4iFcCVr5YtIv
SLel2+eAN7aZ37ngcnx8O6s4kd+FptO8Vf0k8V9nBH1R91micdQTxh0hVq/AsefY
VNiejiRKwhUUQ5yqDSaFxCcdVCxdSIzH5i1r7hGuZhgfC7qjEFSGJyFDJQ2fNeYZ
QvFxdZXaWx/GV3+0BQTNFwgvocjQX6cpB9R1ULyJV2ghGeYicTLZ/VanGPTtAiZz
0sVcGiP++vrtelBwspTTHHqgje4unaxeDzvqdzXvINnborDyPt2fx0TdXGiRyH1k
nVvGusz+v9EG00sEDIiW0UPsrE3Jj2LWrK7PJdXgIYriSQ/99GlkHdVhfJcZ/r3j
+ZsODX5W+xaUn45XtCMnEM+XHmnewcRDG4/iuTtIZfccwjPPdr0kWehr7ivDGnhM
dTbqEZu5fbPw8aUPH3irCO0/k38tZXAM58ETsNt2d11QgMHDUad8r/afvOmweBSu
ScD3s5QcAYw/3YrPIG1V7jamo4ceZ420RGDUPWrISNuGEvumtbh8Eju3WlEFRtFm
a/tBXkwbEa/fzaXg0sSLbtjwJvnkus3ZHa5mdRbC+cPcHqoASXpK2ks8bvRwYZxi
I6N1Ay63B1uZM4onegusE3hkPDM9kr5bZNAwhy/6rcfV0IeZSRNCVneWsxqDWohL
SvqS9eG4hlQMQaP+80AKwaIBeF/mWHqFlb72sqtYusqD8NhtYGFlOP+7U2n9Gm89
FhWxS1u+papi/vosZfr7u8MU0/7g+gwLJuIUJDykK3tvwwVMXM9Bvm9FJtXiUB+4
cSVIEnKHttgoBEMsCbCEFF08nZ86pAf6UogDc11Vn4sKwi1g/JP6tJmo2/fkDCvF
V5c9wG/vOkWIQrfmLJ29B4gwvuvxFoP7SUDO2v1OB2yXCX8MyA09xTDqcqGAIYIz
hW6/7xaIR36l24dxttQLiEBUNzRGquDCHIje99DFZRAA3/mffTi+coP4/lthDMYw
QypPbMPcadDUfnyGvPJkkkKyEu6aIx7g5u+N4KYaoY7YhtwD4AKOOJL8bToK0d3e
4wYtAbnJSuwa303j0A03heYX0qccKBdN4FhVAKMOphMr6N0AuT6L6QrpAW1ztVd5
6uiLmJtxu39ZWbZpyqt8t3FxhuUfYtrdhWmdAGvQvAFJvojYQ33ZaKBUU3X77tXY
dnSy35g245g/U+8txv89FZe5sU8aGi7o58Ha2e/nL9vs7RNMCNIcy3s3BRs4YcCE
sM2L5rZWs558w2isP1Ewwyw8P6ye/apNN1i10RFQK54Oa+UBb8iFyjbmAMwhzLpk
HfcDc3Uhz9eSfQBf4OuEwwGhTYvAE2KAgxONYUbIzR2FpfjUZuf7EJpTTdQoEvBi
HIpd7EU2b8ncFHlPaT4W4Lh2VcepN4oBhWVE1H2XE3Mmbo1f6/3RiwcMSuz4mU0+
iJUyR7yt+mLR9dSpGOYn2XwWALfukmF7FtDqqyq7qjO0VgF1WKZplBvGqAQdP0ff
oS7tqJXT4SuS7+pT1ZmjIhDCqPPKZIAhOqDU0NEVJqt6BqcWE45Zw0ExY00adR2p
PMxK6CKxyHT1IthEUYsTBlBp3J2yNNuHZ85c5NdplOsz9Mzz1MuhpZx4BivytHRa
7Vw77xoiYKzxugTrfXdI21Z6/9UQtBybyWQcbbEp6g03RZrQmKc1LStMnqxT8QKT
rzCoX8S0ZHog+jV0b5sbNrUXSBTCjE5rDfGB0KeRGL4AoAO1Iaw3Bjb8offisR75
mGINQtqw51q9FOYordiKmxnHpNUF8y/1Qnlr+kc8N9vFbsXhjDmYCF6yUdoEdcNm
XZvpNTQP+GwhBzawNS6TB6VphAytdGGU2F0XmyC6grAPCRQlmG++wG7ZQlLU54DX
apRbm7OIoO/01YZu36Lk8ykS1kORLeHMAqBciBjj2t5bWUnqKrQNu0xPYRJVUsfx
fCbyfyt5ETHu0UdHn+kEO8EaZB122DbSanTpZ7QXB3PrpO2um0vLHxUB0j18ttqV
9jixXpaNKM6Upi2EiK7M/VvqcZzxKUdfP4NHldK/ZqRT/S2FFn+Qsbzv9rwnWPvG
+UV2bedj6gpYiLxG8Bm+Uvlh/A9xBwJa2B95QUrTW3KpniCJmKuWra6ml9G8dADu
31xp4nNi192KgVmXZAPwv038RFpXmPZHu4g1BFwVtDAJQ272XaryPAKsVljSUB49
pN0R4G9bzCKGpZqY6hC2laHQAVrN5qjfN41XcjKbxZFIOLhSuoKgV9WjYSQD2TCl
EexEMcPUBBSknzW9ObbVeGFnYIMlfrTYUeJoKLiiDdrwlKRE+Gp/FKiXKBkuXLc9
QL4F1Toz+ITm3elIXM5mFDkQ878vwc2lg0eaXUHmrVV/76rCJHwL/Hh0qIjwlhUO
GCABbRgrp2HMhSufnFyK/q17sgvfMt0qrpXYQI++aAaVN4Kzx/sw6rH6mej0kbWq
/7gVxzpjJCGwqi7LaA8GzV0oOdQLpNAOcrOLv6FzGPbGBE5ocIqaPnSbMP/NCPhX
x4eJdMGttYhZvMyucWKKyqqYzlutCDskxJdlOy5N1SYnb5AsUDNlTEGqUdhbVWQ2
koj/ARTPLB3PyBjNvt7QFzTMO53dBsAH7xWvzENWAaOEZEK2eWqyuHewm9Elc1CP
7fwMdM2wRiliUvTlH1RgtWxQAwBs4uAgRt081kQX72PiT9dGU+IFftOtRhB6eYmu
X1o6oKdnUT9KJDSZlRnXG4AftzWyaTsQ6TcjjRpWXMlZ5ReMoTVE5oBT6IA8ri1O
Bmx4KaLxDehSGrDich82ryLyokG22UcciLSzxpQaM/OKb3OEuE2wHg3ouN2dkzf6
UVt4HFPHNqWi9SDZ9vQjniaecudLgjEte58F/n1Rp/oerrtwtyfyTutRfDpyTfl8
YaR/EKAJjicIn0trIZX6x953Kq7ICCBkavDX6fXslpg5p9Wi87ddtqDKcW5FgLEc
RY/pedgnTdvvwN3f4L74b+wbjCc/F7Fh97qe0rIWSKqypdSbhOsSERah0ccYjhhH
pl6rDuwMtz/Qr1UXkwo4Z2CCjSLGFo5POVPDEAgwAQ6IkQTq/Kk+L4GQeipPqBVl
TB8RLE2Qd578p/B8gssRn00FTfiNAOLKj9eQya2eBwdo9TaQYgRSgr2Bxg3/EEmI
iBJfB3Z2cCBcsxVGegP1lzOg8Un5mq4nTufsot2LVHF6Kk17LoZY/BBOrapmIhCj
GQKIX1cdznJZG9wpB13MWr98WkPkad8lI0Cx8Ibb/FueTRr0o0+mi+wYez8dwUtU
sfq9knQn2ACdsOEEnMgatJFGdV5rsFGNW0EAHrnvGdzTjs4+sFzOsLZWCOLgah7K
fE0Mm9ODDEf3TJ7CEiwTQbaxiN3GQYy1yoCyDfGl0luD34G99kwul9aZHK1bicl5
yKyjaFlspNwQzLyyqh5AuHamyMByaM/iVZI7QrhuaHXmLmMduz/yD0GBrguavBC0
QN4D8SJcyOfWjm6ao9kAWhxAMcYHxUyD0IiAtLX+MCojI5IfCqBUWKRY45JuCjzQ
mbtSLUpJGlIPUcM7CFqDvm21krSYRFpdHOuRRR59AtCHHzgWMybvsKNyiQllnOfm
Po/agMAANYmLUmZgxcSOc7rbv5jvNZMjgKfTi05ZiZUSuWSNmRbwOOtINVMjI+k4
5pGEAcT1YZ5QzGWUhYlNvkFfZS/WEgv39gGxnzL/xnWVouW8WNomYGeffqQshxDF
3B6E+wxX1qAQwaL06tcBRfKDFJPa0isjdVc3BbiQwT+r9jTUhRfiRuU9oGXEWUUs
GqtkytfXdgd7Qg1sM1LKJce77qTOyLE4g+b+Io/lRWhMOkxDrYqIg98aPbcP6eoI
ooipqFv7UsrxjRPqNqLdXbQzJYujE7gypFEx6U0KQEoPgSSbq44novUMkJIQ4Erc
e3v/lS+N5qkfh7CilfjoRXsBR8Ywu149eSj67JPCI5UayabWNPn6f+yora+/Nwdu
YZNL6cadTJrra1ekJmDntsnMSbvwTWDDA3+zhzEiJDVazoXDcWa0YpjikgR4RJVl
wwccAUIPZccE8pMFUVUNoX1EscLPUUHNgbanqFMeSGdDeJJdu/H1jx+AnAkxv7Zs
5FLhD0aarRzsq4ItaubCUtriRjvK16+f1KvPRpHg6PK8OEE/jPE8A/0EiHUJjEW0
eKqbTR+N05m8ebPbQQ2dWDcEDKWwrohajYhdoNZXw9xgHV8xLWchEP7czOVrIjA8
/otf9wqqtAlT+jKz75z10Ao0lo0ocp48btV9bVUMCiIONB/o0HDK2pbikB6J+/8U
3vDUBR2CoLmJ6c5DElFGdHGEAatX8iSQ124oHTB6xu6+9LNd4J9B4bL9XCN1xHxH
sn0RjiQNuWG6QpWDqqdFReBQsYxZGSPM50h/uj3nVd+18mxpP5AdRUaMOjPHzqhl
X08HkZW6p8vntF5Io02n3MmhikqfwYLoQFZPFktD+ulEaNAY3DZcG7OBXuFO9Rk4
v1eltXNEdwTp17CnXpQvzfArnSSdmtrUJM+mANsfsrZqbeFpVZDZ4osT5Rc6w329
YVvKXHkAw9oJ0LEYfw5ngYux2Z+Vf4LNGKbpMqNRZwzUeG3/9hcyMWLsGerOB2dN
SOqjpdkGbADSGlAg1rxJxg1cC6zBdMivGnddu1JTxb3dCHa5W2F1IAF/5auzOHyY
Ar2xJGGfV/P3b+71IKbVaqX9Act3EdW2sdyI6ujXT2kLoV1bE967JdK/m9m3riZX
MfnT1+bOv0MTAEhoBPI+ZYN1wFmDm+/M3q2nWtnLjOCwUsX7TVPAYYSOQvmjXiLT
cU4Nl51l/AtR3XlS5II9PFkTGh1vx8d8aGId5UyDcVoFEBa8+3ydDvgBRK8wdeVt
AOwL09D7jqhdw/OV7TnifZmSraek8ojRRHomtPySNcqNFsqYCG6DFr+B8SP7a8Uu
XWYPTCdQfem1TBZ3boQNfLBZOxCGu/Gm3gCBRY+8O2CxufpXOzKCcNkT+MXauITz
D+XsjNu9AAsREMg8wgt47a/CAs6yMTmwWOaNKHmDIH+qL+lVEe4gS6UadZSsRc+C
J7ZPRpoCe7S9rfw35E96ua2moq5u2ampoHybkyBDW7bGJwfg5vy081Tt4xNxFBqF
A0K4md7Sap+ohNVbazVsfatDq/zSHSudx2lBXdbfl1T42AFF3qa2Mah4ZF9eGkOQ
N8zBndoaIveIJnMaTSLYHcAgDvVePBUD71UykteEgAJRX6wmjsCgAgRR3hcYy06F
wNn5G23Mvhvk1HrHQgCXoYOIlnC726UH5+uzMmsP4y5qDyVG7FTZYp9eloEMPkHG
O+pBn7YimnrUId0J1kCYy121Y23lnuZnn0PAi7A5OjVo78Z92WQ1/9MWWUsNV2nh
YMP9kg5c7DTHhVj6ObyGcjlTPMU67ZYKZDcJIh992TLaEevAGS6lBohQknV3bvfQ
SXO1fOPcElEKTo0eX4Q7KBrpsYwkgkETS257SF2J/oTQght7XXSywUtDyy5IgR0v
0BUOCsoUgre5RhX3f3ngcESrkn7MJ7cpygYjFIZduCwuV679nA1L2rqkh1OQ+MHp
iiNgfSguXj3+NK7hWCqjoAQP0tG8pVkYTXRfWY8ksP5ey+icrEmLQIhEkNfHHWVR
N83X/q/qrPnl+Ro0rN/kupcl7ng8GjJT4CdJuqW/DPN2CB3Xz3Z6LMtr1qaKSALH
44EtRyFzX2qwHdtDhy/qSI0IZH3bQ43MDtI/pgbtoT0BkRssHQ9rmYuzIC6d5fT1
7Qhb2xwIDTA+0OmNL+XcxE29P7Xma743EF3anS4+M2Fr65Z6w5lipeYxmxLKgQry
pZzPW6jKU/qZhxh7dgochyHq7mVrwpPLFpndTs0MzOlkXg/Nb19oRrWFuqUZMAH/
b4zVgI/IknPmdNfltuNHpqaz7cJCZx45gvo1Snx+dIBldbRWd5FwUZeRmcXlhPWU
SzTLZjYkK+kLZpq1jyju+ELEJKe3K8Hnn+NT6fa6m0iOkry9iha0x37rZZxEf1jb
Uq6t88HbiTKyMQVrBvafy7+GmjetL8rFmpotpJBasQDw4Oo+vaKi/PVaRuSH+9Nk
HCqirI2APWMFtGnIImbr1CL5nS9h9QsG4OpeQk5/8UoqrLuijDtxcsGIjYtAFGu9
WeHMXFj4dSHqX5mXQ1vvUe4N5vDwP8hIv2VLEQ1iPIgWU58azd24avcJECNTliLx
ZDW7J3QvjyVdoFTB9u/Ht61wAd4D+JGTvRqzips5Ft/R2DK6CxxKidb/5O2JeGl7
7dk1DtHlRgX6waFKHnfFQc9l/i0IwLoWgkaXmFxboaXqEUyjPHZ2I9AEAPS6w//e
GffV6ha724/bNyq4zRDDC8RX+fuS8p6Cjd5zfXrKw0bsQXnTVe9Y66zVpXyudWkg
PTLYqHRKTwX34VeUoGujJXs3AUxhUbWUJhIYPymTJrfsOdL4wdu9kADt9BzHbA1H
KTNsj3rW4Hwmn2nh/7S8RRTt7pDgdGvvISmYoqKI6Iqn/z81JKvTTI7eUPk6wusq
l+kN7+Bk5Yrca8MPuhYLp21jeNGDiL+ITpyDGFdLhfXzg7WF4hfa2pRmRdcL2k9K
7H5mQAMjU5RCkQrwrB85/q2x+RxJS+TtuwhS5ezgQ40pO4vLMOVxn1xVkM/TbWUW
iV+/wZRNIhsfbMcYP7zuzmt7SstNipt2BFN6868d8S4CW2fzxqNsrvOuIrktc1TP
9J+HRs4HLywsWU+k/uM/lgz1/Ne2nxtzHGNn114qGCLB5Od/XTHnhvJ2z7D8RMAD
Uvy05f7/d+KrP5Aq0LVC2pKhd4JxfRk7cvx4sFC4eViJIv+CXiXh5DE16dRYPRg3
tTRy7tRtkfNagpE9ye0SCtDxQbiSmvRStivVwfneKXSx8n6lNMFtvDt/sREpjE/Q
jGe+9rieDh2nni5jSMYBqwPkxeC3Tl5j8weALNTgC5QzqIjNxEW+/5tGC5Mr0co7
qgAAwluojgb1ddzjprkjZ8TTwseZYhPIaU8Vque8m50hvyR4mb6DFHYVtJTLxQDB
nBYsm8nePqF2oJrDki7aodc0zQq/0uZCySgPCOM90l9r7i71q2uDdA/wRyD0IkPV
kEMTsQwJSLZTkc3zFGHUeFVinOQK249TV0rep7Q/UefpUei1bVirsYtyIl9zbbps
NHSRrQCO2QSHbJdj8rso4VBiL86qralueEDWRqt7YCM+PETZu2/ixQmNUmWI2oEp
jCr7yRfwg+yCbK7p5g6Ze+HLCpYc9h6WgloY+hM65juvf7DBhsrjKF24WayPXJje
Jz+hUxlbc0YdJwE+CSkhL2BXOpqLT37XGZPST0UQmoR1yHRNmXJZWOP5Wsx9sxh1
sIPFjTGCk13UvPVVqyL8JJEpeUqahzOJMsYknmMgo8mcdir7bTs85UCwFTxtHASr
z430mNU3Q/pQ7pMvW/gs29U1sW1iGuz9qK2lAvQSwZdYTqGIVbp7pVDdGXTYvPrn
n2poXtrZ8DpiiuUOIFhNgzg/Tc0IV0OGXJApoGR22tuOeb+RGEj4OoqgC5JVlkt3
wV4eVjtAmaDapv6ZrIR9BfW1COkdE8Am5hYYeJ6pZugUgjjR6RD98CTDe6r8cb5O
/Bcc+NmLd+C8wZIHsAoySPB6FPpb5BeT4cKvDET09j+jINy6MMb6jq5wh17iDgGR
zYq4SkIe3PqvQdib/GKqeYX6dwmth6iL9jjxfnrxdYxc/zOPYPSO7QzB0wL+0aJY
0bdl3ye/932h57pKBtkZVoB9gGPaRz6nUsoDpKQTOXwGtfHKhTwjd1r1ZcJ5vvQe
+3kRaL69lMaXXO0fEGBDphBFeLlQkNbQZ0llAYCBO6WKKcf+1g1wa3InusWfXZDU
E03Ey6vq3rrhBBGWP37ISf9TQeIu14V0O0tnl/PsSF8QA0DXiPKPVQCBiczyDjaC
ygRQPD+HaKdHgWqvOF+b+QP2qmtb17JOZnxzuGeAsZgZVaCch9MK0ZVCbrPha60X
mu9Uh+FCSfofEou1b0FLS+4ii1lG59Ja3mkN7sbq8d0WNLqKsAlD4Mw5djQPSAhZ
cc7lFni0nRNGe8ZA8MI7Q8rHxzzHNnxZQE4/7wJctxFCy7ZdHmyx8MEVq9Z90NpU
2J6V818aoXi1a2krjFehq+IEZKedPbdX3451tIJhcKEn33nNUukjPtM8rMhpi6jB
a1O4a1n7f8/7jRHxqxnqOUqrnzztmx4UqcyLqlCNMbYFtoaDoCongRKKSF2aKxYN
B5AceiHyJaByxv/clansYEKD4qFu334EHKpoIDFbKZ1SMYd4z13u4ZFiB/SdOI0y
APEkok+eu+tZkj2fZpOhjoSUntbJBgWgssGsPpMMmGM+CZGbY2XZM2aAe8uKBZy2
6kYsSbzlMSPJw5Ah8l8xAV+bfv6Ze0xNTXZnJV62DJLKnQ8wM/rQ8Ups5+dqURUP
xXc2AUjhxGnaP7dBs16Du3MefPW1TgyJGm27E38+mvWcfuIOHWDho7rFlW5ZvlDL
drjUY6ASdSAE4KQP9zXOyIw7oufTNKJJdMPaBOzdcdmKjpTkf00J9LTEYyt6gUuf
kfJhx0Djh26DaHL/hmO5VR8hTXVw+WqpLZ0pFSf2+b+yON7Vl5EAIWYPt8j6bnYj
xe/FVCjzGTvPSTNZQyYVwYDQn1Xti0JWXFec8Y3/r3gotfjh4sKBEiHlW/IrbSi3
Bg+zi2BiRRWUI5N2rwr/taQlbOSc0obLlcoCHAe4+B/iSlBBl4xLeapxAcaqeRUW
4XyCyRr51rSNXr7mJ/bBFDxLjCuYU9Jurbxv/IR5ANyjTzEgrYBr/N7CY4uucJNW
gP5HLItnA6p8LvtGEbJoFWHlhA4i3g/U/VRU0Z93ASV74DbKTS+H2IyR78Ni/BYk
MZOkh0NKylhPsUF/AEkUM3GhTzhT1cVNelFwOmd2s9yT6VU0OKm8jr/fqzP9fVov
GprvgiIMhgruLIXch+GyN0Xke4b2VSrpxIx4kbEkvQ+xE6GgaYvG+hk35Iso+NM/
FOdseqpCcMijlLHhMDhmschLZ8taA6ZNEcHz01JDN84aWnxPQKHvbrFAZ4aZoR+p
MDattBMd8urD5k08ewPuHYXIW8iR1xb9DAleQUOucl+qJJBOtufjeGXIdJg3zxRH
qbABtYlsaIXg8MTorySQb5ug8g6q+xL2cyLX4cJoNSVcpHrTbEdrdBPjElgrEjG3
nNs/40sDNlODIlxy1YmIlHznWzVvL0AXxpLiVa3TtdOHQzofc+AxwUg5nHqH2zLP
pQ4m5ETn3t0HhjRI6rl7GJLV5SYy3MOyBS9osFpPFOBT1OB+7qgM+mfCFpAlBRLC
ecoc3DTfaQE4JzO2LAtnKA3fLZ8HGdKQUR7gLScyv36LKa4E7WmWX2iPPyd6H4kO
sOGnz3oyzA3hq78R80lzlc4Vzkc+Mur4Ud69bcIkmrO2smtLgqv0jSKlLQjYzfmf
fxAlyVKJpouraRm8LTHZhmTV29k2fH97lGXpf+Zg3+k5z5IpjSXDFMa0j3MBjnR2
7b4vg65KfjC0UNOLohC5o9QXl9suw3bJJx3okL6xIUyr0+lYTWtQNIzG7aZU+r8T
ZmQT9uyTe91VBSXQJGTZci12wQvKpBDWfv6qFBLfGwnLyv/u9VMlzPT1rx87k/8M
s2OB/dEzYqMqw2+CNraDHg07F7zGKkcrfb7rfBzcudYv6XcKPoAgZM8aRyDh1ZhQ
p6L20NzyPn0yPA9KfKo7knU6KcOl06jH+MX6YTnRBw9W7KSyhNGH7XthpQQLxr5m
gBywoM7+oohk1q+2PU4nBhL2ZuXZw/yOuBGxvvpBU7HeQDUPAXL7KQONMHsvYWRN
BkYEa1y5BA4jx0B4tFD8qImG2UdHqVYd6M961Jfj/Y0+uO3DrvtGxDxneZxzwTWM
B8digbUlsUgsOlNIBtLEAiX1hR8k5mNN8FD5otnnZ4V/+e7EFC7QykCUiKeZn3pZ
5Iy0sxvTIITi9F4vGtIFrh3M5nRJrQDoM5LQ3N4fXTtP9eTTUvG2ISgEL0ihi88u
vPcI+sCIKsDSb8Cpd8xZjI3/VibHcJ+hbK/WBZYW2vtVRFFVeZTixk8gcvHI9Gqq
6SvvKbfIrnE6PWWv6425XIphelfivFF8tIiP2VPybt6QSjGWDaZh21reriBsgOZ1
BLULi8f9VpgHuwsEMwam7cnhXUoOX2V+vf+jnethoLNlvDmzjZbjqtFK3y2MmrTr
CT7S/fHiQrJQQ9LYyvz34IlicT3NoSOlAokuHc0mG+tzAspEjN90l9Wyvdg2JG1w
`pragma protect end_protected
