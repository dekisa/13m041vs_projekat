// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pCEHMUt1F1fIBqrpJG28dGdUprkvRLEc8W228Fmi2ToiG15pOqvjqgh0M/Zdh0xGPIEX/JFfF5Le
0erHmoT0R3SxFTioQEpFJ20tf/QgHjxIX8PhmPZaMjhGd70JY1p46UqXWEldB8IoccNqDQKJQLE/
xElB7eAw71JfEV22mIIDftWVzgrEgTA4tzaVIQ5H8pJ3Dk1fLqpriZmlcQV7lO+dD0rNEy1wzIZx
J6r+cVr9zSLXeE8Vt4nIVv/fYVZ5cY6QIay7/wHGLOCZmyhDLhFmgEX+B2xalmsxrYRvP+fFmwl6
ZFFb6XPbwM0WTpUBPf1m9hobQuT6NwIpe4UpHw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11040)
VRyiQBBiAPPwLV/IMEEEm35jb2ZTwWmMv5XYcEBbDicyCob5U3knhOMwCqDUVksofxvvRi6tGsOo
cNz0DkfUBMY9Vrpo2DpGgaoVX21SQIHOsZcLjsqjx5wAuPk7Zri8YytKEYXEb/Ok4+cjqrASSFEl
8uL/UkXOB7DOa6QZ+tJRJ0Y3hUS9rHEO6jo5eOAokdLEXjWKbFoJOxNpV7mpAnpzGJ+sLZ6WWySn
DPmYkjFV6TTIUwpxmEZcHD8AYpT0Vt8MDeckv8eAQayy8EO8O3/SZ+H8c6lHJRs/W9/fVcwEkCH6
oafBUoY8WJ1QtmDTUmkbD7VQ0mzPl4lUGBqh/VysTdp1eI3/7PyVaYJOiogC54NMh9s2A4k6ZWnb
ilwAku18l2zDE7v6xrmc6niWUnuLu0LIYR8MIqXjeGrpJPLHCf8+7KLgz9AbulD2DO6H0bzA4YPb
SlwejWAJTC9jbN+1T8sg8UkoVp6OuMyG0uSpeHJ/jqd2psTb4+5odNXySFmdE4Ss/qoSxtwSmXOX
CShWNaPA8s3Nu2/euaTJIrheB1zQTDg0H6HdLlbKINq5KitdSDDEijpkHAcL1l8GZYMCd5GnYliV
2pDyz/f49Y9Nm0kBJEIGajjyU5yAtJ9zpYDBgg4iJuXdbgPngP8d0piehjlr9wkakzYGRMUxDGHo
npkp08v2VPqZ3qHDljuZIECLTMBfFOeSowf3YW0LDY7weM/peO8bitpdls8fDb8Pf9uSqb9oyGen
ImiT5en3eYVT32N5a96apphwzqSJ9Bgf/8yS/3no+KfTqMdsS7j45h7DDY3D+YPCIQQuanVBLmBP
QvKhMoQVbYQ8zfv+NlGa6ItPupFE6zrk21j8H+S0GsnnfCvICEPntKHp3SqXm3HlywFJTMPbnRdI
dFp8xgdUWOllwPJMSv35PLLE7xr1wZMkMBR5wTjL2M2Z/EhkfaUQ+bu+Xey1HVsP3PLb6Nmfrgmr
r4GyG07PjF3ib/67SVRt6wxSvkE7STYX1h4cajTNGiFC78Dhk2HIGjCyu4Vqg9DxJRB5d5vKIqDm
zRPYam8Syx0vVnuQlcuYigWJy6G1nfxpwi4DB3f0UfbYtyncYhchGr/K4BOTwnQCdiHIjNe3E4Oz
THL6ar6ru5UC8qvAA5d4Otr3dNXNobj1fXajyKuitXuvrCeS1AZ6uawMgEEOr2Y3cr2GDJ4cR4PN
choRhuJ1chUH33Hel2WLivwXnaOrRDv7uiysBlcc0mWfZ6CB0wLZoWwOR3eu66N8zCBaguaFhyiN
DKE+EaBeEOPT/BW4zgymAhxxouVlUHY/nLtxgHopw7xjdOKDEiVoT+7DE2JDL60Dz41/N5qu+aYt
rDDE4f6+5+vpg8ksFLdWHsXx6dzrVqg323ijnVQtPoq6gM+ku4rNk9CWe9wfZ3eUf7HvxQgb2Job
fxxmpIyzDz5MlMl3tTeEHnvCWSs5/TyAxNPXMqlBCNANwPWdEIy/ZA7fb9hLr8UZsNk1MzQnv0Vc
7CoYrhaF7KP8vy55RorMEhK3mrmFoWS/5h+GGkNvrY8TDKBhmYLbjdNpGDT9apajpX3s1GgBT0SD
F27AO9ulweIYSR7S6V8Z/RfwIJOv0ZT3gHGb/FfuHKWXUVY8ihDD2bv63l8RUu4ryxZg7kaxKoKW
87i84JRhAIrNTOFX8jedn6gK5xroxJ0R/WqbwBP9pfT/kOppJ1w8cn49SmUt2Zg+jBVtADcyEnhh
19fAhuzgvNs7Jg8+ZzbuEvSMMLYmKJQNzoI5rTTihWyahL4fFAXqfYsI0ZyYZwOPOFrMZjm80RC4
EJX4g8/oD8d8gRPPHQXy7MTKKIq6fzg8QVYtxIwI4YLTomskA+kvURjY5YliYGRQUMIt2c6NCsUD
rbb9J+UZBEGJIYG3ezp5+6gKvTeV78o4yE5X8oORmmY9htt7beAsTIAmJAVsSQ3r4ArospL5DHDO
xnC4gRDwbZFDVKYJzUVE4Dd5zwDkDlV1N9mwNFCrm1NaCB+y0x1ZVjpL4wnje8aMANHZp3qnPVs1
++Zyfcd4vqt259VkDh7Xxa3KqhUm0/aNeq+f1PcR8FJp7CoVZtMm8/e8ENNbGiRnp+FTedy78NZI
5CV4Lwn8exlxTWmOFmybgeTwVaSCnbJnv55SRyqrArG2g/afkf7xtmJXwC30RHeBzJjnqOi6HzED
BtqAv4K+TF2EYcTJUQthsT5L/wKXRrvS5zECqknjVNmrkgENFNbrzLZkuuVGj2dW6ySP0unPr1XZ
nvDs/obXgveiZwdnJyc9HilX5/4wC4kp3Ubre69XkWnUlutERk3basvm3b1CMtJZLmWGJeW/9H1w
H7cxzOFcPdg7fhY5GZJYzrbynqggwNGmEPMtVOW5Ol4nVmJKWhV21GdxJSgyb6Z8BFMHV34OKDcQ
ow9wekCLyb0p0w+OsFPz7mAsR9cWSXT4G3qCGQFpCoVVShGlK2EaFOPq2du+KXNvGsZC8i2zrEET
dGESGM9Q59NRYX0LK5WfDn3L42CiOT7b04p2R9Sl7oeCwMuvxCbrSTvy/yf1PSsMoVJ4HHBWmGou
5W8+0oUj8rie07kwRk+8Et5iQ2VfFnEE4gX6IaZ/7ryWdCeeeSSy6Ps8H8eP0C0EKGA+KYl4zoIW
ksZx1D055+Aj11FdLRGfK/nd3AJ9fektgKbFGGxKaeg0Z7gG1HXeGHwqCPvRtk85z/YmdkxvoCsA
nlFVDbIbV5fxBQBPfe5BAJ0HMHr9ZQEB33GpKK7LjaqApiUOQwzeFsopEb/etUEOmvsUGAYMrNXK
eGRrohtSt4TRbtr5oL4AV/GO0Y+U4yQFAFRzpyn0YQnb2xWLi6zfeErLpDb1oyJENBZpDvcOVKA1
Jr5BiH2K+ee1THTRdmYE4kl5PU2p4i++SYgoKKP7lnlKzxrCX3Q8856YbmgcJZRILt9hHdmXRTtD
5lDp39revUMTcira0/6BUwxXurm+YVoGHYRiSpxOZOaSGDETqs929BfnMLS0gBiAVGHFdUN4nNRC
UvW7pkSsCOztTuMDs1saTWBRktLv7ODYbPdBNEWHXsXMwr7o7HvtHsY1W6wlXsSFDoby5CNhgdnv
qcJPso+pPlqO7J3NY2Z4cUZ0SMAY9okmI8g1qWo8CKgRUBqYFkx2R4Xgn2a6DJaBbtHxEpEQgZ5L
hflQ+KZXiTeRQ6R5wIRrZC4iWSLhNdeABdZcGbV8HBGIa/DJMIQMocIgbQQyudvMry8m36l0xfNy
xTk146X5jZMAqGLvs/akxtEpCVaLphwKxm4l3iA3aIE/qqaYrh61b02VZzEnS83cLcIiJSaibRmu
Z4Q3O1aeFTLXA58dL8oDNtg3Q2PFhJpWw1zeh4Q94L1mEL6Md6BAmDhaOMAS/Js6xXjKvcOv7tsL
a1SwZizupZLtAqjXqI3NXBwk0vk0DnS8/I28lDu8feHFjnWS+wjoxd67jydooWG0lEVFND6w2wvj
DAXDs8Q+Vf0unIc6LOVs4pUeMZVc+8EzVCxSpRbB9aUsowsgDC5s9sxYoKwvQKhoiN/pgl/w+Pxw
vTua8BTwG1l1ZAZZQ4oeBPofN94lYMzzGjBV7Mn7z9PkXl9eqliWi1h6a4tRY8lsl65aZ1gsB8Dp
26xotW57rX1A6JaYPMxnxvtZSek2r+LipdJ/AUPRvfM2q9JlF0w5enUQO/aqb7l9r8P229KdX0F/
JzHCMBys9rDyHGrHFFREoKQj6nVocYILniEH9vGtnRkN9mSlGpnSf19VjHmQCwjNK2TUqw1+sUCQ
trNBN7KDrbif1Pi6cf3IIoH7l3rousp4PlpeklLgt/lbf+ybXrjWV83ch2SuurhXed5LeOe1UYQ0
mzFz4GMrQdgC1d1K9EYAOxwH89LQ+U4hq7IOKsS7iv9b5TwXgvlTuV1b8Z90Zteu06JVF0CdsIHd
6C3A2h8akEVCdYHqxa+6fpE0X3PCpJPQ2Ds21F+NPZjxxoUfOeI/6MwcMr3uQUfWrCFGAHTTJnHU
/bht9u3BskZWiGmZzB2n4Ci52PsH/J5ddGr4YABnNyTqD/uL9omW6bf2otlJM5RSDHg1JysZUY+K
JpalXwZka4UdAuNu5qnn3zyezXovln5S+U2u9vEudrDDuW0Z+YiZYsx1O2vNOAe++U7lOUhxJxSo
OR+RNnIEt+BJC1oyOcFDjeaHeVaBPHM/vpfgiVV7CQLcU+AMbbIK2KKOrqxAyn9UZXWeoUkj8KNy
hubp2T2RWi8MiRfa1fpidVpwWQCYFA3LGAdgZm7UNxUqQyxOC1jQK0tUyYnUS7Gj2cbT9OJyTchb
Fg9DOBoLeVHSoUZBJXQHbLWeZpOFuQWxK1xpvMTyECPyW2/EkeLO8WIRw1MlxP51HJ7ZjNDC5oH3
vh5Umg9Jynt1JoMdHi3tcYIyjUSuXYeo0XTQ6LzJzwEYWU4TSDx1O6sHw5h0tlEjs2fFq+7vmQNt
YihtmCz0Q9O4bprjqXKJd/pMAH8OKTCqNpAwFUc4ZwJWwTvIWfoY8TnGWz6FHjZgtIWuQcImJ1hN
XPt9QSZxFkr2u8atGhjVJuXeuvwZo6PXLXbpArMimfJNsFaKN4fdXJ6plVNsw138uFd0eSdSWAM2
aD2zZnxxbIVmv2HeJOg37Q/S806uePLw9HkuP+dJ6XAI0Bf4UUw1StLtjrrrwap+vVSSzIYrReGb
75i6HFcRxgZRuPzkgnZv/X2rPiu6OiQ+FaW4APubKPA0srpE0LXqtMcT3cqrBO6G4n2yeuOE4q8Q
/nqBsVW8IDj56VKPO+iXPzmK458/+22x70dIPqhHJHKEpxbMdyPpnA/Tq/ybWIBOZu7xWSKh3+Yz
+oDXcdEAYIC2hDfQgVE+iLjYqqg2Skd0mo3nMOwqNUj+IKzNHDeD3/r2jcKL7m8ZksquzqBjGv+v
nhCgZItcpUB3tGIJwYPCY8zqm03T4pS0jZskEEFpjiHetSjer8w/qYd13tgmCjMTb7L3jICJyWf4
hOP1/BbQ8wtrSyvotw6SBk2SsoSCG0VGw2D9/NKJijUsyNlKjg9hSiBoK278YnH++rlzZaogf/Lt
8KXSvVTbITE/LgM429CzxZQ/aR3e766bJCz0SNCdm9MM4y/j57KsX/OizTLYhmS/yH7nJHT/WOri
K/2NI0H+d2nK3Hd0u3iTsQUxOdLb3D4jovdsdsB/n+PyWkjVrB16D3Jbb4CFdiXryTLg7S71CPEl
xXS1GJcKuu7jfwuOnlRTJj73vNPTdx917L9vKt18MpgmkmLgpp6iYZeoyKbF7LMGRk7/hQVPLZHU
zQV3pxlXCfZeBIR+xHF+KV/Xv+egAvD9LkHf/w+LU5C6cX5e3K0NvP3jwLUCcQp7npaUruOp+MjH
tNLt1OOGfJXDh50008ygY6VB9NdCGHau82cob/P+DzKNv84Ouk/wl+95yMMbVne1lR86yVNWWqRl
xpfWg3ZtmLGYRYl977jet/jkc+eHlddsv9fnM7vkO6i4oTVjvb/ixTWOZljfl+6VHYPD+GDpMB1I
CD0Ha9nj52xbM4khVsJ4R2m34hrNr2YmHoCP0sriQVNmnvXL0nWklkYLR7CPu0+fAtcplqPPtd1n
19jbmEgw8kvh/OpSwa7p3WGGTgv4/xBBcJfsuruEf7bK/YiJnXGY+PmaywQxPejnr3Y2NG3/KSoz
ElLHR2BKF4SyaAm67EPqOZrqsZinoWQXAg9Wj0T1FNKocaUsQRQtSIcPweQq+s0Lt2LQpqu0F0bF
ZSPAQrh4GZU8bhmaU82/OMx92yBgiTQpsqqupA3819BCtQUO+/Ji+31jCb3bSBUHiOoedr4dotf5
vF3cQR0HXFdeNmgSHn4c0PVAMpbMtZavKYmzCh+vljEOk2F4br1DD9V/tAZMq0bqKsR3MMJFah6t
Tv9J7nHpIC8ZOfZU2K6o9wChPyIVVgIoJVzX6j/AUHY5e9vz++jOceCzsMHwVpX0hn6Dt06XkCuq
70pGgYg4amgOk5NV9GyNSuYn71KVmCq/NhFkSx6Fx7QiOyD73rPN8g2vL1Sf5Ph9yj5DnQKXc04v
2CnbwAIN3j0A5hD1GWHWj4iqYTC69zoX7fqvF3bzwKAqKmqS9Bjy+JXXJ6TGbwwUWWfWvVdUwrcZ
ScBbU0ZnIICfaOazBcrpAqGXtW0V6C6TbdZb5hMf1jnP83X+fEVGKxYVilRzRX2ep7IxnJ3dyRUX
fSLwI6OmohWJ+zDXsUKzdfA0a8AT7EC0LFIIK6x9MQTocNPQkCmEAbrNQTVLUVylRwNXnKtoxcuV
MMeaHMg61FfRg0JJ0iI+/PWF8gQmgazYnChHKEgtyc8z7Cc3JyooZWohK4eANje/7nJJvkOWreWz
AFsAc3UblHpohEMtdCkb4tdee/eOAQCCf/xOExBIbhhfsZEHiveh+yMNAd7GBLWUkmRJOF0jRrx7
3DfkLZ+FE+14BkM2ip4pljby3sjE1/MtMJy4xEORGFmqiKE9Y8w1E5K1mC7YUGoKcqi/e21lugDU
PncIJmhwBmcX84tvFT04R1MJj+bxkybtN/r+0HUFEg3dI1UijM9xp/WHo64SXaAChXSNHWIkgnD4
xU9LCMQQmsWZCF0PZcB2QXMxwPd5F4wuMIUFSwCjyCDXK2JWN2DcVkePYdRnik39PX95N6cHaPh1
8I+/9+rpfWODQ/W0tjQ/7bZs4Md9+gr/cfRS0H0OoUOPkdjWxVhjFQ642SO7rsQHmt3RmacdaC4r
Og3dLyFGYRK5ll2VibyuDxJ9xZg1F3PfpP8RMq07xIIuxfWBHomvj8j9t/eTwEldFl1wGjurTn5s
cay3q787w4iNkY7Iby8I3ie5+uaQXOghfjvaZS8g73pqkaorIC1uakY/W0TQUbT+UGJdngYCAqC8
JXWhv5kK2ri2R5hTMxMcrld+klJ82sex0bJZnuIHfB1oGs5CaLsQEl90SspqsT1vMUhP/BS96LI4
5IMA2yxhTBKvZb4vuu6oI/BwCW7D9ilhZTop01u4OIRxAap+LxpepshxBSa2AhWMvAat+eDyX0g0
pN0LAbEU184vVQlOU/y8QbY8apxNV2Qnv0SnuGRdG2hMtO04i62x8YhDam5LBCUjXVP4eKVzwAbB
i4VIJPlWodsvHNpXKsCD3x4qUODKwjvS4O8bkItR4irVAZSbhy9VSXUY/4aEDn9J2+3iyIa5XB7I
fzMvxjKD2roK/kq3fhFSoV+s8cM4/0ROSHMGmjyMSAgP6uTX6+akdKTGw1ABOoSBnmNO4kwI85iI
k7w1dY9tneoWCHhETJM84Br2B8Bs/2hdLsxC5ualDb+qs9aaRHfIeYvcoI1ZlXKcJIDfXLEFwv9G
QWQz3VxgYjsXF+QDVR0+EXt+/noyIWpZXD+yBEIq97CcWpx46CWauuQsh9c2Qox6ypAn907o4Edy
Yw6sk+NgXmfRT1nNeB5vy763sROw27lG2upqeLpFypt3pzyed9ExZ2lFtuEtqeOTuv70hfygmots
0WApRM+8QfSgGHqDdT1TmQaiSg8jtNdfzCQkmlpOP4hyRfxt/uNIOnbzQ6hwYEaWf6By9eWqoXRy
ZZd1tF6Plq01jpl6T6DLZOPym7RsqaaaOV3nYY4jOul/YYeVfybe1zjf216SuMjzfNHgbf3PjsYI
2ZjNw9ncDRe1bt4/Fx/CjPMqOIisp6j+DOPzpJJqpcG2hphw2fl1OwHlcd59rMTzrkkecUUHz0ej
TeUGaneK+7vlh6ZvZNoda7/axNsM+eaZpyXhDJ3HdLWCWVnATjhvMXfVjXp7ENZTld358fWP/y7U
N5Y/JueHklvylAklGQ0KNz+hssT+oXKs5gP4sQOy1gh/i1ZhQzDtwD0vVVzcIYK+J25xvMeGSpru
k3Hh0i+fZUzZaPOYCU7UQoLMj0HHyKDZyO/4S1gEnMCC5l09O+7czNCOEyA9c7/JObypqCUKxfrB
rD3/ueuw9o2ESBHj0ZT1gFKef/tYKzC/U0VYykmNPN2i3DAZrwWlU/hHZXuJ5bGTM5XJ7SaybMgx
V1wWg47ZqJ0pqw5RpvPvxCOdK7LmfcEFTM/pGISo1g9sWf1fgEvkPPv1WBZs4p0rdYd4dAV+AC0P
QGE50G0HBGE8iA1jKIyrWAZM3BNP7m0R9U/uCkR0PmWoPFxrb0XRr65Mc0hnLIKCTMco+olyOE85
F1KGF7V7vJmfQmpl/3uW4S0mgVRZcEwsfN7jwkLoLBQ2PzzrL0kZekXaWG9ggbqMSZ5eYGZt8gX9
E/k2T4OK+lYEwH54JJL6Q0sweZdCoGZPfZJoPXZwRsVMeP4fxQJfWZv1QWDEB9YJEwzFB5TrjJjl
3prYlfOuGazRGOM606hWhtq/WSC/2XZlVBT1ZesGgVD56bzO1MbODbMAmHYUI8Lrn+dSZBdfh0So
Lenq9oGjPxQ1/wMiCwb3rNhJtrmgrniGV/jrHLEBuyEVPN4jVmeYnLhc8d2Tu+Rakh2cLhZixRFa
ZN+OA/lfl3Wt9Q+K006q6+evURvIaZLPmdaiC0LdPT/lL1WjDywvx4sWW72HPp2CDvqdBz/Bf2Ls
KzCdoC63bnpjeayxdwi62Cy2JNIbg5GbEmKDVaZQp1v9mpLCdPpdl+96uXz7qcsc4BAVUn/nAbgJ
OmO8fbTf/I2KmVszoJLj9oFnaHwMPi4EOiMUTaA3PxiZ2KSTtFSomDbwfn6hHrZzTYFHQB/CBpiM
+ZCoH6ohaXLKgPeCqkQhn2bjnzIJ7K3b5wc1OSbtM1d88RpanLWtjBEwXi3sTxcKmgpEnKdBCkuu
0QE7kOcokT7/eSCm7fDWd3KL6DfRnsKJagqhXL4RqHxAfuj53td8LQcUoeYl8d8OYMfHNkqC4MqS
39DZLmVpML/CiYtH64JGGSRUiHGCoc30wFyOgxoDU+mAXc8ABiXg5oPO94ZMfH3VdlLcbZ5RDYW+
Ve2L64EoCaQyH4mUR5AcS50xbuTGUvgSpfF5Kxjj0FUt1HKiDWKAntqfYhrwG7z8O9VK/uSajP4r
fcL104/oRjLckLk0CU7WrpLyUMlPFb7FnIt1S1VE4MJiWdbwwdIajhuthKoy2iC0c90PjX+9KeVQ
B/GyCSnssPP/7igdS1MKbtuGFhJv3W31dP80acFe/Rf3C8mdBiuHW0Uvxlcp+boFcpcybamk/N4u
Nbgp3HMzDCLD+ibMHMebyICQ+y5yGui9ppkiDbrMyGMkXm52OPakCeCpu8wTeCkZV3KWQQjkKFG1
CgBxT6bXesNaMw8I36hSJc+bfZdb9LBFx6HIAq+U6LbENd9Yy8ZPcjmJE/TmubeQgsKrIRMRhaYY
QBngAT+oDB3fuJIt5eqLdYGeVpZvATi9FOuqBrhSPYlEopqfM9PvkDqu+3IqfJZGGeQVM7Lck+X2
uiw6snPmwebodQ/FXencb9/0VGiYVB3TbqnaHv/a1P4g8mquVQyMs42PWlUvxhZobZLRTvS63LwA
DITByYLxtiUAFS2IrTXjihT9/MIpll9+dt5IsPK6yGRiF3fPczLp8/39c4BC0sq88Tvhd8w6r6mw
xvTwPnCiDDiO+kV/ySq+LhokUHYhRjFJM3lOg1uocK3+CbX7l4BurTWbaHOPyt8cQPLOccQU5zZu
2Ed2dA9lBqxjWOtHlKTvLDJbVaX+ctmBdVOgOBNYCKdPovD6CWTIA/e7SKCTTn4AzANjCfug5y8U
+Rqy46JCQx0ZE37GosWqfR1QH9Blt0yd6A9sU/R0rUoKcHpHFl8V4KmAs5VqOrpPXZti/48pe9+R
0Ljw4mmS/F6cJ8CX8P1ONyN/jzzrEzRxwrA9zUUHPf1xqy13SZr8pcYXJffmvLKBmXMTvMIqYEsC
18wC89IDZk6QPzNgZbONw92i5zRq6YgPhxcOxJTuhpNUXto3Fx930JzRMasKlbuqhrZaIZJehg7r
c7W8+80zZzNUHXEcPpssS06YZrldCqDwPK3NNrB5+Q/DS9hxaYrm+Vt05+61rWRgXpHqC276KMPL
s+4WdCbiQEVgWPJfhR2wU0T8ZxV13eExW2yJ5tGbk+JZ0+GvyDgVStLv+xOezh2uQzYKWuorXSbM
d3+FC+gUPhujAQkaZ+qX2ooBhzlNbtXHjIPaMkQekRjiuaLCFcpjkN4j4O10eONsKnIF/pZQYbfL
LX5pBCmMw+LSRMpBhazYvuF3syY5CuJzDLTGf7MFB11G/lcpHOa2PtWwDW74WGwDdz0NfdGC2yjd
WfyvILdxtGVSe63p3BzzREctAVYgWHdOlht4G4txG0SFitCXzs1kpwRVSr3h5aqmMJlLdahxmkQZ
VMODwohtymV2LZOHipH1OSioRG9eFzZWRcbDuiTywnC5hq0CwRn3X8OjPAfR0UD2P8Y6j4v3rY90
6zoDfeqiKcCrm/r4IdR6duVTdKxlSdeJPCiCkr8N/rRhn0OO+02pGC8OSI8Imy0XABcrc/5k2Glp
vClIl+7Qwv5uNnQcCqsXQXrVrca57oOFHI/7roUh4kVQWx1YMHLWkWKHuCDRmHM1jWsaOgce/i9J
Hfp6BF4pBC+X7+erfV4/8okVLB4eFNNsgm+EGGjr9HAfxV9/UQF5Fd2gsYekn3bdfs6FeGaiVg+g
aU8GxsCZXLqx6vrAgikwGMTHvgbSQxdxyqBT3uFedguXT+TckIGopow8+GZzb0eaTW2tprP/eeBX
R7FUo1Li0vbPiTrp8BLVnsFBR8SXazu4FMzty8WBTtPzznWriTOdAAEThZzdOrsXwtUJB83tOFyn
xro2b/BujDUWpYxbv94qdhPN67RxuM4KTk2TKW3vzxuYjhiaHv7VlWxzTI6hsRvuvq1KjLNAyNPe
B9GG1B3cRooJT8M9hxBwP2WgMLOzJ11rgku/3Z0JuW/abpD8a9WnQ22EkmpfKgxU+vN/WhaivXrO
HDUJJj+zD8abixdvXcd7WT858ENDJDpTbxlc6lwISBym6SOByAu0JwYBBGUSpPsNWXaAGWFyyFwN
NYTCZUviK0uf8304AB73jei1+L74f+wm0V1HrYZb6IBmsd7lYKei6Uv02GydkprXOBAlDrrfhBmr
tnw8Zry3SezUihSVCfuJmb8W9eskgSkgI2C75we1f084oUX+AJzmyiSFifOg+T+LFC7Az3ERNs6o
jyRtrsjag0wXVtF5zTew2/SHSZqyuTjYHiFU1zH68qaEgGHv+FkGj+2hXnZsAfK0AmqZelrf6tTB
zC3nn2LtXhrHZO7pqx/iGAxhp+2VceYbf+9OKBU+F9vq2+Ixk1wDek2OSwVTBCSRVAajXgAx8x3F
W/1Uih+oBrsrTVvJSaeGJyARnMhK5zGvTwZludwgcHM6ceXK+wFRr6hylK72TDnE5KXZc10W9Kls
mKSjVKw/0yxLcH73kEFugP/G0IwQjGxev+aG+CC2M2ueJosdhpzRQGY/jZ3Cl81wrLhCMU2Am+8L
RHMrSGMYqNOkJQXcoPJvO4AelpMhlWsutIFkkYIG4c5lbumltrtdaFqzQRmz1VCx7V/iKs4x3ox/
zpHFO3Jl98yLVbtHeLryfIwQ1iLbeRTfOT512rWajZ+f0JEJIsCvPgJxOEZKrXaLTjktFQ4tpO3E
2+onrda3cg+JuomwsnN2EVu9r/Z1b2wJTd30OhLXvXJyEeO/A9GCJAUZiMq83Vxph8T4/1i7g30P
ZLdemfXiWLBTyJykGDr8+nVy+sp8IJ8+e8MPmQR0OGY8JE/PUsYenVMawyNYboMZtNrsfpChpake
9TamqeducCJO+g2qPbC4idthUs8C6oDWMejzkfDX/tPRzMLANrMDWfXpgoKW1oMpfh0+qQ9NBUaw
CmCZpIdvzCVTiFz6c0yPlCJi6AtsMqUA3jAQ9PwdOOfBsSCJrplT/roOh5FueUxtrwhwlyqM2872
k0Yk9OJcmPk2jwRveAGympWmqcxHoH16ix4244v+lz2HfaoC2Hpu4a25xQ1qQyJv10k9xbRE6h5P
PeAoZV5y3dbkapB7j0WK+DPKTa9POzC9KGcaiyNyThjxwdMbITwHDr0bJYoceh+CIe2LSGoAuaFe
p0VTgiANlBMp0L8oHAH3qaSevrirVeAu5KYGvKcQq+wAtfOJP7c4LwNxL8THagfH7HbbEJ6gj8D1
qGkuARCROTL9JbGFtERvA8cF9sKU/Nu/wiKClqIOGrrGyp6B99RC003AAIxzHRes+3qtAiSqHOwx
+vKV361my3Hu4+PXJUv98ZVPHHgsmvrmjTnlX+IsFDS/jsaUP1j+8F/xlRbPCsChY+f+c6p/fdQ7
I2ae3WT/ZOYPAGriKRlCalUPRdMDdpt8RKHZsaTQ1nCVmGXWYja3dPW7T1gi7U1y5Ap2jEEQDvkP
go9xhoOjuEXvaxkJOj2ADFjIUxnrw0znkK1b74eHUZKKntkag/a6opW+B8OZNm+/3xUe7FB6yGqY
9DvcoZtb9d5ZJWuz8mv8PJGqJHNbZvIj8eazQZrh/pT/2xDi3mvT3miETMYCT9MHZvy6Dpa3LJK+
KbHWxn6PpiEVtHUB39fjL5g1prOwkU6kTyL1608KlULbpch4wfgkHmR5VFvQhp0Ja+Tae64C9Ftw
5zP2Lt51NSmUw4TJ4KhdUpL1gfbSaj+G+ZZulgWLxyKoN3/zm209aZbQ4hYX7+cPif7T7o7pAJcx
G8ZgSs4HcE1W2yousva5MZSQWj2IHaqcOClRf25OtvEiKgtMUUhdw3V3nNwgVTKS52K0QtdL7kd7
Ml/FbOM0KBkbw46wgxOXaxW4HHGomLTAyuyM07Edy5nTIfvqLSepdV8Vx9ED+AktsFFkURebK+hV
QzZwDPEKsoZrh16cwuTCTNWwubT05g88zGPqOw8xghTPK5ZRzVyNf6PqvZT1fCu8lmlqlRYz7GW1
KLyRbcOzmvzMIT3XFGXLKB0JPhQr3P+lmBrIgD94Mjl9M5/a1+3B0xR0BWaLuujG9tkFUHIAJGGm
kJM0rNIEbih/xmk8e4Lh8RfHSQXmrKj+l4cAoULjdAINLlNwU/o46xmIR4TC2hsUXWFTC+zk3XH4
M17h97dF5TWYdjEWMKyQ7JWgYey/Z1cG0LInwLq7SiIxHWIUaDMGsv8L1cVPnaatqkOhU6suPvi/
jtoJeP08Cp/6lvUjC26401zS1PRfSqd0iSv+z3XGsSoB9NHCC5GpcZXYMP+1ZNMI4ngsA3dDe0/Q
AYu+R1EgxJYDhtpFGMuTUoC1wmU2qqEKCfPQ/+wmHCIkYC5+SousO/eIZt8rlroT6J4rjht/13a/
565t4L2uEGlpN70l8cBvjyRkz59Nlp4eS80tKUvSoqxoCQ1CD0ZfncV2KLxo084fcrrpL7A9g7Gf
SMOgKJvRAsP7pAE7DqSUXN6gFk7ZZmSDTQO5siySXc2f5Exkf2tTe0IXl4xqYSKjMhICDni8OHaR
0cLVwqVLVbwkz752qatD+StJP993rHlBpEyIxIXoAr9NuPWwF+Mgyd1TXpVwxqdVTB5ermWLD3+E
29rWzlW2lpUU5GpAm6t1ffRp75yK7QB9XZQNy5PO60UWlZD2g1YOphmMSX1ynx90Z+zfvjp2otNZ
fRI1maGYlvBX8Ke4Ev2OWjYvC8JoxWBBcMDuNj1V5ZDX/Cik+inTOkELhJtv5NL74vJqizhwR7d6
vDBu0xCqlAElBNEG+8dFmc/qCY24X7x4f30LljrKD+Nw/sVRExXvHBaJhQnWVfRnrmTRBBXVF+Qb
pvTzl7jkVm8JqT05nTHEOMppKHd7DPRIlBHa3jKTH2sexnV3fE24p8huurymDEyeIOSFd1ku+G7d
HpDZow2GCUa7fm45W3aeqUbtKiXBoYKibosgW/WZ51S9IJfEqB+I5esATyMreclZMPJOR7WZMxb/
Rs4vLYvVt2QzDP0WsiLxCpTQkuMwe9gtUbx/irOKCRcB95Lj+yWfbObsy6jkoaYxeINyRWPdrQ3I
AbTglKlTI7iY3zN+QEyY2xiDylFJBKDP/x4ODSJuSyL12GoRYoY4S5lDyfLOsbwIVD4latPAnF46
bSoLVgRCh+K7Kr36y5hY+t6A1YlS7omyYJQTmmjizIfh9V+mzi5eBzcXZJM7Ap4iyC2aV/8D70uF
ndsKWBccZ6Z4piZnfHThSHi/zAFtru2e91DDnDT6Lrgk91R5+l3+5BSqgAUfkxt9gSu1cf0o2wTl
Ck78taDHi2Fhs+5qrIEgGmwiUutQ8u1SBaN4WAmbE9SAUPFKz1URZ5oOscN2mtYwX6Qy2Q9jsSs8
SLtdlE6KSva7XHTeIRV0KE6ozrE/WNwIbMrbbbR0tENRxFz0Lus0VbvqE/LgpT1D+JKy7wa/TNzp
ejBrQj2Yya1lary9MgLQXoWBQ/Q3WZnw86VoNxRtFZwO9oCjOQtdkGnZ3cSpq/aCnH2QmeemwgZ0
0UCdIim1GW+XBOEXEulxGT/WkoB0CjOYWa91YuTvxdHwdWa3U29s0Bdh5xH4HPyT0pZH/69RZEkC
sHwcpzUwQsW9dqXvjNP0Au4v0SwZW/p1h5xoV5qu0hW4vUFza8nTHUl/p08JdM6VKUrFYeyIh8bj
YRs6+qPiaO4dGhMV+hsofNqoYS4Z2VLEy/kD+oTLKSGuLCJQSxW4efOx37Kqn/Y7k8CKD65tn6dJ
VTYJ3D6OD3byrK9QxpjDdVhPzR/PP6pfV9VHSQ0y/SehDkH5fQbl
`pragma protect end_protected
