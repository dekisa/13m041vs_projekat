// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
MnFwgv0dlgvnSa+XjBfZgVAuAmM9iajFqUT8ie86+c/5gIPH014zXPq+wFisgrEIE/V/EfZc6ykm
ffNETUqD9Mky5AWziNRSLORnk7/2Kw2nXHwviBgh20tKdlgEDq/0gtse/+3ERN2Ea3XFzyQGLJGa
JlyqaADGwsf58suRtgTFQrxCxw5rlGkN5cl2E4xSWqkOd000zsbjSZQqDpwf2yGQVU4xFYXk4Kd1
VAUmszfgODc1kv6y/O3lt0TDRw0PKaUHGXuxXnIaYJ545XYvmwlaDpX0MRRCh+DggnCsYORsp19D
e906J+D5lXpscVf/c7Cbjcy8iK0nNg3RsNnvlw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 36048)
toDbhdBuoFmLP8V4pD5XlKJJhO04juqHZAtK31W+l1/i3ypotCbUPU/LjlIZtTmPqpJuXUq+CMDo
rKO8HqZSH+rx9EpCdxohG9At53GaOl6aZp7AFGMTAQ07BqaO0u7xtJav6aAgAoPfRvYz9Rs2av38
XfHxE9rI2d9nWNE/t6K6d7HtoVK9ToEi7231e9avJzWtanBrkstdeopG5h6Y4hMiM9d8/+l5Sz7C
0akfLERYSz5/R4zwu/qPsNxMzLtkPOoIZTz3W67jbfkRuwu6uZzqk/D3s6lz6oYxPVhCScMIqbdi
lAnXmWqXBlDIOFeXE+nmorEpA4mULd9GJat/xOXGVBwW6RXG++2xSjzJkXs49f4siAtZLPYyAxLh
X3TZ0SToJOtPeRaubQWEBfx3ALveDBTvr64JnAAPobWJpC1kftlo94Z9V4eIwa5sPVKrckQjn6gS
zhdxqhN1G04ws3El4LC9xnHj3WbaH2oLbND4xzcaH2MCUJ/QyuMghTmpYqdkPyUhyF14fQuKGrbl
R8OjiTp7XjCl4ksR3OhlVc1OsupHU2+50vX/JCMapvnycW2M4iC+ci2FxJK9KJyQ9YND8De5eKDH
KFTudb7ZHGzIX9JwqQIB012ixWbc7uig/9iiQKGiw7t5uYngMheUYSDe7uYsDAt+aRmEN3PjhmgL
/wRCypZAi/GKkyw8u4P3INp+kdFwGudhSBsBQU06uZbdwd9eEJJcsTU5KFWT95RIAG46XzKq64cZ
ygEP8JsKoV0G9KXj4Zzojeb9qOCQBHbP8d0+974cV9M/lEH/jNbO3aLzczGUb+d6RE9A6eWRPEgZ
HK/EiXKXJKhR2c7gfp+w8vmn1XZ1wt0J6pvoNYOwKYDu6/tLlVZpZysnFPQAE+MVbmfHwCtbHmQ9
ZEYutjCuB8wW4YR/+zA8o5hgnqhp6caWnm5ZSx8RgSq1gY9MuHNL38+42i0vqpO7zlgeUjxNQocs
JxVq2KFa+JbuqgIXDagaxFOrsgzb1WgPABomzVk/Kz1DECG8bs1Z5c1nKpK2OdbUDqyeDF5Uakyt
IfIs6XLs9b0CnExzbU78L5ln3zha9OvtTzXBcFDInjCaT1J6OYb3gsReNQ8ZJFWdddClsLO2Dw3Q
ILbIrd+MGWSHA0RAfZR8rByR1GHZQCFppi1a63gYir5Fp/FWw8XiJCubw1vIeGIlmyjWf8xAdquI
IRkBBURV90DYc2RLlApcBNFXN3v7y07VHJJpbTGflNAYBeT7qRfyYeD505c7Xhq5/s4SvYHmOQaW
2f0mzves1/hffxQRwuWMcFB+2J2h1lxzUrYmSRpibh/eiLBfNXO7Bk89FR3Jx108KO3MLc9O5A7D
zxshmMQWAKmI/VKYYjVBWhsWygvPL64l7GsIIx5AR5snTqIDU/uCNOIAzIuQn8tmb3WHvMjl/GRd
5BLS86TRMycwyNoz7Zy3Wzs/vZGce1J+Z9cykM8vZBSaThbaUYVTgkijMe7FgKbDNoPTtJ5TfFx+
Odw4DesAJ5tVFrTMKxiFII2u+Q/pg3jKlov5tfJgqEbSOULYJXGJSlT3GpuuDWiepUZPz5CE6mzJ
9A0rs3LGzJVsPQeZm2iuOY8RvTXY8gFWdu5B62KxhreJLlDQeufbVxtJG8nDEbXBjZU2Cs1brscP
IBSl41IKmT0Nv4G285lyue1twtL4OmP3rCehf1kleTR7nUK8MVS2EuyAgcEu9lPwdMvTUr3zBf1h
VfzkshtjraabupCl68VexhjSnEKSmRSWP0len4wWZEojXKdXaDcSQo7YiSqLoOwuEfagMnxV/Piz
bBGzFLYlW/6pdzh74VJ3SqlYcmQlGfEVhGCEqz67wrDXGGa6a662kjzMl5qVeGhzboqJLuzhxFUs
XWXGKwc6db6I83IIeUB3f4dj2mozjdqvg0ukVoVz7gSRWDWzi5ez6VlOKU+RUJ/XHv/uu0QnQLF/
Zlf2OoR+AAWte+CDq5AZ7XcMnSsZiSa//sjBopK9GFU18cdlKNqdDuCLfgLJeKz/kqsuUxTS/Uk+
OQU9EoECRg1h4Td2XMyPyMkf4RY3pqSjtCCL6LvHzWFiSBMXfGTqt+PwryVGG3dxb0X+YrRnq9NX
ouXjwAWsxhj/k2WsIfMNMuav5GRJ6utwB4WZwbr+UZqch2q5RnZOZq8s6pS3PkcYl/E8RT6jZo83
+sj01oG+Bynl43pTC+ea5aXo0IvF5sXggaStAHfXIxnP/ZLKGWfM9iX+PbW1S2DI0XY7K551DAO4
UIJArlGlbYlmomwDnZVuLLB3xztl9n2X7ilx4yPxgkcU777OE8YcGOlpugqdPhlMnL8VClj0qkrK
1fTUwbpLTTJEWCZXJ4F+/DLFExrwR2eCVOvtP8th9MGNA2QJAXmXBNNQpwnRpig+P3YMziL/eeVL
CYVDtsxGQWT6TcgcYOPwFxa8rteC5ko2Ur/3vwxryGGikGnX4/YRDF3iKMQfUfjExyHiXc8uRBFY
ueSYxb/6N/5q8F+D56flNUn3PE3VxQ9HT4l9ycXKwuwb0gijKO40YCL1JhE1VncNzlAagLFDhuXl
MW35faQJ426fm1660U98EyQIwbi39ANZ6tY7rnkk4RFV6tg4owpNDM9draX0ofwJA1pMKSFfwXIr
T9qpIfblxFe1BGwPoJXVW65AX79Paz/5rJoyfOkv4ur36M7sQaMlzqqvpbPTWie51JSkpdnb12ek
uFJM5IZEupEIYtSuaJAlHsRjF9T/roxANz9gJZmLQiWU47hQHZaPzOVSOozpY4U8xzMRJA+Qii0C
MrqePlHS9iO/FLLFvI+cEBwWq9FT3TR2mvyrPxnAdzrdHMzIJBIpjbf8+VeDv5i6wRabfM5N+hWZ
Seqz20TQ/Nac1ZDtNoPRgmTHGadqtoWSas2K4A2bA2Z02CcLINwWm311JouRsbTCR/uiiWObOMVQ
sIulKQfciwOQm0m8QIYHIwXCnmLrcyqpx5A6xXvEaYWKAycFt9M0jdXEOyyxQo4RI033XbUpRVX1
Ptqgqq427+4nTMUgyQmx+1eKc4dvID4gPIshCpqM6eJxHqeYUztr4T1gPfxHerpPHnlO2Ceptgvx
BI2yqidF4xHrUTc8yjyDcBLrwCRgs2/+CoJ1qeZujFnJ49TskmxesgdoeDzuga/WXn1D/Nje4u1N
IUzDGmms4U2Gy5kPdGesv7X8MZB1VUlo+NpDvTK8nIj8O0ce5d0yQ7Lv8QPpI3WZCoairQVHYuu6
c/eN9Q4M95UEcisSUcP1u4SCHm7bGuPfuma5Yq/k784XZzpcH+o2Nn/orkIIYCHPcU0gbdYcVQSV
Qr2T6F11yuBsnk8pICkFKY4DotHcvV5EO2RPYTqX6oeXf9yzF+EFQHjLUzekMcq1DjaC0Mr08OQn
NjwTuMisG5o7oteunftwG6ZdqcBStVgt/4J1QwPBGdp8rX46owD4sXxG89sv7XTSG0QFK4x1zA6z
btsG5X5bKDbZRXdQUTcMZQ/AZlpURbMccggpzW5RGxIdGLB9lcaz7O0aZunwd7VuqaouhG9fyQz5
NDRrrF/vAeC5wdGWY+ytJM5zs7CDMGiEMVFbVxfxDRwtqjgxlms017WNZUu4MDJZ/JlJF2+eAN9l
dri/Bq4enC4XXkO/9CGcCMENDptLwV3ghx4xW7lhZAe8tNrveC4CwBZfef54xzNj11ZtXKJlVXXJ
ZGc1bb77vPIauIHLxZfABKcN30fUrzoy6nAxcIsyJYqVsqCSh9g3412/C7pgJfTKQkfz3PUr8dYU
Tcrx120m5Q/JuuR12sH8tYawyos8eE6t4/eAOeH8TJG6mG4P69bZWxvMrTeaPrUC4vjHbyWdTQpP
ouA1t2NwjqsJGPTIW/QBl90mO3sqRF5OfWpjb/5ouPtOsCEoILt+mvPWaqtkshjvmfnk/Hi0BRTD
ceuLHwczlEHA+6335JniYESDuA6EpdXgsOg4OAhLp14H2AN8ncFSFLh7wT+hc/wdnO72eBomGp+z
jT0fDeWwagatBX0MhEYDa/WIe8Vd+r/iTOeI1n2TgCdwv5U/cKmVlAbFFJCbbA9FeDrJ8BLRx5kB
pNii4hIl1G4ZI4G9hyCiWKWKiKrSCe8jNqRXN/jW7/mL74mlxLJbVWGbA2/4E7w88lrry2fZ5YFB
rNxDB7zcockB0zIsoZV/6v4DiOpx1PteVj3c9A1twVkTIVIgP9BmPiPVFjzp3g6RyagoSJCkXfpw
qFaHwrmyOIm/g/fryW3y8LXB0yM5zTWJsqmjc8NafLEZiFEGWHGVwNs25y8EINDua0T790paxFaS
Zf7TsknkvpArAVazKBBB6DBMDrqcqP1ab0nLcGtCfsNusdbDsZe7iVDMwQJ0JkOJ7xZBC/gL8JOz
HgPCMuNf8ORTUWhFUKbBwIqHLOSh8+dsTzNZOjVYUVTIyeAh+OYTWB4+8kB5hnIcqDDTASuVGOCM
S/OC1QWaHX8+dBKGv3kEAVKQqndbktKkrY5StSPfakJlwftRGuP5qn14piR4jWTeQR7KHaV7RYgA
3k2lmNgNSVg32eioZvI6Xktf/tBr1Vjyu2PmVCKB2BrblPmX36yJjbYTg6zL8NL9ZJ+3lQ0NKFRs
pz24lCPGYb57R4yVX2tuJ0fNXJz5QL3wBipvxP5u0oNWRkvk5tOFY6iP66zKQr2QGWPH8ESYKQUc
+OTvSURPoZfDRdNCV60U3Q6LX0seOMxeRt4TDLojCf/7yMjpQ8N/e256/5GyphZ4bLW4P3nQQxcZ
exb7N1khRLKDDNHGbrewAvJD2no/yWQNj4douF8YiUu5p8lIvirKk1JPZKp2QgKFqaO1hbg2ZToi
UUI74DxE5RjMWHDL+KoGoUbKkp338bpK+77+IPJBJK7TNFAgFzw/CJAL0iRgAC/IoDScqHrZcKdD
JrCouZDpC8K8CHbHUNrJZ3x0k4HqGlfYtdF8X9hnd8MNtDqA9TM8oWGvp/pK/CV7V+l3rHepWnFL
i2iafivsfNGF8gkv3qZZDqPc+0yx4hBIuBBcpLfWHdz0yfg7aKYCNvYFRctOU3dDMmrylzmQFYrC
+DSax6mul2i7L9yymieBiX+liD8DKlxAKbuzJXJvZJ79SOx4N/GB3cJeVM+6plqO2F9qMensnxdW
MMK/atYWz80Dv0+ZI0mMbCCgE0vPpjd5L4IzMIpeR9EqfNUrpHmqJkINXV8A6loIT0amPYIgk+Bx
vL1BNuv0hmTibxp5QeEnFc9l73rk2hcCJLjXoystFrHBW5ZWtM4m748BZ1rG04XnFGfWpJagEYfT
qaM4WI56vjvwwH0868QMqUhgMOvly8jFc9MLw5tiBYliP72EeaHSoSZdMu0Ym+FkID4ON+7zN2Ki
ba1Bq+MUNeGou9KqLQ7JxJ17Llg6tpKGCmDzEyfVv8BXnMcXDTd1EQEZtL4gRLbBbw0mn5gQKWRN
19UIOZWAFnGM2G0Ak775loqeWQK4cisP6RLLZlJ7yhbbivw/zVzfVVqRk+m48lwrZCWjf8kPaTY6
UZpV+G+ZA7WcZHXU19M/en6R33M9oOcVi+u/SCy6/+bmyOLBlsu1F2fMp31JuT3oFI30PeDgjLwh
vYRjnU9BrC2AtC8fljGmTdTqPnh/OFw48JyFuGl1/rXaZdhowjZr4DUHmEZfHbH2xYTutt0KZuoQ
PG91az/SmyP4LxCQ2hDqfJnAQZ33epU+1piKeO7uVfgYONNActo0sc3BjrrJGNTN15gC2ndFoB9V
LAPW93hivF4uHh9QkrM56KQCbFJaxtB0dJdcgxIY0qehi6gMy9UCWTKnK2JSnuvWgl2TIgp79d8A
av83Dzjyydcgx+IBHl8KhTxh1FZZod+Oxuv0yanr5HvcgVXcRyWQTAmf/THd/WOL1SPnfuG5yBRO
YpubE7xx7FuWl+RIbfUg/gBX5EwGilRUjIaKb+5lh9MDsfHZGdv1ezfaeBN8Y5v8avLKHjj4VmeH
HSTsg83cQ4hcZr/bMMxVIwQKirJvpjLp1WahvFIBLtnz0j7dnZ/WywsQGMj+UfQfI2rF45VrBWL5
DbAdUhnVhZ9KhVBbDtTwa4EB2SIEu8OI0zit6w4UBFHcTYtUdIInSXuYTm2SgLGACtmg6j08NmFh
gp3B7IVD2rCdpvQgj1d0tyvb4RFf/XMbRFZAqfzT7+55ALBDuU2e+OvA6KnMSR/sZ3i/mRuW733f
6KIhGaoj+XbXUBssfKEojXdqiZ01/NTGCZ3xX+Z1fZv3UFtGKlih8PpwqCE350luULvot0Gev/mD
8iGkjqyn9pEAFiM80x9UY2iWb5t6dyHlz4LNC9SozPVi3RJz5NPvPewYl0P9LXzulUfZAs8VcKDq
OWxKpBKRffUtCil6m88GQkpZTj+DdBHAg4aZuC5P/aJMpL8DGM2axJqrYRnm5XxHLH2Dchee7E6U
hRouZKgL+COkitRG0/jq1av5mumeTmuZCHDpAiTLWKF3tJbNfcuQPmbzPv90h+M5aF/2MLswSxZL
1zAF6p9wrNQMQ0qGtpyuQUDDhjMr81kAwQOM2u6JW7+nV4IHHbq40SVasQqovPVrSD66BGLvAdAa
LoIyWFB/byWduQKD72CP5+zOmXL2Z7pwZS7lDLbMyS7Qu1jlUzgiin1fRFKJ4tAJnK0K0bU/+Bh/
D2MDES9f3CXu345D/PJdmTi16iserKVg/iGBvfUNlzQNXJGIkMRrs1hyPxPPqeUq4BDpjr45iRkq
jRdrKQOJKe8DJ6MV+qNkhRTzMTijFltlXYI/LfiJkHSvzBZJz9drcRLnO4rgACLN0zjDniDSL6JC
HBeaRyH4Edqz/aThP9F/xlY/HMBYUcR9s18K5CzfeEBBXoJbzCKZExqGkxXF1CjPWYpIURQSj/TR
SfPpJ+8LLFahQ03f/AaqRp9XgzBG/9Ijb2XsuTlrsNnhkVplqkmECCrVDPY0nvzSIUgJqx3L2JER
nfO6lZWUHFUD4dz66jBqMuHqjOrJAGMuJzy5cjM+oVFe6DwlPqynyuUXlLGWUz5718AgMv2dtjqY
prXReKwvJB99law+DxuWr04Tq0xZvD7EY08OOpJakdE2FsdOTUCzwn4OXTaIC8wUz9N9RV/4K+gk
BhGb6UJLnE7FUzuyJpe3EDMkk/bkdbOYHcDrvpV+m3xKYemMZZyjiSxrLPHLvLB23PBgVKmAcH3H
PHMEO75xSkzdb7CF0GOQmllU8RQPvd4qAKn2aa4VuKRlc4YJDnSMPy+tMqGzpI2LZ6FtBp6n/gmF
K1cajFRoXrnZmTCZNp6rxquzlEyYSFVvEusqcWf69l8g1+ecDEYwLoqCNQPOlnPTh5J6qRXLEfsY
xmTamS/wtZ6iEPBaiDrIOKJ0o7LURe4Jle3XZWTNz1NowFiEPUH9U5y50huvVdDNIooFTfeypnjd
Y5gLtD0w47uVodz4mQhdvPo1rQV9NkrQweeWNwxwUT0vmRKxe/RC6yp3FtjxWIK0KJffL1pIFeK8
jfs06QHZPPjmMNNoEqBfysdVPEjFGvoX6CceoRh5hIOaflAxYv2YCX7SlVUIObLCp48v0hUTvNBt
RakfHhOuCHjM5arC/d8VyVS5uFHS0zrBmsiAaD7wi9LuEMVTaZQW6pSZHc+KYAmKlK+FajQbiqko
XaAc1I7T8xcofwe+Hmi4Z96IdGkP+m4hV0U+ED+Zd1ojiI9Q3sMbidcbUZYX5WuZ78l+uL9d39jl
dgtYD6PNi01c8duYOm8hX6kGqc1XkH9m8BQ9/mKQ3uTrX7A3XidtPE44n+pWTyxs8z3QmizRQvPb
5hi2VNFweRdUJP1Ro0/4k8e5bpQQTwFSTxSgU74qTGvpXOI7JkgkkeRQOlZgZhW+bwshmsFHbGP5
RxO12hEv4HmWI4cUtZEjTbrsBAmgzKt98xC34njGkG1o3xeIhY9oNvg4S0X8YUR2LBjlbkgHnU1+
n8QJ7VtxlfCxasyMVNC/+IE2tKHn0H3b+HQmvky87hHMd1UNHVgYOCRZj2zD2NjzldFvd8mO+4ZX
+izApFSQ4aK1UxDISpxU4ATWR1YPGz+6hO7pW+zDRjAAGah+UKFUSsJp3c9SiXjVQOFay4RCqn8E
HgNpMbai8v2jrA8FkbyLp53OoGgBfzUv9h4RAQ/kd6ZFQcrHCPj0DYFd4D92b4GlYQcwOPwsjNqi
SBUFNZPA7X7x1unt3f0ZJ0VqEOxkGOvPwveQiEWPKSQZo8tFy9KLtijPZ8tutPUf/G7l3EJMBhLI
53ecUI4aMFcTI/nZBVfMf2U7gz+ZhAPe9As412Wm0cJJeNQiW/uM1Sro46tdnW0IP87xiYMB702A
A+8KoqcxCCLtu471TZPYpdno2T57VXQUIls578D0xCwbAXnjnjr4YPE2Pdpg6z7OAJC+RyiWm34n
74IrRDhEPz50SE0rUxNWDPUZZlFWSeNGyQks0K6Diq//DZtpOE73aNuWtD2yRwbG4cG71CFFEVgY
tTXTg999oYGEPX//a2VJVpc6zSZQSL7AnKPodJVjgomnw+kTer6D7RdDR3N27CcS29mFfONTl9La
LQrXGh4e7FnyqfA90+/fyzq8OAGj4BczHVhM1UTd09FGZziR5NTzSukq4ZNJpARVtDsQe9zPLg4F
9zmSUw3E88gAmZUnZXHjfaQcqK/dhVqxzJuAXii+SlKgDs7J9p+8j3mIHLxtaCMXTp538K0cQeKv
4CyUwcxV1wTN5gpHMen7eYO+uY/Kx8rMNmTYCnp/+n9O1j4u/yXXddMHGYpNt+/iToVEFIrXvzcM
gqV3IUTfLvTYApi3Bs/KgQceqrqlLZCzxwkwQ4xLgb8+qw9NkIHsOGAHF9p3DBTapu1cUzN7Hxm8
KmKU6niy1r2WYcgewRFcdP6NLTOXoTJf2MjoS0crM3bSzPfjEdE/nHwyO7ngor1Adt+Of4puZygT
s1uvJQRLYmos9+n5U+BGQAeYW9vMiHMYKkEzaInN+y0JOHUlPxmBoNhoKnosnglok4JWTwc2p+8r
2NpZ9skursuW3JSGGFF+nykzvm396jnyvB44gqkPVyvUppRSdzKeqqwVD+gXG57YVIA337qLnPfZ
/HGMAFOPKwWUsvu8kkLUyWCZf6gRC8aGpIM7k3UEwJZnkeR81PZ/ZRC2c2HGrNcyAnoVIqrKD7Xt
BdnxBSeSA4J8+MNattGIEV7bYZgmRWw0HQQ1eVjarUZ+7USmYLLOMBqckN5OrbnXh/PIxlLBGm/R
vLU49LjvnX9Kpbgdc0Vni//YWFzZlwit5krdNqKE20eL9qw8Nnx/f6SRimbzeL2rgUqTnzakV3mp
V83HvjLNgEF9mgdLOH9K5Io0jG0aHFglhsDynU984k6KvemgUlVuQJduFwyywT0lvtNcwazN+ImB
LmXIZI6KL7BOij2KELtvpeRW5eO/MvdiSF08Yam/GcKwSwtqPRtVHOmNoNjoagP8b5Wq3cySyL3p
CQm3eRNAUjrj9zKQVg7z+TzBobRK+5hIyzzS86Rj2NNIWcp/TD7T0+jDxqyAU2SXoz5KkMtUD4Dr
R6+wdyMFAVh3Vaps4rGTxg/9x5ZyZT00DJ2NjhArQJi1wAcOWzAfGAGzsTvdzLsn3qc2QsO40j3s
ER2uFK0Op/Tf7fJ7VMmltQAiB2MipQdP5muyXTURBTZBH66+kh0SC6jI2tWszk2lX9xRcZx/4t1n
+wZ4dNlQbwaFWvOSN3Uh3dxEkNd+U0A2wyZirixvcU7uf6LAAW4oTwbOX5QcWB7oyvm/j3yFhoo/
qn0Q2wgqDvB6LT+Hz+Om8uZDl413vKe7yjPJQn9Vaj79N9UDkat8zQt0aUU9oVKjrT/lZe3Ro7Bc
G1OL5nVQKb28cZObxjW/R8xq0v+8kC67TsAc3nb9Jfs8zZyL9VedoyrIbFaU66yEz9cAbJCSta5Y
2kDNvAcfnyE2gdtnggCr4yvGKM1clLw0ZBr950bVG9XmzXNlBlnl4yXZ32me1k5eWQrFR5f23BQf
DK79hQidVghbDdQY2m0OkP8YvkETU4Hi9NdHn7RCviy0ejZxmhWCFM6XtO05qxDCBH4zVq3jwwl1
+vvje2qu2kI8F3kBkCxuw45DwKIHnBJ0OBsgKz+qDCZT/x9M4njQOFrQtCJIcrzNcAfuoIQS27D4
kMO9dV5ZZ/cM2PWZXOWwN8jiJx44LrfCuybomAuw058e9u5bRikABfPxDqx64d+COUml7OPrylF1
n+2XVSxPL0Jlf1QMQcibDRc2cZ11wbXH61vt1YlIRUdk20WHrScjRjGSHWw0JmpGdg/SvmxryEyL
eaumFRTEEYRpp/XNxm+rHyunO2g+RNXTlf+AGWqSuE+hXems15tdz4yzwpIGbZtFsKJrEYBinkZ4
Rgjhj+oHOweHxAlyCBM4mcMWWelDqBJoEUbbqJYHJl0DkjDzLfMjbRjJHJ+sOAqYiDQDq2gQnnyv
qQTsnFhuoqnyy0naPrD4mSZlOdJT5zuPJAfPhnEdYeYX4VobnRrjoFtZsV78AzdeQNu66yII/4h9
K7DThddI7OWuHZ3aX2sWO15k7XPnUphd5lu8f3NemhP60CYD2z5a7S/M+XN/Fd9GG/8ZzGDS6Rmj
7KJNDk3wNWuMRHSVQVAFlBqOV8GuPl4tJsgV9RvSQdkxvXSY3pQCwtiLdWeU1rzZTLzQa6Lz03yG
GmlXA7JBOHmJuag+CmIBNzFdoCZEv7bM2jSnEFHneIDilMiesH+diDryMIPjcCGHdsJA50Z3GBYo
Ikhvrr2kLzFMkGR93P0t7acG4+RQx3GYskc+gjQYkNr22HMYb2Mt02cgO3L3NoqSEFjJQEGvTSVn
EWfeUSpXJnP/PHOZejShJb8rKQxJuSigfNy65gOVpaAt8BAYBkseGgtIfTomJC+CrLDN2Onn9VhO
1wcC5mjGPhE78HByD1MK8o/EpYqUc6841rWvU/rzshibZyvNPv6d23J5aFEOldSLQUrW/eMR1iIX
Q66fHIjoM0AcPi4clEMnoMkh7yB8K4cYZ5JspNaNgAzMbRSArTzym9UWk+71IjqnL3ZNjZfx1M5n
yhSJngGGSQ7omIjtT7BTbx5SQor39q3HZipsX68AMgyEzJMIC06qDklVBB4uc6bPiRzMxgSEFlng
Xu2HSU8BDNwYiybtAqaYT6dKcpbF3oIJm4rqBzJNcaGZS9cjD4LdnIRFLSWC+zRxcyMP1hX2Tuo1
PDWlga0uCmTGs5gPrte0jeDxCer5Kw9eI+9AEl2ZK0rjO/6/rTkucGM8RtseFvbGZEzhSXdvbGIq
2vRCw8ozOGZZk2aFu4mUXghzPHMLsHTUSdJgP4ACbf7sJLGgu9R5Ljs+alG2agfV4RMeVb55C8go
axdZF65hyq5mGu3EkEbau5SsEvdXouSsWpEnxgg7GQ6iSqiVB68VncOSOz9V+nTbQena0DiMcxs5
bUdN5evJpacjPtCjNDyirMREiilnOrRasqrefEK+VNxEE8p4gpBVZJkfY9wu/7FbQ38O4RdODvr0
gp+I+M7zpFov9bObXntRreNGflaXKYZbPzoEnW+sMOOtLWKBGYnAP8LBd66vM4P/+hl8msDDemIW
VortxLOluALHUNPzYxEDRl82sVB+0VWYXZvsm2HCexKg7/jvh9I/Ns0r2OTmW2nVnMv28L8B9J8g
IYwpZoEboyKb2Gf58NkeagJONlAJEmPfrPKW8yMhb+UvUAEH+1zrcr4dpgNxR+LKI0yVo4npF8V+
fv0UyoV8/jNi4qwXB1iVvET9hnUibK8ooUDGuAACs7hBbCzlPh4Ci7ljssDTtrqdbr1Z+hYfs+6r
gaXHPgj/++qC46XMiBbIpFcZqWQQFqyl7EOiAu5Lc0nH1Par1CU0wajYGJHnDAFBQKtBfFle7Cf9
g8OsYlFVqZiT3mArjOZdntUHpwZkP1p5DCsKTxkzPm3wCBDi0s7LMlm3A1RsPFHKRWAD83fvHvPK
ne2D3GPy3cXk1s0unnS8pTJP+/ujoIlFRqvJCZJcMsf5394y2AyoAKElws+b4J8PNBfOzmopobE1
W4iP7zBXfJCWTASIkpkrXqXUHXkRn+wpL/kaX9tHPNkuGmcEexMqAtnO/gnVgfGMvgGx/3bYitxW
WsFV1Lmonbi2hjXps7XEfwRDOnArhxTfyVE7WklryEyB3wl7ylVOk9eqzf8ypi8UtY/QpPnbcRw+
D8TUiuBrng7hws+Xn0SYV650VGjercDe53gfCewPyj8JeeFBX9grLmqLq5qXceQ6mn+JVb6XvDqg
24UnP+v1ttULhq4BNL9qk0eFJBTIkQGi0A8zYT9kw3PmbM1UUDNeOvT8hH/L8gwNqx68feeBMpHm
0Nywvd3lHfqyGIojAXjfXRtcvjKoPk7CS9WMpYrrldU/QdG5ZtwVhBnpdhqRjYTu/YbEmNK0mr2/
9X3VQDMKUde+GJggqHMHxXZ0oPKSVUQZCK7mbskjbyPHV3k4WRh/OxA/U3bb2JivH+RfgaBmJnJz
dL5ZChzJv82Qqk5zflblBYUXXu7iBT+o4hHEOIHQuRJFtcVF542ZF5QxDxFxofRPpRihIR9YU6Xw
QFa7cL39agjY4ReQgH+hSkBTZ/TczpwoCoojI1kWFThLBb8quBgLIwaYSu/9FGAMw/76Jz9lG8eW
KGg4byK2GcLb8h93x4VGfHIvjkDzP7GaTrN1URrNn+307cZzNekOukkhURNLQsv/h8rriOBj7PD+
VxboySfr3NNIyTyLrvnBFAWL/eceaHW9zXa+WqjShzCxYMfPv+TDOLc7nF97AZdIxo86sSwKq4h/
ZR0wMD2Jy/SyQT8vEX4aMRct1ZSbC+OGKHtN7BsLEf3gb/QI0rxtqUfil8OuhSjuRMeRl/IaITmv
w2cGUsYeqwgeZLlpP4UH4yZAKmBo1+W5rGyIvagWASzCBf1nGUQbmPKqWltKmC2LcYhN7RkyvtUn
dBBv7xMB9Cy+Z70NxGWYXiiOTD2/cdMwvVcFVgMLqZvYZApLGuLGWlwywfMDLxC/ZZrzEEjYj2SB
Pg6mJG8QyImL7vXjxQKRjIRNDz4ZJdMw8+1R+eW90Roc27fkkK+50EhPJM/MnWdxjKOj/Egp+Cxv
MDj3avBJC1twtne8FXnXlVeWnwz9ECHYNH+Pr24d5VPstEDJHcbdK0T4gQOYoUEhWY6qV8eMg9RQ
4iClsGtE4i6hoSlgrvYdbazx1CUsTJFesenUyKbbDLE25X1Ou6LkOPWveDr2BeosLwqJ319dR+D8
5FTxNEUOxKUr7mlwq4KZumCl3EYZgkKutJBG2jzh/bonmqBEb7dNkRwGzIlNxxamcvQ+GnqSLDFF
mZB7TBo/P1FjlBitmsDo6RIfQ2RvcSqyMI6QPnHRF+DqGhbVWaB06QLbll02a915MzDFNMNmlj2T
mXDY2lOlZJGyqYN8jYCvV7Qj2mGg0ChrsDJydUrA90i7ClPa1ZcROK6NZqHddBBIeKh/KjAdqXrb
aMI7MjF55N3jz+Yg5ucrK5cyuYSMTJ/m1umY//H2tk/YSzxCQt2Lb1msekOTtjcfS60SWNEoSQv7
JLCS5ZuGDY05tFEIooeVbe8LjvGEUq/5SSthI9eFHSRlhS1FjbFQjJ9kWvTOWDpFWbgu5KiYV0Su
H2R8Z9/tj8eUM+EPAjvicZML6zgCl9/v/uJnvVj+W+Ns+A3IjxQTELZZ+2BrO0sRtkivp29H3cn2
5BbMsFBxFIPl8rtmBB5ejWR5S/xJV041Ow7eFEoZNpjfj6IHSKZJFK5R3iNa/gJTGYfcJjLUNpNH
P3aki6L7gLbsLW+dQ1D011YcueasWbJFEtwN7YvT/dCEU50dzCGVOq4BUt6ujDIaqzfoBQSNrfEq
a+DkwdEXZDd0H+25uotOELxZdCJ56SpnYrydUZpD9p5rDGuG+BLBCXqs3CoCE1XtmKx7OnxP3OkN
hnOAfKZKVvVpyYeEpFPEoZJeZepDySEHbnIm+A/smKhufvnhs8/GOeyaUCyPWwCfTJLXPSAgDsa8
gof0LXCRz3LNhrQuXozKbGNfjhhc2dRoQ7fsKphA6mlevGAKpHx4Cys1ApLhb3fEDRwTGvNGaAOd
wsqVw9ziMJx6prcWcShu8NNvvKQQOU8fvXn+KrHxKcOUL3O0NVfBoTIcMX9DgoHpxQK5qyvlZg5L
T4u1/SWeFu8Oih+x26SZTjsRVZLzdbztwbeb6mSjXD/mDalHyE4OjjDPDf0ppMaPd6SAWmpxTdHT
flpvQuC4nvEhlnENNcLC1pMdbF9x1rtzZTDax959z6S9I7s4eHCn2qgTW1SyVIWVjT7k+3lHn7ga
DqIVTX9+krXE4XKOuaO6fhlN+ikp2PjI6tpAsnWAPh4nNTRz/AB4Nh9IcGh69Kv7rX5k+eDXu7JX
wHsA86174mQWtiFDQGLX5sGVf81N3akJjD69dfPvhgJKfDfvgVrqbtFjnCPUmbJQKjjdaCs5y6Ga
X7ZZmWQzmozh1ZmD41V9Z1GbKpF97twwTi1tFR/N6A2N2lNbhkEybcoYcP5FZUUI92qHI+4WgwUJ
56cmK7+I7AGo4qKt7K7zXt3nvJeBd5+d56rXoz8qg469CSrEHZeyVwCpcXb5xJTxrEKbtgzghtC3
xoc8dIvuuag3yqj5P1ay9rfiPxFV96rMjgZg1BQAyvRHeadL77qheNsk+6BDjEEgWhuoZyFXx/VA
4e5yJzyTnj7i1olSWO3DYtTk8v6P/ljTtNghcItFlXYaDw/23SpG4zJ3SKRzeDKxZJcdAiOz2oam
MHQ5FRoN8+oosTs2/4ktHJuHjxukU+Lip9WUwKvJPtO3W4S/KlBEcpJxVENhjh9EWhISI/wfkCRV
0a/2+GAMElu5wnApoSYxy8hVS51Z8fiIXAsY+r2XaOVGkkpJ9MpbmyQNZfa4aMIzVJ0KuTdkN/9+
R1YLilGojhVmi8qvPmon7WPMYpy7+YyJ10WPLyXlNwW4O+xzkOpe2hQqa/lpCW6s4b2kWamQzjbY
P94kVbvFI6Q+/IC1QC4OT7e91cVKr0LOI4Fe3p8U2XUM98/V9IOCytRQelqVp5rD+D/sE1T07XY4
7ueeS9T/DOPTGkB0PGylAGK9KCu2hqgfIl3U6RaFKpEoxwFYUVVO5fBL4k+x03hLE+XLtLepsAes
2N3c/J+a5Sr2XXccRqouKGAbpTChx5zYg/snjsw4oW+47KwKGvhaAm+zQATtA4NPd6zXuTFmWEYP
daudsJX0m4dMEmJy1wxhbRCtCYX3lEY65GaKmsIRZDyZ4Z+b+YA7XU4rNzLtUdw07SQBAQ5NxtyP
arPyqWwnXVNo98HDYRGKVm3WqggXqNydfbuQJZqCc4rnVkRjL0H+24TAb1h9M7KH7YWhWLQLlEff
iSie4uOnMCkAs1WmGfzhcfxnKXzjwzsrkV3y0IU5egJ/hnihKuPyA3hgYL/uU/YaSVXsj4GK0Tn9
ls8x2ac4ZTT9PlFyuySksH1Tg5ZJarwgPJesfuBuJ+8md91y0IuTSjEfF5EZswVRCfVpV0AsJJU4
YDJJyyrPTYQ6CKzDtg3KnXPQVgxEvGFPdZBDm/aXWFk82I8C5YyX7/P9CcYuzTvzJX4mZD6EHw76
otGcDEvaZu6fPd6Yx5XxVZ5C0tWLCm+5CBneP5mAIpNdX+IBXTNML7vRb5zE36Seek4GPW69xZkY
oVg3s4PfvAH2WYVZl18QQsiWhRppEKL7YauucxvPxk5QNHTkGkffnhh1geaq3MjpZW9BwXxAnzcd
NzbMOgHsYqDAtgXFie0tuROZJPJ+C0iRBeE2RXLt80NadXAceWt5S6qIP5xPzpOqEKmpBul/VbS4
0+HSB5pDhIDGbN77RjnahnQkrNEozM5Hnx+1jvtjTQKxyGZ3f4yajSssmKO2o+KA+zihGJjF8dqG
e6ywBlydRWcVO8u0BkwN01wlcj5Xu4yd4fICiMlkLsu4rrr3shBXQLaIsHiyJHv0P0KtM21ugcz/
3WuWWrPa6I1M/6hslAHH6kW18J26y3f6KO6tNjQ3e6NgYvNNtP4QFACswiRTxfjITMtL0bxrx7X/
JBzlX8M9YNNNbo7OSWTlR3nXNw2qmvyVO+vVroBkjbs/wX/pUmEbJL4UUQNMfA1cbo+7wcC0SrzY
zKlnCKIMe0/gLBymI9NIMO9hmdu0+dBy+oSLuGQ0x73JVBlFk9pofyB/c+0nb3pnteaLchSIX3Me
3EUpXqhK5JDeNhKscVIXq7qhO71njSjBwj/Ed9COFGpRe/emaZWhedDceYQPbWuRo7xrJH5ZBtUB
566oKJoFeCrPBbrm5GYg/bDh/kfJw5wy60lQfOJoc5YDLKmHTqjZlJV5UbFlRXCRbEtmKpNvStnV
e3aqthiNkjC1lVh6oEXgXUboUUgMWPvr++Zukue6cJrLuOnXEuBVsbo1jEzrDX59UpMC0tj6tOeU
GV60dra/djBeRLF0u0d4LULUwEAWoM2UlWtKLPfVEsyhlBaqqplHxhxQWWumYjkk2y/yD5X5H5kt
l8CWPvTlfnhba1PTUrgVpL/Ni5e9UoI69ChYudYQGR4iUPxS7+Z1DVG/TREhvCBd2ebVJdgjYJrt
kTErrD+m07XiAjsBi6rcnjFhamydxF2rc3YjDyklgUCsjrobiTZVtLGA3DFnZ9jiB1jt9qSGN+xh
5R39I/4ylLTwJLQ+NvneFJ1rBviO7km44voZWHWstnA/GEGCqvA+d1IBnsY7so7kVnim0LKpVQ99
bnObh/Qce4AI+IF+GExXg8tm6aAqcZKMW7TF1XmX/hq1G3HdUFmpocNCHKC90BDTB+A5AEe0rYl8
J+CnGKiX1966sYCHaJLDbLajg2BPMoFiVuFpp7MX5VqpMLxdBdwsggIDNtH+W2SgDRy5ovi9rC7s
Y2bsu5aS5MwAHpepTKXhdhmj+LyZz6N5LQNsLhQZmRtNJEr24AIz1PbdQOJ5XVSIb67lcOFlh/+8
dTVWm0TOB1wpiDTK5Ji8eHjBrz6ryPyba5aUSspzhBT6slwBbBCaqsnqqMjsosQFtMPg8FBwY6rb
PG9TH8pb1vUckwLjzwlwIH1uV/nnJ5jE2lvmzGrRprK8IV/22rOglnoOw0B3NKXemw8aZzOyhHtx
eyZ4Rg55fx1IVeqGJh8EjU0hB1NPIKqf/EVmdlyybHJ5frHJUIKN48n0HIGxSwvgCxGZQQzvJ8Rb
WneN+1mFT5wT4I+5leIz4hs2EJQHQdzKbNrGR+Thbj9YlPgmibHm2AwwvRqn76Xti45RuZa/KQt5
kt+jdeCEYT+Sq5JTsbrdhrMRffgPg9VnuJnvHnwPFHya0hp24QQxC01PDBSyf0cfZ6QC+akp3gA5
t3vIyq2vo2kr9rQ9ROSONvmZbEeGngW8QSpe4r0IjRSucFIgI5vVxOn32U75i5xl2vCO8cwgbChn
eV4RvWaEAn5oTk92o14cfmBDU2IM9BLIVjUOGVQntJaOWeZShTfZS4GKjh1B4p2O0aU+cR2VElyq
Idj8s1O0vE6csI7m2hWsznwDSX7irNs7CXS8j1pBhCfFBekIikb1TlXL1o5WBSOY/VVNMhZDz/QS
WBCH6Bsv+YeaCMVp28Vrwp/RF9CgLydFsLIe88zpuazrR/Und7As6dfy3COlJUhD0JCpRv+U01iQ
KeSIaNZcGSX0uxmECL4FbG78vtcKruiEE7oWOB0s8kQbApzQ1ZDRDYIpOJj1vIojYhXBLtthGxB3
bsOuLebOs8Vu8u5Riwd+n4Irsc/2otgYqXq194mmwchp0WrTFsHgr96YqXeJvxjI4y6x4jQdanUv
rvFIA70pj6j6w8FzozmQqxtctbYyd5pOowyFrVcnVDyXOSXX4mc98+vIwD7C2P/8hk6vFbLwqQaS
19Tm6OMLTUlbhuQuoMPtbXhxZYD+S9n1bnKisknDQG6xSZ+nMV02yioEKZFpxOYS9KOqcLSNQC9D
sF7vJSd5VVOhg4XCsQQe8WXw4xJxiMFSmMqUfXIzkcXd2ZIVBvOcE5y20VLw88u2TAjqHPkOJEX2
Eiu4BDW67t9N4Zy3yJImEfxgYLzzuKsfnWvUoIdWbO+blxL/TR6JA27hv/yu223sWqNR8Joz2OAM
0s+jfHEyFpl49NIJekNtcR0ZR5VHznSZJGZKazkhpRhUQ9wtqxlXFl03e8A6fVRrUA691Xtr02tW
mAIWsRhMUegcd4M9+xxq7OY3bzPsuM9u6YG427q7RON5Dtza/VcycetvYDNb4wyG0ZGDXzdoayKG
DcMOGUKNBvI9/LwkSE+misJ1Qta5w+sdABdGYY2NgfkbqgcS+wIes7UFZpQN7BO6nBYtUW+tA2C0
61D5bFQcpW5FhDjJZEXTELjIpBWUWULAodSFtDETOP+xEHYp0XnVuJyq8HoFvZWW+7jicbDWo4A5
wlIHgf+RQ44tOT6Kl94HDLAvOWAezBgy1nig7nJ4/2EupGZuvHWUDth1RRm4uj5JOaL9o8PGzW6f
sKJn3zJB/qRCZS7ddV2rySVpQ6PICodTWo6lLPklooBqodCYCuyg14OCAEuNYzWTVw+APz56Z5iS
3Ry79kYVZ+HIK6cxwdBwZ9v5NjcT18N9ZghxVvQ+uz/OFBBn2R3wXaFhzIVvR1quKqHezcqntx5X
qPQqW3A7AT2RG+FI4Lkl9fXplNq0/y8COzmv1iFdLy7vANtFaLFTzCJFjs1KB2n+Bqxl5q4FBS6P
40oAQXKAb92/bNNrJRO3F+OGO58IdlBu/rsy5xrwz1Gojo3GXqSZU1r6kycosxPk6M0vpbmJE1O6
jNzy9ElVuCyZ79kCzE2CzXSIZMZvCXIS38Zcp9YQPyWqbpoSoHWbrHpVHxZ3dq9XB0pRNStegNV5
hkIRi33yKbfw1kyWvtDWwfsZpGSITPwQABFsKIc1OPm/RnHq3OwNI025+Dqpl71W0lsjkazqUVZv
G6i4zIfbKu1TT9p3/O1iSH/Nc/GeOty6cy6+gM4wNy6Wkmqdm+STVLmXY/udeXTLM3MEVXhC8wW9
dqVDmYnpgA37OlbvXkxQTEV5LXE4OJwCJ845a6UR+62A6XUR5kyDhpKLS+sujoMeKxtmr/mfI4Wz
BCl8rQ0ek5ysvy9pNEMRKLYN+hNKws8d1i603P+moBn37YrQpd0Ook//bQra4I16YWjkX9bWN7Y8
RtJxOfSIiozVTZQizpUahkhZiZixexBRHfgRs6cqpiZ2A4dhfN0zujULH9sf+xjDyrf0JOfJ6UFN
vvmCu/JYOfJGELTXj2C5lP0l17rz95UE2xnlNWAuIcagwYlE59faA0sgzZesE6WZoCjmAQx0hb/9
CmP5tyhzoHQqsNTXwarUQB21KMGTrZPGo89ZGU+MEG4kdCAEuGzPTcIlbIm4acyLrbhDTL9t3qPl
DHAuZTteopUDrN5POhtksodiGTu2m/bEv/RCFCpGIPSRwhs5r/ZUmZpEVkLYvbbGEJ4uXNR7wLKK
+lLUcPg3F6tg1L95xyq1KlnKb70lk8uIeC9Q1mUj41Uo9HcNDtt6EkOUuThED81ULi+LW84KG33A
Pnz6zYAuhLK8H0P1wh0SGahSONPycN3Ay/LIPUaFhAsTeErV9wTIC5d7zrjCH6wLdVydIwFIavqB
zfTuE5RD54SJNq77GUevNmT8Dfcd09N4vpDx1A5/ZwYiyZ1pKlBko66uxylclfaIdtHR0rNLM4/t
Ho18+/ppJXj3aoRKKluhXe98x2u6THWP2wHsa3UIh9fcWD6Nfy0Z0WbEZkpVzV0GIckg5In8Xije
/7ykpyy2houueMrYyAiYeIYw1FJSsT4UM8YR24yYLXzv2lGJmqrGEROnh7jjDjoPbmB4cHS8regn
ucQmd14MWeU5sNPvttEWNE4Z63VoS7wRJBtZjYYEDBN54M16thh+QFtVs+PE9CBWHw3cdD1wkfyp
BazAJzad0IOD9xulnh1qTkewGNBSqm8HLZjph6YFjic5ewR87nUPLlh9WSLI4Zq8bQaIwQ+X/+4B
g/4OGVFddOth1y8cImDXsnz+0DOsXzlaQkpYnBvguqqKj4FLuyzWtpgmDKUXYxzminxtk0aDqL+n
Up+E/nxv1QDQ2wRUv6TZ9OLpvD9N4Nb2u+PX1CMt08HjDXRsTU2ubKF3QBem55wM6b0vBuOyg3c6
Wj8mtY2XsgGd7kjQosDPZIxUouZ+UukoJGfV96URhPJoFPEQbj14HFNno5iK218zeNfLAW0ZdrF5
OfeJ8Kt6BT9SiH2fp7zfxa3V0bJ2BwjOpAL9xNDHoDNuxnNBAdGUBg5vKcPPrf4OEt6vKLRx3SE3
mocpugIDLwT4LMXTBF3iTg0PDvaE+/43f8F8Hrw7pSfhI93nhx4HCHtdy5fuX7PaB6qgWzt+yFcW
bK2oR3G8Nvyy6qa/2bbKqKQG5Ur9sw8mxf52xz5+v/TazlMdbDL421otEBp/2YARO7b/MBpptOw3
KDltApVvNhsgLl+IoIQGRrVS76aQdjnnX9fT6uiae6cCkCfp66ah5+5Rr1jOCzEJE9bbMB7QjSQ0
v5KA7iLn0aP7HBwfGEiTlBStrU1C56xcSZfmIq7n0oYlZfCxUs4krwb3XcI+3G5u85+is8rwHNpQ
jXWIN4MKnAiSTa1MA+kR1zXdjCgWI1HICUY/PBUwHt54GhwIK7X9RpPfu2ox0kAVH26BN4bJZxaG
clOgdBSsFZY9JXEC4iLDXUHUot5DDdli4mVpwHitKHJGW8nzyi5QlFPFSMl9FqM+KMsHRTs+mAvw
Mwb1MOc2NQkRDbWctRdZH/OZHrNHaMAVzTYq+nJO3XEtEqjni+WJKTmtP3XtMDfa6BhCAWvqyonJ
udqrPI3b39DwtbZm4xYSZwLcNHNaIxHklHhWgyC8Szp64952tmxUbS/kpCmEHD7nC7I7nrgNXGpa
eLLeTCrocp3pIFxlu2Mhr14DSEFBGyCIRdBPEFkwlRkFhXQHd2DDv7NUgKrXzdexLlq3R5emSI0+
PF9NanUqsVke2e6HY0bmMWbZhXJ8KGnMQEOzwoDD06FgN28zr44GuDcJEaTeR+48SsiwockLd+Zf
Ab6mg32mft5lrD+qbxc0Q1de/JNLsRGJmOcBN9vpFcQTyPJwxEAv5AEHGq3wa9oAOTHvGYx3XwmN
D6Jko+5hxi2/QedCv3Zp3rJHXr4z99OK8F3x1rpuwGD7ad4PVcg6xLTT+bkVUfPNIX7B0cLFmSTZ
KSP1gx37DxCAu0KaujvUitMhNZT8vilN5wls/cs6NXqAJjqDrxFedrPYtQ1CjKkLmF/ekoK5XRJn
ceONcLl0PopNRsIr8NGOZ0eqcVPGRPYpO434a0Gf7MfJc+Ax6YNbP3+HgJ864YZLlRgrbcSQkInK
+ypL8pMhXkhkcy23K/X6oDk31rLSm2nzKGsN+rYRIqcTenHUpfzbmGLvht5dcirbWKRffFJFTR3P
IFqNzioprAn+MxC/rgLBzd+n6F3MgfiAutj5CoT4ZbR2fuBQLaJ1hUVJkVtM1gFY/uH/7dYP1IbL
oEtFOJb7t21QXbPazeBJyqi29ln+Xc6Q/pbm9OaWGGlUN1PG6vGYNDWfhGtyn0rfpfboWbG1oNJl
ShzvmBj9AnugHEbDKP4l4SZKMc1Su/izRgn4lVfoTsRN4G7+FvcyZ5VSuR8EKlXzp9fSe5wmwEbX
3Q1f7UIKDEkLfxcZ8i+X7RxZ9mAvVCTXTPkAihM31fSkUKQk7FqRl6qMw/w7e85CwX27C1gokhFK
A3c+icjxpU8lSQH45ZHIG97BtE3ZxObxZyvH5yUs95MRbRvUy9UvZU3o4Gzfj6jU3qMXntxpa5dh
B8fx1mNW13w02YVoy7AbNflmr0DEbMEFu8zjEoihOmREYelBTqlSPGHH6/a9ytY8/onYOeR6zppo
R8y8/bEaTHY72DMGjfcaPBnsiLE0bG4yo9t5DwfvKTJXPlU2XXyHPhVhUQFFmbT2U9lke/VoiJG4
I5UDOBHpkXRYNgoU0iObuxPnI1pZ3BToyid/fA8Wv0lNM6FV4OdyKS9eXYE5WIGcDq0EcLNJJmSu
9uyHYPN5lIZHhww9vr6Dclo+UP9HoTMYV78oRWhNl9TvXzcM8tmnuNEXI2h25I69M0wx396hRn4s
vbzX3wQjAlsH9wY4T5+T4rlizojMnrzmu/N5Rq13Bv+Cg9P+bpajOnxS8ztc1xJHXSKTO3ixIneo
5VjpdK7UZ5C7txqHHNaILWKR2o7KJkcqK8lZVN9HrEapVZGSXrXplmtPvCFYzYEY2jsmZvQdcLOQ
pKyIFlU6j5vek9QNYzn0FNuIUgO9rDcXurzONWlhYHz7S2ZwglxhcfEK/dnBmwmnikdMymgGuF++
306Fq0GYRgTdQKxXF2lZjMqM19U0hM7xLwjqjOMLLCT7A3MqiDboVxx8bmJ+dNXG1sPXAr9J3Jst
ktmG58oVKYcQUxlA0g4qUOk/oRGwOMISBi7cmnUOy3nTccyoXm4n2n8DF1ifZypphP/g35FqcoKv
lOj237xqASubGVUNJRZ0KkCxJFZGX9Jvtwkjr4PdELN+Z1RvZpucxNTGE7mJASr3vrs8DQ4fKuNA
ktrx5MhItNiEy361Eyy8Fko5G8VfXJOTf+EFhfOM527CtUwgGfsNdNDJOS818tEDottVm08RPsLs
mHpEINEoxcLW48Q88VsbE+Z7E4BV1iSSSbzmHozTA9b6BmZo1hVou5WJ7qmDdYHp3oOnX2rxh0ku
cUwIxLSfni3iKTLaawh4UEaJHG+oMTyHtqPm/TrbSWTpQ6Agqd68SEF4O/Jvc9J5Ugwg+ONJk+T2
EHfNN8xemnaEi4PKNrrii6s9xjtsExwC191WpQcJo0zyzBBDLhBQ/LwH295Ylz8w7o6qdlY7MS6W
A2H2jE0bkRjmeqs7CIDibs8s4M9QVO+Ovyl7Wg+8vLNCZpCMbLlkpVdoPM83BrkqML4Z3GZx/97F
pMnDfgacGTX+4+mEzQ/bZR/o7djqCAfuWiwqlfC518HeRtJXnT299+nRdxYArlwhMjnDBx7BVv63
0R4EXjVSA8b6TTRBWlwsYrqLjH24a3hx1y9BYQ8QLSQQANcsaQrRmRgrk4lED2Vj2St+qlMOFA3A
De2jE+yAXI7Om9fwIUDIlYlBCcjGutFMwE+e58qi59RlX9JB41YNVIm7lQojxwabXIv44MQ/OP2I
+xTH7n4YGiisfjKhr4WfB0p78wuXIJmmGVWf3/7cV5rkgPI55HWWFi0cFwgu5focbEIRrAiJWdqd
1V4JIgIezNN6DCrfOyRv9CwYOf0vagzI2JVgGb5ckhWDK22HLteXgtiBdy613I3P7SQJdWNH0JEc
8abQeGmJzV3t6kGnQcl/0h+zOUJQkExvAYCy8OwvLigm0Jbryej+P4jxQz0fweGpmoTjkLOoblWh
y7Z5UwWxEpLzXHoW5vyzQCV67dccGClzS7AK8xsQ/mg667kauzSp1uDFZOwMaQk+LYq+3sV0QPg9
C7eOgypiVlrXjugWdjyrRfp+jRh2H/ksme4IQYnZho4DMvchVIZVKVTien+5VuagjkXO/2QBoUzW
hVhmGrp0b1/9T/DlCJ8nbvRhVQZE75pNUgCaUEm1DxlSA+fINyUjflymTAboSERx1H1OVLdUOJ9k
EG5oEoa4W8wlwOFed6RYuR5dm3NLMD1qqSp8/9tlOfvOrvujGXJTylTnAgJcDhYd8+RiNcDZ4wwK
oFV2BlPHofql6+vt9mBC40mCcpQXOBDfYYwQ5g7VF3K5FfVL1axcRBg/RfXJgpWGe6uXIsyX6zBb
bb5Rb7mBsoL/hK6RDsOsR7U559FeCfGK8Zh/bqb3ih2dQWKLAJ5AxuLVddyGNP21ersEfLO7Nlha
VsA0jtQConCLyrGe3oqdJw2pqXzxtIUl38ok3XmA6XEMKjjXXs0bZToI3a0AcrJULIUaEuYPh7WZ
17phBfQaPH1xQYIWteM1LVmRlFJdt1KvBGNsGFrwdMOAgbv8A50LIy5871pw9McY1V20olyyjyT/
hoVlYIIz5KAZ3ayBwlm62p+JO33Tb3XYg25B280yPgLNxLP8ekbTABYrjPN0nUUuUEi9rGe3tK+N
tiKOm2QVZGfu9IhOQ+PbsnAiIHmZfKhFZ4eE0Ij/0oUHrs9qetpgLfkYQQie6d0CJxMR4Krd34CF
Mb2G2HJdirS8Dni72I//ftq7Zwd1zNsfL8xOKbFWiuKyuUuL0gXsMY0BKGfbnWkph8HejFWGUVOY
ZsYM4ZH9JcdzhSiJigPr71PKKZ/GWr2VQjdQBebcsKhb/VEGl0A5mPJ8ebhL8e4wMQBG837dk+wF
BG0MJwALPHk7at8P9Q8c+OOeRPsuLDzgg1S9DYmlWh5N92Bh48oInKSq+AvPWSk7s6TrxQqeSiWX
QNCukybi0NxcRVPIaRMSode0KnitGH79yenrDLiIzkTodMON+ccrV8+K4Xjzxzbln8MLjUCh5IO2
vD0zNkPIGy73zTXrpnA+KRLDrpWKhxmuLGYii2TZrFvcF9VSed9taHIzymycYjrrvOKmWbVKOfFl
hZlM6LpCEQx7nhbxPwWkUpKzMde69QOmDmQ/ohuNU9CItzYZaaTsrjnCkV7nXqht9r6lVfih/3E5
EOSlpCo8GD1bHnGxcduG3jpSPosE/jk6WGrdZqriQeumgi0kxb+j7ZlgpQgvEHFhtLBRXAHunE3c
i/RDPWrSljueUPWgt5Xbpr2RDkkF5ldjOQ4YUMQ/p0/C/k6KXd26vFr84zhG7qvreLgHTD7Qsw9/
henv88jdMIXB7K9fHFt0GSbxY2kawnwxcKCMW4b26AObhAdcL4avLEri9FO7anzjGh3O5Wnhg8hM
DkkMbPFTFLYXCQ0lvZCsvLgAMLfDzyR1GY6CKNeH1xR26ApHYxojn0T5Fo2mdGcTiQVug5NrsJlE
GiE9rZ/HpIMxHPwy81VYpQdIlXHiQlslHC3jVKC0H9/Yk5ATA1bCBxQ+P0lmc1DjrZptJHfoOA7A
Sm9YH3HkiXSOWFfX6ruOgZRE61pt9jImgZcTnueB8+45OsyWBQgX5o5j/RWyiGKVPxks8+bocym0
OXhPJ7Kx9B0Rim6jhbFu91yNkkm5uVJaAlLmzr7eNDGgUSigUM3jlStAlC4ox1AVlAHDasSeI5re
ZY/EYzHgcQZzu+d6TJ3gy2a0Qj5KMDcO4MvelEaapH16XQlV155G3r/IRYfI9lujIloPWsKKCoVQ
iqhJEpAj05O5F/XKEMaQMhTOONoHfuxH/NvDmiw9cQpu4uBersSl2yZMtbzQjr9FDhaOwFbz5iOQ
A4Ez+XyNYJP0pZ7wBr3I+sLi2/IbQ5mhaCkCwFASGfx26RDuaYCnuZQVejAuDNdyrGrknCVjPunY
pzj6Z9fHLWFYOQoXsmpQXUSNHV+NSV2A1nCelHRNgaJrUz6ZkLALirEXKez994GxS4fN/Do35wkH
NvrmmUaGt1K0yyGuLBRyMhRdGWMhoq6ED0jMLm1pzf/VWKhMsYLa0QCZbRsLZlASVII/F63AASyE
vMbmDwt49G7KBBJs6YrY5A1kIJI1e/vkOtLsPxV41ixzHzx62Y3kDMCdwsGu6bvmSnhMfQXdMK9n
Ze88Bc3uszQkrvnBoaipU9AhfjJuM3GdbZ3wYOOKyEdR18I+OCLPRcoH24yEONgl3bFtmXc40pE1
qwmfdEMWDS7twgNmRgvqDI8gfn7nu8U4qICocZQVulpoVzqNnKIj+Xy4zacWM3Ts+KVQuMOKwVJk
MGks2X02LYn7Q6sNkiDybIS6AUYicQvzD8dK5UtAmbTHzZw0WNjkiDPZIVR2cmsFCyyM1niLXshz
gNKDXdB3q6cnp8t8MINNk0+CDE40NSRPqM+Fnr20FY/eGgxxRgvhtZPhA72qXpjxNA4kIa2JjqF9
tCOqx+YNKmawY1f7QG2qblDPIeKEc4TwtCbcAnyhwdD5Idi2fc9tm7/mrzPZ+GI3OYMALJNIu5BE
xCLZhvXxoHUlfy8pm7oWIv2GtIQ65MTxKyHMDasQ/yMvWmwWIhTNVNR44i0bepy4dYG9PboXq0m2
kXmQlL80fYZLr3/FGGJDc4ypEDFudbSaOBw5CaCdxdyFM/Jd8mWVq/Qm7pd1FBrFyyahVUZDA2uK
7jdFyHKJ3siclaLFgD5GOSI+Lh6x0TGjqcFsO0y+WKShTHytdGtMEGPMDCsWHMnt6PZIDKOHjkQ4
lsfTrWgOKi+rlvHgFtK+Ob2md20bGiIRijpMteqTWEIgOmRlKqiIqAcYZAtX4KCHdO12+kevAPlI
h15FBbYyUJFIxiOsA31ExMYCsdLXD7DiM+MI7D3KvmTlcEXYD6jNzDP4ZVEhB8wB64lQn5QgxIhx
Nn+Zmn6KGvGHeS8PrvRaN/pJti2EEGXTuW4LSRpxcM2i5rTPIYiasoD74zMVzIXh6ZasUZHBYHQN
GlFqHPvNsxGjXovsdVN8XSa5yv57ZyibrbvHbLYU4Z2krU7Z/wPnPYcI45kPMYZa4hpymYo4o8s/
+DT9p2y7oORctu8mn/IRnyQcZ29twhVd/SmQkj9EGvktVBAMeULuIBXKRA5FKbmZlTs1d8elT6FU
Z8Dq6QqVWvVSXM9no114o7fKui0qqnoTuSktOvEJyRlY8LvbrSKYetVvh5Hof5AfWZ+tMQDaawWP
KR+dCxXeL6E0UtbN/v7tpCSWkc3f/ZD4tmEpGZaEUKtBs1rmSpXkYiMxRjNsQWh2IXMdnSRggy1h
4bnzf6LYUXxL9eBBVv2IEhrBSyg5JWAYxPbd2AzmaLq9YTWDSiRuSNixZM6rPM5muBwfGiqKPGdm
D6o7GrWRAYtgrr1IlCNwNmsGZCWfP70k9zKukxj/g77Tb6Eba7czhq5XchK96s7pNOHCviNQF4+a
eXWTk5KHikihqU/FPE42ecoq5hBw6OV3/feT0ysTXRh/txu9at2mghAtpdlWj1FU17o0TkeEseFp
fA5FkDJhQ0E/nL+VSdS62VDIROKV33QmTFV8hDdvDvVqASpPVIxEnXv7rYNNZCbwnM+iE4opW5Yu
IXDAQZBBHFl2CQ9wdG1aGSYZ5Lvgm4PtOU6eX/26XBXFF9mEekIC9qqZiQLs9vvfWONkXe4/q2Jm
h4jYVIXsZgegRtpVOTzUeHEPQ/c/w8F6Lpn6uc4zkLZiqgZSq+YGirV/gCiJ+XIrCgb/mb+x3N0c
Ik/cFLi4iQsnDtxoC19loyViYy7GVe5Rsx/8HRjn+U7pkc5nS54SixgbDeOFxQx/NNuPBYN9vENU
LiTq8c+C5pIy84y/Jmr0nH4ZaOQyw8mZc8Cgqy0jlTf9JIDH0UW810Z8KHCEUE1JRKaF7ecTzCVB
8mEPQro5o7p0FEOpfdnCDZceY6Ud8wE46viq0mJBx7scBSlDh7aFuKqo1PTc77ZfXXCssndO99C4
OGYjwqRW7UxOrltqtaPgUtfjZkxWCix1jjN8l/pPd6aV2KxVtKcsA1ZaClAVj6lfjodeo6Yu2F2u
1RwL5k1W68q3HkKNW2WNDY6S7oiTIfCqLqpT5xgyxeD4S28JysSAE2mFOTtKMSW7VVadNyxNG5AG
jdc9G/dE7HhtQGKtYBKLKcSqhFYAJZC5jpL0yn7O2GNiy30/kDjJIDBtNQS2u5Bhb+Zn/E7LwgJh
hSGYgG3qrwQEVC2QyIGh0Cr0DN+R1PY0J1RBhJFqxA1zUvAimROfOQd5wU5YgQnjNd1uuvdSkc0q
gol9eHxe/E6k867ue/p7O1k1HY24TLyn09i8W5oGZH4EDQTjwJzS9fdOwDuckiuRFZN0Dp5t08dz
M2Q6tbdNOXilXlDHGYXh3iGwrlthpdRUwGTkqmy727sUEb0ojOjYMXHHn4gpxKDhGKBeCpwDBDF/
nREYtkGv9XW2Y3P+c6ldulO+ele2LTourTC1w6KXqYGD6v9YtHXaLIsqr0wWlEtSRZWhyb2/X0ho
ektsI8j51F054tWu1Ws91Irwp9iRsxTrIZG600NOSbZU8BKRRHulMkjgltfpj++tRMw7WS/9bOM4
UuqrP71lY1rwm4DIz9ppw6Y+5DeAM20vcppxwNus/kYSj4Z6AcIKOtKC60XxkgO/gK+r/hF85BbY
TKdoafVcUtV3JK9eIW8r94fhDlnZKBT8axG0HbKxkFpApocsov3Km/gtJl+WNH8LwoCBatj4ZH7D
VbvmiM41aUr0v1jo6/yXttCpMjKBR9Zm9fudDKbOL9ftjlp8rl3Ahpdf5yhsCff3G6Ip8QXK0bJP
SQL6zi7hSnR19Q+cChMoazOmBT3nEHos2s/LOTRhSjpMzZjDmKjzsupulMctOTW/iW7vCVw9ZUTy
oMy7W3qQ0hyRDUpS9yMsewXtxFpSsSIJHFXAVSXRH91vY3Sg0PoG0F6LRHFecSYlkUc5lphKmamz
BM16x4OEKHr8Izd6eOOqBB+CU90kf56L2Inb46n3kmJrs7Okcd8ziHpXCCZiG3lWYnrsHS7kcvcK
otG1dRQq4kTF27AbDOLw3f0Kz8Ccy/vdp2/mRtbCLS8WVkIiiDsmkGDvDTgqEcUkmSJYSFs/+z//
kzJItJ7DJMSFObEkpcgvjJtgT7wr08/jc8Q1AjxNEof/Icdsg+4PK9Tcz2b90f1qii7SBd6V5xoR
0XmJN6fgwDtckp5kgHLCGUnZdmsVQxqs1DmmzTtbN3BtWQhLEn0HGZJf3lTqTrN/TiSmrtJwXWP2
x6QLPy5WnypI3hRz+eXrp3Cg2DQcGXFwrPP2xy03y+2HKEzS8/MsIGIDfE2rUz6EJrLHe5nK46bw
NhWumtdNhGW0AH2YeriUZG87cWh9bYxU2wW8H9l1cODoRrw/ou57NaMUnYg/P6VfcCLt27JhAsZv
DBUgCxuz2/B35EEjXdtUTri+pu1s3DAOxiujKJl7zJhd044q7DvaO0H3yfzyjP3X5K4OSL+2MvyE
NtKLb+SaOZ0g0/lUrdAULyu1IL9o+wHfClwK9g37e4BRDnO9LtwzplwVk5AJsTaMPBSTpnzfiI6s
y/TegR1k+5k2Ykp16Kku0IZcftTPHwwv6wHNlQhxnmEu7XX5BIiO4wrO+3BKljFCZS1BosZQbEJn
GH/aPxoyPRjpyxa7J4f4TekTC4owfxU0o86k2HFVG3A7dHFu9gJBDfAoOUnTfRdyLqJ2dS3J/pCy
dnzEXzn+UwOaBB1gbabIT5WCQIxWjH8uFEjD3vBV2H1c/05OCnh16bS/uDVMcCg+iBmE86fhmkew
cI3UO7YJtgMMNaqEYzP9+LDDdY4ULSMylWwr1YixMwws5HyogL69V1zFYB4pVddtlrVrpML0Vw6b
lmSWHf0zoqqrGHfIkfdgZb3GVagqtShixtT5BSt87SD3uRl6cnebb4VlNkOdhSgq/l7DZsgtt4B3
qQRzkn/EAhMTPRG13O3MaOqrZwj3zZeQdhY7tNC+3x7k0X3FY57Cuj/cgJZ5x57Ri6FY7gkP+4Ha
sqhlR03ZMhTSnaDgYQSgvyM3fwtUCEYoyNsxccd+0ISKwH140UgyvfDl6tHiwHG2tEh6Q64qLig0
s09hNMMSRU8PAz8OGkSje38elqb3g6XK9D4tiyDf2GBpauIyCZ+lGmgCC/pAROspWKulnkBUCkuQ
4yXI9lhnbvx3DbKOdST/YiUrNcXSMzttk/mYR5wWZwCcTKpX9jkZIU+5BK43VG9kp1+BW2CFPc/c
sfzFARg8A4kmdQa0vDRfmOikJFgBc0LGuSEjsBPKEElG9NtOpoKOPFjThpiW/1Mg4NYIINzcezRB
LhyFOvny5o9AEnyrrUTs8tX31j5jj9FYvvpVodkVhINLc2Qt1roy7AfUjTVIyUcR4SXxszOMtrE2
F/SR6nUsbRRLRfKYoyxLos0fcWpsyJAPMlS0pWkOla7I68Ax0AXzP+IAWeCBPKQ943naAPGT52Kh
dpJeY5Ndb0nmIQmI/Ja0cHaRJqa2U1Cv/jEnwDB5UrnYB3LtTfe0SOtYnKOJvrcO7PHQSifs8yOo
VCDoOyxVu6agZAOUzZ7t442/lwhY+ZlYarvUPNoadnX86i8Room7JLSeZwDHgYGT5cph6wqU8lgy
7xLOjKsZWnqNm/6dfpqlKF0obzp+SmpBt2UwjxLQyWLfZqImAWZe5e1AbNdGmafnNtxq7npr0fFg
QDuaT4mVSrtTH6+YTV7BlrgCaNfr387ndZp0uWaR9c4+k475aIIIJH+VG3zvJLMlR6TZZD4KLq+9
IzXDWXSxyes4xwR9Hd34eBIX6Ez0Lo15+fIyR+s76w9LtJ75eUEEEcyM98PIrKEg0xUtGwemTnNV
/C+dx9Zagws0Ntx+5yUc34ERdD7bPLBNDKXNwoj41EJEnELMxWpEjtW9J7SBi86Gl3IBBvcYRmwJ
lEevlasIUTYBmCuHdtLlNuVDcFpHlC6MaWvvbxOculGSr/TPmVvLSd5UXnMRJnrNs74XJsPzfy6a
AMhdg9//hPQJQNj0YDQAm5PGWigbt1gJc//U+hYEbgf8K1kdcUrnGfEE2GWGZujSeFXP6Op3UFyI
jINfV68GvkgfT5avyVMrgkN8TEsO950aB3IzltneAfoBz/9PDX3GN31WzFaT92aTrSwW03l6JFQT
tCk+/CadmdWnmVw5wSmAlrwybOOsrHSg3+1TDeAdA7pAcpeGyN32/lIg6bxzwoo4/FJwxk2V73UB
07PKfBgI/sJ2yrio/HoqksLRe7YSGhF+vU4oiszj/IGYXYBVKh5DwQK+gYEW/YDt7T8Ue8Qgwbol
2VmdRsSLGq29whqew5eqxvoveXg9Di6p2cTY6iIlnrAkgmsgCijSdWb82FVSAqNe06gNwqZJb3kf
RhQxpgoFkSrhOAYl8G0UiiS01Hc6jagxgXWnKqqfNIs5reiSE6R9xOkeYoIrr939dcf2FegQzQCS
Rggrl4OIM5+nOnxzzz+rnNO/gq9L39WG4ug3IN8S3/vA0jzzO0PxArZKWWsnnNYtlSL+aJ6mI5+x
leQ3MNyVaGiMLjx6V692o+2t1ejtAVwiqq0FJAe6B+fxPiTBnfkp8eF/Y5hEC2lRO7fIa5Ym72CR
gEz4gkFgoRNVMKvSLcddUfGJw9/6VW2ZFuglmbsKegS9+0+cBI6N5/mXJRgv+sO9X+jwUsZzxeid
v55KaK6C5J01smY+bfAWfdXCkqk4Awp3aNIY+BIapVvkA9lkfNq93nX7ZsoytHaVm383SElF/h+z
yn1f/4OEjfUkyUzcNW3VGnBMJLuwMmE32V5e6WiHUF6giGzumG3SIPgcgyu4b+nzhTGPfEutqauP
J3TIqfCJIIWNCt4yEczjWYDwvY13tAzd8bWarfu8E5apeFWM11AUeBJv1a8Vrc8psjXsUrqah6c2
XV+9KqHOF+wxcmQUX3BfWlHvYa8gpT3dI6YBtdAehkaCgOF0MJQT76f8caTOGXzOzEzNGNWKWcB/
Jdi8iwKxnBNvbR9L4m4FWcSXeoTHYxC/BGryIIHk0I47chPunvcFy1TTOKm6bO4r9xps4T7PYGVa
7PHr5GsIsOBFjJJJx7KTRgLITH6d8CMZw3nlOUXorNJXcYhmraYEhGv2NPMmZrSuPoIDzu7T2KHc
y8uzNKPERr28IzBf0lHaHlHsIqQqEFtRroSabaABePRJTUz6uUKLTTl9dzFvrrNbb3lgme7gvy/b
WuyhcJmTcj9lhZYj2FVuI8zkLYfCZUIuApNovYkAdgeZ197lsYhnD0IRKY9noPzTG4YsGdQlCwaL
XK5IV1KxEbaRCodmhSzVTpwyfW6VvzcTTLMpGL6nhZQ2xAPMB52ymmnH8Rf8SoObPXMCrf2ObNnK
BJPF1Nc0UBtep/HiYOfM6isvxMOdKql3WJLSwU/IxxuQ/RS/axJXQaN6rnblCsEcF6FAGayu1Epk
RKJDibY7KquY+TLdGoC8B5ZeC+0JEpPKtZMksvEaS7EWG2S5jqegDYTqwtaMjDEWDoTmIXsZCLZK
ZWjpUHy0fLePDMEoadPo0NysvVQeiJYIkrz/HvIUpwKubHXTonJ50Dit2+PaGfcRqQRb4fBB/bzh
cUayHRGjiHE0Zd59HcwxFye0DgVCnPEXJPaf1ohajXScNFqTrfLa5nKQ37fohjmfcKg6O7j7Ck+P
YziXU9wqa1kznkI7kkZZxcgcJbj0HKPx/clbvl6SbXPVJCTvmJhHOGXzNNMz1BkXdemySf2IUtbO
SqamZ0FqJkw2tfq3riOLZh936UWgAaWNiXi7F8OonqBbWRVaui1BdsXU6A6ZI9GAuyG1B+T0GsAG
bntnRTC6GRD+wKswKgW9Jqj/QaQqHu/WI4fLm527Xx/GUVsgQulFBx1AMWEsi/A0a/1/urjFuQRq
2UtCMYv2pka33ZDolBOa68Bva4CQku8SAd/eQe1lfqNxKQ94sDjAOzeFkJthn6ruu06O64QCGLcZ
W0vMfZMNcrt38ZLZLObykc/cj4SVBRUWucnsx1Dii93rcFKki/5PY1TsTxWo/7DhvUtkMx6IS4P8
L11STeBV8mWJObdjAt7P9BwsKR5aig/v2YNMncAYvWmPhppsUni1v5Q8of4zvoj3IDg5+rkitsD6
crN2/Wnnqr9P495S7PAzq3o9Z9UoHFOgaadaHAMtT8GyfE3rgaBxU2l4NatfW4O1jjIrcwbHkmgz
+Flokpraz6Qw2SAc72h14R4k6GDm8563za9r0LCndMzELHwCrYfmMDv9Pw1vubQjs5pYGzgboXKS
yIW37TQpCz0vkzsqpZF1wfQPc8J1FDDzvk6KjRmpagqHtVO2+6VoYo4iGEfez3sYL2ilLCGJrnza
AucFerONiC//9JxMf3q6TjUT5YNYGnWx+qtEPZOI/jblx19LLHwu8GxkTMrgCrjfy04tQuL4lrkZ
OgI9BPDhZvCqhA8OXpL2AKLEfHQYFZYUTC6/B49fKjAoqCAJQwWcs8xMX/didYgSqlBLd11hjGQy
ZU1/2kpx+IExOGPUdx4oFoGM24i3/SvalLWpPPmkqIJ2iX+PG65+6GXE+33FzVI0UV0mLFqSbdh2
+Fw60S2yttIHP6fZ9fYKT0U9zPNoXF+3SwnqlMOO6SiRZtmUygbwlN3L3kTim7THJlXolznXlpSx
x8q29W0YXNfI93DHLQAKgQAk4mCPIO9YkRa+3ZCYbH9PkELHvHn2fm8ZlbKsfmay59W4bKz+l2RF
MjoS3J+Bk9SYFo7uq2sSZf8sRvi1uCQxjAbO5pxqA+W2RrP2PV7AiWsbWw9k+SI/wgap6TMmLyaC
UfLsV0MduNOw3nNFYfV8ERfnolW/gxSyMRA28+i9tsNGvup5kc0qTqVbSxPW6ow9qRRBydf+0oaY
sLKW9NiBWwkUll/6s53cRSbkSNOmxFKdQHvSg8I5YOn0M05MjUx6xwduJD0KjW9gXAbikUuctYuZ
GhCoqXzAMXy2QRZw2hTfv8oxcq8/otNCFL6Vvt8QHNX39eujZtm+r6c0402XfSNUNk2sJZWDpIoL
e7yez+Ws1LhYBJ0ldXLCtJ1Sjvv4Qc7/ROthLrbLJFqNznQgZyg297mqtFpsiNDH7ZnAHY7Ef5Ks
HSSHTl95XiL1FXXFb09+aTFcpST8uX1iGADGjtwW6xIcedyKYFg+kJEieZPb1T+vFdzzXQgRXpy/
/7IAprq+ruvaqyN8O1Puyi+majFHqziiI6p2CQhO+t2MDHaJgPMCWvifGbbEUMq7LCIufGxh5WkA
AB0uh14OXaQt2AgloAwxQmHWu0X9mYqBwawcEKAG7QyXPgk+mQVLQK7NxaCWKtML5fVLDEIpbeGG
4eaYv/h/AJZk/z2yeWz0YpS2eVAb9XmV5A0jC70pUsfQStubSNd80Ili3FFuP7qDTcVkJ4P5KitL
Y9xaX1trqB8DhMXKWErhyHRZAZaiETiP6MEJd44b6TncVGnfUnvBCkA9ThFnWrxEYO7Gik994noS
a5JQBPyH2E22sokBEQD+bKLCkbyVH+ksSnjzEKGV0zoVb+O601utM3wZPp7yxc0naTpWchggwRbV
Q01zsjEDzwbkUVCsaaCT4NQT3uLQlsSB3Jxe8Owey3ZZmWS3aQRIn8j5lY221wnRmd2JQjGn7W9+
E/2TGJd1DBeJAUouBOJHIZYJG4zGCopRAW+J7P9YsHEuIuVmZOcTnu/zPEsYrmOSoi0YJZivmwS3
eKwuTlDDT1Sb63HC9U3UjLG2LyIvtcEOdMynopQ53bw58IY4QfBLyWlorYaRmZurv1OUC0EONjFz
cx0kEzxo4+JcOPDdk69yDtDUs8OJFu9nABY9KmbSqQagSRGJdcESbdLxkPga02RSHT6yJOsDC7c1
ufjnoGgi7ItTQyYpkh1TESR4yRj8py/hJ94bd8f+cdEOKP8IT27Fb0UvXyvFtvJIKQBWppUk5TWI
1pPLOY3dedoRQDjj8e4zcVaKagaHRenUwT8wvxoqzsQxsgzfFc70OvVRPXoO+Ujq4PqDZH6RZiN9
tC+vd0BZLiIlNPWmF7SZOexqQYo87GtSkcJiPo8sW+XEh5oq8dIF0reOXGN9lO74YpWVvIGiT8pB
QbGLdcgZhxqeqlNIfzC47qSeSch+3yCGwovUIiEMwwDv+qBtaK8wmiqfWz3v2qOtxzFb7QTi9LoG
RVrzJQWNrUSN4T9G5Z6aUC4hJDd/xkanthN8bzRKenKuS0LJKxdYdS7zzJP8sXZlATiltYfvz9HT
Nq3esrp35Ol+vsa8qVxy0M7OD1T91UJEtRt8VcRugjPwkRb5u4/Nkx4HmH9rb+l1/+1Y9/csBRME
fYOdV2q3CqyDPP7j1Sg363V5rcOs/gExikeAyv49vyMtrg4f/Q3m3DZM4O8vb9+ZqJvHhoImes/4
ZnnzgvwiD6eUBtPBjvgVSXBlfFOlrSNAgQGDRW0fxZShDBhv6gNEqbfg3OpTzV4HqC9q3jn2mlHy
hsPxl04ZwrjNB0p8boFkPdIceF8vqHDi4grIuz4hNtcdEuXi7dgJkVFdrZgntlija6cpQcpR3zN9
p0NHoFIYWw6p5Ow1PVkCEtezFu9+Zv/pw4IFY8wy8k51XTZw+XqqgqJcqr3wK7KJBte+/qhFO/FN
Q0SaCYbAjjb2s/IOzqMhDnCnjwVmszAXa0JKQb1CIxHN7+tgT1fGinUj30ymWQH0E9oUCPc6bUaW
F+7gujdMuPk4140lNW45yLS4bx0K+cJirUWjNcXTIyfOKyPQakTy2di4zENEQcDmYrm1e/Jihsrk
mqofCP9/JFkgLaDP8A1TSKWVn7DfF0SOmqh6emde6ZoNWoiDjKTMsMK8GS/BomTorZGwuisCBTP2
t9TyHyHBSw572EZTfUMN4P7IY7X+iaovngfobW3c3QrSM1crOXqor/UDo7jtm3fsDjywkI9UE8Sx
bSBmDpdjRbvoVZ/mMlVoIKR3C7tHk2u+jc4F1eomu6fIL9FNeeZhhCRhl2kT84Y4V8Zo6rw00FMW
spXOC5wBVaIOAD0ITffGTHvC6rL+VrSWKT0feCyXB9K3XIOinkCaaoHUmsR5tiWYJnRY+9PHJZ2Z
EN2MkdLi7Ckeow8LpxyDKelrAH78NlP113ihI0+BMSme3t4Hgus6H3KPmlkg8A1FdKLtprf6DSAS
MJ09lBFAbLLXN5qRBH/ZAMLkiAwkUcTV5zapXh+FiIjLuVT7xt8ou04AZtv2hHH6jwJ1llWaNHDf
2z4J6xrf8BaI8lR0SDMqauZSrQEg/JQ8SkyNL6abO/G5WFWeUm0xLqxlLMcEh/1pw6LTNJi01iVp
N+giGwa3+EFoiUzNsdNtxolGROj6vYh20+WQkutCw+pC0iWMTPzhucTl2/zswlSYvm958P244iJu
V+bqXh2DXyKlvEfzybdMtKGotV8z5a0lKYIQ1Nk+sRbP2N4sqV/M3zZq8MkUlsgdjfm0kK77maVr
CUHUIBAsgFHlO3H0IjmytDnZCKL4HOqEj+l2bb/ShdZuVCAIiPSGpCMdgLqVyPL9vlz2Sbs8/6Bw
iwcLXcUVKWJ0qylU2dr32vd5YFBhTEPyCMjw5MQo3S7Rja00zHj8o3+P7MVvyK+zMICkuVCMhn76
J6qNF82pwQMalQRZMENxdMbPyZGmVBM17O/HVbyF+/99OR82TruoNeraDydNDajdZADXzVFzo8Jy
JIR5xlsq1S+VDXzV3I2KlwFQwm2/a9BtUtul+sLiKugk8VWGc4P4Hce7TT58SicXLEDMoJ7/aM15
hjdNljJW06AriF86XL5G+T1egesH+Qud4/6puasH+0CuwjMXQ7tMFMreroSoBH0hJBY4+4IbF+wX
D0mhhX1Wfetp71n2VXb9Zh/cDc54mrP5abzuqR01xV+VOAY4YNSHqsG6ROTAxQlZqDYBV3yOrYMW
0TcpvtF/5zJDDn6FOIPyO/QlCol6Zl0dLNVjKQSj2QxF6DkUhUuq1pKcHIjpQnE6ovygd3CBx68D
aZbzb/kTnd3wGyCCXsrI9Cuh49g0N65u0O20D8ibi3FrzAxg0rj3861mzZwjEYgWGVhtW+T1GJ9l
RHfoiLFEeSc9vvWk0Ygu0TxR8b990ugpF1O+S4vkO1xAC7uFLh/rE7kbEM/0ZSFzpevyKvmi5uHD
McKzU+QnYLVob3lnVW4MJOfNfadcWutMquv0wZ1atltpDlTKBN/i/zXdP4t5TTSIZxu+s5MRR1VR
fmHnoqLs5pSZktsLy2/4uHhr/y6lZMjdKsS6KldYKNVDmKaos3eqOjnsDVqPhipbfMBvTNbC47cm
VmIqxEZ+MjbE7zNBLw4oLdQvuGeg3iQArofjV/5p6rLhpp/aVSCt2uSk6oY/ybi2sL0UV0xVTdZ6
6myDKmorEUVpl2ue/7FKZd7B0v3ruWXHoWvtsHQwcfRpjmaJxk0GuImhUcNsMGq7V//DPxJfJ07z
E5+zZqIa4wuqyTR8ZBkYZqCu2hCTZTT955wVJbRZAFDCGYahkH5wdBxxSXvK0ctGrdeur43B9Y2f
12NIVGXJQmzK/EA4KCl2Ne3BHIjOuQcP0IyZpqoo8UKi+gvmFBpjT9hT07Dd7ciM5y99Fh/dtSfK
0LFpXsQP86kAzUxn7kJn6ewZFTJEYOsXfkFwFQb1fcVQ7lBDzCIaOYBQ6/NyQa8klM2x5S48RINV
LnswugLK0YA4T0fm11w/GolfFKwxUf2BK4tigHpiqU+Dw8oK4upe07dCd7B2FGgiKO9ZxIddP7hM
yY94LmaUh3nki11k08z+VeZRRhC4LF59wL23qDccBujE6n7pPmwFm/e7TPKxZ4ZQBvP4yxUea1Rg
+Y4isZlTRXVMya3y1WYbpcmTjLmL5m/kzoc8lh4mBYFUs2M0/1fcMgGT+YyCxMnVZbdLy+jGWPWZ
UJvQ9QDkL7AUEPmHSGraT8J5gl0ymUCaKx9/NKxPQNPCpiucqfU7aT4cqpw3Sli50edc9dnGdYF3
x8g1EDGucUwpPuYThujO4pudC8eq72jcuvA+d0zXFedSe1eMCBThVWmgwybv+Ulu314CegYol555
8DyYXEpmYX0lrRMcGTAYKc45PAJkUBnPGeTWVRrkz66AlHRDozU7Shbfzxej04+6rj2DShFAuxbl
EETLY9q31yne+fhlfffeCZ1ZcEgcwclooC3+9k2KyjwGdysEWtbxHPlrs9Nh27MrLaZgqu/vdCPj
u3B0zea9w6nKT6e850m6YYKrVoSOMJVp7z3n1aVLogxFAW2J0cFb5t/H68qj28ZsmjDaqxOQJgLm
g7LWu7L5P18WTvh3Qwf2z1hW0Cc1/Hr5JJ/GyjBnu0WWeOO758GMxuJvpRUpW5SiOqAn/1+10kmN
WNvOgyAqxmWJUT3+qd8onD//Intgrx4DWIN072rAdqENy5cqnG56mQFd4sOv5UmnEY+Olxl/LwmB
fswbhWOTWfPSSf5IDCQnMT52nKU3/a0g8x8Las5IFkahChwvA2W16ySdREHptdRKWaN03DJpPKwW
YVE19PL5NYTUBiSzujemkTRYiLlkjD/nWteLKlh2DV3lokX4T3vHQyrtQsBh05B5L5u6wadWGV3K
nHFgHGtrBw4uiiMTN/F7zccLbHO71et0fb55OCBSHTd7/HK4WFzHxouXM9d1g+wCymPQp+qA9UZD
srfMd/wZ0AxYDPyoJPF5ld1HAiXHHQ9TKY30WGWfvRQ3F/bfgDNUobt74NwM/kf3PbTLOigqojqY
mrnxVtk4ExQNpHEp5DvAqJiNYHUg/kNNpOrLLkUsbfOLvYSJHBupDrhJmbodCnuMG/w9Er4XBLeC
CmPNXWsViLUCm2aTtDZ3XUyq7fZ/3yNcGXtfuWVtIiu6K+LSgSLPOKMj0cQAW866ClqapN2CMNCU
h0dCG7XOSI1YaZE3Szjr3DECM8wz9Pwx6+GsPLZDZZDwpjSFj6RbrjjsQFMRvTrLtwptPBPQMfda
3NtCt1lkHlvczOskELFAtKeDE1gMlpNTVXeAKaHin6QTPz07Dx5yS+QHoT8trXL/kbWpdex7SL4x
J7L21ep4NzsJO/ipcbjAJHoaWyMN/IqwH8rPmXoTTEH6jaiZ+pgwdZ1Lkbiy1gsqjK2Pxi/Vw2Yx
Ef8aJMCdgLR9lAaezjM5TS5gBeVBwfglXJznxwoXEgx5KKgs1R1NXucF/WsjXqjT2Z3Z92NZOSx3
rlv4hdqMMbt3asvuum7xHWfYf0mC2bDkAm95oKee+jaGaD6tNPFRV/ZO9fgY9IdTrYQAF01zniP3
WXoWWdww5s9nhKD3qyEnAGF9o3Pj8QP32owgPZx66/gZFg7BpQotN4FiYyTe6z3nW3WcUs8DuXyT
SdSkx3wJqWCUzcA/HfQP3+6uBmaCLNZjyR2NRMTHml+7B7EN+3Xyz2OQsCvKpwjVUf43VTNJB9tm
dL5IbqPw6XSnD015EMAuQ/7sOkms0I2gz/hPWjPQgGUEF3uENQ56LhxUsk6qEzC7ynoBzOYNE6b5
/d8Kln9IUmDgyt7vTLx4aE8uWL5PGAAFx+H1tpUKOwo/64/9d2bUrIx82y6P9siDHyWkBBtbCN/H
EkN1gboHrugjcryo27aT5oVnM5aRBn4MmgHOAwED4DMeQqLXwyt7m2chkPRZT7kQ2AOJUxk+nlvY
v6BYzGjqECyH5lLGR3bo/3rT6aI5hME3h1KIPD3Y/itwzHfKAGjqsbJiD50O8ITF7IN1wCuahek3
twzqTYG0DBMugCl/jBuPtf6CTnugDSOxwFvZbHr3NjQN95Wwn2dxKYe0SVRLkJrNT/iWF0xXPz2y
wqh6ycK3qBWPi86qG+MRk2WFASFz2Wm2RQaxqxn2X6Ql7jKiAcORr9qRxRW43vPwnTt4cdwD7oO2
My2G9tkrhOX5svG5DibHkRjZpSRYwgWQJ5PWRlKVP4t+V5cFyGkTMdyvrUCdC475g3rBC9GTkxLO
Rni9O2VX3Y5EC2AycLtmA2nTyktLeCuz8UrAIiLWpcKKEt2zdljIk1RYxJ874VxS0Dp0W/Yn4GRE
AmauwTnc8dsq9AEwRnQ1NCFTQTfuJL3QeT0oUbyOpUjHOt8wl/Rj5B1argLUpBU8Veqg9gQ+p6jY
jfYo6a5tX5f7W4TjuMz2Lu4KM+GTZYG+xhq+efeg6alAie46s2qPhiU79YyeZuiKsYolGYH2Wl1c
NeHToGzAInZxSPsH5APellTcOnv48IXxHL4PUrVnLJZfJLvclkKaDJsyNmSkkAQ97cdKkYLSgUEn
JQzEwIijtEXtMtFiLexGX66xMYjxFfE6TL8IlMTUwXY/4SBGvbQv76Y1/5inYMKyG8l9fi+0Jwem
XEHHY3/FxmyrkKG1fmXAJXE6PAUO6ZGo4+nCBR0VZ9sVD/wA3LgB30zDe/eGNeqE9Vup4dqC4c3l
V+d2qYgW/lpHtExoJWqLOtFSAntqwmm790GppAVX5eD/eM2LszBpD9vTCsqWpOdxtOkjVlT4JgN+
KJB0QlLUO5nLjRtS4yY7vKvOWRdHzFwc3PBZfA5onoCQ1VxO1b+ag7oIxUCCZBcznAsw/muBdyBT
gfBtNcTDhszhSx6EpzjgAQElEjGrG/LEfU2Ganu/KNId/ts5hMJVex+tqSYy1PRyArHsJ8N/DRjB
xJ2y92+AyLI4CLuAXO7L06N4rEM6XkAIUVsF5jGnd+RQzwm2PschklMDE1oI06lQfv8vQo0Ds5KF
Wy/njF4L7evHQAmDzF5fw4vy/Yx+FLAE78HSKxOD8vKUEv1CenUtRpLwrYzTjzT0ZqOXIe0x0uKx
b4xwuNcgDgJZWt3V40AvOGBddEkFUhj7A62P1OijIzuwgRuCgdaDoy9hTK5DCutdnCXEn4ckdOwR
nrmXYZ+gYq5ZMWx4w2TLBv0sBxoenJnktu7nK0t7kJGu/z95I1rUD4gTHlQ6mLiZHrwrwg4/HxB+
iBGG6+QZ4xX5W21PScSNjSw1CLTvcPgfI27ugvYrepHXGLSKzoyeeqXik6WhjpwpUUV6ZeY8a9jO
40grrMTncLLVQGVLwnBfZuIzkTPriL/Pe0mzqiTvWgKCL+gCF0xgqmg7k2VB8K8tQeDAn4YlIa99
8WVTpNRsmHmlHQDJJ8szgXScVMn3rRXNO6OYnsZlIlFH+ndsFLY53/Rlwxo/U0DDkG+AvpRdPslU
gQJ2DTxhpzz9MD+LoP5YjyD27qMTL5O5W6G40lf1GMj8BAeBJYO3SBn+HZN8ZWIiXIpbYO5vTjvd
X5A+Dt9TVqQ72+XNVtBVOdBTAOTO1oLc94s6VN2lMqh2SOw/GMSMctkNODxSSJp+jdKLpqBTbUH+
rCzsUj42PlFRq332or5fZs22rYSeP4yWyFth+HGeYGVkYhp6ii2T8pzVkIuxnvL3X8IIoD6mPyDO
M+jYO5Y7SPcpsw0Nk1NJ2O+B7waogJhS1b7Zk/MaRX8r8wSElcHh++kR6kaB+ynHmgeQ5mSFvxKN
cp3QMQ2uSs9C/MAfW3aB10xPMv2Gbw6n+q+rW9UpqzHx4yimIBFATzjqiycG93RSjiH3eUC7eFCM
ZcRzLMiV+pIOuaHWbB3KzQIJvXl8Fnl6hhxu4slf5mxxcEsfuxskhYyJ3AhtGq762QKKTfhAuMRz
7Dpq2QDMrZiKMdVy7vMDVOoMPbfQ+a9fGlMVBaAo1Ax3LjX8bvCeegHOfQOlfpPGvbJpP2jnh+wD
Ia/Ou4/OTQuLpKt1KDi7YXGHws6VLbBs/5jyxIglBwDgGoLg+h7TpvSotlqJm8tsdEJzpTc4/par
Cp1g8NQcMZZ+EhX5Ldb4UBwZhIlkZ+PYBqGwq4nznIcs0eJm3FCoZDOObhOBMXoarRDO+MdD2fsP
2fvJlCvPE0/nOIOBvRZMgmzkr8atiDNvEuPMs5HcH+4FJi+Bjx6dkkQ9QZgm7mqolIcoRRnj4J5+
LsuurGsqQI3LzH5waJB8G0LzULa5CcxzAO7CAB17V6qE1f4dRiU68+YRyGXpHwejxT57ybZB4Ndf
gt5G5Tw3JHq5Wta84+22f+H8G5C1NJzT+1qK/HHxucZS/LQpa79koIgsWDC9sRSz+kjL/2ecen1P
G20A+ZWhcp4yQDyjFMpfyRWU15Hkxagu6c7eomWrRDk6QMpSGuodWyUGhc/0fPtDcgPlxaamppzP
a34K9O6Nu6891gzeh301hWeY1qnbcILMSJbnDpTAy92Rup0ksYYAn3EQaKjvZdhl1OsfzpOPNHHc
sjpYggR69253+HQv9Ith5y54CYicEUvznr3q1+gUNYmt2Vj6m4AubSgZoia5Yodb1HiBb/ST6KR+
2knfwkxY5wVdFduVbu0MK9Fr55OhjqCShDYRaMuP6ul3rl82yISSstY0ImThedZH9eNb7s9ZEW4C
oUP/Fa2DFvAWwt8xPh1tlvPAY5+VIh9OFDgUcsYrvYwxKDqmb1EiYQ5QdVji1tzwkzI7Z3+7EeB1
Le/KoHJQWmMwhW75Pa7OoHi3aD4mDqzAQJi0q1G2kjoYFu5/UYQMhZId2MKZ3425jGj8SO4bbdmB
tqetxx1a5PUT44BOF/dQBN9/cK2/dQ9MjnIQvMOT98B4tepoRuJ2tX6te2OFH3WQprmO2aDBuMBo
xtqIGkW8r28TLKlcOUV8xexzqZ38dhxqQqyxnV5QJnSh7ylcwf1W8wdf0ecqUZCCbdGdVipOD6GE
PVCjRzI/jKI/h6CfEqEmd63VV21FhY2Ou+eLIi/MscG1h0nBMWX6BDoyR8GDu2PDXPJ9eUmLz5/u
6gAtreePI0JdkIWKdaUDXIy3c4K50peCDcDzY/+vEOdLljJCKnHGDbtpiyhPD+dHRmUu94LI7KCa
NPJJ+AzjekjpIjgf0AopaY4sHQRpa4CqO6ZOJLjEbG9cBN5GICHRN5oWvr2dxChSV+OTSwCDpot+
fXkkJcaJWme5GQuWXcF8HKu9c6/QaRxASMfbgz1MlDMf0olPSpWsqcbhJt5pNtC5fGiSe0BpCNLE
e9TQ/dyL2rpU6n1Z34CuFQOrz7SaKPSvhgZUtRye0BvqTsvH2nZ+RyOugA8FSWP6ZjlwEsA/bDLx
JU3PQMXG8gkOdNhhu2VtSKe54tUhNNE2ULHkaSTUG8Jl5z+DAhxjQUjvOXHm/+e5/ozQkyPwzCl3
OqI5ykg3ezA3pJkCBET/21W/OwHOgWS46FG3fowioBEvxnvpcaEUI+zNHQl4BTd0BxruYn+pmBp5
treMtYy8rFqOj6EyKfm0nCuCiIf4PmxdA/RFrDJ/+QJqOF4XUB17k+AirTnag4eo4kRbV2U4qJ5p
lztF+p8gpALzc8BisDqHg0wvMVnNrIhFwt9iRlmCCB9jgO5OsBTCWKho3+PoX88LZnWBZPUWkvcY
z/9Z3bI1nMiiig76inAru5ApdS4E6JjenGDiuRfRZHehZ0/qe7OFfREprf9kHhVXeXLsBRHCSZiM
oMFnIPE771fFFBgmPLKobrbOUkIGNa4dctbmkoRUnsVXnjQ0bC6eMv9rdGbfsz43K18rIPuFmt4o
RbCFpQ4ljtQoZIpIFYO4FDzCCXmK6lB+JY49JCqBNYWppayP5A1yfVDpVvMHqvXRaIya8n1wbdRw
aqf8eJw3v/bxnASPTteSfbN0iN+5qAh/mbsvSawwouNs2EWEUYGwcmJboIcv0aF0xz0MhSAdKm3X
s2RvhygNAEy6lZfel3yza9TZfgO22xbohCr3a7JdGXFJTZGXoFlAbOjUquwBeU9VyjL4k42114sZ
vRaPRqbngnfk8LElKZPFbPpjb2D9yUCE0owFlKIxumxxu0vyp+9nDD2ogtg3R1OPbBIn2LA36wYF
vXQ7o57DJr5s4dXRJ2cdURR9ebwngORrv7uy6GXBKiDCHIajVwHrF4UfzKTBZRlvcNI9OGbSuTZO
s1TNAPNfdkhDma2R9xe8cSymSuiP982myjk95SymraBGX9uNFTykcjQ0ZLIfqNeLk7/Tf+hv9JTT
sGlyZHna8DqpTKDpkb91Z6iPdrjZvB+CArNN7rs+YChgyg22o6e8X3ghLSSIjnw/AEHut7LHXF0D
e85eh170aXna9p+u8b6o5oSCSlanUD8HxVGj4H1YO8tcEWxlVppk767MfM/skET1j32VY+nJecZx
XfqEx2hCXD7n0cK1VGYrVwSujmYy0V536IG1dKJVJSdaI892HKl2lP34m0D8O1MFSY1GQjo7U57V
aMUu6l6yZD0D9H5L60jaMIlkQUYj0wN7H49eOlqvzE0wMg2DZ2cxwUEPW4Zmfxf0HPxcJ7A+Ui/l
26N+HyUyiQGg5SCYzcvt5tnE2/CTNKu9Xf5hDpB6utx4zTBcotLL+/SFW3zus1HrjjzN15aGQ/3d
c3Oiqpc+19J88d/pCkFyJ7DFNG+skEvQwVsehyLpVejYty2zC76PjWYP4J1U9g+sYsmM9CCgysf/
R0rq+mWZr5/pqAVdHXoxVX0dShgMzRXZIE/OAF4K1dWV9ETKsycrlS9hP5buHWSEIAj4HpVBgG9H
PfxuU20IQQzSvdPxL6J35zvcEdgqaPF8F3gKIY4HxtYspiJD9xzuzDolJtRw7XJ/QV/aK6faYOqq
o7utkhfMw0ShWyIg/BcB2EbIBjE2Z48HhCnEEMgi4+VOTmgi5OcEFRHDeZXa/EGyKietpyCH0wl/
FqIfqEDoHQRpP4evp5TYl11lQg1S5fjVb41iOF69E4vvC6/QEx7sHAI3ctiO5nWLmxRqMONEsvc3
6iefCs5XvQD/WXIXedWkweJbfL+V20cVeYMgRW9f9uYsTLA7mM3ps0+gK1Fh9lDQ7QajdPl+PTJh
D0l8I1taGg8YSdsC1V4HAGrrgCEydJIfTG8TBaDEj99x2+5IaZb6JQ61YdtGlN5XX/bnrZ4xrIvW
8sTzfx5IbYBf0dj9BISCBTa98WmD11ThmzlVkfNvFbyJhE8+LhK/kwXRnCUPRMKBOUs10cBsn6/Q
HzGfKXSioLL0K5dJGnDDg7ZfYquyshoIkIW+pBzVkMIMk5ovQpaQMsoZMQTKmGwQ9tllKCyZ4j9V
k2X6Yp80tSmmojmyYrLjbOwZcgDKADy8Ae6V55dxYVrHfha8Ls8+i7SQp8I4kNssbvWK1Q+TTQ3F
wSQIoVaxvpkIsl6ttp0nmCb7TvxKkJVI6Eedbo45ev1JJxTppnlY10vgUjFyHkUJ1LXdgSfDWv4P
FjAWrwJcdDG1JRE6FHW4JZ3QpP4THhEM6+OgT9U9keoxrormMEz7E/7UlXzqSVkgy/htxHhNSRrQ
AicFyb0AU5VDOLt/IXHKRtZ0c5K91CjLg4+t+yQmN14WLvMxhv31e3AFqB+Ue4F98EYXmjhKfkGh
l5VjIVNcsAkUd9tgp+xPh+TTcY/VpXOD4Ube8wdZZspKb92C7AoLS3uyUmeG9YJrAgkUSMtFYWiN
NoqtPoVd3UGhaejHGvj8/wFNFlJFRifTygryAkls6ARjH2Cpf1BvgmNxqBUGfxg1YDUMZYhmeHkg
lVPodH38UEi8IeX9UQq1qg3sI1Z4LtBTHIlMYnok3CqEvzd54XkNlUcASzdQiO4iKEKOOezUKDDi
90WEFhEXfLLWuY0WT/kQ1wWB3ul/PZGB9UwDsLSYlXij+t5r8GjBsWSGCCezS+wIECyVGPtUZW7i
B6dnGG1KAH2lGqQoJlhBXbul6WBgrDjyyPmzUISXQ2Plsf/kPCZdSSoy/nGOKicSCoInOXjql2Tl
o0W8B8rkt0WyunXHcCl3qrm4MSbQz7CpJbOeDxsdSApOKuAmC2xmAtb9PYYkbrrL36p6xqir3iMV
2mdL5QswqsJUH6BBG2GyLTcdQ7bkJL4eeymxuaBzLY+vg82uXN6g8RvGH6Nvza3RTvJwCzIIvcdj
e8/mwKzGDemwF5ds4QNOwKXVaayH+aRG63ToKhqFqzf78S/RLCk+FSaf9EXeXScAgU/ftGvF3J93
LeQlUNx+NjNIj87AoiATiTKOuVYQD6zpgz7AAE5gB0uBn3EnmK2NQDzzlRMv6Owq87U19oWSWzLw
jO5Nx+AHltLqRVn/5wUZpX1gKDhNjOxamzwMlQMLgn4iTEKh6YQ/Vb9don4MxgkaLGV7vJWqJKyp
SZVCzhvfWw4xvjcwv4S/tnj39YYqmHiP4JkpkSfjlnhelqs4rEsGKSrqtK1J3lE9ranL1DEBnjjc
qBhxS/LdCeIAVXdJpv/4smAJLfJPhy5NHdVDElFQ+hT5a58YmMxT23hMAUMaDc17JpfgXHY+dtKN
KiG2hxv8AfN6ubD6iR1cYfROhqnYpvrODgbH8TCdZOCiAm8CKGW+xVBO0n3We3y3fAmG41dx2H00
Qqxruv9oPncOKRkmEdlbpm+tlRyHn+eZgf4zkMMA33itHLfP5yYSl+FvvxhbAxC2AqUG51GpbM7z
hC51wr5xC3KFpJkK0BdyFp39fBjFSznDBogF8bu5x6y0JxRCI9yPG78J69DQoOPhtmt+hYhNlJ1V
ebf8FWoYto/U1De5TmQQub0a4rfXCYo1+fcSDZY7DvB/yHCuIFGnXUoDP22KRaGKym8kQhWE5dSK
iyMbquN1aX1laDAPaipC4YeyDnHDE/hJ00Vxv0i8D4g7WKiCpasKMhx8u9Z+/dROh4//Tzo7s5Dn
kP2kzmASZmoHRF5AghehvlOW1pfX4kbHdnEqJfjXzN1B7bbCIG2CjJpDpkN4d1SjG74PH0FW1UYM
nF5r5EpVpg7LOLRxJx6KLYsuSn9ismc70urtLLG4/S3qf4sQqj42hJBs0mjiPFE99t/AxDIYFz5A
1KaC7UCEcK2j3gPxQpEr1Oj0l4cBtka7KOIzO5NQvvN5MB2TH7fhFhVOnsF6S8SpHy3WJ8ndvanS
6pd0E8Qf/MxaB7BXGjeu4z63IdbFLEWNLdntyKCTwX2x/+XtqVlTX2a989euqveOVSBwH7456eIF
3hyThqFVYwCcmCpbaueNJwWiko9fodSG0H2Gecj90LJsgqxJlZKOvWQixYlTm8Dl0I9RQzQK9wKz
aTLrCWv28JOfXCyMqBSyUuTy5WhB4u3kAmrHxezp09JJFQ1FZIASS3rVVQPZqy71UfFFJTGWPso0
bmjlZX47NdO2CbqZv6ZWUSNZQHozyWPr0WazLkqWZ7nI+RGUkyqpthI4w/7w8J1qFSTmz/wn6Y7B
xyQEywKuprbSzuVm5AhdLwX6o0hKdbg3/wZYSQeaQc0QgNqNeN5lYJXRijQFF2hGk1SP78fc7ZUY
PRZTYMAcDmBtgoEjWo2OuOQmuys/z/cn+B3YRfUnZzJz1DexsAYAofJ84zdKjxbkFn1YgOeQUJmz
eVTIjCW4JO80gyLZFi3/fhwTVp1qOaHeC2u6j5lwM/TP5bCFsyG0xwfJmO0zmhoIXosYsPeBR5R1
9M8rVx8g1alCoxgJBKCI3cA7V0BJEnscDpMwca8dCyr1tHmH5OhNXQsMf55/4+Nf5Pil+5mgopf6
mET3EFqikQa+wQjnue5e1Cr0u3Ju0kZP48ofeg1qA83iztVfRlORkclqjex7tDcVL07mxL8maPMJ
ZAc2eTBuQZBp1fOQYw5s90k1YxApuw2d8ONxMMgyK2h3P0eo+8zYBuyvKr9za751/UX1n4LCcCIi
6DTPK9/F90RI1vGrT4nMh5P505i3pcqaousF5YzjNhURIZQ+xeJuhxSpckB++G1ya9+EZHZGzYBO
DbB+8v5OHmuMOpEp0+y5wQJiB3IDRytIf9g7G9/jJ7XWc9RlNADENyJAkUqmmXB+wkwmlw4wgKrf
bw9JZHXltbgFmnhpkvl1T0sXVqmBGcnheHwsA5DfxJCV5bjXwe1n7URfgHyIEwmjpRuVbYF0v/g0
18Y2lSl4TCwxO8AHSyW1+NximPKSLOsvOe89xvSdrhSokx1d25WCXi8Iti0FnqtQKRxpwmJxAX5Y
6laOVOny6d1HFkz4zrObG9rL2Ag+laWkRZISyE1CVasiQkOJiN6QtBIEdgdLMrWUFOwYPhBio2DO
Mwh483iIgpSKzpon2sMO2QKToW/aS3tYjZ7r1QApvAOapFxBeymoreqFtrvVn5GoOeaNHZ8k0mE3
cQQ7hfEoP9B97AvMwfsANKO0VSgS3IrATlrjcyGINmLFMcI8KXWZ/lkbLzzdKBslV4t8H1MFeSzb
eDDzKyJ8wjJ3q3nAHmz5Zrp9xy3mUOk6RlpgG+nHpV4wXv22UzuXh8LQ10QcC4/hItmkgZOK2Seb
xHCnMIMAYOm8l0KCnfa5xJPvnqa4VDw7+XNVrKquqqViNspu/6blcY0xDCdyHgL2rBp5x+jbQnQ0
nWXMfqc4nCRy2MHX40XvTO1T1DrnnvN5ORvOZqY04wSnVV5HR494NKUjzTJP8TwU71XvFrjzAaJ8
AyAvEpPrU5gILAccFXKYTEHeg2rPdChPeu2ZX+qJeIjOePfU9FyaRSO5Qw+vXQG6X5izIv7BCuC5
KY4GEWfAYpkTi3034CWVzR1OevTucGGq
`pragma protect end_protected
