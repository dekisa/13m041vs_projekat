// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:29 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gidse85poVsO71j4IElN4Q4po/ZJR7CF15L9s+ckKv/tY31TtJ7cTL7sebgFFqbo
MJrNtGBoOWExxROFtILPHZNHx5SDys6OUP9TunUiYu8J7EmG/72ThqgSaYBb3Fmk
q+kHbqRyO6bdlz4HSUQU2MAzd9FaG94ERJ4fLeqDnCU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 55408)
rAkgqL4xgmYEFV/CF1k9vMS0DlDu/woCJyQELTAKoDz56PGjPkoMnQ6uHvBwEMpk
BuZVgRkJ//FmnMr/Vjd+zgoZFXdm3qGf5oHt0OI9DqGko2SGJg6+erGOa46lmIpS
xQvTPyqAFoNcld48cZkv++0nDSOLEc8yUNt7YXPTTjFmwnLXCUgqXUQp+hzF9r9L
eDdCRxexhD8RJhpW6F+t2tKGPManFuMxIf2Aq9Y5BXHBUaqcShQDvpiW2+Z75D0p
stxguFqSHcQjNdQD/+ggU7OZ+pY5kjM0G7TIqqU3AL9mfcxbBBCF5auq2s+rXD9K
oOVOos/Xm4t4t1xjrIqUi5lD9dXr1LtKpZyc8clDGi8itAaSv6X8Uykj5a7xovyT
RhRJKfQFjXLuGhWyfqj59f00sIu5r14lMUuu9s0sc+esdzGkh7shidLqTh1T6z7p
33DRTh8P61xZ5oxX8iOtnNqWPfqRKIA8CCJAagDTonFHdBI+YASttt00QWjtpMTF
lyNX7QXKFGpL8hEg2lCL8BBtL6ImQqCsKrg1mEiOr6WVaPp5+tT39XaWQtAG0tBx
AB/lsiHEq8byYhkLULUHSKgB+ZkNgIaAbyXvmFxU1jNhwRgyv2RW+K1DuZs0+vNg
PrK1RQI3bYpbCEikw2nFX34DmcV4Kp+YTJkVuqS6I5ajX6UXQenoePkCg+QYxwLJ
CihD5DfkHZONWwERis1urUnPSPGEob3VZc7qZe2Bs/d1XOFrKum2VPKNm89Mw4PY
XY6bT25xnZIOtRS7ebQ1TLJwHf55LZXjjpYJ77JhLDRRLMm3LexVvrzg9JIqLW7P
QinzRAJ7uavrAFqhC6FDxfR7VK9yP+QT6lknp3pjeTUg/IntCSUnm/Qdmr7cuQB4
beTE6kXZLriMjG3aLZi8aFAzdSm7ilAs3eXjbSAl1ZxpKdiFGgsa2mqUzwuTzaFG
d4gDvBNb3EIG7dC10wJ3N4xS6T8YbXPR9PyQ82+sA7XSRbEKT69ACZwPPU3dFiJ2
AbXGVyd3eJjISjd19Lt3b5z0mqr1fyzl+j3XjZuq8UNaBI4BKAEBKF3Q0RzFWDBJ
zTOZWjk2z5z2OCqk1rb9+KGMekPwR/8RXAbLTPqN1ytOiYOIR8kXunIBH8NHYHDN
4XyQT/3RcMP7dj1K8SrH5DbQyRoYv/0puX5nUEHR5TyzCN18gB2rHE+0iw+R+JWW
+bFiprPebi2I3mn/yGQLx5G4j+qsOdrDSV0qx+x5CJEa5JRfhOhx+5VaCmrjDwxu
HsDDvVUYzFtnUJ9QZg6u0uFBVEmdHkSQU8/VF0+v9mRsIytrF9L/yMdmsRFpgpyo
MwzF8tbssTpoVw0tBJqXPx/JePiqoRp4x1AXZQOQXNEcEvmLMFrU1HCiYwLMGbgX
5iWCHMR7d/6OIbOcqvKiozjUNtg/PNMBeIfM2uy0QlCkt2iYamOpvwNEtpTbqxHl
8vKUtbiUJ1R7YnNDlTkqIs2WansrdmC07hFCgIA9KinFiZRtIJMh1bm1U8k7UrqJ
Qc45JUsju70J6W60AUXhjVIslFX3prREmjWdxMqxtBQ/evctJ8RK2PkTNCIikJJw
onTnmcERi+JJbiORCZRUw9T2H6ZpmmU/1LBVsv5r8tTVirA+lcdhJpE5wprKZbtq
H/eGRqtFXB8nNP/Ea9V0+7O2GAquNPfA+l2EqPZNR2a10udN8K/X6VO7odRSM2Fz
XKbST+xEQhessfN3aYZdr1Hs+JoqzdVtB1SLGXMYksFonsumjt/2LfRCVrSfed5p
p0STJN7j27vNIkhFISuW2X0C2V9vm8VaDguHjxc8clompnulHK2ooQU4RjFH6mkM
p3B9hXAB/f8RN55JGpXSM9CgVcq8P2GwVm22LRUlBaPlmhXdDTW1FZOugqVL7iBw
Zl396nrZ0vmj1jLZlPnaIAWglaQLb8AocKG7AaNB4K8TM3YjVf9X/UxQwz7iomjg
7Nyy7fY7jZ5pYOSY7qekN/Oby/LlxxW/Tuv6auEE5kJZA/78nnX8dI97Dw4igrZN
Yc6An6z9ghd4YC0GIdYejLi88IPmLKgQGvzIymqC2Gnd/tXjB+aMjd4Duml2nY/n
mjc2EhNV3SJLIspj0W8Sb9w6ycLfdSUQzmF/vywLi7kenkBHRyMbULQhpiapMzPj
amb3LjeHMW8DmHVswtR8XHeyzRI8G1VYZiMGrzCTE6heAMwNxP84bj0/Dgqk2JEo
X8gzFs6gShQwmsmIGA59FgEZKOEG11hz0TSRieFBahYHHjcSTeHtgEnM7qLc7sst
x69AyJaLXg7IYD80gRcm92hb+YWsLmQlbq7e3hAMBMxXmTDE/haZbXUKduHgPSun
Snpp2Szjq2AKl9Y3MSJNLGVxpIHabmgIyJ/tygkx1TkeKaF/VpqN7VCDQ2AU31D3
SaQn7HRf8C7X+wtI6wrIPerVSAqjsLPCPHVSUAwD22CSdgedY/igeLIz7nPGtw/v
tLw6LkURyUcG72jsnm0KJfQeu6H6JJaceMEsqyPFjLRv7eI0xixF9EhFSF40YdON
3ufb4J2o2hVFwrnZdJNiQRS1El4pP6VEApauWI1eI9E6gmJa+fxA+HHnSaG+zlF8
T/XCzHCNpKOeETFvhXGIIi3Jiss1G2Pz9UqTP69YrYu6p8q4fOQldJQZmgsZLL9L
n8A8VlYKK58Kyiw1l4Hx26kxhvGASK2tRJBRaEbLl+9orZyySc5OzSCXvQkkY68J
YUQ3sj9bALY7Wk4RAr8XhzRywAlvkgFTUSVkuRuDk4GGW1tdhq+b76U72Bhtwvh+
xSp59llUnNbtQoc3Mi7W2P9aofyTGuVpUvsNMlNMnK8XGUEP3jaK5e/PSbGcs1PR
OSVbd1ahzuufW+G0pAIcQ0ae3eDjm4PGaZVGgn74MWKfjqO6Gqkb/5sXpP2I3QX0
+VYPtSVbn6tdsICoDFzWzvf8bED+sKeeUA/nMx23vCAAQrZm/7Uni/aoWURrfRja
h9/syl/wO/QywaG09naiFvxqIgs5sgZ/p8/7sORmQ6c053OJ/2t+CtCr8uWeNxQt
oeuLKj1y0NEBRi6zPtZWKCtri3teH1Deg/XrS00jLVWHShhLWk/AMeR8dFjBmu9R
nE/sFpeJWHbJQa6iw9tgxnAoKPaMHylWIba7QS/K9ih0EXHQdxlrwxGj7CwZo9ow
u1dt+Pe+tnqBc2L9g75yc6RuQ+XqcKnlHVyfKJ2VAn+wiUqwmtYuz4bmgBuph3d8
qbGaFDZ00/VwF2KnINTCjEgq87HMVwfW+Cu9nHQ1Tbg1vk0Hx/mvvVOdKcgXxmqz
wfF8NRZ1rLfgiYCQrYf53/YOImZw9oC36cPX/4WEWbs5mg5qwDXoxSGpEq2BA0Ic
WKzQtNASDYUth61HpEV/2g31zGQ3F+29zXsBo8hmFR7a/QqaYh/kQve9pItO7bKD
VucdfOLkorzLTCjVV19zDo3IBniwdYEN4FFLZRbPePwnw/jHuY83lojF63DmDbfe
9Oe29htZdy5hWb2eZBMIimT5fyUGnnFJxH25HzJJ7aLIVSdJYUC/b/tp3Q6WhmHx
wbH+g1Wi6W8dG8mQlw/bA770/b5zNGOH2VPpQbWNGLoP5lPkFR2yNW9DRlfClcWd
vt7OLg/aJONWGf0lS3/Q2C9BjoNgxy20g0INkhv0e795KuM+A7lm1YzURhszosxO
UE4SNYOGnJJ+IGOAi9ZKFNex76RPcIW3Vc6Q0XA+XqnOwPz1uh6Pvr9DCL3nlraW
H56efgUELrwhDBb2mbkS7QuTvnNoRFvJ2V2d19pF4bU/p0dV7jpUoaHTqn/8Hxo1
5flWrTM+f4w2L9Ny/NX3BUY8OBYwV4gsUL61Od/6qFdl6ePv8JGOoM1bd+Zp6pUO
X32WNt2xjTqcX8ugtI3e+GH6F8yzRaxV7UzIMkg3UFNCR6NswUJQekIKMFjHixWJ
NrjAE9IyN/IXDrUeYNWz6yGpWDDX/a6bZLg9D4jEOhFFL9wVC0A3gOCiZGSojY4Q
zeR+Wc54OswS6Wgh4RE7YvWGAUd4YZ8AZKNJjXIJeIvOgng1/NXQ4yquvUANQPMF
RroPNzcKDU1kBpvA1tAG6VX0PS9OysP/icBAUwymiG9mCln/zOsH1/YNFIJChUiN
00rkXNFKB5AHIc2Q7snLbgn5GF4kIdNJ+8PK83Y07e/0vk1rqh1LMc/FsKu9IMrE
9Rb1BhAAyKHsX6UI0BXSQA55VaOq1gEiAxlbqIOP0RqMHWzWVGc4ZfhWqU/3bQbz
DazIH9AWWeiDFmwyylCFjZQEYJgCo+EMMv6THUtnF28XgRL7DHfvFXCybZcudytf
LTJxHi8JUAnQrAQQ8+sVHFu4X7v3zAnXZdgwzMZ1jwf5vlLwsQjnLpuQ09UuQRQN
9j2gfvoLQV6AVAl1nKJC8rlC2DZhHXxBs0BJAOI7bWhbT+b0ujy7Ey6iTBWqC77O
rOpzrMOqgD+B+1hxPBdu5hFzGCG62PNJnoM6Nz9mI+rye0Iua9aCCwfrUjL6Bhju
UkP3iwjbvUL03hLu4koSTlV/i4CIA6569VUew8yZFo/nj6f6+7WT/DNN2vJSPJQ8
7f2RtZwd8L7WhnYsERv5gj+XjLoj5ygvtTsnPd58Y1VIMI7nV/hxVHFOAbuwNYPw
WyVWdCMhbRuKQeclBShx9+rGxS8wz4r+0Q+e7kRgh5EvOilBzBpx/tPi4fgc3iiZ
6f1KdF1ZdiTalHdOGacFwdmz/0l93K/xrbiNJlpr1JoxGpEtippQOt7tzb189OIT
WrKOQr9YMZNjKF9CTnywNDvB0aSAeNgrQiaEG9I8spcuFTrvF7BUAmO/GBHIS27d
ALVG8auG5j0yRgmQlYF5DMOwzOTO4NZ+5ybOplsGWZwnzhIHu93WNk6As6Pp8xAw
P1F9pcfvu0P0ETb7RJNHX/h+9wTt6VATRBwvMtOPl8cikTcncGJ02+b2uF774kBa
jJGw42X7BSMnyZ3WsWKyfAPZEYO/2+Lj0GHSet7umkLxbMSeS6VsCYzCLicCktaY
CUV2hqZ38K05ynptkNvYROO9aTWHHmJ1kIQXhYYmYiC8tcjA8jj5wiQ0Um9xlC04
Jfr/J3YlYGnQsEbIdv16HpxBlGe9WxAZQkLiL7kFDvqZiSlteTw2vxx/TOaof95/
KYIlf0xhsnJAIE3giZZCTm2ilKDAfNbF8620EnKFDsLQKWkVWvgUDUm3N/An1FkT
fUI9B3qRL5EzF3SbkAPnxpPwHg7bsy0vuTa7ZvWZfUxUsS4y7O9E3m7KTIkLS7qO
mPX//9yVnA5z1JL7/qlcnV/XxewIAR9KT3nL2be24iCsCESngeI64FdRw38iUimR
9EBKCP/ihw/3WDl2ezsY26uUVjM7cIyt1fjwnBoZ4I91xmZl13W2RNKJz7KDCKjI
xlQXTeGaiCR2tB5VYBfkn6xT1xxPyUMVieXsp4HJvf6j0yaBs350kJHhbokEDguc
XtoZHi+Tb92a+12YSirQwg6l6Uwr1/8z3YWh29jcx55ihKZRtrKK5IAYc+U609PG
o64jL4hRqWzVkGEftWQewmSYxSirjEui/dfER1Y94EvfId7HYSO6RDVDne9cgX7M
gh6hgRgNd8cYdBHHPXNphjzmj8GILDyFYD4nhoqK1FOAa8nre+ikYjXHIEa9bAiY
3Wvu4E5/Mql+cbheXvDZCEXMNJzG67vJm3lEKSEA5sJ6dQyOVMjDLgFBeMt5cpKl
bSrvlYfjrCTBKvpH7O9S0OdRz3/EhoRrq1rmxB5Hp7KBKSARUHrteJ5sNTYVgMz8
fa7SiPn2cGBSFcQk08HgGJM2njB/vBd9cyaKjJ663bF8STPf7j6u4n8NJ9k3k6Um
aYnkpG8np445izasAXpuszMulhQn+tsn2xC+0zB585n7s1GDAxoMMwIoBL8v1RKl
zsKGV3H3nr7VuPRjbtVU7GhaDGSMM/0jZE1oHxi+jZeZMMoL8D6w8AJGvpv4ZpAw
ZC4f/2Uy79+e9xl3aDmQlkd6yH7S/pJjvv43eS/PwsHhldL6OoncQOIE3ZdeQcqJ
ys2evaZoclX8Emy75rMfnQ9XIHoS48Ks3Jr5wHSquHn/xQ9n+ofO51hnjVp8U+BO
CmlnXDSuBjaYUAoqbahsoq2poig6OPid7o6tKO2vBgJWGXnroXRjOtOc5OoDcnee
SBC31UdLS6S4UUWTvWcbVrw1jmIfb7u7ma7FSPo7Qw0r9xUliMr/TQtVkmuZ1HS7
6lK6pNGQLsYsYtEojHeNsvMVMKXcpukgP4eZaQR1RNsit1VZzzSitP6qQPHdVGZI
MQFT6rvtTcvnF9NWcWdGe9P9+PTUDpkXJmdTcfY2QnaM7ylKHV5M/u4bvRD6lpaF
pPAzMzh4/fC9vOjdtpBiB6dR9pBGKbMsroIa/YmRVJg2n3cDyAKJpwE1WSguPrvG
vKH7nX6Gn5XGdI+wp3RN+KC2OcRxNChI8EzWHGY30ogeEVqgui75b/aGaiAZBqMn
Ggq0RRn9rc9aYQNgfY+u//RL2IlgG+/PVbNPcfXUH8ZyuXC8fBGSXd4nCIF4otFo
ZlKtXo13ngLAf4UYgZx97160hxhQmJU8gIVsnt3dQns5WFxTDJO3RO5cuXctl6oh
26+Ps50rc0QH+VeTR8Cm7JG0/8qMAsUnRtnw6jnRRB4PyCz0BV9Atc2qm0EityKP
rEOLx7zlwoVTetcvxvK14xpNRH3+3kJD4viNtuoBv1dd+zaiEMsQAONRsv57GMWw
z2l4Nd9so0lLlohQ4jjjRFOF/L2oWZ+xq2W/WeF6QtAG7h6PJZCSi6c62yCeCnHd
RmxC68jKHq9/3dkQ4B+5mCr4Khi4KoeW0xX+MXJaVS4ry2luOvKVzogo1jLCcE3H
xLKHRLkgyqwaEeSVWeqQqXx5dW/i46h+NGZBe5K/ke9mmfZ16IbOBWqxL+o3jYWL
4qSfgL8Ll0fWuf+2+wfH96Nad/8Z8h1tamadAjMlBr0GgGaYG56gaWLMepgoj33n
UjuwJ1JVrVeA3XY7Hl1U7Vx5GyXDx/skXQ2XkzftDL0Jf4UNjLQIcAP8sLTuvfx3
1eJcIkNtC1nWifXxKE4ozL11xFPvBjTXC0vNS4qw8KJ4tb8K/cRnzE+LOsdHarDx
j4j6GC5E9vsr0u6Oaj0fbeDiDvjc0achWLZITI65wLAAxcVifc82KERF1+fP+/A1
h21OEl00Jzg7iosNpCeZicFWDvaiqZWWfxMBIX9sCZoWKmCVQ659Yp8d3CqTaP73
HknH2oen3qS/kQfMa59pCeIJKhR7ZQN4WKACjaYse1W0dza/CrPTroHps3WBhgGf
BwHO2M2lNUG+q1WslAME+rWziL0dpasnEYcyZ1zXNvCUewTre4V0gBbjVhDIHqRj
mt5JvRYls2vqKn8Ds6Vi+OktjwUxkqStUfhYGSSyd0wJRq8jyIVd9EHbbQzvnzug
dnUEaCIh2I3cNQYt5bx4ZsYaCWxL5uF0Bf+sNhZrwxKFgOc9V1rKHWODpDFt1TNY
75eTi2RJFGa16VAqO6WISgR8I7nEHSD1+s+jTjiQhA8VPPRtIarswjY8UlvGHZIY
E5XBOnW53RC98ufGurHf3xtGCqGkz02EP6pWVJLxtktc5tbMavdAc9WDsR6uV2Gq
j8+2t3XH0s7NqfYAqkK3hbphpDJsmpyhO7rargMVcc+D7We6lD8JwOmEcGNTaA0v
BjeU3D/wtlcQy8D0zUnVW1R5DyF9k0IOH4aYwg2VIm0sl+cPTimzKCRDu6ahdJz2
TXm2IN9D0UvTRY/FIdlz9Yi45xN+rL1OD7mt936Yf1aBJM/0NnY21CFGu82JUtsN
ramQhRNsI6iEXRy8c1iegFhlSp53X9vXidM1WTzKMKaOKFdPEPRjzGTTA02GhsdY
n6ILYNpxl7KV57qXUuKyAkVzMaN6FnblZqqvLRH4vOSmYm/EzjT9PedcbG2nHHZN
NYx+JYcE+vRzP9g7GNdkA6dwA/27pSSUiyH8J8Im4ujiKI8pGOa4YvjDb9Tis+IH
ZKzvR3YTWI29CymD9ei9Frazf7hPJKSkZt99ks3BY0FDMF4XQwZgZS1Puu2js9+g
kMjIQaZXjM7WuEo/8pQPjWnRb5thMNHuOdfrLLUTsS15n50VrCvY3ilMgsjYoAQe
vtMl3G1HnJMITqRiG7ZtWtL1gz5w9VXtEfDVjfzz0iMx315UTZDthiq0vHDxcIBC
du1Z0QrgBmjrASgZVV+I7Sfcx/be8Lp/ZU5lMg7K3e73zJHoq5aecDDlqpMuu7fH
gTF/ERThh3fVnE5aeV4RTlUQc5rdh21ds/FmEv1jWpktOHTFAw0p6u8+Z62JAs+F
ZL6A/QRM1Nc0CR+6LDZktP8bI6ziy2wVSs/6lkq0pC63oS7pImh5Jgy0aSUkptyS
0qCitaGlHc/zZ3mAfrbhDNm+KkNNBVtEqKPcstNpeg7bS/X/cd6KfHJtGxQaJBc7
O1QsG3anIm0QuZwf7HTbTGnzTgYFCIcJPf98SwdQgzS9vUi+bN0WB6Tq2pjwB5ca
3/9smmJBh+EZb2tXSnGWZQiZ1N7QnN8V7z0rdl4sPMUbfyDWZe962OmhKVdPeElL
VsaekGLMx+Su1QD7v+IXCkA9mOaJ/3fEXs+pn35r3n4WlVPMTDbyrrTAnanR/KEO
ZBDW9WXlXwEBiNT2cAXixnuW0KFJ9wD/06+NTFweGoa3Jg75fHqveR3MXH4yhy+D
nxU7IXDpu6+V/U9yhafEEH0Iok0NHgK+hX0+/L2wOCw9nAb5siW1i9OLlSV/DoTK
zp1b29QTPal05VB6tPIULf/FGaw4LtqY2QzOeGHv0XX9xv2u8mtBBgQosjHyYjxA
sMoacLO9/+g7sOF04Bpx6Uzp9oEnz90TgpLk2IMbPHPE7tBtRQv2QkM+9txqXTjE
llwp32Z8mlIoMPbuz3UGE72IylHeErXAnLHm2XE7AdtAZMIptbsJLVoSQ2gftlc2
BrT2TBV+uVjnT1WqgVStEzK0IOd10v8SNRs9A63PKKDtkXk9uvTJVjNqIc6LraSU
42GiNZiE2i+QmJRhM8Wj2z+V9Iz4gdaANZ+XgEsXio5Uz/wpmM4rMIlyTMyMcvM/
0vsnnJ8tlesvcUNq9EyWl6ETsK50vomXgfQm6FRuAjwILTIbIHj3+xXUHTfmhqBU
iz4aQdR6TqY9sj1xzr5dA5BrW+SEilygS5i/BzX6JILYOTzFLkoDL40M4+B2nKAi
tdK466w/pYanb/pzjBlBz5IIO1BXz81WvaIXrAzN9ZLlyVEPpSJyGR/lr5Wb6bDK
CmASv4KsncW9kfhEnllp8tRmlexSper+fb58bKxBQSr55nzdoya19BMPZPSZeHvB
Tscv0n+MbFztVMqtSHKCrsZZLhMHl7zgRMW1DmEGQ7B3Rw+XlIvNugUV/2bXvoAm
ODwUjGrlPyUlZwP5l+NliBAogukyhm05U602ZtUV/ZVY6Ndq0gzbLR+6sQBlY/iO
ClZaX5cecZOO8vKA7fzmlVMkzd3uG4hdzWg4RFotnDVGZwuaXk8A3jmGWlsKlJGa
P+cfsTBrp4fuxEVy1CK5pqopMzxAH1epZCjjh7ujdUtxykheW3PSX1yxlysQiQGp
GBY5Oo4iH30t1+he3SOBYiAKjvj8HZR9cy6s+VvInOEOdN12Nee7Wb25aSTaDhcf
/13vtmSGtqDtwSB6GMVKCrrP3iyQhJfecW6dwa5CsAzv6gCqUnD8GcQn8ActykRa
nEzys5xE8lM/bx+dmfPwFJ7acP5JKAzTA4XYouwl/W4TKbSjHOWl091GAsA02u8I
YmB7RQfIrV570Nrpym0b9FgVFkJeHSxoL0tsj50ZNl97pBuTv5hsgTvBQ+jKQjNJ
3ZjJbDjbzRidOxaQIYpepKTUayEBmjWvjgJz3Vh4RhJqahUarJDKo1fIH2qtA4GL
m0Yc2pKxLwNBXXXGNry9RLy/gJdJBfacWNvBnufxhTh7uaDhgcgG6Ue6qUNWnBiV
jBk+GEvQxpQeg3GySzsZTm0AXcxcqw2UuwR0pFdzH7iWNv6I3fyhqGVc4rlDs0Ij
cXYuVTL5EOkIj7yTD+zeagWZ9cxvpbeB+ai1d8/SiIi+266Te8oQKaXXdgOSsAqD
2qQy+Q9FfbJAcEoon6T9Fhhg3QrNoAH/kUFPOjQYHVDtHyGMHQ1oxMBtrJn5TUtL
Kc+dxHhsd5cJDNbkaUUAodfTFwYMYTRU35dtj+6ryKWPYMwOB0KvnPkB5+1p2rSk
3g9/KNg3dUx6CFwbyPmlPyaalt6xRaz9OJXZ+JR5Fz+P7Rxai1pLAJSpyLmOzmK0
N0ScRp88kzKl1XKjQJaRl6LB8ASt9IN5/RlaMsCkqltJ2jfy8jqChkT746RYWonA
Yn2lhwIYf4HVHIwSr2rBEHeLLEj11jPDCWfhT4HgdVFvo8xBDi0KcHhteZW1q6TJ
InHzweK/bfaPj+/BzCHlV3PezKpBdqd8w8UASNH9bZDvJ/lh6AnMasadi6pMra8g
lSxXOzKA0i9y8Zohp4D5H0O8mfn8aBDOALxq0iWzp56aKyjk3HBowS/bPJe4T/jT
+91pI+zCE4SgTDrcCnLt+0dxtud1Bmcee9VOv2puyO7racEQeuUp9dx3cb8BZmcS
BB+Te9jNG2Bt5EvYxA612S+AyFkvIESFdFA2m6yglraQd/qfVI+xQiSuVCW5x9VX
h7+YlzglAdWQtVndku5FNNgc/ueuHPQqZgOlziSe/VpTm+lhxdNyPwvPOa5yXK4B
XuwKkUAd7wDgm4UpiUj/teUJKwR7RxpqP9yWsUCF3B4ahI7W0dX3+AxESuQ2H/Mf
avvKW4YHIgMdzTidU7LbYfKgp1aHZoZ45aWgD056bLE+/fiMdv+UOxWWKVId8FDg
3Xh9dNn8GqRnUs8ul6t32DAOx/9QptON26sp1LtiEKIf2GzhFUKCxLrz1VIVdHuH
dv5GABh6TpOgP2jFx//e9qHBHiCw32eb9hVp4zwFegv2SMQ2q2KVyH2yOlHZaPJW
H6XM79Z4PPj7f/m+SGVf92Gxb76LN52JF463qltvEHEw4C8xJBnAZbbYSZYK43ja
WvsM+NXEd8TgmXs9/jaMt9ICL5NrHdZY3D3RQ/toBgaOXtuRIfB1nKQ5djQUvYji
9bJBX5LXiQfYtdDnjmdK7MMt+nnnxaOUcslhjNjPPh7eWPJvQ0x+gEdAcknC2gAh
AbXRxckNVieKDUKOUcFU+YIMgp+GFmqgDw1sErLrtInDNKGGAJIFekHO3bLI0bMi
BGepgxDExdvPK2unsPjzrgd3aVvNkS9/3pG/bXXPGB6eb+Cw3XeVnDiKm+7WO0Qb
FSm9AADHFoVL2Gp6pllUlePsYd0vmxXhU7BtV44E/q4VqIzjcvGxDW/RfnwdUPpS
Q/sxcpbQR5335L2SJZ35D65uVU3RCQ7hoUDbb6epOMz0bYwVYkTR2r4WG3D6YF7W
FuCEpBOMb85J20XsVvXsiMEfRBKPN4JRAS2U7h+YNeM99Q1HP+kTfHj3IXu47e+r
9GJl7LyIpJROj4c8WFhqr2fIlk+KNhnVXDHTnduJQYZY2Zt7MiXWYwZe7k+khhQE
0rTCMHb5yczdU5fn19YmH7C15MkQ9jD1NNJWjVAgmq5efwvLrfFhXxjCJDUFoeEU
hGaQZeTyezvPV3krt71KjBfsM/cX/AsxmDEflKQEjEkks1miQqX7gtWPZQ5+6YuV
MkBN3TsBDO4EBLrVHkooTR6bFovlm/VKotanIJkjsDknXCuYO86Cl+CZhM5iVyDi
dh5WUGI/6GmE2+5jZb1hE6GtzqThzjzoJobsdHr6CuNLFI24o0nb2SS0dLrRv+9f
kpoEb4fB4ExRSXTot0XPJBtcFXDGixmOqKSqSCZQTwUovxutXQqdf8RwxHPGrEUm
BbIAGr/Vi8Ju9XdO4uG6gb4EqTc9M7wrD99IZDqUW6Dkl0xLpJpiXQoGFzHQh/cG
VeoVk2GrDMjsE2FoKWGBWFIY170t7NZ2TnMxEUfb7F/DTzO0v8FML4uVPW976aH2
KuxArcTesw/CkWkIJ3nf2Xn3YuoZt3XF1aogX08t7hWW8YEQEY64DDvCUf+orwxQ
UuYQ4GmwvpQOvJKvVUi/VNiYS4gif2htto8vOBFNlUVb+0nsIgdZuD6yxb18wEFP
sC2F0kG++VElwGFktJadss+PW6YzBcEKUOr+ksFMLzT/10I78fWGj/2JLKUeIIhz
v00dphuQ6NOyBOPca2cObEBILggYIc1EYToINDq4p+jtHEzGoB4vWKv6d++8Nepn
rw6p1WaRkoJytkjH+1sujYG+RItayG8OcZ6wEqey2M+JoKp6TsuJHeXXUDecGaf3
278RFU1vA3IXvCEz770AWus5Br7NCVs9qDtCuPjNxCw5L0Zk5qM3b9PHGVxL9ZOb
qqYaReSiEWi3mBMAGyM1hdNT3SkUainXWQCOIKyrGYGDrj1wnMfsc93hDqRs7vea
WqVeGqr2sTDfFSMkQC15oNE0TPo9FQIc/Uh/8V052460L2R2SwVZ43HoaE1d6asA
EQw+n44umpyML6h2SiCUF9h4MmMuSKCjfE1A0P9JoTPni3Ck5sIUi/R9tRnmZC8o
JdxHWVaF4J4KWqtOgGoqF3MUkSSSWHfMhT9Lkbw7yg3lAJRwQQUmkYwxMfxk63uq
LsH8ai1BvSvRmv3/DAqbU7BERiQfzHTNfobXEDCa4nkHEBdCNufrqQNHTd1WTOba
3ePDYu6Xof1od8tih8r2pBcgHJKqbgS0zJPapwb+OfnXy+zvqeoxV3s3kpejNzHt
taAEbjrcYsQ4CuGwgQK16U28a1cKHz8dJ6IImAiUPCCSDJD0StBqEbEXtUEo0qBO
hdCV6Z1s8chlPCe14DSZne8viB1JVvF4Ewotr6KcRc3r1bqmerPtX0kEijODQSeu
3jpbQjo74VUqYbDboAQ6zmPIg2TTjBkjexz08OkvvkMQuVvCuzvofk7kJ4MrsWhR
gtUV+RV+MDIv0cc4dKqF0mzqU3ByJk2qTxRWEBi6i4GF1w+0QelrKsSyH7zbXGDV
pDZv6PNA6xjOxeWwv2daZb+7G4CCKP90+h3MKaDpbAHYRiC7b7BdaTtUgh7NgoxR
62MnzOll9PT/O5tmf7HEyvAH6EXPxoevkdFcqr3vncPkBncx2xOjJ8VlPPewG0Ib
XszYPDsUSzLVcywwL7ZJr1EuyPQ1pfKSMIIcQVHujZQqSMjDM08/iVw9QaJyQvZs
ny788C1RP+ioH1eqqXD94Hch3Xmd9OD4MpSmAvedeMkmpuozWaLcXVkcKpN7Phvw
d9fBtvmTha5T6SbEEIN7ZKh3FR6z3i5L+i9pd6eN0ladfIwid7VH+pNFPO/6uJit
jaFHU2WAotxG4iXBdMzA2UTF4sTZi27jxSXLwMH4dobcXHVxrkPPu09Q/UAUbQEK
Esit/Rqg18eVQ25WuPZsTnToTH/DHLb/x2RW2RakStSm0h4yPutTeQ8ZjOj6FFx5
SOuRMtylla3q4iikh4MVhrukJTrxw/vVOQx/GgXxD3EpW5JdOpcXuv5pRi86BUiO
mAIjI1ADOPw1YPpS2phmaaHTMjt1L7JBWlaDVMK63KkvA+EzmXo7rhKQJODRihIk
3MAESewnl/Z8syM2+kBRczAqGJEobsByBw7sE/TO63/JEmAQLJ81Jn90mU8bYj/+
naWH8qItlH6uoEG4qUDqA7Br515Bt/Ytw/4ajoacXAYwIOgFhKPkuSs25V6q1qJX
mA1zmOaOeHIJ2Gph1rx8cYUs/1xMmbjMoDFW3EzPQA07/jRLBit3WdfzEMCD1MTl
ugpTaEd7CTCMtYjGOS1OWHPxCtsmj0ExCzAGgPwAFIZJ9bQvxL+v9N+AVl1415Tq
5DUpx2bOAjCEYN56hk8WvkZsBnQe3LXgWEM/1kEOFJUFEuIfM4cPo1HIyWS7KC+p
JRkMBA8pMbQxoyRRSRFPo4SIbTRB4R2+0aAKRX3FhbTCHX8Z/bq9+DHSnjG46U+1
P1nlm0hd8/f45WaC1DRmwps9XEguaAoAW3K2EUf1THCzgpe8eY3IZXW/tdxjc6Zh
HCfUrF1FyY4iFFd5sWBuyJmHxDRcCkuo96XaxLrYnqr4K5G1zxiAwOXw57zBKEVa
VzYMySoV/rg8h4YrzNqNqchPkrAy/Zu4RtKQb3KssFO2U2F+I5nlXj91T/5/8kKn
zM5ykP6wzl96JOee9pGcctQsDEblIG5mcYHmoPoK8EJFt2UTv+ATwnApqpeF/bss
XzwqXTVTOkWlwL01NXqyKSi8qNQkFWdiomAGlWHJJpRhy1neTKg8LLYBRJ5/NmPR
IX7NfWGShox0x5EX324iz9C3buncECY0D5tc4I2JhVm6/IbuhnwWsD2dITR/UEEh
jDcxOqvPY93czOWC4Z0o48tPdeD+NIK3iTPvJg+8DhySYZMTFRkJK5kzk7xMPb0L
83UyltHP1N6zagE5RqfdS7CEV7+ieeQzc3R68j6LFJ3k8+0h8C4Ok6UTvioA5nJV
hz9A4NmKmfMkikegUiE3vC7BQfetVcDwNSwNcWwA0BXzbDUDDxnToacbcnDA9vyj
9x7aRBuVIOBWsLdVi5C9Vbq+oF1iVi+r5vxwF5nSncq8XiUoHBHRlpJLYCGxCV+w
OY5S+WB7fBFBCie35CPDpkyM85dSZwPsk5+sDZQztYMecw+qi3P2JOlcPr4aWVt6
iw9fP0DGOoDeeh+epW0rKT0V+B5pt+Yp15MPnMqQDp4H2woGV+Dcfjx3mQmCakeR
rS3zntpD8XyUnNVbJ9JlvhBEJD0Il/63VBQ9LpQsS3jl2fP1VL7F3rFDTW/2/65c
SB8VIlWPb86ieP3aKMDT4/B4/J3Qca/kNWrIMwD6VIZjhhVJDNkW5a0SH94u/yjt
tyayfC9gA2NqtOqRBFo8RgJPW2buS+5XI5adDyOsEHAA8/dtdzUSYqcGxVAHXFNC
0pEJ2To+G2xZsiS+zgWErTEavphTNFYaQWuUom1ObdrLIBaYedjZ4CLazRWWhK10
15sZxfBkT+qq/KaXqRxZmeSI0I3QqY6da2/TSNiQ7BdN4cy3/TZfF6VHt8917TjE
f3BXHAwFRUYHYUks0rhx8C8CiL+JaZ9JnUU2PY/006cI58c+Q4ZpIYaLfv9POv3u
/QwP1+EyBEst4WIkzBxKt4LmO2zAgEvPFoeeoqU5ivrOvay9LTZxUOX0fljXqDl7
I3gu4K//XMnjXtGTqlWz8CckICe9AWHI0h5USME6PdSJY9h3B+yrKTMXqRkVCztz
3+rC5VBphcvG4siI5lzoWidAA9KFCQF1F1x4zbVa+Gmh9V/xh1j7v7MzF4D7vJ5P
meiGDmhozu160w/H07FkWlspjV0xrUhrea6yjzNzZT6MfAs/8j/oFWyBOUOsQlwn
HhTS0gedG1QXQHgMPUjfCZOSj+x22V+1QHuLQdeOvscvVEX4aosN4DveX+g7xZIh
TNlV8g4PK0qZLtV9tsFR86D7q1O0xcvsMM9gvudVWiqqap+kvgVwvwptWTHS/ziJ
8QcEwXswNvql47SfObsCpAnVc3sgKfCNFVeRDrmKrZXuy/L1q4YHVA5f7wv2/YDn
QBajg14hFINSCQ6UYhiMnZYIqeeOjO/n7oI6Xoyt10d0TxxVywlunLcQ/m2X1Img
KSSFVg7XXhcQgHQPpzlup0MHsCJBJEVG+0x6cUaggZKAL5bWKBN+PvjNoaQmZkGw
AVVWIbVuY0I35FZMIJ3XxELe3jjHEx1D4iGq1dr+DfPkLc5hdVJu8/p6wCsBuViG
AkFCtHAbaKiDCfrhg2FGYI3N7zfJoei7mmeS6LTz8Y5LuvjDwVjxUkSC7rGdZfi5
GXxD8WChOVAc1P3oUBTDDZzGrwWhLMU1idyBiMp7dOWqVvempzyjtPdmaZvofUNU
JZEwvLmwFoL/zsd5v8vfEZsueFCXYRFaEJB54517IaCrdN30xwbKQ0idBuMX0rTr
jANiq2T1xz5HQP8Mu+CSlN3jJP7Jevcyou+VlUvICMlPyj6wS4PBnZgtKHRwnCS8
q5/SZWmjji+CXWeIprNRG208Jg08x6q8l2WonWRZt09LMqlybz6jCWuIFiGemhIb
4OtO9CrEORVAeiOkBeirDjf9L+LGJvTSvgkFjfAvCw4n0pp2LBK0CBe9NM2/FmiA
7IhpdN9h3gnL5yIDDHgqWGh3GtwlZcS6xsBom2B/TbPFmZB0cpcOR0CJo657hf7W
uj3QHkzAaDP2NCJ0JHNmmFix5mETCoxtgNGX3cJNQzxI79ZNaOzJQ0Hcj83gLgMZ
H0GbcuEvQ8pcthfoif7V6qOS561NcTQ82qMUcC3MOPlsyjUd0OgywXZnCd2Wy8MA
QUtzeCq8T/YiZRi8ToLnicRNR10ccm4OJ1PhAKybbJJQqWI7D7KcaJarMz3Tfpxy
EwucwMiQIOm8uvEMu0fNX54BKnFaqkfOBrla4CuwRVTCoCkWzw/HPHets/wIjEhu
1mX9ONobnlidOzfl205kF1ywAxfIPTxFfUl1khr4QmGpgVO/kaVXHAaMj35GQBdC
xC2lA84YEvRfqy0+t8d3Rb0GAGfiPJt1jXXf+zS+wiL+rYgeFfL0ER8cW6fMw2u8
HzAX3HIJbfOUVSmqtCFlbkiU93zXNRmNVZvIBtia81TM+8lDOwzwMlgj+/c8xM0i
oj7mtI5EpXUCNwZd8fCH7ezubKKl1ZxXMU2NQDoO3t2Hpx0mLJtqv8esA6UnyvMo
qKKpl4Ncl3nANdvuGDeVo9/7WbXAoDpSzAB8paqKiQd83u4qH/lE4dFQNkCPSDe3
JkaXBpZ52ICFKQmLKGoQmfL0TmOpDOWt1ROnkzDqdLy6zWXIAdlNFmiiJ0gl/4AZ
N4StafOcPMOjXla3PjW30EEkNoSwR6PoA560H81XQWMgppgHLVMEKcHoyCMukJ8h
bfYFerP2akaQ7Mkl0gkSQFV/C70mFDEyo5tg4zfoC9UwMvxAr2U0lwmYOGBlxC73
ph9xVN7BcX9yUr/Ay3/Fhz03suoxXqgXrb3A8hHn71fxspG0WQVcr6t3xniVOV5h
j9mE3N9KWU7bknf/yJW/RigG609J9PPdapRfWZzJhoddJAeawxoJaYHLiemayEgh
V1IHYGC5rmPNrVVOoYVyg4vRk4wnS8b+qPsSuWaunATNyK2Cxro7kRk0K2n6aeSX
Io8i4GxJ6yW+eaNvmJ27kxFBveH/oxK5LXJUGpENKsTa47VyE4hpGUrXAIjr40Yc
dZB+NGPOdbkHRO0V0s1fz7atinfIeP+27Pa+aW/VIImnpYFhta/MkrczuPsCN+RB
WGp9p7AelRvvzjzYggKt/mxS4kT7fSPfxUGrRRr5phdzYh/iqzueaRwmylmNwbjm
LK6MDR9CJV+IHJxCb20UQgl825HUDPA4tZg4LZqh3JljNxCsB73w7K0/wC4jqUrz
uO6IWU4f3hboduDe+w4zw23GFpVg6lzWVUrk/oRIrmvJAkg8leKTdZNVTfMqhyuL
BWHyJaGDlLQnZTUlXiSnr31TVznGQ7Ta00fM2vXjNeURiqUVlTyif8wXdJDW3K+V
1CSUOxRV0BIKXCGFZ9c815/TdUF58XTlSET/3gGaDHqjOlpyrp504te82yCdOwHl
p50A+ExyLkeWcsOpJvuOPaji/A8w6+C0ZBTB2j+52DLrYIa8rWTnJ20Ll+aX9nqU
NRt2hr9u+yo9BEASfRh/hOqow33HcPhqHMcxxeSpdOTWspYqTyH3SvztazJ/0Kc2
GKWn9DF99AhWBmDobOx9+BYnt8TKz3QZiUBb/wtOVOMV0gvqSbANadaOlq8VuqNy
uBu2hMxK7OrvInURgF7blsNJJ3IDOg+g0u+aFfW00+nCaaNHB8TwU5vH1MVBgux0
MQEHQwgYX6mGk79EurkAHt1PsjY5G00Enrum0T0A9hH+/1q2Ay2mfWveAB+A1Tm2
GHyZDjyCh+cKh1VxiweocE47X/Wmeo70DLcAFn+fVzGt2fthdFhzpEEjjuCCTV5q
xVWtcqqNYEY6Bsb12rHH/6n7iRMIpgHchDVq/VkYmReLpxwDresXDXbBqj9cnidU
5n5BNnjfXFGhuF5Kn82fRr87zfgOcFLJ/9hXCTFcuw6fP53QHOXp2wUQcgQCbdyC
SAntlRbr3Ft2D3m5nBzbgAzmeJeCi2RfCI7mShtZXDtC5iZO9Hh97V/pbdwPZd/9
AyvQEwEtYwSQgdCqHjWJ4Qo4L/zZuO/5Su2DtumxNE8G2InT40r0zoDSKLf0VFDD
qoldFuhFxz5elFGDugn++dyS5QozGL7+c9WC+onOV1cjm/3aljLrwP70kYPR5NuW
yl+zHl5HjYUEH1vNh4aqo6Uc0YlI47x/AyZ3p8a85huY0gkwkZGbet3mdDNt468O
MRhGB3Az3F6AhCvbaJnk/4vSvy3M3Mdl7MOHPLOkjnYpACs8Z085HuEZ4CLGHH3l
Vt2V/GSQz2FZk2nAxVTHqf+aST+rULcoqS2+vG8gUPFkkl8L6o7jLvHREXYTpIH1
LgSk/NCKlmsdcBqg1TXKDREV9xkEsIyGdMKUCPxGu3fb6T1vtQ6Gu1o1/7XHm3bW
acLf/QvpE4mp79mVYXqq2LqdHHIcrvyuYWnTgLFrUaoMCapL/TpPla1zHgfDP+Fd
U9SmoTaUuXLZQ7gh4sgdNsjQS3RfvvHjZkdn3Qb/Tlr2OD69PZ1OFbd794ClvwjR
uZgtFl+FRaCX1uWUuS3oorEFCryAmNy1QLHF7RZy/NSDwZH8WOP7xAb/OjmERBq6
JLDcRy4MMiIkDtItDbTGeSEUsmmXz0JwKo16gAbsir3JbWGXJG0tYNraEdDfk6KM
BFU5peZjm1GAWxQ9uAs/F6rOJLLZfuR8rhbHB083hcvVNhLL8Nsteu42GKOHcIbQ
SiQEe02FedgCol8352AZF71+qOjvhTulFR0jzEcfaOCUXZj1S6H73azJJ9SG67Ys
jSJHbWJapa0gmDOgF/qHmzBFYlUmlzk7c00K6FPgjEz1fvr5q/psGiJayhBZJtJk
NQb3bLTzRAguKhvjqw3eUe/68G27a1aCvjO74zg5Xg0veONAoTMbOqxGqJuWIZYT
HDjSizrDOf5yghJiR+qd5yzs1DZtNILWhCuxyCW7HAez7sLg7UfK1k0IMQEtMd1h
8BBGUsyjop0w8kOxUMXqEY0zokQaI3liMOkHIZaVyox/DbbmIGfXbdMrNDO9D//2
/rh8UgnKN2SKrg/w1wCdMYK6sn8LIAXRbQhXR0DghDxbMVrNK0Kjo1lqlNIVCK08
qVjVoCVEs75VC5qGzDqEdLn9Osi3SYEkqvVykBs8q+Z7pnxIPtdojuHiCMc5CZS2
UdnavAlUssu/Q+3eFxIWKA3pN++yCL+gReYkyKhwZbEark+rWoBjDAzLMM2pvvvc
vOu28U0uoADGnq8fRz3A6Qdh+an4dzNPioEBmGOTK/aH+n0Zh5ess8X80FGxWW+K
3wC6W1Mny4jtrahyRovoJ1QaPjaGBkWvGOKkC5+UNakpdfC10IbQBLcZZgLtC6P5
b5sxw2kCkfKF/QPHG5IdSOQeossxd72hBM/pYbXbuJEbsQZ7V/njIcmgRbk49SVG
mzFL3YVoHH7b3VpxjUt2v8EYiVhGAhDlTdQcCrpByyasHBpC04/m1MadrotiBkCz
OdT2eI0qfmW4gCxnwFSrVVteTCkGncvCoxZ/leC/a/w9CgDg+TTnaCtMcGQNS9HB
wA0vSBUuUKf1WNbFaX58XT9xV4zHq20wpUUGU+YTN7h2BrckHpgNkUq5XNL8O3Lf
7GKZ3pDNV6r3CEihZA01AlSaQ4kgi5Fmg53dBjybdsRfEMHsqWVNHHvOEYDww2CO
W+7ptyyUOTlSQ+U3MctYjrUqdb1UdOxP3t3BVU2rdkDxI5qTWVeK2uNginGBlWAn
oEtO8XwUb2CmWRNSDKUmZhHiWWH8akD6xfOxpa0YcT2kmyvTaXY+dNd/4qAjC60a
zRwOYsQgcYnO+8WO/EP+lNyL19QonP4Lwlxvjxv73XZgfrMZN4eRe4uYdslhZH4f
EJYkhR+uNHmlHBkBjEqBE/UNYA7BbLGvtmwLMy+zH1XU4ec3XX/Nr6K5AN7sY2rX
PsTGq23F94ME0kMyn3EbilhV1Qr3LmP+JclGUcbJK7eVAKkFzzHpvSjq3zcFabUM
VpZ3pVqtxMsCsznZ9BGBrGkXopXpN0M4k+ww9qc6Org50mGjvD9pWwXv1zDO8RWW
43CqOdxnYNr0FyXaplsakOaB+u/t/VmLYabhN+q3fdusAAEjJZFVpUR8VQf4Uk2b
xfdb4jXtmgt1AyvfG8KqgRNiZUnwgB0MBu3XOlgTEkhg4ZYC8qFWZbqPvpAJmRzm
7bddwyS0d/j6zbNGK3LAgOzzV0PFMy5k68n+dQh210/oQtmtXdnx2mEs2WnJp+y/
tjH/k+UT/MBRxe5mq1HkPnY3qR4SEVsSQw32ccfykFHLS50PaHH6Bv4z0bxiK/yA
73l5JJmQh6gspHyq3ymIRWgfHXZ18ejjn8DniZJMkDWX/0va/KCdDU3k4SxEO9sI
PutqMuyhJCIcfm1rtbbM69DWjowQoxcnY76uQxWyFiQtt98JWFD8/e6eKsm7JxTb
YKv5aUVshcC74RJcE3849d3hBwIHWH89NbP24ZwKkmjxv93aVZgb+S/JZ38U/dsw
DoxDl94UGVKL3f8qb9dkm/g09OhArJJdpI86D+6wCZn/gMLzcUE/qyuL6rdMRhYE
6k42yvFmOCKKIuPoZBM/RJt56T/3m+KMwE1do25nFdjZJ3DoTUDUtYjqlNjwEzXO
OWIazbY3kh24KdtkHky8yvddhyw3/H0NdSRXW/wS3X46xN17aa26fOh8U5KwV2Za
xGG3yppaKdYu5DoeIk3YGPD5P19WefHfw8bJpY/2gGI6WomTSuTIUhjFHK7ZPJm6
KD0y3PmP0QSLeGo9wM3EfqSW7yirBKwmaqU+xUV/q/HiBYnH1N1FuTUheyw2WkE7
7vfUoMcfSDFS5VDlpKNVtrnwyDqXVgYomHDtRolpYTOQ7bj35LflL59+9l1y8aLp
Fq+75ziDvVj4YjGHthM/8sgcJJjaB4RMpBv0AbnM0o6jyR48/avKvT/ecSRDisUC
kXN7vd/dFD1cECVnGKtOGcHDZLFXySQC8sk0l5X6O4iRBsxqUo//HDdokdHAfupc
rUY4ALLbbZBaL+aAHxG621jzDLSGd4PCq8dpxZtwtxWSYIAJRsEwAXzQsT557zFv
plOOrcXotWZfEwUc+DBtru1+NPRg4CKLy2OJemsbfkVoQZe/ajPFfumkWDMCbgjs
mxQaAlHYPOCAhM6umBcj2JegQh5Vbn6A+dIoHn8nWFaRJbemHDt/iMc0NqNE0cmR
f8TbS/ZkdQsDlyuRL+USmJ5AE4CyhiY33cGVIPdHTdnrTKOsYfXiaorfKJHSoAsI
83Q3Z5awY1hdHcWAUd634USefEu/xfSmeCEdvNbLTsX3bJEBttRNqbwMlyMSDygI
Cm4v0+/64P708WZUBYzBxMdEYRq1SW/sV6avqr3+i64qzg8zQM6emndExlh1NZHw
L7HpSx+d8GP9KziWzhT3teXqcX8JvZth66rV8uPCuI3UAbveT8h6MNrwSYXnOYvN
KQ62zwwVR87zCW2GLeU5yyuFm7PraTXjlTR5oncS9D4dXrGVKSJOPOQaRbXCJXvR
M9qKeEuuwi/s2dkrWjkyJyyviZWVO62Nk9CQRlzObbftZMVbwsJm5lFCXtMj4it/
urv6l5EEuQj09Pt3lelgrCUo0ZTwLmlwTY19RfecbUK7+i+Im3tXTQxwfHMorCwZ
g33yAynubNaTOJxQ+Ct9BxAJ/rTErokbV26apTHgnWLxOAkjSx7wwdG0BZXmNDXB
BvXGJzEF1/Q/6hwFFpU7C1CZre3L1aB4i2uxlY41EFkuCOXpmg7ynLke3TAqZJlo
tckZmKTLg55/CTQPuylmsR2eEg5kcfLRqHbqONCKSfjUy/7mjHpvSa+z6Wl6EOrI
ZyjY4SAOWFonbaNrnZXlEeqUX1UINbeLGK8PaM+P3NE3vrtwunAvgY1MDqG+jrEI
JY8LJkmwXfDkJ2NoS6T3GuisDGESI3HRelOfWcQRm936Xb9rRxmAz/VuPUtO4K8b
/70mlNSBCf9+1lC7AjZ0DHnzlMrGiNOIjJr1x/cODZD/B6trLnFn+9Q/1fj8lmYO
2V4vpuWdFmmcQ67RUF2YhHIOE3xa2pRXvv7HFMT2kksa8KgmSctz6/zya0x2WMEF
qz1rBENW6VyzXLVF+z6FdJvp/dGUsFmfWDyilItwmQnaU+JRnIHsG4sgbCf/JF/E
ZkaciAKvoy1FlJNW05hjU6tKEgwvXbbdAc9lO+saNX3Y0Nu5DiZQqxfCfc5QzKPY
POgLF0oyt46XiUItAIL2Qq+AuZ8Va3aixtMrzfdOkpmqPIwhJj7FLkvdudXie9dO
NRbSvPr/0xIEQ9d6GIMCTjHeQHSzxiXEvZTesm7Xitydfq+2qaufQbDQ6uuEvypr
jwF8j5iW5YJr9ROWbagCZK64DY2bsXKFNmC5C1aglgQrsmiU8EykTPOHreC/n6g2
JrsQRUhbqP4onk2XQjGqaPalBbRqBI7Kg1Eo4dJPTtu5ZeS8G8vJZP8VoJTffsjJ
QF73TwvpI8Px7YfcOudpVVdvoO23noTWeOrRLP91yuhnmG4D33bBkAbDWYsivjwe
Mp51fFTyPEA0Pf3XvR30kenyhMgeD5qXlMmTS3XlQe8bqjmzqDG724OyHu7P/fxO
Bt80/fMsQChWWZQE9gfEwCFlo+XlzxvN2h4VGNV3Gu9Jrqh+iAd2kGfXwaRgBwKZ
glaRa6wDWJzhg4Ze3eiN3WpMW1Qk1H3HChFw/1Osl2h+qICj+QJRzcBVFeVJ0/Dd
hdPRGPj1X3ayqHF3SAA02JxUeNRHB1Po9c2xXvOBh+4DFyEe6worSjTUQ4OAyR+o
d0vetnfBNdSrqSQwYDNjMwXKpYebUWJljz0V7itVdham4R17JakcwaL+cJz50P7l
661YjnGtWLhLqsueja8nH+VgPkb7Z9pt4KAWinCa9RrzuBEI9sdgVpUg6QPJxfYn
ziDzw87FdGGs+MfdwcKCUZRDTBQMYHN/cHSoRVmXLb+S1nMI9TIWHKWGE2nbru0T
whXbr1y127JSRlsXbsaTQrt1FNxzbFriCpaCoNWhWYxeiU4GhcLjlKCnwTiJTh0B
frh3yJh9lbSkoygLr+FPJu505pDtt+ODxRqRAjOv/t3YgdMyVlltWDaKNF85rocd
MPDInerYmMlgpy/4Izsx+0K+1V0tKD86QyuFWAYIv1AouqN6ztzgOEoEnaV4nLBu
0nZk/voDer8TkMt9SWG992s6vuMCOJvX5eP12NOfhQSKf9dvXUPPOjA9pne9Sr1C
itsznTozesMLDgQOTyUj/Bb5n/iUC2DohCS3+cL4IN9Z4DN6k7Ms8Vvi6EkazaYp
um9FLtacp6Hg+b7dS6W8Uyr6iUCKTyGunIHA5/wrrLve4TP5r0qAFljr4eLdzQcK
3Hox5AssXLz9oXHBN/RgZVjM57CadVmSSy787PO2+0ywkBFqCKXfdREEHK0IgiTh
05bgBq+tvlvPIhP/Vq+G+qlfuE41zwAaLeEpvKPmTEv1bmYFx1Qpa5GWKcVGppk6
o2C5p7YI6ug5Ub75XDDHeW2o9xLFvQqZYaztAwPao4wAybTriU5c0xHvLd1vx7DK
ODtFvX7tKEdxdZGAyOss093LJ9tYYxLog3RYMuGyXvsdkPiGpwDQf57OdMMuUjCX
4EuVC0Jfx0JL7LWyzXxpFn8y/s0G3KJ4n2FAD12qzq1mKyu/ngBd3jlkhq4aILDI
0YRXVrH9AQ1voEYjdqjUvxaxXJkLhp33SXZcuj0Tr7fiyh8XWatf4EYIvDvXkKXm
sF/7Zdfv3MHSDrYATTRR8zo5oEaa1FStuAuXNkZRlQhMQl3SaWfN5vfwP3dveVoA
2y2YEO18uxFkmPDCxMBWRkEFStZshR2cWEtDPHPcWI0vxEXNScFwXA0fkuHbknOs
P8LDF8CFRFBrvA/xwjmoSV/gQfMZ4uLqqpJ8caL2XX58arwbkixx/iCDPjQV2uqK
azULdjOYisAhn6MLnqbwtQHptxL+AmRes6hnrso3F4r246UZ6rPma/iY1XyxOve1
By2JDN+K+ihTSjbV7zsnJHF8IeWvacOwuIT8aCfBC2+T/tNBaciop0x9HJtNIZuV
xdInqA92vY65zB25EhTPi95cQEqXcl7KqN/r76CY0fjMD8rzF/dP75F/w6pW4trC
KhytxyTxigVPG9j059gMO0Qu7KrBR5Pd7TXGbzYZABpKpMRzEsFxMu8NLd1HIAev
glsDlyuNpynFVRe1MgE3abB/M3I25bWUauK4AkVHtVR4Kk9qHuSTYTLa5aE7k8ls
YEwf/vbLo/E9WoE810A6c6lpZjAmyMH70WDxmeaTy2zGTF6npK7xGT0Wk8Cp9//Z
Xed8BtZ5nFfhSUR7QbQg6nKlZ2OAn67Bv1+c30Vs5BfvmQDeeK9SXuOb3Kqw6xe5
XPU8J0L4hNeIDBn1nHux8T0v2Cw23sXN2/PlRUsH3s0SX+GYtykRvvFg6y9ONJJD
RcaMksCnKhsDmBAJ2mJUN8yCFK3cLt22b7W5GppM39WSfdBcqC8k/YMCtHj9yCYL
m4t7bxBSNEWIA91IJ9+auy55nTFJECEBkPeVVgyedXE33gqZ6bdKD2q+MW57kIpR
O2mG4s9GPtZqyoreEbAw+9nQDbx7UZ7aC3R+pT9y7kDsNc9FmWOLgr99/5xQ9O5F
bOVdo1Q6BuuOA6fHHnUKjk/00rVswyJd4PQHl+eNdgg6tkL6jn+GHK6TKqQD0p1F
8G9c4DZSAZYgzDikg428P1oC8pmJz8L4n30EnGdRByFse3FMWqoDHXIDYZ6NqwBH
GbkMxnaKSCTToWOEgVZnn/pBSx5BHWFirVmuvuRab+ihbTYEQmN2k6Em/b6Mlws7
YTKGkuX5MSI0sBN07x0yatmunFz9kokbRIU1WirpiX8QqoInOSYpzLGWzYQgo/cm
5g2Haetgtoi7BEPhUY2O2g1yC8Ds+FqBunwTMj2FNAD/P6asVP3h76La6XVfKc2b
lznLMeXYBymh7hIjsG5AIvI6G6F44EEAvbDGo9qDCqoUc7ZMQZL8Cg7arPTKT33c
5zPoa0dFhdrv1lfCotRQdYhqJ74gAoanec/+s6A9Fg9uC6CBxO2oLKvf7ZzGHywV
bmc/BeeJ5M71pNvpzfmRy3jWqCkbFJmNhdzuCovFKeFBGisYQTXrEVF9HIarqn6J
69fgqGHGKItOrvtYuePKqzpd/RfCL00STmA4qma7bSqGODo6a7zcOAKsTn9xGzhS
xxPMZpbrMlKIR6YLqXcLgJEqLRkGp+s2fW6GvRUujj/FKsOGqy/B8dcHdxx6Cmrb
oD6M4tlFi02HnUR16EKTpMvzlbp6veaYKoEcStbP9EvltB4osPh9FOjdrhbwtku7
742WY+B/3XhjeOOUr1RQsr76+Y94yAjQjvmj+qFNYgNrtLzGNe6h6qe88miPS415
FUGQKlEi8OPIT+kNLvt7CpB1YKDw5pRvPYJWon3PP1iozyUE2BDYUbavfyp+ytL7
rwuzSSAdsPhY1ByncDABAV1w2Jk4GUtAu8qlBDoOZ1wiHJ5Gx7ZcfWj4R08CCkqD
+gUyGp/HZ7G512UHNyHaT83ybzF5iOFzTJta6a5uFWMSMvFsUcnmYywkPqac/Fb2
UVCNIrz2eQRgafu4sBwP9c133Nl7f1EqqjPqCmAvroEFIThiVCbpQ/P7CBpmQB0Q
XabpB5ZBCeAjVGG1L/cetIpwIWL0pD+AkVQObAJSRWwH+SwrTCsSR/Cu2e0Pnqbx
0iNQoXL+3O6D/wevV91ePPKyKhN4rjHkBhZKmBOaP6sthFuA4i40stLPYee3tGjs
zmRn3wJTooeLrz20pFNRCqPCHaIQZkAAv6jknEfJMDsrk2tu64lgEfxMfKJA3ffx
p9KROwM6f+TG1Tn0EXOKEukuYvMYB1EauFrJltFaInMpPnyKB80r2Dbk8IpgcZJr
Yb9MgKQYFEmzq3wplqmoY/EDeUsKBCrdjsI45v74OjIfTmPp8286rIW37Tmg3PTC
spv/+B2yyqFRAWx+2gwiuGbWj7iLm0wDoLv0q7lhr3LAcuz0shoTl3m/FWjhxRfi
S0S0tcctva+B/7ArQm5TMLBM5Y8zKuGrmUlY3vjGXsC1CRAW9uQpzm+/nJbs8Ig7
U9ivr+nHIK98piBp3e1ZLncB4mwIbxCMMfynYWKt8ofV7qmYbzhyGBkG4s3xAYyj
oTzu+s+BnytWMUu9+I95SU7ctXoVrutLlL3qZPsfYVDS2IffvlREcbXe9VSzn3k8
5RylggCYb071BUCioi34h7/4dFMbqbdS374PTVRLEmOIYmHxPvjkbILURALw4b+Q
y7vNHzBhPG/UTkPr2toIXPBm8iCHj9d8KPzz5pHG4HrTBE/7ZOWYdiPdPz0jdcum
ZpDgM6kUIlkmXfrRHZNnlV/3Fau+7IqPBD54zSXkAtJdDhWsnTx4NoWA/2aUyH5P
S2SUtLTfK7aISaqEkdDAsSdvKR7Ze6u695d35IH3n/dVSOJWcKJovW60gWYEiIZ/
0ZrJkBbXoN1u0fyhm6z1nwuxoTC4P5wo5j1jtABV1mB2lgqcxzEFplVzyxq4/HDO
39xriVrLbRLTim4dFD91k3K61Ol6Jgq7T3EVlPvJVcGdtBWtUJCbd/D4/A8bT7pY
qqZUbpA+Cco7Wmxww7DZMDNXn4zjFTgLmS+eYblAArocWPmr+BEoL4/4ICQCg1ON
TBRUQIxvbfiT7CdDYu61A4dYSsBvR6ec69UcfLu7GtMIlWwpv+9c1QUwT4yhCTei
SYfzvutiztTnW/daRrS7kD03sli7bB/bUfAfbYhBj3+s8XPxgo+tr05ua9RM9rup
96ApfiVCH7onqeIpkYg5SyV5ctXABTxfOL2HkxE3SCQ7LWKsm+qonYxhMkCM7gUD
Qi4hrOHRe7zP2Ca79nGNXy6vk5hgo8sc0amekMoUGH/y+G891I4fwlV/BgYBToG1
yrTjbfiE4A0EUSl1MDQUH0nSmtI3kvEVYi10sRRpfXufZMu5CsQIxQsoui54W4Vl
WBUWMjPFCcG2s7HD7r8Z29qlSm1cUIfbHW91VgGqv4JtJPEtaOKAriHkmW2UCPMH
kzYFT3bPrS2RFQJqDD4b9xA5HipCcJYVHdkhhqZvHu4CPk91AlQTUsUlTj+S1ALV
8BX04LxROb2/k5H1RTHCS+r1EZV4b6UACuCogoM8SHkuyIXuT4vJmXr+a8CEirNb
UTCTPofB5FagrPYe7STCw3/FG5Vsd+7aus75E5gYBlYimdMlMlpx26AqHZRGAK/5
L4mBIwVxVuZj9qV5gmaqn1ihu/I85PRZeieaPwcjov7LoRRJAsIXK3E7qfrMWzFI
Zc7IIZSOMzKMfoX1A0waljw/Mfp6VefbDp7VqzCubchSlDygrOhhMbG122ntmlct
E705hamxiHbBG+VO6Jn3fesTh9+poeChIQL4sGthNZxb6HpNE1ERhj2awpMZgBk/
5A8X/cqxtn+qdYXGhP//zNld+Oz8s2tc0mVpn9jfNGYcOAswzY8RFpW70xYPPQ5h
WSjUcRdbuK2AjIwfvGg2wFYwJomu3H4JsjZvpD/GvPhN3XBP/tooaChgwHkJNCl2
UKOSCoB14kL11pAhrOhr/7qbGuU8628BOzU4nmGZTDeDHDwzccghF9Hy62nmHzyU
TZXtZ93vnYNZD5tGDF/h8VuRM0th1XlDqNQHcHjBrBkapJkpolMJ4Ot+LeHId0mb
2+K+okIO76wVHHWYVIlq/MfjRqfykCi/p6vGzfDlg/wwZR0RikCQxz5CIO2lMfWu
1CAw+HM6uz39n2exv7+pyltm4S2PPAxQEDR2ItA7ozkPZhJDIyJk75mxXjIdGyrr
j542D974s8HaggIOrRSE8o9ukgJTpnUQLIwtUpGNBWEHXhtsa3r+kaEw5H8hX4QS
2CgloBaHatsi3JGF52DqLtSIi+nlPf7dLB6+uT6kGAt6PfTG1lbNQEaXRNvplKmv
D2AyHE64Pcz6hzpUpQpL7Mne5iIp//ZDwIdVNW3Z+GiqJIfOY7Y4HCCJk3x+0kTc
ynJXsdw1UqlqT0lw3298MkY1DKTphRf5fwQlmPZ6zqmompwceWu5hUHnq2PCwWFE
LyV4Tkl4gbHP9TRLcsO28Msx6oVISHDiwt+ph0L7z5Zha9Jw5txAbShMrY5WbQ+d
PqwwwCoUX5hjw0gdgAM2pL+vtrvNaYx4ybp6/jxgx6fIq1QBENcym670ttfzsNMV
GpmJibTPAMQllnzUro8DDCMk4adsBnaDsTpcJY7/ixpbDpvAZi8nQOYsETKqCxS6
U6kLNADpuWo+wjti/weHxPWoSOBHIAlMeoV4m+w38jxi00nSrsVECx4X99MpuYgk
/GM9nM7USFclFBIPQRvT08VkCCilr7+2BtN+5PT2Q2g0zLUUouIK/bpENY3VdLEw
T0VhSonHwB/A7QyAjOiwmyi1v4vbfnnEbxN5beXyb0/+RkI3sCTZLurCEmE/jbRe
m6YD9vCzJO+FCyKuPrnTofiX2O5nJfydHESonUUhLrErX7bgQnCTUB9Kl0VSogm8
XZSCbh1h0S4CdGKlsj4mZsqHxA3EJiEwTHQjefqN9lwmBoMMyurXRRBYybTJXp9L
Xmdh2QsztLDkdERhBhJsURwEGtSFUKSrECMr82z7cUbSm3NHsR3Weas0PUQWe5E1
6v32W4C2ZpAIponWpxBa1pqJ36vDRZlUnQpB7nRowDOXyBs2NJ2LxKHt72nE6Uc9
PRh57oQXuVY9CpH7g2YiusWt3nIx4aXXOThtuPaamT3N768aW1wjZ+7lB8Wiwlqp
3yt/+theytIvKCW1VF9c9KOz0aC7n5uuRcPpcWSuU7hLAfiFmdsy9oJcxY+yOqm2
zsNq1XzKtTNFWEf+PVDjfdRiaSpVOkw3lwZKbbBCBy+3LlzCiwmd7Zs1kkh00L9+
q6fgFwdIxzHD0F8rp68KEhhor77xZabjRDzG0WVz0HXf/YZLn+wWyo53ezrLrJMQ
19LH2VuF3ywqhra5Q7L35689d4l6qDQqNEhTB746j1ONtXpzXadfOhCMzZyEKiEP
F1367NEzBgBu2Pl9q5BWd/GWwT5y4pQ+3yyioqAQsFNAFUuG5QmGtRr2uyJ3awhS
u5CrpQYgfNHB/5T2eM13CEC2S63LwrqI3axbYc9KXGPY8JriUxIwS+2je5t+0dO8
NuzRW+iNRFktHEK6JqH0UUEQD9O2oClt8i1MH2Pq8Vt4MD61o3nJfvmQLjbqPhX2
HyBJ9H/Vgl1X0trIKLNwfhN9VW2oLDEzzgC/WMM/su1XOyuhZNCQ8he/qgtsXIvK
CeGXiIi7mOJZmCIg4/3qdJ5T0PMUuxBIwC2ta5s4btCfGXFwnkx72PEUOy9OzIiX
ODBIL/UIsiTPBZYQld0LscTJdn4LobK+Wqrh/xElsDR6pbY27qv5xhqN3wNdoYue
4ODXElpiniJnWr3GtQGYSiWLCp+DWSjgYP9dGmkPx22BqgorgfwDnxJbJo3+iJxC
xl7eL7tOHR3APaCIIF95oMWILyzkh5TpBjFwjmobOr4hjEPnlMDsLKXsH8DLmb2F
VD2BFzTcYbq2UFDP2YHyTPy6zzqIZHy+L1XXl8BGBaoo7N8a1HEkc2nCJEAOMc0Y
oZ7ups0WZRjPdTWcbQUqzak03rBmbsb2c17XVbXUNU+LuuNRUlZ1x+ePF9FvvsmI
vTKWI9y9NfqxSuekbqZNctcJd2WoEt1iDP0iuhYDX6xdTl8v5jBugiPM7vxI69o9
Llb+WgZQ8l7Oh2rb3K20nLh2tohje7FVn6VdNaz9TmESLk7ntAaV01QLkFXYptja
WvpME56dXXPWGEumwp2LcaRYRYRS0OAMorbCTWB+i58l8wZWTBydeZ3wyyiydqAf
AqpnbBQUKluOM8wNApVaHoVosnEiQVAuObtOMAVG3dCyJpFJFqCTiggeUUVVh4x2
L69+H8EWR/g3lEdiaJunXTERyIcAH5F0R61NwQO+wIbCGDtFskqPXSrbQbjQ0iqG
XtNMDC3fc8rLL+p+OF1f0n80EeYU5Vx1OidbKOFmCYkL/tyGlIRDLYxWKGwFI+Ik
A5XBXmZ/DLcpNng76jNpOALl3LQ2x0NQyPTVMnPvSduGjx1qrWhUY29sk70JXtgx
nOIe1BjrJbX+oqAsSpwkhy49nYBVpfKzsDmkQdJmVoZ1C7cZwbiwoYTfx/hL553R
UYJBBVVKqRxE1Wn4uxTjaEgBD1VP8QZ9VlYZfFy6gS+nNZsT9nw7jZZAxi9c6/mh
y7muRSOGHkerLSUw4DqorU/ka8t4je/08bFTJ+0NsTU+m8UGW0ZhcRi3i53S5fJL
RxswyyqPdRisVFzHCjjVb27LclxWHGDXjnzdON6mBdVBkIYPmZLpkTJVZl8FHmrc
//oAGsJYJ5YPvp21fQskj2FBhDbKrYDWlrcIFnbTGt/l1nn3Mb1Fcz24kSs3VLyx
RivDP2MPSGHKF3NBbd4bHe9tKrEYhwtI8PO8eyf9e5zXIohsPcz5CMYAp4VWS6GX
J6NZoNvBg+OcAGOwvH513e9dAPDB0FfpHaFX5PH/QTy2vD/W8pc3vRfcGIxagml5
o+tBFZxAdvhiea9l4HkxjyvZzrBmFYbKQxAay6wxFILoqEJ1RwEFCAImUJllzGHQ
IYlVV58AOhQk82Q4Hdcd/H9TfQr9TAH5/kL5mdnYnlwUVOmUx6+mdJoBQgpROOkp
T+azvKSoHSQLk8hqzs4Ogqg3wBy2yl4mprYFQNmByJnOKICPjR+0y+XkHUuk7KL+
nOM4LPuS1DYXzm/7i0SvB9u5iSqgKGWWuE73bXw9r48sABFX7BFTgEhVGfmh/YZQ
EGPCSqtLQpB1EGxvNahaCtahdzj4/7j/hlY3ibN8H3o9JfWt1jzeM3DEQsnD1STV
EnJEk+QP32tFFVgCglhV3H+uiIjw2wnd7Q3VDE0xnGKhFtDNVtOUXRL4N4/E+9bJ
qGo/JP+mhKAkDA9sIH8fpXnzhD/rkD46UYpzzOcz2+7TSVIjOvuFqxJLNDs9mDZs
dyfFVA5kaefcVpWZBq87/pJ6Og3ewUbTn3/SpKMqVLUqa7EKNxtRWKXfxAx7gO5W
cyg8w2XvPY26m22rid5EftkdSGx6A4Ft91DGmBpkjdwtFMnHqDI3gFOZ67rPLY22
/nDSwCwESC77wlccPN/U3yo0d4gTj/Dp9/lTm70LMvQmFvOKB3e50qCp1SW8OAdS
nSHRYaKVRMI2HLk9KKO/u2IPKUobYFpYFK1+ayi+kagqChkSzyxnibTsn3msAIUS
S05tSKO0L6vfUD4xO4gNmOrctMQQ5I7cyis7XkCWZP4gq4RhjDzPJ3shhhRH/7hA
84w7E4D8YuNEWC3Tw7E0n5bw4fe7/Gi02F1MhOXRVvDn8M6p4EvAb/cKkukObVl4
6jbPKYqZ7owG7dJ78aszZTp5qUiC2m0FSJVxVPi/Weg/HV2nwjcMGWiGgcu7wfZ6
LOVFL0uL0d7CvY3Cta0mrAsmGDlddfGlswIbdEL19CW5cJlTjarOceJjyZQz5PEx
pSbiJdYyHIpGpzG3qaJDIeaL66/JPVfXIsyPnZ45w63SDYxDjWijRZn3f5AXnxAW
xVeVRfHz7/mn3/uPYGgqm/ebl6diOuvtPYEKH6XR/cS7ju8+HldIbe+VyZ+YJ6a2
fqV7S9R5WPbzB1RPAlqG/b7Ls9NWniY8g7jFtETvUDYyXDyEY3sZ2QZNbfxcRvzg
m38uIsEA5e0G4ryrShvnIHIqk4bYJR7RTOgOU5NNk0U3CRL+lmQYvtQndwOmXSUd
LPRXGEzwUCh4kk5rJQGqXCw5EW/5bWf2P55D7FLBbbyfHQcUHDratwSHuiCNM/In
vf3evCtuZ3HVmWj8/YaURtt5J0uw+jfru3FH4XmzDKo+Ei1Jq5F+etaujWEvcugk
AC6ZwqmxGqXyfJCYrHEY2hZtVr0/B9UX8sFFbqFj3wAuJAbTWZCk3BYYmL+2xinW
omZNdFvBPvtyH0MaT+jdof2n1LG6bXaLG0LcRz2xdgsijUyHU8eqY11UxQ+4fsLd
EX+hc1AP3s+gbVJBhDOwrfWzZq5TcRyT4tOTLFPnAsxMWtH0FS5OvwuPrVwqoTin
GMZwKk9zlc3inyb/hzGu8crz362AL27zZZ7/9LG97q0ggITKe+xApQg2dSTlSCKf
twmX+9VW4PlL6sXUgYyHhxpcxgSuf6tJQ9YQuO/m1gayr/ABQufM7596aOu6hpW/
AUwWYRj0Y2jTBdn/LNBZhewisBxhmJttrNlEd8aaxNVKwozG3pZtKvPySne9R4fW
ENFWBkWuFnZqipU+NFJbUPd8ruN+4VSPW/b1DiWC1cRzEXim111cGaRU0swZLBkV
aVsKcFS6euF7wiDWs2EookfLCTttqz6F/gpT0NYnrogTDjtZMXFo8qFGQsBbfwmf
cEC+fNMR+hyB0qklGCv6Uumkt0Q9N1Sp9MM/VCs5dK75tZ5CTr5bu7ZYTJBtiJfO
ucYMMzJq76XjXFwf08EqX0MS1FebGWK0wn5Xbgn01DOHjdVYoI70FuSyU4zMVSDT
bR3HixB97JyhK9O8ZRdtx+mUT6Qu0orwaCUFlqgszsBioS9E9EpuCrUHXZd5FIsW
sDuQ04o4gSoZubBIA8W9sRuHid+YXNQX4O5565+cANeG6YwpUyqKoX4Mfmc/q7U0
dxRbig14YU6CrWULadYF40EbR/XA6Tpn7vg43cTxY1Y/bjC70Nw769LtcbyUuAfn
R+kYTOG6IRIZIXqSv3Dzq3WXJUpT5YsMul/k7NjIJ5E7lWTCttkeYGcW5IRPSmE7
nqzYGAwJu0H1v1f1c2cr1wDeH3xjgOgLfckZlcCwp24x+qzLzWTw41uTQEXYpomq
oMirYpx7FCLPVOgodLrWw/6Nd6ZM9Q6DVDtxySZTr0x8sObqYyyE6sN6aFY498VH
pHRM4kPwQrte8UJuiTrjLxtLwi3GJgFs8XIYSq+I+0RAq50DmiDUJIw7xx0L9gzT
URqp8Edg6FqzEhdSEPFF2QbJmCY6RX1WLUy9OMV9c+oxZkbZMTepRr+tD8H1iEyA
n9yzlVFWcGpcQtgSkDxZGuQy4VdfGFfWrQvjFivFULkIoV/rivD2d6kjXLHy7H8L
63FXnq00ZRdEl+ww9gFYqNah2/DGBm3zk/eX9LgsuvvTzePYzJ6TF37FK2Bd4suS
Lqn7kH/aH8ryuLShfRB1XSidoY19DA0cJVvOAfJXyYrhKPN1C653dPppGEWJIym3
eIGIXEq4CIHxkWc5VqaF3p2VOdga3wFgWsSmbJHNRZHYcYm6wVA2A6nTe9Gr2SXx
9T7ZgHSiEiMZ35k9sRd+bKoQ1NUUr9v/YoXp3PWnutA1iQqCdxXsPUb7xA4exw7T
JQIHUJbSpnXwg3gBhlnwoE2ZX7yzj6GjVO7hjvqAbqmMvyDa5zgBF2BPZaEda/au
86WKDTprK01LrPHmzGH5Zk7MOppdHOFo/XMO1oXgLAtKqLMfZcpv5VE068aCeBfx
0ihzkHIgfpy7QkgjasblGaKPT3E5PkgPu300JH0t8udBQJnZITiIjk6YQOkf6ncG
vO7mDISUG1URgdeaNxH2UGgAdpR7ZaAZ92EdwkcDMn37iOchlMGCw9/FgnwhZkPN
qhn+e8hjbdiHRVF9Hi+oHEQaGH+BfK9xJzLyqSaDHyoVlweeo4vWUS0EONOrcoOJ
RK96EKZhdfFL5YPSDPly/Rq8Wfb3rL3E6DWYmp19UH6S1etl+9jzmzUti0OYIfqg
zNzF+YH4t3cpkESsU0gs96bYyQgxDwgcQaKOgFgyX9hCrU9dOjCdbF8pM7ECLa9F
L3hMrD9h8BUiItkSbiRtyMsDWwKzVRUHXtUJGtht0fqgcxD7qdDp7cXFmlXttQ0s
0v9F5avCqRW7jnLysCuY8Sw5l7k/h0ZvVDxF5JYoKp1Iwa3JRShnT7c95+tD91kA
WDxx+V7NFWXRSF9RyqWX+wLV88L7FCTIvy7ympAPy2fN8GuBvZEZ7k0oaQTKPH+j
1IwPrTvi1KcdYFJEniFH/NnNTC+z8dmEX97WYoHlXS801xDw9wWtzxL1F/Z9qN+Y
b06Fgx35DzbpN/MbRkoccpc/Sr6ND9/6pvjhVC1ipCZiWVP8KlIBlNYMyDRUuk/0
ZbccX+KANgsPtNe9b87+lPwKiAiSvqBECJGM6fye9/vdrEVkp6Ar1TgrLbApN7jI
Cc4EPuORRYCc3Kj9UiiAqA7VPoZOci4KF1Fr4EoJQUWjz7/dYBBwWhAYKY7F95Nh
HDYi5aQ0iZLiTYk00+iTL7yDTHU/KSk9GhLNa8+UB1ucSRnlIF802Lx9XUlIWK0o
E5JLqNWSredFvgJC87arMJevxWypdkMJ3BvgobykJLCA427MNGLIq4Vvap9/JwaG
NWTNIPBHmM5c42V6/FXdOLJFWeyNuwL4yTbaL16/Oux2fZWefD4wG1rLLBpq4PuT
mDMU85e+i4hsPwLpaUg70mPnD8neuxZyh7XjoVB5QsrfGNMXLzz5Td7PWdTJbVVB
4IazUPYcgzBD1df2Q3d8Xch7qtTGE2ENzpGAI6AieTsNd7XPruNhofkQDNQGGgnJ
YzWyIJO/uxGcY/wNTUqvaj42x/INLux89yx7wEwrUcuShoB85tblCI+YvxrC1TqQ
kCJTK4r99sW3TvV4N7Hya5WnC12C7RZ7KTDVgQ+0dC5sTOB8l9kyreSjarY0fWlk
ENIDpxFofWNFcTKG0wx4nF1HA8LBEuiNk1VaDYEmLVrhQJ1hLzGp6TIo6OQmUC/c
JxYiR33xHCkN/5sYZ/mNpaxKO1PjMtPIrFNsStZuCsqVlqmawBPwaKjti3vE+hRy
FjlWUxtKCaJKze5GMCmkR1xQucMWuW+DhvDnFgMwydXqzr+JsBnnC5CY5QvxW7Pe
ch/AP1RgFeHtF3OaAtSHmlb58jcWtzQZKLdO8pbhlVD2b8wSQuiKA2/+jGho/6sV
KZKWExsye6LbEcRwQtTgtkjj8PtG74XmXJPAQOVyWDvCHf0I5AG0BgY+5+fSuSDX
wV8I+6dP/k61xJK92IgxlnVhAI2OSufo4XY9sHK0IP46D8r5wUITQBZ4ijuQQb24
FwroLccVJUALsXgb0s2UpNcAXvZkjhSYo6KJzrFVq0INkMHP5Kl8Jfq4vo+yQztN
PpMMZPpSXZ3ec6KQWBljXHW4vWzRz1ie+o8nyi7ktOqYnQg3VupK2WPL81joIfBR
4xBUAblOTv4RxjKdV+JpWQBt8IiAExiGAUlgJP4xiqNknnsaSgKlfPxvhL1d0BdV
vnd21QTxkBs2pAXxVxgktDcdWGvWw/EfFyh4c7eu3J3AFt7IJDOKP8Y9vGlNX9eo
ZtzlfagfpWkQ0F//1knxkqumvRU8D/QP6Dc9sM/iZaUorWcUVCQxEejwNg1KpVaT
7q494NVg8otqVKEuXEsQBQKrgmJhyVqIa1bZa6JXT+lV8H3Gb2/hXpBxVRSwbI6A
VOhxXPAg1whma5GuU1uPw5HbKtzKehX5etSHhi/hKI16TQ3G63bA7ak3ZZBtSJgC
IfI4B0sVUe6cIVKN62LiDjPaUiMkJI6nTbEAenmQIOOlOLC/VdcFPdwSQMkxfmlu
JWuty9ztfOE4B/dY9JF47TrgKf40E3Qd/3whDOsamwl3ZsRzbwNe7OmrueI7TS6K
+9YE8H8H4qPzk5OweOD6Xds8yhjUXEjcTUNoHP66MJAbzvbGDZ+Nwb4TMrYCumjR
WeDvj4xvYJEmX4tFZZB+e9eAQUwb9cMcTOgv+cf7NMIt4fJi3KKNtbXCe2WJ9TPg
/+umtLFKmBpsyKCLvo8OZTZXcAfHCvg40nWSh3KPdK5azAxOC9WGfxlH9Z9yrIY6
q/l2dB+HTjiJfjHrh0fIbOJTvhkoNyK5H8RSevZ1Qcp23+1f98qdEh1vqtZDHE1r
aRI9joNDMU/5dk0Nl/wlGxO4eAMQvv5jgo+QhB8qXldh6MmE8fzO8f9WrRe2HKR3
+7AHvBVIHlzdv8JuoJzG351VwAH2LgrzmwEetQ41Sr+F7MiPWOJdUO+f+/Xh+cHr
T6FanFGxSh1FwBNRrmrnhHZZEfxQf5iF1xTLUsuAc7uesWpzqOZ6lUDcA/jGng0Z
r8r6HFBbe2oLsL+u5elW3MMYsYHkbKTA275jF8Oml057X6atGbhNLRiDy+NyqpVL
ep/c3O6Ts7Qz7vbKEJaI3CnsuDdpkNQtAsaR6+BfuBeCeCYzjnSlXxpVRIUgAYNj
RBJjPCmqRK/liJKG96ZP11Uj1d8FjGZIa0DivAcT5ySF17LN4Tbf9v0C+/eMJ1RQ
Xp2LcuLCmIuHrhDu+62Vbmw+020ZMTdomICW4PJ/hcHKiVF4ZAaiBW6xvSERV5cH
j5oML2c+IED7AsKkhV4ZVRBJz0Z7WIm0SYrYkf6a1rROCwqTDr3aN8N2t5TkkQe8
RqC3vT1on9CBeYd3qSjUXavSqJ//sgWMvTz3jEMj4gjJ15NqQ1cJl4mUQVnn16sG
zp6UHu30N0xboiOPqHuKIdFv5VxyqXwFqxOMuEx0UkofwzGZCssq1LkVDrCBuhJ/
d85ThVbuhz3dXPeWM2wzA1IxTfnBNKvQaPZenudnEfmJWbdW5z5Sm0px6s+YuY6q
EkTz4aS0UBexl3LkZo1a0N25Gn2OLrPsc4olSlRG0wgOLpbpx7XjP5jaHUyoEncB
aG/tONCjrMoUnys5uD9ZHtUowaAJtyL+ghMyKiMbqd9+F7+fuPW8V4ZvxmbdQqy5
cGd0Xy/4/FRLzXKKt+KlGVsH13kZI0aTkiXAPNeyUi3rcaOE9xw6q0hMVqF/DFxK
zJugSLWHT+/kks5oWmxfBrhgL7zk/QTCoLlVw5RBKVCmN7omH0HPneP14LmJdOQo
WeBhX+v/KJvVw3ru8S7JEjQ6SrvW88xhvDMLlRCquvcRPdjORtw7Sr3zy+oOEpdS
q2uyB9tAUNoFvDZJPowq8zaOFc4UJGkEuYgR1oEfZwyUjsLiyEnsTH//SAtF7PWZ
B1Lj/jmxk9EJ3zua1TjR3jNEImWQMPbDGZL/68iVXzgSsSHI6B2SKYoXA3EDhViH
wGuxTtqrFTotSvMwMaIhKu5LjOW1zls6N+Mxh0mVP3dwvxMyFxkcPGGt4SN8SE+g
LV29JQiW93C8pMqnIgkIWQQcS9cQ5DHuTuiFEwjZoEYpbg+8mQkV0oQmx8f8ukrS
2+nFfU8qu7xdDPN+ZOF7ciCwHpbyKiUbu/+Pbs+ecjfgzHy+ZHhKmJDs9xn+uZ5i
7uBBT3zJbjPeqTwSNBA8Yr/j5+MZERVX6dsSsJ4wfKzcXFUUwCnpK3nO5Z2W4GEz
an+pkftwbB2smgKDe0tZxTIapkzV19youkZmXpTemrRF3GwZClHz7uNhe6HNW0z0
D2j7VoXE6ZTGGl1zO9iyL1o9Tsr58ZPhbFGeEnTWDuroTvjwfL7jcbhrRpJJCjqW
RlLJElcer6vLfd5N4yxeh11nhGdQlgwemX+wD4RXzo5EBGcpQIXofuM++fLfPR+l
in9MwpP8VPDXnTuNW0rDsL5XravnqTSzPunQsfv0QCl74IrvAS4+PwhzrgxFZZrv
3usS5blb+zjgCyDlmO6KDxmuiwsxLhgiaWoLAvBB945RPvHAUwpM+aDK0KAxhK4y
7sVPjjQvTuQgE7A+0iSEx3+w/VVp2vtElSm9GvlgQ9PcNEPeO6FxGj9PqGOFps3l
MojOEAPdIoQ6M6gq5CAwSHHKOkNcmOV5FD8fuN1QWhBO8QJxCeuefniyCxMP/Sek
CLx359h+hkNSYwWT4z7aIbYwFDL5Ssaz3MC3kinnPRENGWLmicHwu4DkQ9lVX+5r
XUu9vq8pPqvyf130B4QxomhvmNxi8B0dfRL/6RfYmW4cgbt6KNXe+mGY3U3iiiWu
iAxDm1/rmSctykzYq+CZ9AJBejDdnVspefg0PF4icwdguV5ERjACwbaPzrumrtAN
s4T/d+9Ja3DvY9sMbCHNKl05stk2he9/yWvNHgIZkj9YhVdNCypR8lBGj63U+UQJ
QJwZIfJIHmyNb967dXlwr81Sa8PhnIlNupJRjVY5DYIBBeFXjOOa5GmykI6VS/Xa
vnPg2yRWCkahvT6rY9I3sYq574qa7IExPSWHD8WnWVdqrRnShs1fg3Yx3Mwym5hB
ENgoAnnaDmsg4WkrcqSXGTJ0OLElCESEZY8VGJgrTIRq3PlIE4O4RSI+xzzgmP4O
LeQ9DCu3cHp7qCyS9p3wQKL9AmpevEGv7Pdg1qhCp7fvvuttmhfIshaPDZvcFe1/
bg2dt377yS+NdMfbDFiH5rypS23M+FB1OrFATSo8QdSmms2av1yKd/x+LW0Y6/7y
Iq0sy1rt0cL8dsMn9m5WwwfBUbn34jwRKPCX9Kme77KTZcQ0cltg3jPvKMSe6q4z
JoerV9GkYZNPrj7qHCnJZOEuBLGV9Drd4oPKeWtlo//MQBdfwXC+Nuk/zxgOmbJd
2mKOOd53iuCfeHipcMaNHhm5aN79t/yRhEKuO0dx4onZBRpawa5jlBe+RcnLWr9U
BdDgCzQc4/8oX4K9MhlyToWTNzwTXoG+IhxZCPhFnqb6OtvqK3+09TX5grd12uO8
2FOxdJD74uTDaDsiNdFqzwMb3rb2YPZCTN/S97hfV59ckc+vF4/7JCk76C/eAyho
AngP3Q++msXFDeKt4VinLMfYF89qHngWSI113dbtadQqILA7JsxkcQGhRPILVGwH
r0335bT7hbdf2W3E5Cj758MbJ6YKllWap8BA9Jm6yfdENsxdOIfmCXxNkXA+hoPi
Jqbj8lD8am2QcHFZx4ALRkJm3uVYA0fll93CvEfGWH59bgGLSjfhpdHMO4qv6u/n
u8alGQ/I0kG5szZOPSI1mZC2h483P7L1dbivOqOG5ywhAIqCprj5fbAe8eTjKNO6
xuVH6B9j18iDEAbo9GsRsmtEKgjHMokZKyQS+Yh9G/SBrHTa2EU/BUt/AWi/MAgo
xFvm85q9ZqE4imEStK38UntCq2LOHqrj4RX66G9gl5Hpb+eb3pFQYTRJ/flpW/g7
JqDq1ABKLoEta3La86xTgPlrNS6Vtbhve8/eeIDr5pQ/eNdfaXI+PlMJovVettQ3
lGA0UcSBG8YOxPlrhZTRUEOOt7UIcZqFJyI0v9sT59Aghqd0wF8IXzb/duuJ4nu6
5pyLE3lfyrYBQQXQlLxlJPUn6zzKWqen1z4olJhQeD8Nbr9AyyXdqbI3sbgLi0ik
z9D39Yyrj4saFZV9Wo9XPNXe5A/hWq0sK5TPyEhj0tmFlYF02l8dCEBjpMUn2OmJ
OC1MlOFgK532dGZhk6PFQ7hqjm5XE2DsZkPq2U0kfzQkEaiDT2Y5eQeGQwrYBQ/E
TSfBOg/9NhfECHR5mAWY5P8mtBxhVXrREFbypmx7wxSsl9yo8iHMP9z+L+NaW05q
PFrnh3K4ssisgUsYlzGblTm5QHhEgFcT98HDr2ybhxeGHHKTEtZJjq1Xwt9fIBg/
vg1CTvN+2YnABNWgpuYklLEgzwU/hb8rTeHDRhsFYYpgBUBgLisLZBFV9TH/6MD1
Xh0pdRTKgbFd2V6xWmYuB3Sg3ahckF8NDMd/+zqA7qmxFKyuZsVHY2oVvS1vhkyz
EttQsx0U7Z04lQgH9eFjzZKWBupjJk6sr/e4BHnvWkJu1cfiAkfU3pJ9Z0Tpa6Iw
lnMG+XXZdZeh0IVSJ9GKng5lsTbxtnEFWq8/0smwPdlF8VIBnj2QZQMRIRZHsH8E
ZDSRcWuLp/bOAp/ABHbwm5EG8GAmR38htjCeIohmQmB8jgZgsYx00OE0dTb94pF9
V2CjKJOabA1SCDrovHgSQ0jcr8c08/+TTV0KFzx3KqhIi/4EZaZlvoVQmeIJ/cWy
ZzE/cMZ+1gzB5QvD0hdgfmFP6tSEbm+q8rZkxep2ezoYa7hcM6fzQFi2EBIbqehI
MWsWvhqmLibWnBBGYBYYqWixEjKKKgaEs81q1oD57/mGoylgwrIa0g6Vr6SGAgTk
MM+3VHSRMSkAFmDkkcKAoZVbYvCf5aNpU/5Qt1bIAfzJieS4NGLS82aT+2qPGtRT
f8DRUiehw3sd01ZqyYVoOX6ef3Z64KVwLqrfyzuzuNKf2FMMUKr44VXYE/Q83Qk6
WB3qprOmvDfsBWtMxCkS5VdfojDNNvLb1/gds0TggRl9UY8n8vH2fFSa0sPP2Z56
AE3oMeDUTHV9C3BpksCoLV/ijSQLF5Av3UuGp0BkcomoX3SepnYzbpu/k5d4hHCB
xeDDwKiszEsYYuEUhDH3Xpyd6gx2Ojl0KaP+7snsvewzf+ZtbDhpM8HHjZZMhT5T
wXSGQNjHW2AoBpAq1Og6dGlP0bKb7Cni36tTyM6aU7IU8BJN8oZGDvtm7PA/2Shi
InA5ixTEAFilNQEam5BnpNH4T25Hq5GdksZBEJeDNrfy6csVTZFZG+zin3ZK3tZn
lFEoRXa9x1ze4tx97omCA+r5PzCpT55nHWoi+aeWHY+Vq5z1jSXqWHBaNgeks1s9
WRpX2vBUN172G8IKrUGXDBLkuE/gM8uHJV25tB31qbENwJBOGtPHf/Lhe3o4CmIc
EeCmuMhXfJYaJ8vG7fvDJSMBy7v+gGp00LL8AyjtTwmOyE4TB1KEy7dKy5kAuyfH
HLo5wggmPV3ETZju9cksfhzhaWrk3KYjnc2ykWVuOUE53EXHO7Ml2e9hT94Q/TSV
zJSdU7hTVPCrTkOelS4V8tCFAyPomVjqWPp12QbiuO5iDD7dnk925vg616z1Stzt
ams5cNFbdAWjyumPC7G2PH2Bhbx3Vn9eGGK0pRBGQB3EMRHttTukS9FX6w5EaIWs
KtcEZPLLOkEbWiqfy70GmqIZ9FYhE4BY0RgRNN994E7V1Lf71zR76cekw+NlF4uc
dRRmcbHUzN55KNf3oi6m/gmOcwN3a5zLKEwCCzG5u/LqU5U0GCfBjllFV3ecFczg
ZPL3n8OTrDIvHZdzeNctiVH2baRPvOFXhA5MSwojRJ0yJClrUIcFihh1vNwDn93r
AcOzWQnji0BBD0wz9n8rNrELgyaIFMJz2BQdDpHzUqmlfF2DGEPRFJ+PPinTKPTS
gzkHIzgIPbIPOcH5fm7QGrwOXBjYH+Wh1KDsF73mHs/1s3Fcz2zXBFmgcspQ4qO4
1MVtz9fyGI8fBlEs3sXk+wj1lYuqvjeAywecI5Zo/ua6NwANpSCg3wGrGOk6iawB
80wSrCTGshYGGQoWmSShLehW1+Qm0SsU2JxNmEYKzu63SJlRQ/xtDWiSiRxhE/+/
bk9Y9uTVPUm8lgnYvkxbmW6Gwn8N8muoH6Zv88koVd0u9ZDuBVqBhw6Fa2caJFdL
FMSY1MfDJdEoqe/p/OD5agnzEzaLgwZwlDnIO+0z3Lklg+v80414BWAuBY8eHKkS
p/ulz6wWvXoGasik7A15puNXJi0HuAiCnJkhF9i4O44NjIucDtfAO0onMLGw+toY
ljf/Ziuq0ky9jIdZvsB0WgsL5SZtcUIFfBHwVlSAyYqwugpi5BoJzVcIQX9qgyDZ
8Pw7ZR8fK/oHHLMp5p52oriYBFoVkghBxVran3/eV1iBFH7KvpRAl/IsUVVUeVYw
XZmmJNV4oB9f7GUmHSj1oW4LSMTur1SnovhFI1KKX1Ar9EtSlcnxmMiMGF1cd2nj
i7xEZHIFEkdjYRWztkmSdpF2gAnFOn8phzKnLy8NC5olRGFll9PpdWLsKU4vM1VM
/iPzcW+fdrRrk9AQ3CzFK0CYuMTnI7iILtwUwanhiFF/+aUur0gdFnkYMAAglROV
u1RbxZNfubnbWwPbEz3cxYdah2+nfDWpV2RTk80XM8veEDeNocGkM4V6rg8g68wQ
kW55qg6B1XAmONQPRcUI7xvLt60OUuuYTleFiFdUCypOvCa2HYAXdJoElIE2GGiA
sQ2tuGBrzEyaPxv8HZVpJGZYwO2UKZpE5piEuOwD3cBpFEGoBmKCqyMOlU4yKJ/l
pZuq5SuWsUjxM45mwRSlVjWXMxChtHR4M/wXJriKnJBkM1mhkIbRnIGF4kPtagdp
76JDqDMkmKFUnHvBPbY4lm2LaO+Kzny0xviFpFlH9RTnSedZpYhrc6+FC4nr+PWT
RDQcvscXjcNheqbfSdSxee7FrWKoIzV6nPWetu9VfSPZ5DHnqLAU1+2HYU5w1VLH
dRvTjTLBfHCPio1s80HXgP88Ul/91B72UJ09ib31ahmaocJ3i//sQi7+Q09GrKnH
5r7JntjQYyTCW90GCU0kHX/SRMrVEocJQhLG46gK03N2xAvt1gRB/TCrwXR686PF
RCkSI8hFl+K3SyA2NZapkSwedE5uBdyZC3mT20uFPVXpCValb91q4mW569GQ/7Ch
YtUSQ6tA6PNxL4vd3llVs4yWQOy8Ny4OmpzyAZTsgxR6jRgecsorm+ruAnOZecLC
+sJtrQHtDNvdSsz1UBOzaZe4O8UjD/RpSlWnoafKy0s23eJjNuHqhMySJnJus3V4
Oba29gMWAq3odKzmY2i0PgYGJRxB28v+PvBPMSX3NpnR6KcnFmR4Edhwp9c4S3el
WeIiheBvl5rjvq4kjSm40SqkxHCYImjBsePqqD3bvBUsUZxdizyO4sp0ArPW3LGI
J1wQYSNFCm0PDAiDgBtZu81MWG80Qtg58u3Y1T4M/HvTmjyJjWVOgSGSWk7spjYR
NhAQJaOn2mxcmOw/KrnfQdTe5TfABC3DaW4yDHulSzns9AgKzEC8CcGd4S85wm6V
YAd5ShJ9OJSKenyLVNcQAONfIz3Y6eUpKabvsyukiHi0T+rDqsqFmg+8K0xU3QBU
uBU+rNfj9wSz0V+FTvD53sHvfVrxJyUKhGrVrRSYI7A/eO629jlADDz0Mi7S4wxK
XNWL1Bs+WPF+iZC9YEUm4lV4LGsjQ3syN42EWFuVZaJSvnFUtuzSuzN5JJq2kSy9
YEQ3AUcxqcWI9yxDdxccBoJkMM7zeNXPTlTaFBhTnGblFIlYmpeQv2M+q7tISmng
2pEIxmC2dZqpdUHXmA4FUL2PKhGCc/IB20QLj/p0alSbzUZkdKvWDvPM8rSzRFqy
iFFeEYiHt5seN3kopt9XPEyqbP4ZSK9wa/nsWmTwOukbGkAeXJD7U+yVLybO5MVe
i3RpEU7IJreFWEfBOBkwBiD3rsp9/nLAEBVAm+TbreFUPMa8rrzR36i+qa8yuzLv
wdGwg952m/ylylE54L5zEql0lWl7DJmuw9/0kcyKo2sn1U4D42YFtZUy/HyxJPfD
eD2jLXVNUsJLwJghjSjfsG/uuPePEpYn0/I4kK3SzbCZgtLr4Pgj8i+YoAZNhrhj
1hPlNYCpFjGc+XBcoLi7q/H8wPS/gcR+X+tljXyoJIWE7LA19BMAmKBpq+Ji+pcB
u5aX8nDcS3glLVrSjlqqVvqMjAY+J/zdaeQtETlc15fYK3o1nkfb1j2Q0NKWzVtN
lzenDvdjd8p7Nx0u4oomqrXkba2W6EeNdYP6vEbLtalKON44ueHV1+ZyEdnuuPgr
DrgkvN9JLx4akP1nZLu/Hx1TAA3StRgEmzYHced19r5Z80u3SzhbC9SE5ThJCuv4
9lCo1GgVwOqNzu+Lj+jlDlM7aQ5b8+nyvtXKyWb8PhekaG7MK7vZ6rs+ipb00Skr
EwqgpVeht9G5Pms6QQhJJ0fs9sBeRApeMKw5OVqDlKC39c/YR29lm+9LAXeMGLBn
+jPGH4hixVbPl23kXQcoq60g+1rWwh1SolJR1QUNHiD5+eYXanIZbg6KW6C5x49L
SnwV8WZYSPko52f9/8NjWyLOYJaYApzd5N6NLcCc6rJXFVqnZN75Y2XQwWcnCx+B
+n7bHcJJRZsslIVyjPvtiYjM8osbnH4+oVAbQq/j6zBj1mbaIcOZzWBJpWB+7Tho
a6anvOlrSHgJ7jPeaiXBKtSbTPEjHe1hO1Tko1kIxdA0w55eoIbrzsS6qdPvpjjn
WUIFwnS/usn8bDKQOErx+bQ4qIJBHwC3ev8oRB+2jOdkCu1cnWGkBooK+69CF+Wd
WEZl4LA+uG1AdqYpbw7uwB4hgwHDjhuz2kHLHZuTljT8kTy3Lu2WY3Tah5jrfxai
3vvyH38sjjRdBRe7tBWXu/ZZv5Q2k6cNgFOGyaEZoYbkZjEYcgUyuTKQVaKQgXn2
JX9zW/04+cZ1de79U9YJvIo7/qme329fCqcO96C+xECgdA9JmPIi5vZ8rv8YFJwN
VhB/KAESaImmrP5gW2EWwz6O8AaxNeKj1ZX7IVFmTpAbymO52c7lhCidVtNkbNZ0
aeq7mwCNYvdkpXz82LcR+s0FhgTNfwhLHMIvV4h3GQ6/tBayMc5O4RL1Rz7ArriS
/7uWsu1Ftk6r2MlAwMxVjbkHuiSs2+urW0qZOVthhPzTZ2lLtxhI2f5SbVCEnkGN
DVmK/8q5JSEe3JM3JzsT8H9FaHal9Q92vMuQfZWIxeZWMpZCLF9GdE/54620oq/m
CXESaP/Ikz/XM9IDTdASG9ZRwIiYrZuF20gZGnXFwUoRl9/4og8kvaWuXSnegJB2
IHOhn+Gbh0Js4xCEjM/PJThEob0nOKuBpzhJkVK8pivH5HBd9AfeYhajzCZNAU+N
N4Hmcc9L3/sizp/Zr9Efem9TOZrOUpRLZaTVZFFYQwikBjf8eufvF4lBISr5FWLF
oWyIid/tryI/0K05W/VuOPyXWPoLNuwO+kL4z5yBGMt2ia1W76nMN+iHqOxKtTgB
59oFqKdnqnWT8Qh5G6+kjcsrdZP2mOyNsGiZ4iyTDZD7AY/zkEnCYaBqDsEG1O27
oZJOy1EHB8D0hL6OCBu4KEL03catzXSjB6zZ5aMFQo+xhtCrPXz/h2YRM3Rg91nu
YsA140nUqXmwTO2/ikArQwgzA08j3fWmaqTovB3wxs3Rt0Xm4bwcLFrsrFwYdkGO
cq0ltKHGHhx8cABtVg5cQiuOhJUueNMJEbxmRAo/b+5NUKfR3fkn4QXSVtfnhamU
ohxy/XtuGqZcv2BF108YRO3d6pnbxAghdgxJBy3yhE73oj1xFTfiqFPgzj4eKKv8
gzKVzfZA+0quAz4LdPjXKj3f2HG1U5ey17qPw0thOmV3Ah4qyKZNzxWzKY2hvmnx
i3oCE44+WIuw9qjXvS1vzaQFdgZes8IpXYZdPvPgBS1mVOc27sUhiKMdGpksm6Et
Yf6DNPMR21PELLb9XNXCeEjIyqDviqsaDr6/V0enTnNAKNSZgvNb32R4OjKIO/pu
eKoFPvWwMKGrSOyaeVNnKw7fTnSP/6g+Hwh5qZQgune00kSFLrqe167Koz2/0UDT
uqi4Yx3y0BXx+wxRB1k0QPej/MXKjDo08epV3CHQBnCEm3LqRRJ1Pj43aqhs/SwC
B/aIKJwS4TIt0401afvqd5CLE1lZ+qj90MtA/mFcag5l9S65onSVJfLyTmWayrDO
xC1zdQfR3VCDFr2sMhNRHX5tfddZgK6b1xP/mkUPtXMzmrPKrJJC7SRaf4vWhD3p
UN5Vc8XWkuyHkQ1v53rYyqVarVzjkBioMtrkUScXi30RLXJ5s34J5Dyg+/imJypg
vfsqOk6qN8hhrcnOsB1KO5DILYK5bBGecusBu5gksZunQr4am/ZeZ+wW9+xYYzfp
llqnGBbfSE8J7oCqrnseEIfJlQgclJOmqRJYN/RwL9PVWCFHADbqnHHM8qKv0mHj
ASw0FFiDx2JaAefQTEymDUwl/xhP116QKNsuUMDeazQ5fnc4BkZ3MRO2GhAyUSyP
yVSbpl/rvRbr83wwxrVPZYy9qZM90JcVrut7/0u2rpdgEzAHoPRakwEVjymagDeE
UvR8VU8rzmKDrz/LaR9Xeb2b/KQw1gLzaamdUGg91kMm1lqnhKDqXxJityvB/Dco
D6HIm3F+hAxsw7GX8pihL1CFGmpHyR5jqQ71Lt+Cz/vYRb0Pi2DCKl2V1rA0mAAp
Kc4/BLfuih1kd361SoswhWBGQPRgxLziJoO41nDvnpdneGER7m3sp8weEExjuT10
FlfRNfWkurkkLTU1cFBJo2X/1zwVu5jM6QetnSxNpVoDP/kaX8sFle/eZrz/zZZ2
wpZM9FYxdgdTFZ/NtpSjmmFJMjHuygkmcJtIy+fDZHpvwuD9d6G3gdQwecUiW521
hn7tfp1lp0Sk6WYozWTyRoTDmm7ZgjpaPwfR6xrJDunITBC+ThgooqI3Q6o18W6d
dtkoCL8W2qypDXQnp8B11BcPxcLuqYZd0xEmPZi2WtM4Ku51J1KEWXzmUKiyPxLS
qQjf2tJXnEquPfqqL+kes7kS+QOTA3v9xm1if6UHhEXI1KIk2+Yj2PEwlsDIWqm/
UH/zZFaZ5VxIUUbUPRusr6ykpYYOxe2D5btbBt8XZLpzcLMgihaOZ71NNWw5BRXx
09SnTcZoSa2RHUQ3xTZH0f5r4wBrcTgvfw0wsGt6K4aZ73A5MrN8Aj+RdLBaChmk
+U0+r8iYbCDdIs+jcB5/QyOhuJzv20YAGAIAN3PZ5+3mofqcw2uiVRr3MoGIpQxL
UUSpM6PoElbzujyKMtyIg45SoHkhAWGqViy4JpmEvz0rjj5Or9HxYeyHcVam1UiF
V5UZD99eGs6y2U5klpbhJ7uINAKzcyb/fnuLd+tDFkMGcIwE+Q9qk63gnMAgR5Sq
kXS0FUlVyTCYw1H7/aMPPpYnhY9pEOfFLHO5D3+XX6+wARafQlsgQq0N0Q57KcIH
VpazsF7XEtizOSaXOEz7gaTuK1K4y1r5IgmWw3l7Ivw4EHzhVGF3Fp5Zkm0NTRgh
YWzVPPNim1tGZOEw8TGA8O7kRHgGiqTTRdq3nV/RDVGJUAJR74CKgtgs5dWgcp2D
G/eElWBY/eRmncGwTx7dhO7Dx2J8sGqNIPZVNIPjk5YFQ7/4db5jgSyQGGszAkrB
wCbpLFlrxWZrtanIkdsDgKMqFsnHChgBy1rcJffPYcmRL2pMpSzjtgNf2WrL1HMq
7d3vXda2MU8tbTJqfhuQ67d7An3e5DhhAMHfSh9kE71gvLs8fCTwaMXQUjUKmq+t
dMHfBQ19F7TEaDIuVp+4bgKeX0GnY8eYPn8TSRbOhPhBxGS0to7LZBY0jScT4Ey0
GgcW7nzIdJAzODmGRRTpPsdP4+E55X9+n1wsm03lRbrCpVsexOlsnFw9Io2vqN8p
hhXug5I4zD6k2v0ns8opYFw6N1OCEItXaz6YWqpT1N7HJwchIUo1lUcSWKoTAx/l
DxRN2yraOgQJQn0ZBFoPRsLMMUFzSyQ340zTxnacOq6+HOTtf2+1V6E3egtGlzpO
rlur4ST7j1oPKeHYfy/kQk1FwUCr4hM2IBCp5TDrtlXcj0LYV2ya3oO4e/7G2NAN
AvG8QZMBpAjeu/gfBaXnbiIGUX6SOMtOn/xBw73bpjfJFMaWjteLO8Rwoya8qofD
RhzXQMXRbAcwgrMbQ5JdzkMRMLKxumaFBxRRaYE7MeCRSXL8N58WwZGKkw908Eli
Xgpf8BWBSMp3+Ff5ibkKmYGgvswO1BCS7iBwdNCM2Aqps9L4+LICIdw8DbyO7209
Ni5Uky/an11JtC8upQoFSSz5v6ramc6iTBaRyYFO7haGv0hUkKJO9r/wjIJYrlmm
OUmpQ8UQl73ZtHFAc40aydZ4UHHHSCVfltQxgUvt2uxWayi+y7PBjfDZ/MJnncJP
+cKWou59ckYWAcla8QHyespOJqxCjnkBQDDo+87ziVC6aPuzhuGYLrPI+8l5E4sF
STezf3kBMz+dqS/bmI+gBDPn/wnJ6OUS2Ut+lhZdMGv7CsV3PDoM/BgSGniaiByN
usoFRS59AF+jHKVbX9XGzhMBDQWaEZJuY9DL1+/ArJftt2rmAQ/rWhu7nfmaQqha
brpEdCJ9BENGbAu/7xniuwf3neAc2UWmMy9SRNgnKDeifltP5OfLx/BpQtIRFfob
YHUbPhi6MpQ6wArrRb45ZpOQg+DoCi3wKGeumDavj2A2OiQeyCAEW7WH2yojZooJ
mPEzc6FDKh8nMhAyxo6ld3CCI/5Jwkso0C50kG9U2QbWSBOGc+RsdF/aO/dHy92A
PTxogr4frwFY/27FqUmXS/lJFmULTx4w5rSvvKKLTILJUN99Ixv++djq08UJYNqh
GWa4kZnRP1gj63XruIOY31jB6bKuVMoRNJ2YcqrcEPnYlqXcNg+Pg+0o0OO1Kk7k
Esae7fGWyBrDeFrJHs87ijbi3mmEsdbdEbWuXB47WYXGBTPE/zK4p5dHLlMRKVsw
6xOKsgWlkrcDZ0wFlY0oF5Ezy+6/CXmOKEhaQk0htwuxGyGKPMaRjtfDof2BM8d3
ihYkLhIozxEvee87+CsWvSsZAkuu33f5M8xxmm78LaBjc7OBqBPjAGnZoeEB2zUK
EXQAxO6nKBTE6vbdnoIumfIlNJL0nsYvK24xwMllZm4wDxFoiNIgEMyN77YUxHnY
ZbBXtQv70nY4QNnxVtDr6QAN5XibqDRYC1V0fPz/PBhshf7Qdpb+M50r5JP6QQ9Q
TqKmiQZQrnvgrr6oat4YKvJ6ZyOJyNOmkS0niqupUQsswwjdSNcnlLa8GTFsSJsa
50YmQulnRptflEC8IQZFHRCSLybR3q4ppeEdirKBlcxx5MEWmtO9DFE+KpiZHLLY
0bQm1HzwXJ4Z4d4I/R9mqT9FCkxVDdY1j2+T1NTycOjAgSFKAEHGJPboeZFwNKkQ
f380kJ3B6Ur0k22jI6Js/MD5C5E/nAd2YkMTlq0TZ9x8vBJMpd6sH+YiM/kA3Tlj
wD7r7/2SJFrgyU30SuSIi6BOubRXf9QCu0RIFSUGIBfBAs3ZsZnqla/C9kWEVCli
Dc1TFpw/v/UEzGd4MN7nwMlfChg5UcuCqt4iSkMxDHLcXTGaERCJA4JBhbqd5Ern
CSJE2+987A8fcf2rA33Rgx3qkGEzv9auUpKnrBBwUIDcEOzEYXKHskk0l5xlJYyJ
lXnIyYuUOuu/igB8oSqpFq71GwtBsKm8Olq6qnERExBibxsg/rtmwGO4duOFoxW4
SurzEsSYzF7sbmpeB8WVs62pylPIgDDyLq+ecP+Kwsjq+fc5x1Gwo3cAvZXou3JP
bBzJifsMNG64Fxpw/LZ/wa1Q2GD1Db4Tm7w0y8SjSxaAGElayI1JVj1+d/C01FYO
hWzMZzB0ZtWel78iYPJGyhE7iKOYZBdI6y1O5GJWcRp4+qK5Z7dbKsamp6U4PPY2
eFj3QZPY1UPOfW0n4fJh2PCau87MB3kXBTSkaFyf1ml5wonmeRZXLUC0HfvVM11I
5rPZ42gvxVuK0O/BUdDdbkYORZ3iLbaNm7Gv1AHnfmOeZs70CTbUI9amKgWdGepw
GV3n+WMEGyxa0Vz5KXBLaeDkcXGjq00u/0Uq2Cgy3zr3YzVlJk7Vv/qzoVlxB8+1
rHIQCYSuVvjGNSh/Fdx30KcXsjmJgJWcRa+3hgGWwmsQbt4dffhkZ2xsRTfJaUnF
fd3hiPjFEzq28aGyjU+XmTgGYkPZgYpdaVMd982tLcSod5d60df2lj2aYBeyuDJx
1hSDQ/dvy457Zk5XM8xoXyScUpveNUEF4fPyGwonC8ocRxY6X4LWK++ypFnzQ3S1
BGpV5qUG9FHIRnsYnp3bAZYHUXhUUwL0YiaVX5MF4Kpp78CmDGdG28WQoHgrz41a
KFAY+DjAjhF46xr8c69eYQm+eZCUkaJJWkY63yBHY1xD7av6Lw3I/YtEEqLnVleQ
lhzy/kqXwrlA/RlF69NXfM1cqI9riZUeVp8ShAReJPfEauPY8yJnD2d9m5ijyOFo
Bx9daogmPex4oku1599vV5yqd1qR9sS9MinZ+ZTcrk8Xa928AJOAMtrA1dkqZ0+t
XpvQ4ShB2e8PWMTK5OOXRW7A57nwM66GqUaUS8TWU34+oAkgX7czpv6xdsMxzZqX
54+hBsglPxRhQLodCuoTgqgqh6h/E8rDgAijgMMKxwZqYZZV6Qfk6wCXX2KkQPZY
HR1+DLh81+PHSdL3ao8dtulM7eEKw9H/fUeF/286t1Xcagwj3FPVTJlFPVvGkx68
4bZP17JGuMlzLEyukNaOiuzACl9pBMegBtHFZVD0OSSW3Ry0DR16p49pX1rqbVkf
uQGwM9Dolzy2+Hz1yiUF5k0k42YpIl96PP99rXMy3/6yxyxiT4oeOJQ2PXog2gJW
d3F8ja2YkYOYTvgjXgKgy729holRcQB6ax5mlr+SmghAoTPHmux3ny5PmNe7k0HN
ZtjUNk9iC1yJdsj57fEkVjWKcFpDOHKQd98ummcHOS8GaUKROh4vAseH2VweHn9e
xVwlsqlNVa5Be7pwiIZ1eltyxLeEtXb+ZHyZQiYHj1iinfxWHQvdnv1PKshoHMgX
jEwryqMVq7dT0+ypW9b9Ac7eg+b0nj47jmHjw9sqpEZ8PYtCXmJS2RnRniH2lCVn
+rE4z4FSH+bbHXLsJTMr2neiIuqpxywPCEJ0gfsk7v2OQmuz/qdm4ktPfYaUreud
UfI347os+Yf2c1xo8Xg6EBvC72RxUg7s90wv2j3qw1dXuqQ1YifYQswp8Td2F8ge
x1zkaboQ2oZuRplybALfqnl25TywWD3qmy4ZC0a69qDDha95U6/IPOnnn+yt3nmW
kiJA2m/riW/lRRySATAt21Gz3XYSfOj4xd13JwNuFRkH1orlgeCe7RE+f9KMCxat
TXxN5xqlFTBV6c2rhAPSHroEVzOgQ3zeIzBO6R1YbePj1KCRE2Bh6WLla1YpT8d3
BqMmcW8tMOYD6BWBaHZz7QexTcqh4rVq56Rt+dcGuxQWFel5sL8UlUJvyRE5CLeJ
a5NTqC53Mr+m8P6aVgrLl6z1t+E+PCY5T6fEm7z03y9n/e+ckyBITd39Uu7G7DdT
oQBw2MqHrvGBN93YYYk0Suv930OEFCJJ2wVdBMRQQh1v3/nRnFyGCCxPiZQS8/zD
iGYi/m7ceFKpPHCB2LThO9qkxviUUz9Tk0+GaRujOckSZeOX3wz34/CciqD7JsNg
sCC9ATb6m6bAzgAVnadOYHUwfsK4z/C7nFGsPyEudWOSAll3G9EHuRBnwCkNKOcS
qGavyYFGwvXFI0m/t3fC86TR+InorkoOWBQZ/9wstcdUuuVDNeobtTsGtueSthk8
Bgzl3QhVpOBcpK56KFBolgRqUhHLbrpp/CSmqKwIKRi/wfLPclCqhUTwj3DUn0v/
vD1GgELthcdNSUzQ7h41lNpdRll8jpn5R/qXLdZSsSGz6r3eSo0Fg777fxVeftiN
kO0ahPg99D3uh+gf5+cslV6KyQjmhluznFj8RZMabqMlIr4MSEhgBIxeVrMKyiv8
rdcWLrdk7qWugbnk4Ob7KbgKlTOogSP8/zkT3dPlnrDP5ohCmgS2h8sfqKdjCdCB
pYxFcGwXzDy4KmuKvA3Ed7rdFFw+ldVSAqtOO9k9Mpul9Em11sLZkdRlygFpk0v5
FVKGKsjKqAtXY9iWoWHGw4W4RgNj6GXQ8iMzzU3FabGodgQwxotgQDIXdBjCRQ79
yFuiQ05aMBA54jdoh6yOduAeixMSGfWez0avTjfZxhEVPn8I5IVXU82WcRo45SPa
cSD91M0R3q6pd+GXlTfty0NZHYNQD79J0iP0NU9l66aIJIhOCqTMdi5G3kxXx4Gx
Z/7vxNM7rLuWP3r8V9NXyzV75oNGiEVbAEEAS1SAXwzXfjzDmswgSKiaeFVYRGaN
XsFKsZUlDYmcHxetjNKBPIwUcl+S4XdT3ErmoUbwblee+gk434iEfe4cLrzVvhVM
vfpfy5kiEeeR5Pq+thds4rlSFNsCszj5OrAs/w/lp2Qps6fnJanpAdzmAt5LAL8A
Rt9hTgnRyMebqaOJCnNyb+D0M63yFio46EEL5lTsPUexzGDXEwJi4HxJ/Z3oBk1B
MGFkFSX9AF8nNGutdszftVj3WVNKQb74MdVb59xANoLlKjKs2BgyQ33MyPM7pzaZ
+MD0vKfujNq1RPfkfGPypBjwnZS+qksGbDjkfDOHJqDFvQmNuMtDXNgmblU6tmMN
kRn1YKegaUd68V18UU+L5pQBymlIIOfyEVupc2AEiO967xyQ8dcxhVpDgyTLSo39
SOKguNbE4q8eE0s3RIAFEON6q+59c9rltFlMyH6l1vYmQMuXTkUDuI6SwfNRUcbj
kKal2XQoNzp3GFdbvbdP4TCqh+3J1nc9QJoCORTKV/cPXcHzukC56fymLieT778d
qBBlFJv8swJLC5Ouv9jZzpaLaQZaSzmYHxsHlmnJNEOdiHHyYDPk6YO7MzPcZMVl
gdOsULlzukIGYTXaJNFqfUkhoTTVgVHlPEJV1bwCvBnjT6mu9WND0Gu1OA9YgaJe
CXK1tcWXN7mbKzWcIAD0Oabw56cnm8YkXEoydI2JpKBhX3oCGRyoS5uk3VCeqnBK
LyxRyY6nqYY2y21I+TIgm+FFTuGqIobicKApk3CLN1rbPV2EyiuXnvvk4pQvwBsz
86m5WPpT0R2M58w14c4uwNXZUTtGPJF9NwKQ2gVqLnKnh6Cza2qf1VdELURqCkEt
xnvMezJT3PY4LswT0H1P+tvk4MvDT8Z7NnBcUtqphYOZwlsJTw4/QrPGrPo3FaY6
AKUMEeIXtz3mhZpV3wyuUNY8oyCMvnSb5KGSQDvu040Z2CqTyO8HQQWrDCRF+EQU
6FQOEoKgz9ihNJYVG3SiBZwd6NpfUpvj5O01fOXIRrs9uZRZ6f6WV+60i/1O8kZh
gkSaSNMSe66Z/i1etyNSr5l921b55okUHNXGbgNsjhhq+ao9JSYws54IWsN7txNA
9ZgP+qcmOMXpG8zFQ156t+r1rVZ+v2mTh5+gl1AHOm1OJ9EpG7N2ghoKd0Aqi4lD
KVOGtpQCDgYDNufElpEYhkG4EwQQog8+tD99tyh+rEvxsp/PMTK3G6M2Btz7/p2s
579M3hV5Cq7pXGWiuBlQpG7aqbl7vQrwPz6G/gbHnKQ/L6Wm3leQOv/VAYrQxI7w
cEOejDuXabrfZtp8YZKoI//Duwf7m6swBJ20di2z3wXf9c2yndC20th9+mHbuS5A
AtASdkBRI/8b5QGQAYj4l/4xKmw+BggOlYPk9f/skZtw1oCbbVBsrSctBhJeBSCt
wH1WiWmNZ6yj4XOLzRt1gWeYKnbGy5LpvKm3kDjWv0z20MPD+WvPrn+L7kGmAXoo
FtZ5iM2Cvj8WywwN/Q6eL9L4+5e0Y4IFPjX4WBwa7LrP4WAITzy7MdH6qO2bs//t
4fl7HHXCcVsXMzZlD0KV1+xnGWPoqXB6ymELLyO/8xJWQ+rLIQqzbTwQ55GEi+5m
d2qTLY7HMinATvs1gGPHNc6LP3LjwDcuvaZLzUkrooKa5ClPLI8Pwtnn5U9CcXao
+TUPxAdIHfrKVWwbuQtG9K4mu43HXBuvoki7Y2tFBcqYiG9mk3LbmiU9T94lSpRl
i809USSRxrK7EM5EP09qmWBU0mRZCmeqkvt3iUWtvRePzRAgHjWFfw1Qj4+gAgKK
uYXhhQmEhi6JPwYmxs3SFVxJCHbxnL1wUqMeuDirreriACngpXGuOx0etpkFD6Dz
7++UDYPCeVRIQeLQ2XoImiGi1ilD/9wF0KLgpxH2RaYE8uJEKSAqoCsmhf0BZo2K
8EM8Ke3PhasSlZ4Cm93wxQC2wUOafeUc7vr5aCmCYvdZhBzCmdL0JQLuLVcw53sO
Inl8jdfkCmP3f+ShhuzWydpO/EOW6WNaVyt+HUk3HUSuJbWMmtnDT9pjWEHgFdEv
pXSz2WA0Lp4ikYw9kRjivpZGnvGCjCBku6BcZFEDBd22OSIbfUNxqhwEiQgVdj7a
wpTKjZRrWZoDXSU2BIOLTNkcQZ3QEt/aYyRoR+1W48fWWhlRIQEkct7W5yUCZaho
U+67XrRyHeVM60P+WXJqZlyiG4rMHjnakSRk4ciwnWt5bwtNiEn7oizGBiqORtx5
dmO2w01eGAowr9Aji9fa7XmMTLPtH/l1aEgu1ZUt9qbUNh6iQ+JOuHzj2eOBuGf2
TocgZ520zYy+PbcyIMykVLdyJI/RIFyX38IvgAUpG04brQjntEYcNyupVECPJhdh
m3C8hO4gkkqkIb1bGDVERqutyQ/EAEEjK0f45EEu1KfJwtoGKFUl5nDuap7EHYiV
RYonQsMs3NpnKQIuo/d7Ezn5pjnKTOUPia74BI2ILTcUpOJvLwpZkRpj6xzIIsj1
4+o9djvZ5QbA3lr149TO6eWxfMLAanM/TVIlD6ePW5xevS0KTwUqMfQd/QcFASCj
J7tpZ8RtRE5oS/g7A1KLkuZLA/AKS3lyMkv9Vwj8MrmZcwvZnZbedpj79w53ee4m
KPbDrRFXObR05DlGVkDg862Tcuf7OedfeWy3dFPfc/Ca+pmwo7/k7maSVo7kQP/z
/EhRcMNpUndCXG0wh6gVREWWzc6If1MQp4V09JSd5iQtZHKPKTP1Fs65acScUSTu
KlrkQ1IZ65e6JAByjRl+Y3zH09vBcOFtznr8bKFIJ9qkb0I14vPlBeuQUmUR/6nB
2O26urDdYwfowvh2uT5B0NMBvjaM2yR+V0ThfH4eGG8vZj8zHfvhmS2uKS4f7tF+
wLCytcB1ilws9TXzC4vkB59quXasyObRTTFK0eSyBY0hRh91lgeVkVJD43PVqvdP
turs6WkMCQV48Whe5BJmB3KmVKzlSsOyJn2hG1f9gjNGJ/nmwmG8KSYDsdfYbL/X
4MS/Ht1YOHeLxivizkcvdgDU7tFj0Vv9bNaojBLgBQRxd/QPCKqiDIHvk940BQrG
9QuHVFSo0BO5bw3wF5C9Mo87htUtQj3mSfyjvkWs8tMBVxj2tmTrbt8NlZ6XCmMs
PAiHq1How/T+y1TpwjtpXYn/jPtBKKo3c8fhnqpLeLnZJ8yiGsa3KZvW8y27IlYz
V+e8HF6jaFf8JnJNwPcXer6ITNVDQGf5KidUQ5dNsZNvMkWjmskbIvRhCItow/TN
5biVWicx+mVvEKLy3VTrR+Xnz7+MoDfqpIZv1WJkYJCrKpL6OsHpMzTIRaBAO8yk
c2IGThShqlVjIW2IUfphcp11tyxoj7/0WbjET+xjUrFcYjPNl5Yl+49Xd2jgY2NR
4yjwD+zA5gSi5XRM7XJudLUZlWvuLeiWRe7VYqaNZfD9iVt4d11U9squP4quF+If
5npd1SnyQam8pl6RED3QiiMaxa0n7z01E7Tg7/82twEg5XGXpxENrZruh1Hf7AvK
nxhnsZOfjOMrex3gATLgZRP28KeNRF7bqXwxt+BlGX/Nc4vLiDHWbpKc390JCLSJ
61ZZepJrb0aMTGTUI6ATWboFofq7Qi46U2XlvGcd7V37K1QY+ltPHeZ+TDMUUH5H
PSO3lVTi+9deEECkM33Y0rAnxPbKA7a797U32N3lWq7mA54tdgUBAA46e3dObYcF
N1K4ZOhKIiVnRvmXKyJ9Hktso73eQsVVNdMcAJJ8rdYs6IfexzNYmwds2B1VL0pv
3rDjrFcE3hAGtvY7PvS01Bv+vAUCpmvsYh5Fnlm6AzwTyzaKtWwy4i7J/etZxSFd
8XYovIfF24VnL0LrcOeAY6jyyw1D6O36SqSzM0PL93VfNUqflT68X0GkmAjh/cx9
6mbmd/BPj34zCzGXqB4fc+MOiwwUT2/EjQWpAscxNmxxj52e4Eb1jacDzDYSQSuO
kKM4xJKzVxtjx6Jv5V2IuhTm3c+8wHEwTCsO0ciguE8ORhkWyj0J5vRa4flvgRr6
585vP3jaeB0KOw6hws3KHl8k7MtKYjjwns43VyFUkfKc16ptBodovpqOqQyyf4S4
w3qLPEdA/vwCsR/hk6aoR1iPKqB8+XoIzXtnqgBDvYn4llYcprd1hR1T08e2qDJK
Rr8wQ1re87HZF6BOCKoQHKjsc4oLIUHCk3d2BTiBtTCzEfzSh2goIEXSEXPORjrD
cXlo+2UvAG6LjfL27QCpo6yJIhi2jTdk8J4VS1m3+diUpJqNsjvhf/sYzYgVbgK1
5+bIzQ9zsHSiA+EQomkpz0n9hF9E9rQSVMtSn1P+ea3AVXNw4oiQu2eZ3RNo5OzD
p57uInJbI8KGfpO1Qn/PrzuLCixs8EYQiYaXV7x0guJiOcspAfeyh7TjRknKe4lM
nKYNJSdjMKK7lw38RnmXDDvMBmk6o0Pd8gWgMT8BFGA7QDQwqulH/3Dx+7YYaUJE
eTn3bxSlD5YX6YR4qXLr0IC+kzmwdbaSDtJvQr3FOrHUuGvUO+hOQipdTqhlaKya
qntjYaUlhlvB2CsQaIB+1bclXuBZQBWjgFMzFxhnDYLrr79HjxljYCVefE5e5zLC
IpLIjWZmoWptq6zELcfxB+BKJ+uR/bjrjRzxQil/VhMr4lh+NbencGCV1Ivnutu4
4jkcbxupEKb3LkJXztflcjOYmpqRksuWOtzdPDce4u6oSf1tqlw1CUP8ukA7WOPv
jfC7+BjbXhglSfXNH2QSJzztalcjY3eVHvIByhzp/yAlItMz6tXK8nClyiAfCv3D
CkD8ChjG7xdXsuEyhLzHBotSTTSxdUvp9jfiVz5QU11dVMWuxqG6rxsULhdLwgbg
sTqIIlMm+dZpI+pVMxXO0V23ri6rVeAONSBn/hc0xLeqL+WVlwJxJIaoojPQiKWM
lkYBEfOfd0bQagdUQ2UT0zQE698HRQUC6sKC4JfNPJvJN4qtluv4BThRAbVqVtsy
9nkphFPXMB9IMcHCqn8WASkkl903Mb5L4vTvZPgtXkdyQDTUnCeabSpehgURWVlu
uyxGftRJex8ONeCYep1NTbtM5TXH1jn521taFxcWGhMo90dS+s2b2lP8lPplvexb
snrjJEO8E51dyZtTqcs8b7xIxwc6okwWIbN/Sn1qZu7BOx4+Vb6Xy3Ty0kcVEai9
dyg2RabPAlDghUymFYF/3gZgwZP0+zpcYlkvtQCOlfclHhknpz7yEb7XdLrXSyx+
uq7EqX45K3BWp/S2aDFzjhLm6M1A5N+i4rXFqaQyR0IYpx5FQEc1DSgqibJuSKyF
y75mXCAiDM6lTDO+qPY8y5KvAw/Qr28LJYDet51GyPNOix2IgClU7lHIxz0gjdfl
26tQk6xdjwEAnZOKPmBn3SB5gvpaHo/BPbqy/bo+rT4RRztlmplWRj2Cv1yNH5kf
+eq/M3Ruc8nsxqWb8TI76SQt385bGR/Vfee/IN/zc89qdtZIwKodezE0pRr8lIrK
BiZW8gKlFOl7ESujHc/PX6ALxwCphbysRE3YGGDLxwnB4pmfB27YeFlALoo4Bf/v
qUkko5sko8GB/lHgkw0y4FoPJbcG8MCO16QZNP62pGXFQWvWNvawhIXaJmcnzPY5
KkN84m2fzA13riNUHsbsH8A2CS9YkFHBrBMjpg8+k4VMCBqOENjdEU/foNC+ydjI
3UcnxR12T6fx7Nx3B/PV/Of+5FTJ4EalWABLtrICC+kV9uCJV81p+ybR6Ocpi4m3
nlG1i40A5PHioDQUFpnmXKFCTHft1pMtENxJ1avX1jDTsRNvn8Te3aN1CTTKwn9u
Kc+yE821bJVeeCn9CKI0p8Pj9jj+BYfe3ZSQF2YRLD0elO2WQF8nM36upvonmIhC
AMUlYFqZNVWSSYHcXthFXXMAgTFfF+Hy6Rx4EKY71v4lD2k363VpbiLMWBZuVipR
UYAEW5hhUZXYSDhPsqGIc0T1eP3Ry395XtwblXUUzF3wzA23BgF05kYQ/qAZuAAT
JN4tCoD8UJuhxwLcBEKoxfbBG/Y8v4DBgHrLcC7+1Z05z2wkxFNRjjp+/UPNlTrI
3744Dbokjvq81UCp/CrDEObb+U0SuTslsvrpKzd7pDUbaz7LmZ0I7jc5lyOVxs83
xcbfFfF6IQbtYRRyzdPB+nGV4HXsq2n6LIy7/zEFqN+w4OjAQfyDz4cQE0r/gNag
HL11NJooMlfuBLxQB9oXAL4V3ZXLDlmmhkPjbxT2mqbgeWoLTZSY/ZYAFhSdz2pX
aBXRuWhIhyAV2s42IyuOHZw125pB5rdTyF+MsjjlujM2lglQM8bb/wMIHxanxkBH
osClmMMCBJMP7efpF0qORskdMb2ATYTG05zhqV8jvHuZDEwhAIw3kV5ZWiUQvpOI
BQ+aSTTT4lOj1HZ17lebcZDWq6hXERKIu4X0RkfnwHJ21G8ZJ99oh6Z0ZiieDx4w
GcPsMvSbt2lsFHM1yUUi+SxfqWrekwzuLGJNs1YqosBtCrh1fNDrEpVOQnsSmSqv
xHdW/Ep1RK1piUzDq9hcpJjGXiYzKM09OwRW8hdPF/LWAbCugRpJvhAoRqWwT9FU
fJxrUbfYSWdJiyczjQ5T5D4O1PzpszXdqrEJuVyRvwAHD/vvBS7NQ9teHSem+ddt
knKfmhHk6rHpejGwmdWLN3L0v/G6iADIPR323faTbq5T8XkEKuk5ltxcbNOLMLzK
bLwyMPxmUQpZo8wsr5tqmjrhyK6CeCBgKkZiQDuWUp5xcq5yj6J4FpWEmGtIbv1A
SiV2xSDsPDLE9OXiRTnvgkfxZI3jA7kLOH23m9JN2khiPydeoOxGw1nC+cNVToam
cax4QT94QTT3JeXiLCDmspl1q1wdUVFlAinbUgAxOxEiKst38X14GPaF6OG15Nd9
1VrILtbDriTHaX+uray1xsppBVQPrNBluVMPorK2DbMvpjjZXt4kNHI8Eb3GG4Lj
6kfcCUyuN1NFwQGSHiuZQINMKupIsqP1muapuSHzfOSMd5a3U/+lUOfX/uOKRpfQ
3zTqBnaxB9PifWg6E47M4xmOy2A+AIWhmMkhsajtOPDzxYMyHml1K/uaRHpQ0HlT
i5U0ofB6PSGFkkxsQxAjOGk/XwpZD+WZRrqXRHFxwBn4iZkXyuAhyhw2bysdjA9K
HjFY+fIttM523IxbYlXPW27JHo5OhTfJpTxmuEhAhUJmPNK7Dm5Og11nyplD2Kr5
TePlszht/LRPXemp8Zdzh9m+c5dbmICNxQtOeGO3ToHfu3+mirlvwnaC5AgMjUUg
icjJrEylk7zErXuGNhk17h30iJmxZ3ko5QktXmQ1tA31CZJTM0jy2BL/tFE0WaNM
TOkoTFzOJhDt78GQ93pgmUL+t6qZcw/KkvHLceER5ICtzxGwOdcTIpwkg4zkQ/OE
LauGvijcWz85rDFLlAfHgSPPni94CJqRy3i+IUf0rGsAFkgZwixcVZ46Hp43kSKR
H1dmN2jh3qSu8mmuGZpN5jYPIwEhKscA5/j0TU7eBZritIHy10n4Kqkr4FmcuaOe
n1kU/DzUfup28gVcRKDpdpH3J5/d7WpFW9XKlsL22fsORP8vfLJ+JSYesywt0Sci
w7lx4nKZkS4gNN7i0BuiAVDc6eDMReBMeVr3upGJhmYyAEXtNIGxQOT6VGU6vtZu
QTrErooc7HeTssGxXvmvkZTbFeiReGWkLfTG1QIQommh+4Rl2LQscuMeDO3niHQq
QEwLjM2Qy7lrru04qQlk6U8uV2SkgBCo7xlmlvQ1B8eG0zX0iAzoGhC7/VtmJYOQ
+ph4IR+3+EkDlJ3lz+lfgz4iaEIh6Iv0uC7x18Ie9EgrdWiXYNgneAUc0c0OEatl
ZFUbPyywwy1KuwSXZfcio0fpO2Yy7XfPCdaiB+WoVe/ClsOCJx7+n8jObCByQfpI
FlDEwDej3DyjWOE4V/3ffBMp3w7gEbN9rU4Q22A3sS6mkiJaP3Jk6g+FR1INjqiB
nQmom0mxKRT45RQ/4XiY+Clv/7G7PpThVLE3l50ysUV4hzK60yhniogljCvgzJMe
s1rl/US3Ivdpmwd28c1S4PZx4pz+I3jOqDG72hnU7ww3HPoHyFjxPslLc27mNrYj
iBGbWFkc2IfyhdmeaXTHIQUd9GT+tNtOJ5rChxI1VyMTNY3T/mJwLdnF+O/F4T1q
54lE4cVXTeGWf4xC/huOXTMZPdSWIapWTfdWBajNtNQDBBKEQT8nK/Vg1Lf3G8Am
6ocsgJSyUU8ABJikrEOnFdGbEC9U+8ih9xS7S3ch71HSmCtCv2STbmpXHgpKJfKf
noGuQJDLe5d4G4jmTTn15KTbWy+LkXLcowLGydQ0DobeCy7SJjnF1522IIDtKuSn
yhQzWy8s7m8rNss7S81q7jch8oDidppLW8TkLFf0vP2MnQfrtm2bmuE6K/eS15In
APesFf1k3UI8zEDMwOPf70pCIkRSHiqJuiLhUklp1FRo+w9LDpneHbn6Ekm0Y8lw
ays5M1GuHqxizKsmPEkV5zIUo+f5V6sreJO493fWWhxDPzknzAK6dawZsGc96J9x
hWYvgKC1weuyYKF6G45r+a/yj0VKv231+4k0NchPFyQnuOkojioUMQ4h5ZHnt+O4
ZuIC8njSM6bNLAYFoYfl/Phlbk90qQbsOAw1uhxZ6Tam9IhAdq2ZF+GVx9KHXIrB
SEJsX63sEy9hSvd2Iv03MKATV9JxBAr2YORSezwcd4xe4TLNbVG/XZXVmDd0fO+D
nkkTEbIiGGoT3ZgUkAhGggFElZUjdpX57qig7F/Abd4f+75nDRgh2fLGAR8ZotSe
Qbu2cWWhAHiODYr1TYNZR9mp/Xeu4gTYE9rE8UwaFsAQhHXwxAqrMJB4Wd87V36R
ty2b3tZvo62jkYqJbT7R76JSvS7KE1yaGk0wu/yGKGosyVYvjEeBa+Pldv1887NZ
81/tX01L8r53TviwOJ5Gj5CgAblKqPXFGm6G96pXe+OsNdhAIfVvye15xkV7lgOk
a7eSSRfnIuyPGmDLaYkDSgXkBfqu9c411vkPUTYmn5ynaT/6zFPkzfrpZlF+TWp1
cscELpHMVL+WXRqRfxuK42S6usj/iJ8FLdSH25/5G6NiBAWneMkURgbB4avVNiV1
6+JZyciIvt5ABTxVnksZ2VICd9t+qvhlt0zEt6GZ5/x7zpzzyRYA7ax0A9LHH/jr
S19/qn7WY+I+sziT/4l77IggDWm9grnKOTPzbTrPWHkvCIatHZfBnEGFh6mxyHy2
xxaA54SLy6ADK+voQUUsK//IapKxW0WYVmE31BonE/OaN8c85EJ+q+BnL1D0vDXQ
Mrn7EXcLuI3mDTC17NMR4j2faxtVIiepnXvJb4Yynopy0NRKABR+EwOC/nCHoJTn
q7yCeWITtIjUNwS8B4HZHLCXBvQQsRsuyuyVuy05tp5H12sK7/M3ID+aKZ5Bju4s
g1n6gxP8ZTAjVSCICiSKiUn7mY82BOOXAM7OG7NRXPxyE+AEBD5zAJBAtKpxjSfb
zKdRrZ+rO9usHQV223xaQvy6I3ad/yMta2UC6pQeCc5IO88Y3bOdo8XulMWaw09L
qxOlAnK5cwmL1ybqPvPga5vkLX0S+8laTadieZfIbQVBB90qDN5Alol5zUPk/XdJ
WLLy1+bHK0mhdpytGd2WDE03fRN448IdKhbuM8ngYj7u5J5yyOvvhSpgb1fTNXXm
/Gmq14eCur56RRJlpf3ujdLPfF7txirxjftAlBtTPUvcCPPrhTI1Cqax5oib/Xt2
0tjHeE+FmWgkPo9a68Kxm+anVQXeFYhTNT0syV4A/sGZyoCo+gXo5HaAkBQVwNzQ
r03T1XoiKcp93LjFDBDTlyWkVlb4j9DiBGCRzlNAlarR08QdnxhBC3xSLp+S1Nfv
rzxOx+oDebw34Sj6aoBSTJF7EscpXS56Am7yrGZQeSMB8aThPtfdwR7eo7HTiMGR
V7eXNp0olGED2R+Kpmio2GpG8Yt5OAAfuCK+H+bkhNJqnTLfuUYx4150ZHtmUBvO
HVjJsT9bWJoplYlS72e6PjKUp35zBeg3vThVumYFxMjP4D0PSovdmHyCkf+COSkW
EmuZjMNW69T7FaytEZsxpxZGeMNdgotIGAEoYuhR8ZDCH/0FGT3+va+Sr/TDfnAU
Mb9fPy/kkVlOgHTGtWFj3NKIjSu5Hgr9IpOlCDRhlEYvQUUHkD4EoT/fMUdRozlt
FroUMtsp2mZomxwcwBBBdFCprRrqrQaHC5uzuE0JsLH+gbxouik20yE+h5oPBlX2
w6xxnS/IS1tKsj3+TZcJi7CKJMMYuQErCVyVdT6v691TWMI/ylG83SyJVzY33VC2
foB9LDVa168qrVbwBBsct6oUD6/t+jREML7INmncdr55UW6iO2inwBd1YmHQlf9/
8n1ru4D9MSId7x6kk96GkbrZfeL9YyZrmj3S0heMf8MREzQCOyZaAbyN0XQmUwUY
54WPZY1FlHEajWDHIUIYVq5FPZ8FMR/PI3JKjlGnwjo71mC/8GqEFzwAUGuJZd80
+r1MyMTDGPjdeQWwbyMTXh+8wCR7jI6RDMiJ6RzCQ7uUN4uFj1hxVFbBTK2rMyRS
nFTVHpbLN1xWqCdO0fidoCzFTUl2OQ6Gv9Kqul2MZYUdAco0jR9k8/BKlUnufS1a
ZYrg67J2q0lXMUx3GYWlNkoFoowJC1wo34dRlGPpedfIR0MBtaGjIQtJryWn0m/4
KRH80JOT9DeIBHErpLQA2vPwlhOEei/G6RYGuWhH/i/ZW36jTiM3KjhuZnGdWTpN
ATgXF8nayACrjjMY7W0ar/hMl2gEmVPXCU6bCkPirKtUotkGI6qIhltEPQIlwKyJ
uvvX+0M0ug+bl6V/xzhsWjfVwzkqKcP4wRhx1EPooY2RT8D7S+tTdUAZPySqLQhs
s2aNCGoxXLGZauodZ7jajayrSzaCA6AscubEgLZkfpDMzfnC0KrRkxvn8H4/J+Hj
QCW0Yf3bJmA5fXy3bl4SkiOyKGF7aGd6Ynhm4/Dl/wUfmv+d1lccDVI1w3kGD+Fu
boVeTWb0szIXhLT2D524yzqH0Cr1OGHzsVoMEVzjeo2/ofrPzIcHI0yMvN7ogzy+
jPWSMu2NtAu2o40y0rGvIheSjE0toKCNE/oIRRnpqUGc5DelJqXo6uel3lSk46uY
IWP3no+LyOTvOiF/xM5c3HSUcBPbqj+Qp7UYezqIK03cetz3tsW/MxmYXqMnowla
v099nbetC9DyJfJba8mHc/8B83wdsK/Kjg0L/VWyiIc2xzujfYWbZLJt+UjGcpCW
uJfOWM1R/yGaP0xZFv7Y243xDGzbG13+ep94wDxlFPJNEXAkSp0raQ+9afQSIqFW
nr08h1Rec/AlUE4mJ2+TQLQSbnu08No9WX23ISQZdcleAt5RBVYXba3jw3de3dqi
aHe/4JxSWQI99ITg4KX4kE1cVBI0H2dUAI/yVkAMpcuX6DAq4vkzHQiQJoopcsmh
+uU+9BTBXIwt+3HvlSBJOUZOFvQouUm51H5ZUXZK72t0IV40Z+tdH1unLZaNjVD+
h4gsAkuE4D42K/9A6Fz6HPw8ympVLEpkdHnHB8Hd26DRAcmx5nxSrGWtoPCGTvc/
hZ0XCwHxeihS0PeZRCo7pQvSklwqAyTPkiap3zgAjbZonEGVkXgEUE8YM30o2Pr0
YfW6E4r2GZ8dRkOZ8Q1jV16emS9SB7qHek6jygvYroq7E550D8fJzVYmSCRiTagY
Z+V2oxJNmmQbIcAjfMe5NsfJgaPzy0ahybj5R+j8H6XZon5xtj31jt7O18PC8FiM
s+t5oN6qWIbjhiJwWjzlQL7nNBDdaaMO8YG6o+lLmXDAAhstUoMbg0d1QGw3uwL+
1NpJ+gvTD1YOaPN7vyXaY1ZDL6habKC1tjiHBjLGtqg/WwyT9HOGjUSGWfVhvIre
j7hq35b6Qz0GzsCpuoXza3lgwYSqRCaWHyqVeMcfWZ98B0tQ+PFJ4ZoFhWP400nz
PE0KkDlgXoYiOp//sOmMAORngcOyPDkTqqJy6+WjqHTN8xk670xKYo9uu49SOz8i
weuYEpgeRIfcZyTo19+WRiWsiyj9hukgCYonSNwcSgtUVvVnGpeUlemFCHGDlAA8
x9bCtcXAiPU1wR7fcqHFMSNXLbePrrFXvHPb69Mb51MFkFyCsRjn/tCAadhQOai9
pfkrP79OAin4VDWoMTwJ58hUd2UYSJuz0b7zoks5VlNLYIq1e8nMNYZdPv5T4TIi
pOtxBJUI9i5rozMtUKCphwmGkQqm6SLauzpUjjwtSJNCcS7SJrnLkIHHdEJl0j38
UyW/bw2xU4nIR1TWVDY6z+qcZwRviD/G693j5QiYksqGJxOc67PSmGp5ZpHSs7Lm
UDtYVqluKUHL3Xj87yaa0DhOXYlSAJGkcNLPvjozhI/tSmQYWbVjKkKMuypcb687
jTa4VBFe83Z2iQ1BGgdRH3lwJW94zp6RVHd6P2txKueh5xbY1zSSucqkVR2n+g4Q
piIHW+w3M+ABYBuPfsZD75ep/d1+dDHPc0mSCpnT/8EANSMVcYz5ACuCNEgIr3f7
cZwEF/Gr0dUOpJrtmwr4iJi3+DQfAjQwfH7+4XJ0N1PrGO6mY53GLl1U/kn0Psjr
niPntJq/Kpgaehz2ZkQS5Vq/t/MfIORhBnaHPkScyx1NT2D6O6N8LHAIapA4SkR9
3kYeJH+pit9K3JTonpr/KXjfWPSgiFpPlsGjLg2fYxUT9XPKa7MX9wPKSbCXU4BC
uzRkUO0xdhuPekL1VzL7+zVoPYMc49Wj5isEYkGzmRnnm/bE5yZUH+Vnys15CWK3
TNuakNsLScBvMnblnAq7cIvI/GcNqHKV0jbtsRT3c4jcMjZAUdKFOtYqAtmAr7SI
NpbIrCwrSKqw1GU7FDlCZrFWKKkq0tJKScH9YxatT4xEc1i9AWnu5r9GEAdapBBu
zlkMAMuL2DMUBvBjGr+7ZjgACHOuL88K0S7clttWe0Oau8nJVnHoRoiN46t6pSAP
u6khubPlJdbFYThU0zjBw7wtVjCWQVA/eaeCX8ymp91PTRo/3sTAX6haIwT/y9Se
iOyLdKjFeTgbzjQp3s5vwX5IYjYiJMSrav+58Mqa/VknrjEuIyewkJLTutSHMI1n
E1g/yjoEvwZZeJZswD0DQfceqpcHFP8+UrxFbTWgXxVMK2fxeQgc+cQbvpt8x38Q
zvGEf/Ia0TzcGKmbcC56TSyvepo/5bM8vgLzz2RVlIkvz7cESR95icB9PjxDB6l9
QifVS/L7gPoLsqGSZJxHkcjygg1XUWKWx/Xr6hEbcQpTzR6XRES1sM0DxnbzQ842
O6x6yZmA/dwlWwOYyRM7W82jGZOmmT2ZacOHnjxRUa7h22HZqxSs5ww94d3RIWAI
LD1o4qGRCaDSAnOSMfq+6MrhT2IWXqEwpcTQP3UNGzT7gJaBKlreeWnR7UI8yfrf
owvZ/ezNnhKgK+A7MmwxPcLduZv2P2HsQiFEDeyHtPAwXdgxZKyUAeyKjYkBMKzC
icun2BNnWFEH7sGk/Oik0i45DUT03KCho56Av9oPcwVnIxhRNjAwzzafF1p1KSS2
BznvKrZB4R9nEn+0X3T/i9J6qIwjnMkTa0whajoGAb1GdWgTBYZkaSloZh0j/YrG
ugBayxjiypk7f1JIfCJLD4Fe6xmaeaQsSLkQ1ZD2DnuOy+FjA5lD9AIm2oXMYHAK
lBVRHPSPK4UdVQcyCWFqzNnCcav+COYsXS3OROz7clnRw1g02kf1ZQCCiLx3PtIt
S/iJxyamUyixRuwPOE2TbN+yUKw1/pP5aFTCEqBOyNKrOAPL2EFJjWnZbR+1W6bJ
rTuR4sBXdT4En5nk2NkMwszaPJnE5D6sYt4FwSpV6Rb+K70M32AlthmLtU29N7sn
Srfh97zwLHyYEFbImozASI9sSed/Y37bckdCuJXb2gBCMrnbwfac1vpclKYLUB+i
JKrOtgu0U9BTZew0qI0inCKKLKIcWaBbRB6ZrOLlF5x0Xw36sl0+jytrl3xyehzv
P/Cbx3apvSG2IESmAdXP0zKFib066h3YWY7bdYa23oE+qq8M96KQwsaTegib7Aev
8RK/9WQVoDW4w2zth+a664rvJuPFjMFvNKZmsmHAE5OyEvODf4cqGsPt0uTWaMWl
0WXADYmIlOxaNzqiifnT+QXHefX7zR2HT8GewWtk97jLMK+grvQN9qTKRoKtLSve
Qet4wIewvZ0wRwQ71hirc5W7G7ra0BId6e5VnrMnUvD1AVcVYBEoEKZ/H+iL6Km3
DNhSJTisdtCkMyu8JY2ZAxCw+ru4xcdb3kqNGD6SiCYFBNGwYG2sDdTe6n4p2GYT
V9n0zor5CGiEIP5nqnR3GeMzkDdoa0hsm+tDVqMvc2F5cCLBL6Lu8ZG61RqiDyEu
kmMJ/6fAr1o0EWdUnAet2hwLaA+WuQMdLG0tY0a4anXgXlkiGp9XL5mU29F9DTC0
wFQNhZzlOqvIXQdeIoktjkbuOT1nSThevmEf9AhE1AFfcMT74is15/z1pdUllD8y
iJCwBg+4EA/loIkKHZei2C03GHJiT/XOfnBkAQPH7tJXhCIxEYu91QyGH3Ti1alh
UjjAByrIgL238j9l5LGunSRe7oJ9wt+QTUcQs3jvZOwEO4sL9bt3jZPvY5Lx0f18
OLSxGWQjAQSucy+sJAN6m7dVQ3dMyfvQapDtopf63MLrL1oCmNo1aZ3rmvTvupNv
Ed9ycsOxccQwDgY+7OwTHfdFdbhlmfsW0fnWaP/msOOv8Lx+D5tWeOEaGDPgwA+o
WKPnCH6Zkn/KoS2LdUIITLyDvhnSsdA5ShpcjvXwQFrpSW9CZinsEkmdaRj03+xU
4UHVEgAktLdnwCwIBfxmpODqnbYBKr813hZs/aN0bd2aBmTLuIrm+b66rlltRRBt
gJxPUd/Vqe6jM0qrIpy+nXJSx9eo+Ex5VFZGVuePmuxeDKkT8bz67u4QtTS8SwAi
5r27q6oDboWOfjWlA4DydjHKi43dGqr5kM4tuhNMqPtpG5EyQQEe6i2QWHVnTbD5
+Bb6CVrrEE27sThL+XkG2dsPa03Q3ezTkTmI2ABBj8TmKF3yd4FIlji3s2bDEPNw
QxdZcOo/SetWCKpDJclPorl/8U5vUwnchL29Cx7YyR6eEgUZe4CdWDIgWipVj9Hc
vTFV8+hV/6yQXc/hldLTmyzwBHxewhroGF0fD05/GX3YhMYUe2ghUnJg33jjb9UE
gwhN5tFQl6dqr8Uo4tLo4yj+oe61LK2drkZGU+CNW1vHsGCW80YgiH4HmO1NZKbx
1GOc4anFBNDtNCLAOhT7fuIIOz7LSiE9cd7w6u23IZyNuR0zbsYIcQEejR7Xnktl
i3sDDy9ty6Dlpt4U4yGnOihdJY2yy+qMeASERlemsHf9Tnf55CJrld1POwksQlrU
lFyP2o1jaVPGnos1XeLqx2fzhSUmJ3Fnq8nEF2eTbXlrGl1OCJJsbePRpVKkgQPL
znpk5OMQwwBkxTapVJa8pbnBnd9AZ3tH8yP4E9ZDtqhXiaRR5yejujPDSupZFRfC
IlrAjRzOaSQCU5VLtYsaCx6EGoen0s5JIs8YLqjCfQqnepiEWkAFdQYxd4deeb+E
WU85fPr/DXkFX8BGW3JbQl7kRSsHYRPPGckJMAIJ+J9CrtetuvP3C0GuG6J30gBL
MOe+w5pqnj4QK/CylUxaJvU4uDPRSB5QRqnza0+cm/svK2keJ/t61pnf+xvPmqrB
rsBpabBj3VxaDmCJO11W2n3Pb2xQV4NyySqazig7KGZ97U1QZu04rvdG6ZXpLAmO
TlgNVFmHBhnb8kg3KwIwAlFNga1Ss4P5kJ5hZ5hR4EtUOWoKpsZ16Maf0CVecSdp
ZjH8ydgQ38+cCMP+xCbxkaEwjmi4A6oCBQw2Bo/YAVbsVseI7W+DNP8yN35lYB6w
uetoaUNItoAOgor4t/SFpOiZOj2sXWiOlK9jnyh/ItkGsA6/5vSEboo51MY6lxFb
qBypKEYmyFBwrEOxhuleJQ4XgxT7Ko/qGjqwkHZjkeBJVigLQArcqciP5O+j7NNH
933B5kX8vZ6WhQ2ZC/135MZk5wS5/s3curg3DZLjJj4bqwM/euRdFxfnRfE+zvxV
a/ZMQUzn7Tedl2jjvEFC8P8Ir15ZEhKvgu40iMhRRPKJH1ds5t2g8OvMlwRcrChw
hdNL0e2ASvyf6kBW6c0uq2scOCK4DBVabhAEcG0m+v3vGHiFNYzezrMsk0bxF80s
ynLYk/mqyM0MYXMOmqserplk4Xygqz0ntf+BBq7aLdHwr9Uaw2uux9v0SKdrXnZD
zrqnfxkegJJZ3jpjVdSRhTi/96dpucW0yq/w7rTlC2lZSUBDTCgRq4BemRMbEISE
JJJV4jHwRcACi/Pp0XV10fSmxToEPyn3r+Qwu+XZYCx0QRgWWYYiHZTx8Mr3AdSJ
h0YhF3denV0XvN/ji5FTYeg7PL/Em9Ly3iMW8WYjL29L7ySOmdlnQP0wyrp2Hn5g
Hjhe+D2dkLeNMucx4ugLqcaClsLKQKOjZ0q5H1Q7z0aQuRjRb/GhV4AZtZ9t1tOr
WDpfWmJpoGlGaE3BkHdMRZHEY/nRBLVdnFeDj9iWjrXiUDC81EBJGR14lUYW74rh
hywz/F/7LHxMuVE5zqeseJ54luuW2AMF32wvzPFYnlzBxURcqHQvEJMyVI9ZD1DW
W/etSqDRYLALNR/KVgl+TAXTHfZO00/lxKFN1ALEYTbauJCboslwg6pc9GCLM6rt
U5oiy8F8fld66eue//VItNuXC/b3wohWY9kiZDRr2A4w5pBpnL4DzEZlkiAY1Lsr
7gIPmiaRgwKr7N+Nzpfp+r1t3080dTpAWuoiN5skPxA80z3XDFhm3a2SMrqsWTv6
/OPM96yoaF/jsEtX+DoOpiR4BfU40Kx7rW337Ds/0NiX6wDBTfDTPL99FE/K5+3c
n6iYD3DPXJwWKn4F9QRlSAF9oOXmu0wosZOfqHZjn4LMggoREGrzaqrk4PFW/D6c
/WMCkGgNxEC8vXPE00ZMu0JMBH19+YNGY4wFc5PLjXLkP5VjLHMOftkYiJdgca1L
w/WCQmGJrC0/nB48X4A7+QD/6RrLdS1PSAdrUavrnJ9cs9D7HeITzq0QqLCF1cDN
XmgjqlhCi9Wvk3hL9LDiLPZvAlz2wz+GXWWvXqbt/Sv//PY5F4hz6/aZUZ38Xuwu
nXUWbZHYsJ8Vj4vlPpa/+ZcGiqAdAcu1FFkcEiTlbVMPEX4ICc9T9JCnoRwu9v+3
kVpwKhh/prO55ft74xIefNiVchlP/Fi5sSdjnq97J1ZFumT0InbNVtntWljRRV18
3VnIpFT5OOMHTG+LroXzdBWhSFnRwnvFjUIyVwLtUVniNpkOqmdapTluyqzm4IN/
dGBhEOjGoL4K5fBKPZ8E7GuzwrTiyEfM5llbd6D66ax8w5eEhWe2CajySwhH08DB
n/1rmCczJ5XyEo7ORs3X4RWoxuQuuMzq943WykaqdEwP5YoZzbPuHXmCfqQ6e03L
JlbZYXTQYbPsOxuSn+a1uMSInHXCTJzAwfSnkHoLmrTl2MXKCHN/UBCuyNJfdas9
jPpcnKjhkynTLfP4nIq8EEDxUqj7ogLemPuZ+9w/XO0dAduEdtwCkNYC0G3llAJF
ew/7mMMWWqMawbOTAdLqZOFvxbSt31PAzCk41UvqgpWr2sjYM9VHk4Zn6IskCfkL
bWEkipaOPnoX/xFsSiMpFYyUw1lS5U1gja+tgRl8M0ZvWEbGmbQAJn0KPCS9af5D
WWIivEKllDSvwla0VrsbPpAF7DSjuUtSWygMX2sVmFPtOgULdYSJA7EGqCXi4WQW
6kohuOYz8JVBmb10S0qVIuIKt/9puoOqpt8KmB13q2XmZ/OWIQMsD6SnBOCRD1xd
plIX1AJGL+JbVqYNgOZAeuYusV+S1wV07Ks7XPrT6p0ybnRn05oM8gpTT4z+12aR
pRXphWEJjHGEIJB7sEPc4TcHmnw0GzXoUXgwFN1EtoqvBGkEehurCBhBroPS2uxH
itXz1auoE1geGXGla/NGBwpw+/R/EtmZvAxTAmVD/FXLZsLk5YZd0SfXW4K+DCpN
0TrPVO1zhTquntCeSXLrgDq7sYgK+ZcbEnlUtJfAMbaFcl7lL/aYjp1XYXgveQUT
e3pBNhyT424g3enAS0INlYyBcGP8SdR5BDMWdm73QhaQBdxMRo5qBwGtS29PwTgt
Yf+6+Krp38dGwxO+1aqIhNaLMcvGPYsytrqEcJvo2mAKjkx1MiPrFD51KR/rJLUz
IYvfcUyxmn56U97qK0obtgfYZNXqJHDX6tE+AatViO/EE500I9BE1aIsJd9UP+sz
BFWBRIZrNA3M5HYNVtWIXATmIPbjSJlc0xQak2bTBlFu7hGy8ybT/bTcR3b4Zvpi
I1omHLDvdVR4C9/BjUxiPcCztsfoylkOOmuG+OaO+O8HxHjGBPFKchpI0yxGQ2ez
Lu8VssTIMQ/rkT0UfPOwTB11JHaGQVdFtu6iNt8CN0BgwlfMdhjgNo+i2S5mUQ48
RtSGcRUFlHjDN8rc400y5OlrJp6TMWHRPVHajLeYXYCxw+v4JAtN4ryYIjugvFFa
GGzC+q68x7+5B+24CeEq0Zb03dPsvrFhcp51qWuy5di4pEozTYReIj1gkN4SpL7C
KBRKBvXHWtiW1OHobyoKE0iI8vzVw3ydcPir4uUfdxGT7E/CRjgsSnvbq9EcTIvG
O1OpuqWbGzzrirK44hNZ75R29mPstCO5H/r9yEdmQa+JyxcBlieC2cQyd+xtAFNu
odUtldy1rNMJ8He8mu0Sx5oqrjnRsTb3OGv3CFEp7tRPQBgkeYVjREQKAWhHq1iZ
KPFzN+DPbJx5deLMarmd+5I5hPahOUpVHIHZYydAZ4h+gbddoSBcmlHcKkAhHaf/
4dgFwU67kYfWOC+uLixs8KG+VbBTro50rTIhNyojmmiJyUlpeq4g/VLgzccQdRo9
jWc9E9a1EFbjRON9N/9XpHOGxjlxYtzaQK+/B32CGy5FsAmDJL7Akehb1Srgqhmk
kDFXZyJseU8abHooEmKgdGW6mB4eic4a3QNgF1eW9cBF1cocf1jPzsUMcgfVCVxb
WR3Oh+dJZGaXmZVp5BPjsn5gueKyhOG+lmo6B7rgqqR8mZbKhVudNawcSM5FilXX
Mj1RizFOEsAzpvTO3kfVQUb6FjXE1XWR0UibQ1Uo+MVSyoYM9fwjsMqL2uwwjpl9
bdanKvlAoV7NuXPbv5MIsClJeZ1h4VO4tgjI9pocF2AU1Y6Vb0s8fIaJlJZZivta
edZ1zEB7qsiY9KJthRmEjdCfnVCYgnqbfxpEpuu2rp6dqNeEyH1zdSCh4mcNNf1p
XOvSnTmA69NFDQkMbmJMBHifUb4n22OVFRzoVJeTlSu097FDV7FIDt20tK11ZHNX
VJ3Mb2I6kp59EeIE5vQ7B9+21emSMmk6DL4twVUrfsHbWlJ6B6KD9a2q4nbQQmCO
Ou4JdO2p+LNzy3LqLh21MRcu9XUF5VxjFpXKwhU44NTO9ooE/csLx4P29ARDWhls
qi2IR12RDplH20QG20cM31h7bu+ux/vNHuoSR32Yg+ZvesL18Xcbjc/lJd0MyusP
5+Gzsq2OWwfA/o8JQIL/I4NvdeZhm9x8nrE9vStHQTrNbUNtLCwUVt8b2V+tX5Dk
nKB2lKOPXyhDKnVYSAPyoaFkMFJxqLV/UW5oFCaYio+CNCgnKMVBgvj42TNJKdHo
R1+S0XTpjpRJN7Zfl8vDruHonGdrID85JzwQC7gUVjAgXDq6ngWzXevqgzuYcw/Z
kZIJDfYLfGctpS/EBr8x7T40GGXox4SFKN83Op7MOUL5E49g2geghPFzFf+Ev367
JnIRmIHOUs164ClEg5TwOoktWhOTJhJ44l62cNYTr3ScefP22cGvqA7eWwE8Sp4p
jp/CRR/+uSjqagTe+Uv6za1kwTQVgid+X+wcI2yZaDAvR/0e4ChaEFdMt0yLbqoZ
fa294YTH5gv6136d2QjUHdEXCEkB67Mpn2OGyut0bELDeMKY5DCovOF9nJ0u1E2h
RztuMIIfHNrJFwrLOGSyfVAkaO1ANrboYt2jXZkh/r4upWNrlAH/67KoSPGNdYgz
41vwiS/ogEHJ2AzCZkgIBrWRULMDag9978CUngHpX8JUbnTnG76GFDTo705W9GjD
ZvmEQKXl8jcrbKK6Z+awW1mwUAgY0HJ37vIhUH68DRM6KWRWZ6ap/P5y92/F2w6S
aeqQnaw0+4WmS046YPigqNzyonVeZpCf5Y7NzGatkz/S0SEfrDa2jOz6erSsikYX
gaJCtrahxV8zxqML8xw//NTEBOrt5dzw5Q9qW4ib8g7zp6sJT3aE59kXJfAQU0eY
SuWcBn9uLyQeE3zdLJiLlBv+in++yFnc3OT8U2XAKgbjHh3FdAnvQQOSgsmiHzR7
FsX3loqvjdB4tHHIDESwlWQU5njADIWMxxVep8Q7uywb0j9d2ECdEVmwkHZ82ail
cX35+aRTgsGB2M6NuCGxv/wZvbFv5YwtKCKnhRtzppKMHhH3M2P4eWb8r7pTr62N
MP448jzi3iXum9/xYQ//5rY2XbOgV1bTL5rOF8By4BUuOv6ZJ17z2CD6HiL+26bO
HmTJB64YDrnrDM6D/i06oA64qUGIuGA6sCnJe1tIKvj3b3AvDaraAEZFRh5b7wcp
S4iJRFYIyezfaS3ekuctmpMvfM58J2w9BYswxOg/LnipUMqzhMAwrGvaEJ0kL+5p
qgspSSNUVvtL5d7iUi2DMRqQ6VKFzXVAnUImrBL+PQn+QbMZYV7DcSd8TZxWl9AI
nQ8CSIO4sth1UO3ILGQgv0xz34je0KBVPYEHh084X5pNl6LSvM40Dcss64GVDucR
STn55UGJe37+qFczRLJKkMfFf94MoYwZZcldND4F+mYree2Zz/qk1B5nKNmVafuh
XKU3acjwrU/1GYrXGhpBltuW+Ga6rlWgl/K4CL394Yu4HIC54e4jBc3feezZ+qJ1
5tGVh1tvJq8FOS5rWUELatrAdtbZ9md3OYQT8NGjeTSBSaG0nO+d8Q3uC0peM6UE
3dVgcDBH0b9NMJqH01+4mznn6TXYqsGwzrzjC335yWEY22pyXzIGUQw/fBqIxO9x
L86cwsQTLa/FqKnEM1Y4r3M7f98d2z/PxCPeGLA4TBc6DrDAHJ/6BD1uJO8+pcLZ
YR7VhDuee5R0YR+7otxHWPo+T32y3quBxy/7qw/MbEvEpi41TlezGVZ6wbWTkCYP
PyaOIHD/61NJXuhW3icyswD2PPxW1oEg/skrXu645eULWUAYtyCX4P53i8P3ncEp
sEIGGrNNoLVgcwCaAm8aF2K2iVkaLTIzbPlb4CeydQXIBaiLf+2643Qpgw2AxbZs
kFusz6TZXpQYziCu5WGzFtwnrc/C9AhMfOmZMTGcbZlk0bNCYPi8xQ/gvK/i1SBb
j1ghym/fvwFAkNP9OWzU4MiBoTLfxc5nWQSkBw3/ABOBaPhtwW3+0ZoTb4qMJnLN
4onNlTeUUParX7kBE7w5T3rtkSf3nB1O/CtKY83eNBzSN1nGdI2d6ZVtbWPyCRYv
poMovtA7XtNBORHMO+Ft7CVWPRuH44W0iHIsWtUmt63tGRt0PBqMig0NaJLp/MXV
iViKbm7zbbVagHlnoFFn3w==
`pragma protect end_protected
