// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
epRZSfgteY1+kZ81AyXnGTHBaM+fdKnFNYOy9sFKDXVQYva6CIx19Ti/RWcSUdZMFjjA0DbbJIKY
FetEt8RZFef5OvqNmpalVUkprvTC/LAL2ckFE+AYrks1KcM4OVIcxHnQOSkXzfyINyXBofggl6lm
rujMPh9fCttkUIQYEkLTy8aJzZHad8wyc5KO+7VTeCv710SXUIZOe9/LuSbnp7+tf6TAhiwoEzd1
/ufekl85Y/xu+0fhO5hAE6vxuFHFl35/f9XsW5ttvwxoyhqyZZ9x5684G6QlgbYg0ET/pVvtKbTp
8u4ncyb2uSPbAjYgVYM2mOdqes7TZhPPteb8Pw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 55328)
zxGTgI6sbDCAv0HjHjY7OiXR2en0gKPe13WenGPB8e/59LQ6Bxwxte9BwQdRb0mIBP4P6mZoAY5e
nLj9K+GJQbI1X9IUzCAZzeYktfgwN9b+ouVgYnJdBzQquOmweQ4JhjXr6nhBWSiR4XcEJ47sb+C/
ChM/Wgrc9LRM3B6Ky9YD/5DS3VJY6hgCAy+68xPaDCbapG+Oo1NjrQu+U+xewQaWmlBttcLVVgOz
hkwq7ehrxgl224MNl7f8xjyIpWaHToL8vCjsrHnB6w7PNmQsm27UeLGobQfoYKzJgT/gvEINfMJa
AW3UlxUN7G3J2puFpSVIC/sv7t+T+/BAiutjs6aNKVvd22VJU8Yw5Br09xuvjC1/vbwAbuO44uZt
6BIvsRMgNqL73xZUt90yIr5L1/oSKMKEc3QGGp8AK2jeqZ1/Q26eu5eU04GJRQ2v+iVoDIUh9NOF
haClAB7p0Yt628axLWeIWsEe5rT+rYrdaJX7cmLcyayy4ufFi/mjeZXKHVgnT1QsuYJgia/TM1O3
4G7lm1jCzn8ftdGYo/syW5LwAbSuY7pNIj0e/qQtHvEx2d2XZ9q4qeswC0CrMEqKeQIMsveUKFCI
ABmFGWsDX0p+nwIIljgT/H9mPK6RYF8hpHd4MVZmO2srloi2Mj6lCLxBpTQ2dRuDRnTGVpRVpADU
A+G3hx8IfjTcwHHG61rN7yx8QH+BUC519AA7em1/HhXfJMHw6afSGRLhCvFJvVoFijamm3taLDcm
SEiaVbRpxbwF/sZ1KdbYTQ6WLNOWZ7uhFTNoAB8MMUEUF2LrTrgLOp0n2b0cSFX91r6Fi4RH9b4r
6nMQh49eAyJGieyf0g9so61/0Iy5gDXlgWwALaDQsDAr7UWdG80bubS4x/hKF1cFgFTyZFu69FOq
z+OJ510l9AAzD7OujLFTLh+/7obrU2RNIZOAhv/0fNlMo/CniAWsew9O86Uwg+/ZxBSn4n87Blbo
aOuMDX1Giwm28XXnSme8x6ThQnuPVnYcS2mWn57fOgPQgiiU5nfuzDPPpbZ577w/Dx+zMYRp6jTT
H7YVgPQKQ4WhZLZWqNAVH3v+5BRvsoysaeGz6nZt7LDoBcDvGKS+6IhhGLoT4BZY8HRPsDC5KdIe
w9SPLuKI5hMHCupdroZsRhZpj9XjiS/gyXYIJFmldJyv7uW7o83Pzm74x3lUMPDCkFxmPEd3EyTc
MzX8LuY3O7/pUKKb1JGLa29ouQ5XLndIxCWYa674ULWWwqyWpuoELlCKTMhIZFQjH04PHDdOy3IH
BT1S9J9Wt3C5cShX5kMpJ+5FZy25hZ2HfJDn+nzFwWvqrAJTPxsDEE0g2V70Pyeai4fyiHh/psm9
4ZaOILRqTC+N8uAe0FFFvTTq+E0ae60RdB5pEDjXUUnF92EHpvWj53S+ukowBNLkBpwaSCJ/GR19
e1QJgH6mKnfW4+WywsTEseBZTvd+m5aXuV/d6udv4vUrVHXUm9Q42x5RBPmRJ9BbxzhktikWt3ya
HkOTWStkQU5+G1ivYNgY5eMJVToUEHDKjXoxYmkdqN4AGdNBFpytP+Sugo7P5tCMMl+Xud8GJ3rq
cMMIodF7kz/hE631VKkLQ1UpH2zmzRAb1wN18p+UuIUkPgKIPKjfYupP0bFICKUI3TX6/1JI7M4B
MY4/Kh0i1Kta7czW0GGWMWP99fGMyXn+PKA/NdE+jjPuyiQQQFzB0z3g/ja8qvUpU7OmaDuyUyoI
JzQBf6u5RkuFemllxdTQ7Nw9HMwvfp2H+nQOKWFFdL+MYcPn7/uv1z04yI7QnDBqiJmdMEWZ364g
P5i2CG8EKiUffiKdSq77Ox4hUoDTyc8cVM+46VYSdg/Qd2SOA7iXh3gxRxNhlRxf5sRGxxyzYhen
SCZfNo7lMoojplAGvyCLUBgBsdtg+pg1eJabydoyEVFP4qPWBfU205uaF1fDu2DJdVIOfOsW0eA1
Ky3uVF+T4bSoMxKvXj6qvSHIi0N3NnEy7iPgPNADpfuOVDuDS0Uli4Y6kGQ/yG5TaZb2cZjnzsMa
EmFdYePuDZnoEgoV58ddPtQyyd2jfwoCgOS5dde4jTjlLMFGaQzndTHe1GK8I+JRHfVr+JB+z/hy
efv5acbFwYKMCxqGsyGOqPA/+Ba6q7BaSuYjLE8FN7MgCqY2c82YbRzdXKLYfoLyLKcFTa36pCeq
WcUDRCsy9KBAwbHSefjf76Mu0avGdW/YZxAPgl7xK6+8ypJU8f0D8ccq3DbrWlmK3knTgeyQqsWV
RNjzQNL6baa9Fs4jCj2Q6jBVh2LmsFHG2TnOaPl9kCQa/PKwjLePihoaVMYiTm0bMMLn2j2Oj+Xl
5/r5r/lBofZWmEsUMLVzVYXzY0S+HXwy+Fq+6IE4kw7KgmILMbLGviuY4Wy4w1F6bIvySKl3JSm+
/K3Vo4FoQvhYTHwVeqLAo4cyxd3C64642KeC2M5q+MW7005qDUFXxTLUK8SSpIGGfuup4cWqayxT
F+QCTUKIxQqtKLPXrCCULnLzf/Ogecn0ZggagxOjNcaBlbzXc2PCvdLvDvh2quHyfWQdbufQRwcn
AwqGSElM56JtPr8+jFgPFwULyj/TvanU1csbPvTWY/DCpO9ADzVxa3yTZTJ+l5ugcJ0CHwcJIBB9
LLt3RqU6hhlxNv6/NAIUxJs8o0JIXZmDOfR1Zp5Au9MIanSx/QndsvC8NQWZJOapXGde5ckow4SP
0FV3Kg5JcRHA0MA9jsJrT62GaBGF3v1jy7tEUhg8AcSeHUs7M5bShXhLwRqf7GsJP5cKC+Tk3Gmh
/bxWDETZqMILylaS3hep4TDSzfzsJfmwE7R66IAShTJD0ho55SsNsg7uvkjq4WtuBD+7mbqqUbE0
XexXbIS+oCfmifTsnfKuUooibzySkHIZscckecfmcliIOi7zaofF7BVN8wdu5uydlwMjFA4EVRKl
9BhDGrdVCZ48lF+hjGja34TZ/cZUJE3cN0aSgCfX+IIjqke9kX6FzAdwPmfmPkyl/ibS01XT3sTM
fKjnwCHNCZ4MS2NjkHZVM2g9Bn+liWYONWo4dNQXdMYjyhChuuatYVu+0wrJSQjYAFRG+nNaN2Gl
tT8AhI3WaRRAcHqxXOXrorxU0IbqyT92N0pVea+n5Nka1rTAY/f9PDStJM59wOSXhRElhpVug64p
deQGWQhRoYOaHfwN++afo2esIIpxWUmLnXmQDMH0GnE6VjaNH41eqJPqWAu5jDJmM8Au+XpzBOLw
Eh1Su8shLPP+I9FiYc44TRdyMXTlVvy1mA5yDSIrjQjoqdZRnBmICTMg6SV3Opm3sExX8BPthEL+
YoPYtxMisuFyqLRTZOjtXb+OW9gnGcN5H7qB/ln0LuZegO08+lcjnkuGZw0HMU/D88YvIzR/NOSv
7fjcIiLAvd4eM8HGPgEYfbJlrLAR+vaJGOlc0SQ69dAicNMgAWN8wm4eNIo6QO7IXU+/y8WysTNh
+yyHHXfsGwXss4GM2XbiebtyUzv5fLhbpWRplFQ/z+a++dSgYvMWzgDle/Tutn645TaCQsmDGyxg
o9QwX4wON//8jh62ybMeVAs2NCRwJmrGP5Z1qO1ZW6WKv0dg1navqtNOPeHYwCX3mW8lgECYwIs1
STpnkoHuaATJi1dWTiY0i/aXwOxMIdlAZ+CdRFfPt4sB5FyxwlooO0UV+c525o+FjhH/8Dxl7x56
kw8lNV9xsrq/ml77cx1rWnJP/S3WVt8nsIKYeNrXlC/SxNY5gpUCoEyHE1RJparX+mJAbxfBf4iW
4cMZjnsL/BBNCbmd/KOLYsXXqP1t3pfWu33AwkDISxu56juo/gSZRyCi4rOc+vk/vDiQzKbWse/Y
Y4Y2BGWdkn827qMjjRjfpNlpTHwkBLy+2QyZyJZmhat2wOmpYAasBIGMvr+13tsndT9R1L9HH2A4
4ICbRadBfBSF9vKr8PZa4HgvP1HAXqOolMnrtsPH9nhAiIMDfl73O+EU1MEcKZJD1oDkgi1rT+1T
ZDhao/gMZvSvAS1ar5dQ1qkD62uyIumu6dCxdk924LVjzaNh1NYfWaAfe19s1PSVhR6CjNxwuwlw
Zzh82N8J2HKkQYaE4ZASFYQ92bbX417SSSN0wF75B6QYymMcWenN9Idc3Ob2uWCRkIidaXUfKrwA
v4E8/rYQ3QRYfEowgUQw6AhltaAAh5P98Vyg0w/yumIb4fcHyTHls8/9vqGTvCyh6rNmjbKWQ/rb
tApuKtJkST0Zg3oqSecsrR94zCne+7/YOQiRyWBROF/duvnwn7L2bTZOs/WmtF63wzZsF3AL52o/
6kAi+boXGr+OBXvHRRvoNANmVIk7/r3jwc4ahC2RvqAH+Uq/qqKInOjK6D+Drkb1/RKX4yRPHKJk
4flw6EFF43awnJeIbymBdLVguQiemHQ7aJgbgMr8TkbNGJUw7uU2H/eSNDsjD2CIuCCF7t2eZY3a
dqJ4VJ27juNTA+nL1zXCFjOa2gndB3IIT9Z+rSXk4TUgo8yEJXNhP545b1hLa25mvd8EBEt+5Dwa
GV1heINy+YJO4RsKjB2NmVjIqOpNI2IuyzNLQ3dsBOzLG2IgB22j7z8ZEkTlchAzoZtPBoveMJL7
m+maGxRv7nEGDdwoY4QFooJumRxRyBoMAVkBwuzzZA9JI/WE+fAY5/7jrx8p7A1cL3QTWrL15/o3
M8KdWURuTxQo2nW0RnJTPz3c83AQHYzYiEoJsvionSciEjxQu6RqG8fjcKHtOVbqYXnd4fz6G6j0
coDUWd/ULqChvzuS4H6wV+49v4kC3QjaIZS77g0WYo7R61QYy2qKKb1S4pOqaqOMW7cBpP8z2DKT
rXoVpEF0ZaUZ/c9Cx+V2WMf6hi538f4kh3dp4PunzkZdUpsIX/aAJgMyngVAUARjMUrb0dauEslT
JN18USgcj0WhbPFv3zIoBn7hajllNyQ3obwMCxuU8S6GeFm64I8xjopTYMzdAD66YYcVhHJeDd8L
D1TaMOVYKDKb/On0hIjRdywFi1j22YUIqPudJgj27vv3Sp+k7RzCJD4udH1uUvuNIwM2aqzydrGM
b8gdE+YO0YU7jiWfn08GLbQV0SOVPfzgaJlx+69F+yKjDKcDGdBN8TWJg5M19AHKciO703L/tJ1o
934MdD/YK8yQ2PRQglNqK9Lm6fnHXqT861ifUA9OKXNuf6CtarTKrkSXKagIKJeeZcBISzR3WIGz
rb3pr52mWI3FvTB+xDjU5CYhSwGwECebIxv77Lf4+RE32XiD1Du9pGPa6qo7N4qUDW7HGIFF58nn
WulCU+Me42XkDMyurrIe1MDxUaiBD2uhKjhG60uEYMWtJJF+n/ulXlaYCXI4QumP8C2xwzpoGXCu
RMr5fAvJE8ul/eLPVvZaTZivR3ycOq/BpB6jIMfgYHu+/ikn3qzSCfnwuGs62GVL9FQqL2qZbtdO
qTh6k4jXIkkdJfsNxO07y3hFWZK1BKyTom6zqLRbj2pw3GeHpYI7RFpINTQhDu2Uc0hEJ+n3hAOo
9TxCHAgJipk2uACafTTUDJSZQQo8cpNK2LlVdjGifDkFwQoRg2AscvRiypi3G0a2qoRRvyEUvcDT
GQQ1eyHs/eDcj/idyMSty+RsWnjNZGnnWeWBKyuGbGXVO4ncLsC6iKbXnTUh0ZvakpS6bpjgxf/W
8bRSHu1YbQS/KKSVXES3Zdgweq4AZ/TeiY3w41UZjxUuEHHK6mbB8sN8cpT7SiCoka4pTmk/enGO
5vh0mpTTHH4bSujMtNlUcbwRlXkuKXm1Oz3iFj1ZVxoZlZdN7gxOI1r4ImcKeW4bMfVo1+ap65wr
SPA1feD7xetR4uuVGkOHUiokOxRTy47kxIqPVk6A1xSnEdHua80M+y1aBTpeySCa113AepHRdMSK
N7sMTWkrIVTtcD2FUrn6+OD2SHW6Z7dvpYE2vd1euMO0Uw0qWrEGeAroIKq2+1cGe9+eibhw8Hnt
bXsS6h7kSekWKkpUHzX39IeaUV5vPTDVE0McenNPijTF6rC9/3Ligno/K1oVEHrd/0+lhSR2kVqr
pgnZ+yD/wV+GW0nI2c1ZvY/IpoIDYYlQFxvf2ICUPF/C00GKZ9Ia8YmwzQZj/07+sISoyxPDFGPv
YhP1huAcYIUPgZ9SEvVMC0cyotD+VVvVm7bYCkDmtnBSjlfwuPeXeVRUYo6X+Fma4zA1ub7JmIqt
e2N0kbB66XCeBIUGbarwZbnMrpszuZem/fzIjnzFhVgrEEVSnhS9hQBG2RVR9Ye1p9XtIuhwRBot
vfpSqaO00NEKPFO1wLJGAr5opN3I5gWkgDSNjY5G1rjmyWdkiHrgqav6tQN1KD1zuM7apakL+WG8
Tfn1hNP5mSuLvAwJ0a33Rt5u0tkb3sf5+8o9ZRoobDYImvu7PwwxHo5VeQPJlisum86UvWzVr/Du
ozJOhQGSJI3qhm/+YcE/3clio301kf5wlsQ2k8B0DACu7bI8wr1fqWKRWhIYcP314DlTsFZ2+ZmV
ylxMbncAjPo3HdGeGdHmxvPTTz1HG+mhCTIy+n36InF55/E4ylfsH70+VGRW6rWh2mmKW+w6usaZ
2dGmDwGPoN/Eorqt3bEjhh75rMQqQctqi2tcfpWejCO9xHaccF0kKqsKVAzmNkAZa5ohjji7xhCR
Wlzn7YpYXBib5GTSJOHbe504me17EKAsJl6T2DdBeR6eHOQdnRBw8TDO6oELDMji4fPoCY5Y6UiS
NkjPlwcYlU5g/S1H+SKNGNv8v2jVFlDIuj6fxekZZYy/ardJBmSRPWdu1PM98qQuuH1GMkNF0Gda
an5Y/PN/1zlJPDANGA88GYk/4ZoJ7lJ0wC7Y0vLqwVtdizgs+2WlNLzqHAruOrPHdkvdCATS0ZXR
+z6xyoZw7LyvoLw7/CosM0oNj5i5ysJ6cbTDO97sVzdMuYejGnzvr2uBtaStlG3AECrg8qSB8Gz4
Xa8xvyrxdi7v3S8lNK51eoQdb48bOs28vVeQJlGCfql2TTSoHAyo3iHlAqLj/FHueLkOuENvPb2W
HT1Fn2aGTs2sTZYc7OqqKwIREf1hNH3PX5YxHcIx/pvHfmrm9gtNXpSKAbYtx+TF3cLJIj5ObpK4
TAX/DRCXWS8WmXe24BoV3KEALnxLDFFgEGtLeOyEtKfbfde2sWDnNFhCbaiGu7VIzRiTImcI8gby
MbyueAzpmxyuJSu9Mf9GSimRIVYIa8wWaiJzjFZ6rzmLu/vKFYTVvXtVGnEA/jqBAforhn59DYUK
ywQ2cE76Jeq8KfZLwNk9jTTCQm5OQAl2sWCfHCi+Hjae5yUGjFYasLCNp7nEszyIeHVtJGGb7DwD
i6fPRDx4FHV1o9N30WdsUHzxFR9f9qpnglLRpW10ezpWo7h5WBakio3v1cxcvwGoJZ3f4NKT8oQP
N4xkSPPWlX8Cxk2u1FqNZuyYpSKALeoJr2zKsbinMMHw2DaNKy2//tYtHBQNNU8pn9QnO0buqP68
atOV0ni2l7EuzOZ6BDnwIEl2emzjO+Zg7X4HjVItva2aYwcyRqMAsG61u3nPKDf3uxA2ufnvfGsQ
MLXETIO3GMpuy8SdqzNOJMdmCz5LuD/jrCeRUrfO8R809+B/mNXxjhD5k54xTNVWpKsrnbBDsDXj
dII1jSp5OyEsRunmMPhENY145ofeRSyiovuRivpQHSkl6hUHHYoThtPbqj8kx3bYW1NdesS0UOlq
q0bOCtbQB0PDmQLMgqERNXSYmWXYBp8Z/kTc0JT4VHue4JKtQPPv6TVB/BCCqIJltWBZ9uRFTOaT
SPtjfUcLvHnSVgQ7dTLn2K3PWqRurlCDWLcY3XSxjpWuaV94mw8MVwivO6GPgtynvMEZjSk3TM2I
Gc+0tqXojRwcHw0eYqS/1xEQJSYO+4X62vuYXT7ha+MD2wBsTxI3A7QxE3XHjtPUgMZ1uIRqsL6u
PbDvh0EOYt5CKhHfniw+ccGm6m3FWzWJK3jmj8gb95zP1LEGo4eWBuB+emcjBPnMgL/XZT9Gy74E
ulvwomP9tibqbX2Wls9IpKDsNZXRdlsM6INuBI3WpJihGal+E4Djbvx2pCgIBK7F9GHCbjobxZf4
P8DNCbu8jWFqlgS7tTi7bD63ZJZEHXR+PMyzjPgEAaP+JpD6+F5cEtuFp3mnKie59D/SB0m350jI
tSFbDJbAztm7jAq9HQeShQuznUsflBEx44U+zo/0lq922k7e17sXh7lx/xDndWcvJduGszknZ+e0
WuA+1w0SfUpWKmJQFFK3MmEzd3fyROR194VI5IvugFPQPNqgjP/bpVDdsYIXGOhJ/TKGC2kAM3Qu
upFlmO4zkZ4mfzV1DCv96satBKHK06+R9FysKEeMGnB+iaa+zJZb3PnAuAvKHJijfMxHTNBTQWY7
6wlUUKYvPdzycJY+TXFusqXtCipS83/9tphoc2+W9mBUpCV/4P9dDNT5bWcIP11iFHGOgHwlNm+r
ZBcHY7fcVZfD5ZuJseSrVMQptLHm9ed8UypcIDDr9ni6wvV+0S5+pu13whB+mUFQNlTrN/rnWBcW
ZFAF3Y02NFMA6F2CKdn4WlODr+ILfVrR8mcNzXRXJJ6N5y7Dl8GOK2WkaJLlxfWPsHwVUuaGZE7+
tGTA9VM7LwLMjF8+xn0P81uJdY4i54yjxbKj3t11w4/eLKQOpW4XoD06opOHFRwtN73HZdTNhkjj
AIEViCyihAH2mcmd7JsOOxLSQPxmCIC3Rfdora0KCsvV6Rpx57c7AwoH8pCghZ6bZT8mN918x7lA
mW1OvNMwG2XHuKuL8JwKuX/n2mRhYel9QoKkSrU4bNLDWkoi8Tu8+fXlLryXjArJjY8eGykJxozS
WGxdI1wvhPu/UoaEuu+5yvB1jKX85MAhXu9ihg6t8vamzvRH4DNBm87NSCh81B0RgWyQufHqDN9o
J060e+QZ0QojnDZm/KAH6kWKfqta156Mu9MXqql6AGkRJ/woukp//yXIh5+GtHitDKoc4sNMaJKK
BmOPiW33mUPxAcGYjqvg6uKM5xAaaOTMXUXH4F3SQ3VnJQb3ZhdhCGthDeJ31DOeMiTDFvVKN6Xu
1pWrlGzZVne0TdyeleubaXnN1qsZKsd4hdKEKJELZDidedAs8PSmc6CaSScA0x8PiTOAH+WcWJfA
6WloZAGd20vgu2l4dlaUc9WWhaXHkiMtBW+VbqeauERT/ksQ2XNMaHtV4BFsM2KSMfFiaQJZqjzK
iR5wwrWel9snWOM+Fub9FGNtscJmzfUr2zwIGZ1xoU1qmitIku6t9jjWb6Pvm3YtSTWu4GJzXE6A
HEc2bJU1BQ48MDKgB8CAzZgf4lB8fNbez+H5kteaKE/MtE2L8v1ipUoNUf4Jj/9NUmggBCq2PXbk
KHjCBq0dx4giY4XrAs0UGZFJ8YlhA+lb6cd72jfXborpHvAqTWQYra4wLpEBgTI+U+zYJPUtoWoW
3RDH5/9W7p/SpbGvVV55VN03w/5hCCdmmlm0mwyqbzjn+yti61tW5HzuzBcxy5oSAXFBXTX40uvy
xEBVTZSURGiyoYr/om1K0pK+Va6ydCj5HnlqyxOs2Xe36w8LjqJ6311SQEqbsVDqsf+EVgbcDKEe
D64FuLQkT4lnCisoaCUcCd2yc5HroeKFtNnSI+Ano+8dj79AKwTZ48Mc1Id1iK0ciy5RLAd0own3
xGQdIyMUxRPSh8y+XuaVfljqgBoqJkKjLB8KKFAfLivAv4EY7teNnJa7/S48dST2ENE3/NnggTeT
u6IkCOXJ/iE1cGO0lfMrfcU6DqxnTULOmsyNu01cqoDeSbvUt269smeAtP6pcTBX7l5m/fHF99UJ
UYL9AauLTViiWmyath1RNfLdIY7JaXrnD7v+AFoqczGxr5+IspwA2rMyDUqLEaZKNIWsiXxVqZgg
AlFjxJck5wZE98tiCJcL1E/MeBU4qRzTMwX5hTVUsRA3bBGKvcjIAhjeMLA7IFIPPhdYOQw4nHkn
kgqEjN7TiVPStOvV6tPu/sjfA6BsymGDxOhfr9Vo3KwZpmshL+BY7lZusWN+0MtYGUpJX7s9GInR
X98oa3lnuXrucsKD0uF8ZBudDBzCLbXduzGxRYld268npLMQLeh4MDOv+Wi1DbyYMzN27wzBVm3b
OmgzohtA1R2P1L/K1Bp5xLqBBav/wDhBwmTWDHzalEsL9PTx20D8OcUiLR3W6+VZ8Kw6jjWYKx8p
CFYQAPzS9ufb1C5fiPdByfneh8Br2TlMkgdnmuhi1JdfzJyemHJtxi/RMK0xs5UHJlQiHdPYdfQH
/V6v6Pv5oL5qOXRjsjDvmlaU6LoV5S/ek9thqJKi5ZDPrqZwJ+Gci9HRdL8Bcz9Lktdpb7Nep0mB
JRmV5eErYd7MwLpdzWzSIN18CBjWbomW3Yf0VDrfJlgytAMt2MrQ04PVgAwRz9VmKIi9bO387eBk
FuHMUzolruyteWjr1fYDtWrt7OzUsMOSB49E4WjhLoyFF3gtDzAZbptJXFXqCjOZaOV7bwvCA/ie
CeQqgf8XkWBgvXOxtADvX93estyEmvhl6tf9Hq0X/O5KHOT6XFeUawQ0/nwC2HCqGfNiI0QB4h4o
bJZS3B9+DQLrovvol93wMpLD/EswSyETGUwncw4Vxw5Z2cq1/Sg9DXbx2lsX8FsZwCqCDll2WWrd
XpZZWTgqeKZfrgBNKYR66ONte2PH/8VmRUU1LI1kI63ICnI369gb1ABkTyysdr1NQOWYLO6mW48i
H4Ok60s6cPogkoB7ZBhYvWBlf4LfU3lZBZeENFsLM6vx1nSLCScOlv3KDKMqNGCQ4HnS0QGrSico
5CmVzS1ygr1Wod5/J63sYJVhDAT0T+SA7wa0h51sP9QdsSGWM+B16qlizbgvrBtCvawA7II95mHg
OsZJ84ixsyICnUQ1AkXQC9gweUM8zy5Ww+suPkyfRtwzcXuNtjSR/Uy6ZxXqK9BoOJFJOQBlKASO
VTOcM39/V+vyBlUhzLU9LoGNpcs273R4Z3hebehS0BVdbQetA8oztxt2SG/OMQE+P62dS64f1noT
S/+0MN4PszRC/j6DxwmTVTI3FPwrJUldYdUbk4o9b6nqZ66NvL1iUTiwKBHdsoPTFfEKyQ9iTUul
fRhKtAsPDJXVlV4qKxvk6jAlQSqA3UJC7c2bS0o2JDYazX6QCWzdZKrlWhxjXE/RAxNZEMkW9dd0
+wCE/nHZpiGJ9jLwfHI1N169Xx3glV0VFVYTwJq7HhFtGsFwn6oOb5wkL+ymfNzGGZYg0ZxL3FJ3
OX662WnPiF2rb/JiGv6G8+rTKdlaK4mpKZiQ8torWbbR99hYHtdtFqb8OhE1Fn5jeiID7e2hHXk1
LuhZWfdEExekRJkEY3djZF7Let1ocRtbYH4BM4+xxxqBWqQAAQbhBB7GUroTSZCALrAyMIfO1bce
xBri1fOSYcBWYg5/Db7YXTDWivSOs4sF6ciI4GSxcR6IIGx03Jzdw1H6vNkVYUdZYCr9klivW8FQ
LiJ5Rww/UV0nCX614xITCcFpnY2ZSk5OhOuCc4w8iYcqk+AO4YzOcr6llndSiibwndl1KpWNDlKy
9v6ofmdYa7Cb1ilptSW/HfHYsH4uIvfkaP4OYoy5uMZOXAjzs1RnxnTwi5aSNUJ0OpkEbLl9ol3X
YbKl3NPBr18jWQSBNKZpVpd4a8quL74ALKcBKvqyGlDwzOMnYQf42cZWid2V/Y1uWv/D58k447RZ
w0Jia1vNuM0LQpQU2JO+Qbo81FUPiwq979Alll1MfVLt+UYLRgEE6LZZapIX/BRiOYHxiwejcuLG
vXw4ofIf+akh4hQsmUGQ1ir+YEG7KZxpueLQus6Aetkmy/Tg2lNvS5FYN6q8sO0OUpmRPR6taash
B90bsNakzDFhT0rFmG8UP9zLgPmpi8nknFRti0bgtqS6MW+areSF3QEUFVybG8y++nyAFDwDiXYC
vAMv8cGxjQhfOxywA5fh8CUnG3n3dMnD46G93Dd5az77jMrlvFJKoZjhKFHINGkgaMhalfdgxcCl
9IuiT18nailyFuoq1LdShqS0Y/PnIRm/eMGguRrJKf16j8QjPRl0+x7BTPQNc8vpOzChV/pp8ixu
IIHsHYl9G6m4C7eEx7XnkChCrrDeRlv64DRH/cV6U8L2bXM/Vf8HISLQBVm81wL89lAAIpQR5ODY
aJXYzjMwdT2Qv74v5nwz2mq4uOmSFHUnyjU7YmxtJydWmWKg4etC+CaUnwpPjKxYDfCYChYCz2Na
TiNwJBXNDMSSGjGA4Nvg6L9RBdC2vs/GE//P0CM5DXgeaNcYND99CRGCetTMobncdSI0JZLUwfgj
O7fx8gfh6z6ZidFyBGfOOYO7BWUWx6ZDCq8kyTf360efsT9DmbSYaYKJQ7qa/Ymtgonxz5JBnjGq
ulXo7rdzFXiwL/z60U+4VVLq70ts0K+RMxT4YSRmWmBW+Ivyg/XoxWgCDCcrxGzyuuCu7aWo5u2v
EtaCfRTFT9pdK3Cl4DRwPTOp8slGXwKznp9vK+zXV6WzWtWTwCl/RpTBZ6MWUpWPB7aP3hhVjnhN
mRZXrYB0rhd+CrX/6ssN1YeB3Ys0oLUOgv767gGuUmaO7V8EY9YZIygaw6dyFDlYMAXFnC9fYSQi
/ANc2ESc3zH4VwWGXmX+Tkl2c/lnY8/yzwYf4bl7+vTqI6VwjWCAza8mnO+7xtBKurRh+BZYNkvU
R5uQ7uOXsVkj2Lh9JQ088yJzUs32nRXm4X9UoG247tOC9oG1CoPiRkGebl94a1RCfTLMGu0DdURN
iSL6ehEpkJCxYfFGRKHJ3JSMJ4E0jc6/yUA/l0/dIuTqHN34sKhD2ZAgRs8Ql/PyTIwgYEVX28Ju
+aqQTs7wNjqL6iPKWGPVEDSamFOAJHOl09r4eu6JcglzYzpgZJR7CioPgN/FY4yc03vuThmo8+0M
xNUDoKUGQfMLmBeRiZNhpNWxocePWd3jlG6rLT07FYt3WLTTiXLEqSG2h6D1zQlrrUEindFQhnsV
KkF9Qj3H5owFHjBil1+zMtwxV4MtlxaI7VojpkuhLrpLaK7MPCZppuoQhipIQnHl8WqdM38G69Mv
K7zVECU9R5xNVF2ha/3eZhBOlBfuGGS7UFTD1qfCN2ZCMUeuiDOYnPuiy3bwEr6rMRBKXHGHrpVi
+OAd7nv457YElWZH2aAQQfqLjyj3iqQZVIUI+t+4yrLIAapvKqooghfq4h5ju9p29pphiXiFI6Jf
hz2r572eWMu7IOpvtyiA0oERtLz+JxU35uagyTFUMl/kdhOimu3NNWOfTN+sT1qjipvw/YduZaSa
Sj76UdBYJ0gmGGouIzJHdSbhXdGKwKNlEDTiJb5Ly4vPRzAhmkQzF5aIvsvNbs8XNi9XVbDsb9q+
6qQ91hwPXhoEouz/yn1fR8Of/gL0Ojjw+2qEa5Ng77ewDLRI3ZJmH+548CaY2OkzzEI7Bb22/CyU
1yp0AQIApIGz9lqpI0jyov15za6DFlmsz9IQFGRaIV07IxmekG0B3eYEyC+s1+TvgOcGceE72TDN
zufPX/nloY/HOE2bcggfe6Jol+/Vmxcv6AiWg4IshyfLg2DyVZnSCvuSJZvDBq8akcOYFuSS2eyN
PiBWF4T94Tn6Q5syw0C5v4kktsAzQ8k0c8RnEPLD5Wl5QKqBf7EnOBVHrisvfKnKfEHEQizOfI+7
fzbDNG8295j3vC5lk0vnigH9WS+n5poSaqSuOhOzEtoXmkQje+nzV2aQ7vaEzw7uJQK6CDO6E9Wy
HVKwThEaU+j7jLHmRmz29c7EmOKHeli75769P3HkXTb1OpSXB0FrygD0Uz+liGenhxgMgQjiz+rB
J5SKx9ccd6Y6PrDm/vQ2BmMUsP/pcd2Ryfq/jwXmS5b67lfTQ4FGEBq0JbYK1+B91odYpIr32hGN
u1RJl3xmdXzJR3QY+5l5JuXZbi2lEAzwKUkVct5MfzqcOyIezkTfFvIsfamnj29cQbY8FmVtWveD
KeXfbGyVUkBm9K+hr2yc3cGH2YgCHBECe8LNGo/P/l420nglVGEFBGoPQpdfGMsNXFpiwtVmfXtT
QEymFB1h82OcvlajHKfOBNnIbPJhu93ckNwr1n/czo4a4e1xoheQ27D4g/mctYQIvMF7XR0vvazT
nSZTey1rkNUo48rW89hLFf9Vqom1m41/f43KxgyDBCTt0FBYcB8KmTIoEDsN2u94lNcGTV6nTIg4
DlA8Z1RJAAMG6+zh8gquv2D4RQfrfJHKZNplSAsn9Ev0R2Bx1ReemEiCBb/YzSXkAOaTFbZqGICD
iYAdONlotIdLRr5Y6MxT0mMAlnsP7d6j60Ix7zbWd99TUBOpqpxMSzyHzCLICORVgUzsmJmfs6ty
fa1MueEkyas9YhD0HpARRTxJcIlQhKKOo4zAHLdfCTOsWkYBfQFM/kZJpoLekbwAjnVpvSEyCX8C
ktG8QBnOR6W6BDJ2sEIdGE8WowMzuyRkEr3Oh/qS1PU8RptBH2XT1WLapjpjAeYadf+3GNEKymDw
w3HDXbE18sA1JMccU5RIdkRe+lzA97sSXxHIVDovTD1HVNtlITnS9hhfN42I21eVPO//E85cbUWT
G63Jk2w/wo/zvrfr9/eX0NKsL+KhcIVOOeP5YFWgLJZQZ625Dzk4gegdOgSledoQ9rs9d41rmZ0a
7lUKHoEXxBEF2ioNii0rdNVgCDu99y44ME8Egf1PpuDlYg+13KGduLz97Ed/EmFb8C951Q/0ngSB
A2hHTNtBAuwPwjLiCnZ4bXddfiYo0nOZB3RV/5Q1ZkwLQCh8LUXQd0V6s0/+9qL2qkoQU4PZNkK9
9S8V96te13vMw0ujTtotC8VW4UiIBAFQla6t2j/6WRAbwWmm0QYIkLICCTdRr9SQppHfBvLdSgh7
bVsaxIPQchTGwVDvpT23fflG44BVlFmweDpM/RDBXa5a+qVOQyYuJegZsv8mHJGG6zvB7YMiDLbe
qKy+D53QYGFj+a4sfUv7juAIUGC3WU1tgS+gXvbkA5ujy2L5RFZqvevlMfNvabpDPuEvbWteYiZ8
RB/iEWm9dZrd3UFHvVgqNlJT/EzX1MPKsGfDGf6BGmIqtV74JwetXJuYXgVW5Y/cWGnlljrkb9Us
THpsyx9LprVBaQjqQqVqL8Kjkc7Asog1sNv3GT0RtCuEzNq/OfHPAtNdqSsGmVyZUyLsSdzsncTP
4TL7qN7VmCZvPR59NCTEKPgoPr4mYYk0sVOHoYxbkfAVQ5OewvJPwR25bWx9eO3D6KoODgQJUj0y
rBRABFEzJTekiucWEiPmfTTb4QxvxeWLVLvO4zlPwQas/fPKD1hO+LOTyFh0rKEZ4m1V+uhjQg1C
dH/W9HjEF1JRO9FISAdOIqFMIlfpLoHSlJvuzBR6tijpfBNH0pxKYmZWZei2Xts5WvNbHNr30mT5
BDaEtKHWjKeZZMX9tvg9uiRySZ7+j7m0FdoZ9lZpP3Cdq40RAWh6dHpXI3wdz4XJ4NZ/cWIoWf87
Gj+PBJBj0iaJzSSjVlop4687RlUWJ+uzVnaEmQZb3y7cgfBuhjJUs8B44MtkaDcvRhztbwI9/Lqf
hIChlxpVGw7izfrJxm6E8JS/EdfoOTFIknuqC27/ozl7naqgQMgXfsWkQ/P2llJXXMG2+nAiVE7H
gg78pdqE7aqvENXtcsh23hrMUfsAMrGuvnCBIQhqRTd3urfO5KfQQ9n6NXt5oxX7K8zwB5aC8dUe
rReY8cAGwiEyR1YngZZPPFAmmi7gb6oKMWZ9Gcejuyt0yxxDyZIYlyMY6Ll+7H6WbTIq3f1CxbIF
DFBs8AG3hYliyzo+KQI8z6WlGHqqnjnj7eSjiabN/MMrc8svEbEBCc+MXlwZP4Ro/6ioZ0OtS6Ha
sM1HOBEFvBoc2upbuHH6Ol1myO6zM45oVKSCnIGqD6l3sXiymyhTlmmJDmpVTb9hgjUGbs8f330t
NEITfwC+VwsThLklwCZCmbzTdmcrGSD6yS3bAEo/JB+O1PtWuyyUz0PigkLCQ704VoDJB6uZ7jI0
tRKwTc+ILCgTuBtnlgL0K+VIK8fHZkLThC26Tfq6GwVJUYySTNanwlwlvdMOj0EzpXdlMQ1pZMhm
UJVz+AKB0+NDNgglHC7HRYhQwcDM3aM6ENAhgBwQClsnWgSCT0e/7hTzsCdT2W8hogzXpL838ozu
JihGPfgqCyHpb/dHUMT6QUY/uqB0mVbIuD8+oggssr+tRZlsEKD3TCFPBdldaY0mfDqLmnOxFXq9
M0Ip5OE8tXj7emlJMccTwaI5g9n+HbFBzvihoAA+J7BCeUQms01VpDPyAqyLXRoyJN68R5EZ33AN
Uu2w0OmOE+bm4t4BOgatJrov16XWSW135x4lW85Zi0BH6KgqWCjhf2xkh8F4YgYBJgZdEA40N4pt
dz63FpJ5Mh+rmkVo7Ch78DQngQa9u28EyuQCx78H1Bsc9EpqFSutxdlWInJ1CgA/aud1i1nbjAAk
quJMzK7Rn4t1BkY3pifxTjXKOWXk1cyeYhjgLXvG1ZkDQ1P3XGY0hRhP5dbhSrNf8ADItGTihY/p
gTEzlnPr97iZVMSQ3H5YR2PPr4FTzGH+dO60WLnp8fjM0T/1BfULQCmGz/SS6xiOQDhjbTNzKjVK
VloeoqXxiUvo9fxaxj9EgWF4uIUnAegrz3JxiIxAdDqoEzRUpaAISyQ26rqc8XHkW4sXElNgyL9s
nVkYMrRH8EamHWWnk29aKE8LuCgiM+jpFz4JxtiTzJtotgdOYaI2zuYomSY1VwT3zXBaFj5ifbbm
HMaL96qdHvwYQhob01hUeuHX0c1vQSMSV3U5XK9kmo/M2nDvzMXImP2xKofpebCEkvIXHkn1BVNz
SvpTbzLPd5V0r6zC1V/XAjcoeuri8zouUAHGEChRb5HMs5vLzW/laXKaXV09Lb6cQGdZUtHLgaMR
j53Vi3ohqv8wl4m57s+cxSEMafI2PSazyzh+iMKFM/TsCTVi1bwTO11B6cWJpdv2fxcInJicreTB
Kf+sQ8iZHCdB5kVpblAnniaUTD7NJO/gNFYEheiPmPQQtGM+n+K5wDIgMESQbJ501w1Ph7PlzuKx
zW2JYNrqxtCwRF6KrAryy23I9bVJz+MqUpzaory9bIPsIU8qvd7mOwhT3jrpnloAAZbBFurfYL/k
iZeIUVRHP4ZTe+OvOaIfmOt2bmnembulmkJXgzwbnqZAPq8+JwnOzX6xLAsqHEh/nwKw8N2slWCb
BqoLQsiOPTcFW85adR5C1WhwGLRNKNqxHcUF0L5YzggjJkHyGLeJ5ZI52Gpjl9SRDEgnw683BVCc
0yPhDP8vQ/ZU/AbTw+d7YN/G0T+3ePV2C4GebkGNXy0ajrPi9M6djJ5aQkroUsIB7FvWO/gsk0dd
6r9SqJVZ26dDE73KEVlJ39y0sloqhj0NarzwAQmrouSetfkn/ViPAVDVcHkD7cWqOIwgA4Ca8qdL
uTpjnu8uGxMhQIm5DIdbkT6HKa/ErgAkv2V7F4qtrpOMNMRZZiJKB1/eJMByUit4vaV5fz/EygJw
qFF+NOnuDMwtFCr63e9tt/ol+SGpF12pSmNEbCKdthczi7aiCdLjl6TJRP7tsGpurIifw04wAoH3
QIHnPPGXTqiEL/jpHwn247UPhOChYp616XSga6kZRr0Vm6JNBbn4RpbCSnG9S13uphrfgjGG0l6N
aJjhJR6LdD0jAklQ8Re6SKdFSzCRI+Dw35ACH87Yl0+f8sc4dIqwGc4ZIHPIQVV0ziKZkQTzIO6z
t3Qaaw3Z6TRbooTzukczY1eTO0oiC+wn8NWHQ5H+lDyf6yxOR7o+aNYDWxSm8Y2x7tLWnykYMoRf
O7dRYnXf8rAt4AyBnyzdNznnOQ/uA4fNlo6dwWMgg3efTztsRb8rxzOaXOg0z3ChOte9h0IEQnrO
WOIJEZD5+k3m1yMz8f0BIftP25BScAt2IJwAlVUdC3UH0w6Que8TCzUxMKufTzwG0ywnyeWVhngL
rsK4cZstVq5Nze/1+4K1/4g1NNlDhPdK306Um90xBURWC2RBaDoWqhnq3X6Q7nK5P09dy2ZH3PSa
3309/h1IgVytKROoh+i7xOil8xkatPzH/P/nBnCLZGJGUJkepmkv1NNtLo91/o9yNTAKL215w6hw
PdBE21etZc8A9ewWY7NHdkvraxO+Vi4Mf+CL14enu+jieCV4Lo2bWNrE+wQpcgJEz0xRAE6dVhp5
DSUU+mWRn8QJo3iAw7BGPD55g9NFOjK99r1WxMPLKA52eqC2x1pDF3tXLucQVeFaQb6wepaL7CwV
7Y4q0poeEX9O6I4kkvFl4kv3MF/4vJdeZQpmHPr5PHhwqCrgaUz7+1NkIclpWbayy2EZLWts9FSU
vE4kcHcasfwBb8Fd7ACFaq/9tIhmCzHYwMNAkmtpf0jRLfaoDddIgO3334DNOMWQBu+j/PucBU+t
mecky9aXC4bNd/5yzPJyFV0thyop0S2M7LkMc6E2cTSx2f9P8U5bhb+9OnNaU6li2TwYyxMpZIXX
XwkErQdxDvqK2DOuYdJ+ijtBm1B7BVGj8RVAAeSGrm+gEbp47q4jt1J9nm+soHKM9GlMEbAWuHuJ
QZ3QhTRUpuCd5XT7KKMZsTgvQGz27Lertz4FHnnsQQpYRH69XpuIa8yHzl43qJ8snNRPjIKIErLM
lyof1wbtDqjyjlzQ8m8t2tDbfjDTmwW732E5+DTZ4yevGvDEdLAU/o9w3c8XLQK1YP1+pP56y+dP
YccC/G7kgA0aVlc/hUb8Z8mcwaSh15lmD8iNtBYgjedYld1zsqCzt2OnGv+rRfZyl+7xzqZbht2h
LQS/dewMwyp+irF/HZtr9DSF5tpgt9QtYkAMlUo4he7dLG38C9DY3MB9O63jbKdKBDkDj329PyzK
tmDrnlsLdCEqjouhFXWEnfwdlF4VDQtv5Pp69dI7WxXO2wSRP4BQOsfzxwm3rn6d0r5gLfKyvNE7
2mL2Rr0fPINSpAeM84xd2bkVGcoWfWvjvlLCQm/pY1oey0MBmc4FC2b/WU6O89A8NbSZYDWXz1ub
a0pURdXM/cxS+lVhh+zRRgPvZ9E6E0WRw+q15UkneWHqMfmw0Co6RWJQXWk3puB4hDuxqxc9Pzdd
owtKM818S75cZH2RllAegU3QOc0rYbrAKgib3wXhNmDz+UtKiq6PkS4CuPeyRuaKzUBUY9iOsg5J
rSfBHZQXKevSY076M0DvR7AfVuPulP+tzZtiE5mIaTXIdcCX8ap6SOYtsaeonbcV/AKqffa33IEg
eYLWbjzNUGoCIi6vze95Uv/zVoKubCeWwObpmIAi1KmiFllvufzQNqY1wQTkyi0meR3njBwK4AQV
iejAYaR57v2PVHlBBCjdGcEbagcAUkRRBynwN4MmSHYWUH4WWMUjr1ojZJx5acdEFHa1tBAiZHx6
YASRkswpD2tjv3yyUWx5VOGdgCA+SI1HAFQNR7yriLYJuCiOw8ew9QEZn5NROjxnyPr9gd9gnKv3
2GaEnNTzVU3C0W+1ccKL+g2PmeHYnbkbupXs4BHHeKr+hldLULvOuOPIuJxdrcoi347uoz/TyowO
MwlmDCVBlX95iQxS1ND6It5sboAg2893JCyO5FtE8W+PEUKeYRG5QsrWrIB18k0umElbYYaDeFgs
fYhbdQIp+aTbGn7kjSblVR0FWqOMD+CbNuNbjXn5+5H6Yk93KeQM3TGrgVY+g5B2k2YASroC83f3
uaTcB3J9bwCztYyOWI/7SJGL7ZNOyFAj3DgFc3J6MPOVbkduTy06NvpLuIhlBmFTW4ItOslZra2n
zh6MKFw55prKy7g+/ddqHx0e5OAJi+TzV301aFltw73k3aTsdeCn8IjXx+JA+MyChEPY5MlX1rfi
vJvtcCH5GYZwUlQMDSLCjwd5BixoVwuBOhHKc6m5uucWHmzLQMQwPK0/HSc+cogPrlOEAVw1erKe
1BMDO9uWpYYzeOUJxs8dq0CysZlPPJeGBeL32elwrUxIwdlulbNxnS1Hu1xc9Km81eFywjI6QUmW
9ro7nWtf4hRrjcdITFgxMiQUw3s9fEV5DnDbmfcdgvmJnpmKH7l2gmFsHvskjlJmi8uS6WwnLGII
lXoZayy/EnBJ47NOYdEGObX+QKD7w8b0NmDffhfCiijm/vmAba4bh/vnzFZpjWOK2d170i2Zokvc
3zIOm7GGX4rPIDab45rDlnlwvFU1Pm3QZn5pK2LWgAxbRnApTZ1gd11FZFnJBRrmB6qkAMynjnCd
ogfaFZx/AO/IPGwVEKRJpLzscYq84wDABc9pm99WV0Y3lNHKGgrwC1jYCRPx9LYFe0o808P/CVEt
VRHvQVicQzHbwu1GvjAms/bbHwWA/q0kk1V+qa16zGjeHCIa8Vy/belCPKbtFpJlGACTJsYJpRsE
Sxvmkqd6yPYIE8gSeWzid7/QqqBTdg6vW8Io8jhUR3C+38MLWaJE4cDXyzFUGibXskU7TPWft1cn
MGmLml3jr5CTk00f7JDZ5Pv7TZyQ/OLZ/+4tN+sMZci0MhIsR+nQons2sAwvvS7igrSMNHKoy2F9
HT3vsJjTeavKg1G0QWjz2OIIn5skrZqtD7GCsSnQuEUqIexfNUOyfzbIfUh3lrUSmvqar2P6TnG1
wAla1m9FbiJrMu14HYpi0mBCfWi3VAy+/9Rk3Nl1kPWeMmp7pI8yyqryNFdi1wUdTZDi2e3IZWZm
+HhmGfczuAD1esPka8X/yIUaLpqRky3hUnN4fJV9I/hstvJkth6shzEgeL29LkYerUdVi2R9jLHY
WsdraU5atVPS2bCO6AsFQpBRusHGWv1oSE4q2MRshbbuh38/oCI/uVySFsGfwIzzbFYCStuHDgHk
alQv2ZNZEGeIDZD43+sXNvvWZ/wqwGqaveXh5rtHMZ8QSsANaanaWyRnDcL37YQ5HEE/XixvoTwA
vpnlMD3s5bJwOyHFMkD9h0o+nZGakz2BBINyEwBdTOZKnzgaFceBFKHB7vgW0a+jR22aevGeQr5X
Ll36cAZhZoQaZE5W29KwNmh4nEgDSSMgSLHKQb49FwgK8qrLlgrfnnPneCmasrYM0Z5boGkGmRTu
vMXlYCBuvVXrVcSJ9K/UQY0RmSb/0ioLkUXMDkl4in5Jm7snHq2NhUT9r+MS1aqI23xUTxLioQJh
wW1xFz3/9gs82DyAPNuLeciVOQnVUpGCFZhTvik9Jv5I/vFl0sEitzmxCkk1wCTNMHyDk1uA0lx+
pJQFuzpjoJFZyLVz1Xx0PjaS0VWefjsY5Rf7BLgIAvwxyMB4oZUVad++xlzqudOnuVU4i9uFAoLm
1hxwU948u1lsrbXWn6rXH4sgq/S0HQX6rWj+kuPLDihjaZXwuZGmqBxV9+kXt56PZjD10FTXwAuJ
U/R3U8mcmE7jRfNwJhwvZdokncpbZmZCBSAateWDpdPMJoxeq5d/Vx7tNIDhk6On46Sgni6sAJHG
MyUV+bsFEui+FAjm6Daxdxefdl+vMYqlxJlcZxjY5W2OscH/YvC7VJ1eGCuD5YruloSKN4P6hW9g
Cpzyurs5Lk66zBut5JU0107jYG+1i0B1VGkHMFOj5H71jOOiH9dXSIUCaz6AzBYy23FD4w6O6APs
jFobvGs7aqLa8AUa9DxkZ5Bjzboir0CVJXzIRx7t9wSjJaGaMtcOFtMuplT/IswdWYPC3muQmXW6
bJ6n1jwz0g3bXze0PfLalhrAuq2RFNFgzs4gQj/KF6mJqUxZLXbimd279wOkc5+4qW4K7ZqEumkl
EXe3JPojKn229c1zRs2CmrBvLuaGYvO2sMDrTiwcJiN5vJcN5U72fSE2q9OBDNYNjCewazEhdqEM
bbXRa9N24GT5QwVrL/GS575Aka2tLTwWze86IMeH2dfc3ybPNSVgedmNlgU4QzqVdVQc4dWRm6Sx
6hoUq69iKqerFvzNbvJPEQOtgw70DqnwxPX7h6C4kvDJTQcefPsfhgC3/3Kf7ERxAVIPHAjTESHD
LIBIv+eJnMAo8Kn7tPlwbziCBo6I/9cnenzL+cMnjv/pEzcNyw1zRE+jVxWRrLPCDH3kMHbmMIPI
N7VoMiKnC0prNVy85k2X6fqMUeuBWhrg2cb++M64cHUFfRKxe0n6dkE2XNdnvvah+s74rYy52p6E
G3ATe/RLgYAQgqATzaqDcTg0Fq5hk6IIu09Swl5WlLkCpuSVDwnOsPJKNV7DSYDROibI86E0L//R
pkXabbod66H7lflImbJmjbg3OXuvvnapAVdv1RRkWdCRxBVZ5Rxzoifl7QiZ1gQhZ2M3tAkau2T5
j49Z460qMcN+YZFdC9B6nmkcq2QXMbRDraCUa/yQLLaNqFHazjmKQAGy+YIBfdBFBQZpAmwtC+ts
xUS0HXAtCSvGejm3K2DSkSEmdKcrVmQ4LvIUaCryo2ZvMOMV6yVDCmJqQkB2/IiIQ/KGkOhGoEp2
KKkifPGEW1UxT/VPNPLbithI5CroNRGepd7B7NYXezJXl1X013SvS/L0t5IcnpfRd7VSuDFZ4FEm
twBsPlDhOwqtVyF29o+qyPkY3N+gPa8frvYt13VOn0KyorDsQKcSXpsTCcQ21ZCcj7xBXzHprSL8
p5DwnMSLXLuuPn4UWheJ0Fuynxfg2JYvCHpU200Yn81FBErcb7L2UQcfWbxxzOqQM6tDAhfTWUj5
U5sh2VUy1Hq0S0awvMD/xA+fyNZXy1aRxBhI2gUK/rpm9qcVdefKk5jRxGeGOUzgjpdPteUlLlqb
Dfr8ORF1i9LxqFgLM29jDE5yU22HpALWyof2+eyV9YV0vvt8v3HY05ITozfHnJusyXMuvkKctjkg
uLGutnuBG/xGFqjPFM2ojRHiPqBiFlxCB7Fh1pNdq0/FMTcEDC6IL5e4x4/xM1gP9VP9O31tGQU2
QyTXGAfSudesKHE5S8jQE2+mbyQT0mxAAfuHscm9C4jTSNSZLCHqdkTcbrSsBNuNJWW7TTB/1ALT
jcS7TO7DRPhT1dxlQyg4Oue/lKa+Lm54NHU3K9Wro0c7eZgRhQSzCipsltwW1ZL8t6xaMPrDpfAP
gr8WNvzXqES6EayiEuNIltsT+v77shXBq9pYLbX/ntjjCyCIBbbFqFrHrplIWQ1ALxv/v1J0uXJq
KIcvyg1DfXvaIEKQuzsXejv9v3updAhN1K65whtNidJIMvS/WADAY27nIPBAFSL6T9AJCymSIIek
41MF+ZbCUtnk2wr98bj76146fhouj5T9IT+ro22mZz3hsR+Zrj7JmpmJfjQSvwvAxHYL1p25VHwS
drDplDLv5BSWlbdjY0SBF8Zzhb6w+HjXGOGHqeSfNomHWm6JyJ1tw+SibzBo7DoPpRNlP0vMhoqU
lRQTzJONEDf73WCRJsB8bU9EWjSm2unfMN7b9uCHsLbk2Cupn55Z6i3ufA2T71FDtpdW2UVkcdDx
L8E7YdAO50kUkCI8ibZDw0CPY3Jq7gmcWh56KZT1/kHWMpT9rid8kwbcG0ekq2Hw/QpI9+HJToR/
Rsoc9ZPradCGxDwLnP963GMVYKx79Paww9GxZGqwZvasHTRPXfHE2ha2GcP8Hj53jt2ImOazWzEc
lGhvdOWpRa+ohAmYHqOVrBtfjoUwAQ5PhY78uo8INazYCxIyNR31+LXOib0zY90ayv+eCB44sdSI
7nuWTnEr7VVDK9xLb182cV6WqT2dTlB8dfw15ej0wVj523U/taZh2ul8ZP9wQWa2BHfsGF3beIXA
NpHzqPRw6C90xOGslRxZUHVmJLsWMqDZoEXM4Jw8mkkSkdUzbMlG9p5rmhH6VJnn57VRQch4OUR/
RBj5D1Hfpax+fsWMLZE7uFfhbNnAWkVFD7THwTtWSQis0r+h40px59S0FQzZYlQ267C0eVs7tJif
AM/9aB2bFxgiDSG5RHQKtqNpehLBdHdyzXMdh0A/oP+0gmETEJr69hDp10/qHoh3P9yAQkeRmKvE
aMIS1/7ZW6JhPbrBddBfhy/FW3C8D7/mE1WF8USHeWq6QfruW+/GnBXCO6OeogLPSjF/3h5x8Wgd
I10EAjWecokihABMBR82hQlYU0AGSHyFBuxXnOpkfO/O1QJCDlm2o1FNIOwcNlW7Pqmyk/LiER+w
SoQ2BojXqL5Llu5+nHSDkEmjMukZlZicGyMjfHWodQyRTM27f5beB8tvDm2vAPrwefoVIugRFHCS
eVQ0jZlSGSPJRmvMDlZKM5vakO1mjdEIGg7kM5i/m1ng4mp9jU+QHOLSCHnqZvh+fZMtKH2W4mzy
O5W4qXT5UhoJGixGbaIc4ZmNGaDBtOw+Pe5KtBgj9C0SsWcurP4pHL8TwYDxLKAnzZ4LkaB0rMDe
DSv6rMbZN4xeIlf3ATyoFIScyaHcynD248agGdBC96JFHdulUADO7khgOB00vXR56vqYc8CcAvAn
y5cIKgTQFUxLMydZXn6mSXgOyGkjh+ReebKhxLiug0nQwVYkfI+vCZehVzb85OE0vfwhWr30fNIJ
57q4A7Szwp/FpFaEEyJ73LRA8hV5soYeaquTp7c6q+Q1x3wci41K3+rK7JrZaAoM5NZsgGr+ar8c
Km1+Fcf0I4XgqVVtaFbg0da3rTFwQuuP9yenrcZZR78g5oOIWQJj2ZD6Kj3QH8qDV1b2MSiPN2Sm
Wy4s+IDkPu/GzRGeN1VbhF1/IJAkZNCQxppJuHDddInU8bgFdg8Ol2z1z9KjHqh5p2Dguvt6cwpm
2c3i/U0TwOQ/UEFmRwgkUseBzcHXlQ4NsxDX8IrwSVuN5q3Uusj/sl1MyCk/8rxY2EfRApU6nnNT
lyADUYCLv5jI4qXPK+iY4uGipua7u5aCpM8n2TbqRchUk/o2OBJqYGn9t67tL63MTqQ7DOZrVv1c
wCiHkLC0ckPu7uLgNQZab5hm1npfeXzu13E16tiyxuIF+wSY+t1ZQB/MHtJUDvwJcXk6E10NJEHc
t97NsQjUreDi4Td21QSoukjw1l3rAzNseuaewWuRLN6qzsy2sKuz7Uem7x9gkTvHSH4fjtF0pnlp
YKKxhkPqVGcJ5dg4sN+GCZJRfQqTKLf4b1ufIw5+CF7NmsXW8q5GhS9CIvclMQF/aOfkSWVI6O/i
hO05X1tKSCeemBesYkJhTF2U8H1cJxRqkUGXJnUl+o/XQASOe5/iF0iFvo859cClwvBat/WWP5FR
/hFFxYSy/vxiJOxSvXM8nkhqIkPm+Ph/vwaM3HtGYyA2IXbDAHF37ptY0OB2gsYL53OAkFC76uDR
fuCbJMMYHRfJQwr6ajxhNSyyyfhvgx9ssb2igiPgvZ8HbOPCYLgI/vHhLP2+9+K8Q1PaAjVCeOXb
NRHUoYZ6pLYTrZ7+uJegv3PVcTPnIAUj4DLmNlcP/Y4oFExK39JZYAzsEj6j/OumzClDoUoThlre
ctGbsebKdHgKuB0Mxj6rKQe97cIG/UaUr7HPcejF0qZ7B8GJ0uI8aM5AzcVXolL9Ki+fDdVfb2Gb
bJDANY5e5bq9N1WT4f4h+AZPpNQCVyJTDH3ifScTAsBhLRqyWpn6a5oWppWBIJGARTXO4CuRWxs0
m7SnbpMUUv18Gv7gOhRhnhL6VW17OWO5yFEGBF6EvPJ47zKkbOqNBhbRrV/IZj6FxnIBqbshciAw
GBZo4Morwk/tCmdhbwpjTb6ypfMnq6IlGo39h7TJfBKal747xpg3JHBEzK2AmlbduZsQBgNGx5Z1
vqrBhbEcRr0jtvArU4EQA6ZWvaaE9JZbkFVOPosxYQeKnguLnbpZu+eVEfbO+rekcRrxLDX562ow
sY/lGv3Ycxaage0VvGD+kGnpBtYfW0aKWAW/d5vS3nulih6lOnAnjWdxTbgHnDNT/nydvUEOtKrm
caYg2p1VcFRbm0gsA1RQuX8Mqc+SRkjjBxrtYLN4DjEgErYpGdEjHjON4+HkSuDhzv+uwrKxHWzh
1XDZT8ABhu6EvP0qI1TVq2gINOi5tlcX7uBEdQqKrO/Rm9TiBBvpr4+/mybQbJin+MNncsbVRO4M
xeO0wXrLfzHIAJc+Skp1pBDBcFsUu3OFyMgk/n6GK60yuyQD8crTKYarhJpp5gRFTsJiFFEiNWrd
hTRiVzyn51LSBtcipUEPn/ZhaMwfZ4hVzP4DL0kSv9wqu6FlMmEsp9YRSh/wEvi9x/OqgZc0B8x3
/Qgab6eyEYo+I4Q10hzpsUABbukJ2gEkiQR8p+LNz5AIkjrMPKl7bpVEJYwr4+ZhFVv2meHS4QyD
9eVPnMV6P5ITEjm3zLBYsNTbXREcynbUUt8OxWBl/wykeCNFLjRZn7uZj7sErjsNgA2vUL1G0P+c
uL8KkRoYqs0G7EG3dv4xNhZbqotRpBWrfhBV9rp1fyfC7cfhDoJpC1O4HKt8tBRIw7tVtiJkUjte
oeB5+jALbHtC+NawdaS3PTUZgmWIlWqH/7p7QLsHXA53NbMk/qD1c6025SHbnqzSUkLswnmRFRJm
DrUjVdSqBVjGVX9thUIlj/nGj34U9C7iuPYGfiRX61RG+oLm238dUnxT/kqaqHHDarBmAuhCRHqY
/TwM51K7wEUc0PUwY2jhgWc98r59wcFLjYvw5HpMpsl7h7H64omRuqebVJ6r1QOsJyzPRGEgxaBw
0vE9jnA+Wi+X7qgcm3HFwoYAuDFQmy1ijxTVO7rlkBZFqEIfnM4MlXD7fU5pP5kZ8FYooU8sbKRq
BbIvK1+89tNuwvoOz8sbVFVHuu6iLyCMfRXndvno9PmuKzKh8UuBOKF1SdX04cNc5sljZDI3EoZz
d6YNUHw8Yx2T1yNCyjfbltD/wJoTcHatAH7r/epqYMQlmlR8B1PxcKE8FFLjx4tao7PTd4kmOvG0
/1RtgfuD6d7IvB/t1p1ZvSZClVeA8fNzoy5KhDI23mrjLyuzitGQiY9dQQLp5pYqPDfq8MHogt3Y
v7FlRRHYevUxyLnzcyUinR2SLZeXFQFq6SO9p6mAq4fINCUcakFS3K88jHZNsiDxmgYVOz+WsD2v
NLYjB9zbsLPygOFhnbcTmUwH15accsgnkRan5Lr0oqgEkIJ/7W/zFL4TS3E6ArmUbWUMp4ZjxSOC
XQ0YKhUQGeoYkOSTnvKxsgeNcSJBkX7x+IhW/lleAe+NTPmlMxkPPOtGrrY2NPJatFSKrk2Ie/Cj
b6pniV4y36isBtwCNCpcXZnrBIfNOQhmVW2oU5crmYIdGEYdyXVjDJr4biK+xA/zLTI34Y3y6VvF
wbmMEmf9Wk32BI0DC+6QKiZhd38B57h1bJdbe/8O/+tH2w4Odo8LEI1ARcP6ElJm44cGrAVm0tMw
Nyaki6NRM9pQA1ZXIEqPUaTBFljdROpkBqVUa5U//pdRjNrPa65SIeeSp0wyjqCY0gFCK56Awl98
UPEYXQT1orE6xF5quZCYd6mereA9z7Q0SeudYP9rSozLK3/WEMX6u4hRvSbNXa4BMltMga3V5pwJ
voqWaFNMBhVnQVxuyZs0WRkX3tWZXXslXZvC4kvaxesUyATYRhc+UF78s7tz3/LsxaBbC2Q/pCtQ
uOYf+ze3cD/3jdbsv2UCFwFbCNQmsCptfGFxfv91PATfjC6z+/xKzB2si+gjowrIM2Ph620LL78x
c/uWhKZxjzQvs+InsfOHqYz/i5lPDb0DsgquBsbaT0XtNJXw+Ow2OqPXSI/AHRl3vJaTwfz9m3zQ
NMflkQkCI0IXU+S0+rrAmzqh5bddpf13Iva70SZvFKJb58m2Ao+obU/e5h0sEl9q94ybXhHuFv3s
h93k5Nj50MKitCg5PZBk3SOoJ9CFsNykwxMcsChBe4udnRI3ETZtKyJuA/m19FsNn12D9RxQA3gS
MTuIIk4wVePHs9H4Pkd8PacA+5wvfWNGYygWKiebUmicUVMIuUEx9q6c41sU/QlfwjtVGEsyPZ8/
TYTuhF03xKf0uY/Anx/FaTbMESL0r0eF/nEwM9BTy9hTrqfYDik0D+aVqb9I4vdrR79/6eTfnJEH
P3aycutL1bncUiE5wPxk0vtr+yUtkaG6LFbrtchZTUb6NWLHrhotMGyyBs/UwPaosQ4m3h/BbRcJ
yCWIsBBz4US69h0wMWtChBiokcJ+UIBdPpb+C9yOM7kPEMEtT/g/Mi/A6Qwgpb7o7S061Ux4V7/o
Yj6SeqIMaCMLuKPMZhFTjKiAaODtFtwq+mEEQZGXxDbm6oWsk0oOQi7snJ7xtg0VOs9LPFPZxTSj
YCL6RPm47znrLl5fsgl32RIDb/uXuMvE67S1FQ5I9YvYOOiRd1T7vtazL4XtjoahyWRlLjjowygk
4thwSgzUxSKRatTqhsrln2KCy41/Ssjora7rYiPHJee2P6iErtzqpg1X3mlIyFBFUDi57b13KiLA
FSMODi+WvwCK3Y/c8wAAgzdOGFX0/9bfMgasWQDILo5YbFVFwNQC2225dsjNLb54JyRUaxzdj8Ik
7Vc9xuPn8XQDf2Ms+Qm1WKarzBJ+TyVWTk7FnFbS1F+iAhTQQO/bky4Nb2DU3E9fuHdIuKQsCDHX
XKreFA5dDzGw1Nt/MtjCmbC9PNk5xjpiFJ1aJyCrbaM4SF2YP9W5L16GeKwLShn2MuORCIbTe7ho
m3ny+BPgfkGhEKUVxHafWvjAqIv+VDhsnhFV1lVRlEIbsCKHotajUU4AFDrXyMHSIrmyDA5vfaO8
GVVYbW3aLO0oFHt9NjwCHgq2TYEwZsdYuTxFj0u9Ncby0uqQRhVeqieJjG98IONmn6XPIpTqilRU
zWHsREkghRAlmyjT1zXI6K6bieUOzTCE0kmb2I11roms+kj9+Zq/zT+8JNTgL7c6Iwmm/SyyuY82
ycBWAEKf4kljVX5o82ffjLFf2OLchUyXRXDTlS3YNyB1MDRO3wDB3Y7uoZ4Ct1eCTPIrqbm0v4fg
G+vblb8xsik3eI+DUYro23aYRk4r+TY5gOsHK4TsefC0jpIarMVXLCaDrka7of782Q/oOwA3Ns1D
ZjdVBdixoPuAZzjyUVwJ/z2Py2sqz8Y/ek7jq6cKyLDxjL8yd3c8cx/aAcTUOECeU4WVSPoBGl1Y
dxRzJ++MrxD8/gGg8IRGHUrthcfreKm+vfy2fN+ykk4YYYi+0+BJ63soyWxRGN1CrQnGqHwLaQTe
n8TYMhREgeordMeX+DB9y9iLdZKhInivrDGKaNzJVdXHbGmZhtWXNRojea/q5QpgfxUPPE1eVFF9
rArEGLH9NJnDJ8YXq1NllMVBKhnMOaJJweT3m1mcw+8vy+9b9vDIWYkLVaaTf4V1PFmbB+9A3OxX
IVCeWXmnX0Si9xZ48bmkeIX54sBMoOd/jTkMpbI0tpKlu5AGArJ1cw+vwmQP4UfAvUZVKb3Sr8sG
2TiYZ2IAy0EhwGlk489iEWDSzudVX0yYr9+M7bhtsHzfvBL/n6YizOOsHrkwfNLuZInhks3uGTtj
f+7VVeqN9jG2n1nOW0d5q+e7MQIziCHHgLTVPgba1oYH4fvG9lOzSU4aR72TW4dJlm1bT4cPqA+7
pe1C49nuAs1y/EZ85Wz5n8alkZzUZofmnA5BZ4oSjczYzwQN11P5LlBhWUNlxVxL/y4UL0m8uitn
8RBJ/fde3gUEA+BBG3ogaF/fx8y8i18QzmCkzTpSYeojUQ09VEOaC6ej88h2NDFDgDVDVPo0Bv7D
vGcOnilrjBK7jFPCK1dMoi88ZInZjbyCT/YXIp6+pnf6p/PHJtlDhd+kEBhp2eVbyHe035ETWkIe
TEhWHVNqfl9pAkOTvobUpUPFx8Gaos02SzKjZW7eICLhq4sdb5wMEPs85P2dyfrSXr9cjbw+m2k1
V2OTlHNqRMABfbjK96ofBPceK7F/s6X3c1LmPxfEEg++ziPaOkswbk+UQusE0vPWucQOD50WHjx9
j+R+d0YQQ6pYSLJ84p/CKL91b9zjVy3MDd9X+BqAT8IgZXYNa4l+7rIru2uUtc4ywIqINSfDjvpe
RJDagYVb6bifq53mi0yspScc71OkH0K2eXEjcVVGE2N0jvkFuttpsPxGBdQPzTuuED52Co4/sQM1
mmMo0aSUrNZk5aXEv0hYN7jdbh/CmvyXdB5sUO0u0BbPdpMKjCmeoF4nFsDQQ2eur9ABYumh1hX8
OXnTJvWYs66av9Q+yNSLH4WFVbizhgK93GxQGLIfPUGJehqGKlVEfF41sWAt5SoJqd9W7NcIhv5g
i6MplPNERLE+aq1BZL+SlTKTUZg79JsKuXRSoWOs5/MU6Fvv3wMUqpC0ZludfU+CaRdzlRR9fMl1
xpDxwcdBKlsID5O+TfaTWQOfSksxiXGMf9SqyySYoRR3a5IZzGXf1CPTO7jM48Y9+AH/JrG6MEnK
g01w4XoJxJ/RcFNbk5H91F9wvSnlYK1Ra55UAR4hJu/8v7+h0xvRdIgljN7obPGh9hJSaAWbKGf0
LX2gEwQ0qZvCQNl5SYk9GuV8rKsZQMkwXBKh54lZDDTlB7LmklDFfrrJUWSzFZGXXDJ8ub86Yjx8
dwYoO01/jU188HC8nc5Ql9NMNXEG2U4ndHgO6M+A6T6b+dvbgmKsSFzGFK3qWoqXdd5ZaVaWh8ws
ddI4j84qOg81lVRnfcrl3yRgrUjfagl8HbUhZuJFBmDR8mVIHHcZKnwI1jU+uaUmwRkBPKLfQIO+
u9/kRc+fO5Xgxv2hkFPwYbTnSOM0RLLBRcI6OtbiMGY+lzD0rWbhSyuO55knfK0HIs2mMWuET/s/
m4NlPrdXoow2jx50t5+nb5w1od18yq2O17LOT0LQqCyQkEO1OrhWGd3WeZh0PYoKNhH0MS1z8swB
/QyIEpWXXd97Q8DRbC0wpug3zmb+Cc01h5g7R3N1T50KO49Xk5mtaRqJ4KVs4PNkO4YaY0JVMo9x
8DfCand0whxd9Q3tIGI9QYXkV+doiPXNMJeNvhUdT7OdwkfRQav4B2iMLOQR/SUF+sg7uSKrBQdb
HFEOYomD7b5EWjgKZm1mW1p8ttH1BE9ETyjp9AM2UsgwWNa/fTgsZccxfyhTvEiQGnxWSSokB5JT
2YoWiPMUAs8c9mk2QWUcunS0SlbHNhxFvBJkU7ngmyf48ODAsbFGrStifiVPfz2hJe9puX3iUdFY
//U8aiODEMsn3ZAelgfE65Ng7LTQmBkyTtQgc73l4UFUpe6oZLnv30KxC/I+z6aeoZbWs4x/y+Mi
tNuvNrCZdJtK9aPaYd0CxE+Brzvlm/diBRQ95D5BhZbpNh9+6S1GsW79noigrFJx9S5oZ4HLqAXi
VAcZc8vvXV2ybUVesVm+LMb2j2MHPeYsJR3OzX5+By05cDS9+5Gh6EGeaatX10Q76UX/pkTYAK6P
5A0TO1X9zUZ01QP2ld/iUI7FaB+CAr5Eode3hBAuO16HP9VCIO48m7CVaSs/K2lqe1nIoo6b7ahC
32KamF+57GAAtOmnEFes4vusrzHjpr4EHKXF17qV0vxD/nEiEKhvoGV1n2DSzNu0VzjDdv41xCTo
C0YmWWz8Pke3lx9Jf0k6BuniXL01tlaTIDtFM6mLMxHNjWa1gssavpind9bZgJ7Qk5pdMvD55ZxL
BVapuWAjK62EiQDwpp4Zbgs2C+NhpnTLVjY3Tz0bu5yDPoeuTula2Ja/tm5oDpSU4pN8riH6hTkw
yzBv0BkmSgB89DvFAVkmp1eZkuI412wOCFgeufUqV0Jn/nZj4cER1UZ08CUnnCpVRWRu9nzEnz1i
Jy0tlTzfo9UuwXN19Icon+SoGoODVriVCFiab//WYdS5iPmUmgQ1a8JgXYAj9lpRkO6kHtCPuO6P
1bQ8RXeiuDBETtPBYvZ5ySRO5VnjzxQPVoCLIyVJWYnaYno3DwTq9K6nWqWns6hjxTkDMzAXTp/4
bEFNhz2pI+RRPaafZ/QOxkgITNw1zPmdntE71mbLtQVwLDaUNLva/LsuIu4M5cPOWRsdLA5qgMbe
IaI5KcDgVhs/7K/bf/Z8PGbAC+r5o57U1McPddKvRXmRC1FkOg6Pp+n8Qt0JnHY8bWa69NtNiyGc
C1yT0SiX4YjZyK2xopwqxWsEHCi0Tbfl7sgebZ5fPOOPV4i29J2i+CVz4u8LRSEGWvAaJVEGZUg0
No8/XETBhk/17LZ4zqN+NNa8vn3Fs3kTr+3OUnSfA7doGMuGUlARSVejAqtT9w4X7KoZKng7xbfx
P4zPUlHoJzWc7Y7Z/LPqk8igIdox0pmIb6cdX4AbrrjlTrkBPTIYIcf6z8cI3g6DTr6QFyrC2DT1
ZD3qWczknJNrNDjI0PIpd+j6qVfz3dvb86D92OJ+OISJVG0BeyvbKVkqTIqwiD1LgE1wU77Ja2cf
UzXu1XNb3aqjojUDF39ywqX0i2j19XWlmdcpTRsgkeSX7xSVpSfJeOH1NEfD860ASuTCne5/suMS
abcF9n2cudrok4vn5CORHM2D0lKjbW8ZCsRsTW9HI83wed7jVssszvFMMgwg6x710S2XOgAjPOyW
Ty0j/F7cOaxl14S1pqxLEtHeo1vckl6nXBEgWa9nzZicO7Qg3ppiqujit6L9QX+WXFsRrRIYFgT9
Y1WbnWkRRwFpnnW3WhxGeNczWhPIhNWJuyzsys2pWr9Nfbjlhc6qL5p/P9CfycEgJOfkj3ez/2/l
Lad1pg4HKx20oU7Fxx/MKEqs77LQzxpw7XXxE/ILOKq+ZJvr7BvZUIIla0+pkT7qqrT+kghnXTXn
aF6YnBY1wC0MfTlzG+zp9DC5yTzG7tczPLb6YkFhtPHm5OMugN9aWvaHOHh3g42ftjkz5kZ3pEeJ
FQHr0Gpy4uL3LH31OaytL6K/ex3oloVI3FtPKYLgIw1g1lGan3vOsbIzKvesAt8SeSy8jO/kKRrA
qeXaVnwUAmRCV/fsTjvj+TP0HmHiIJiK+TXA1Cri5L6vkHmA5psxwNCVIfycChXxVkQW09M6woCX
q6+MheuAXVBagoenagotALImiyibmH79Ns+/9B5p7uk2yIz/UsfXX+6325yNMzuuVAluaMKZnIy3
fy46t555Lc8DWkiRmDs3BdyNirgz1u3gBqaSM/wCYNQuFvpNIyoCpTN7R92s9ktaQf29L3amWt9h
c/52a1h8fHVVAkHf/k3pfj1mfhNGGqrOyxfKqI0WQdP/CZqrPqI3hh20/8tyl/8IUYCyqt05ahgj
UC5X0nUykaizMNQx/pxncNn/XtCBfuCadE6IsY6uj6Nvg/jwGdEG1tEwjCih88UPQt3sVZpcutT1
iP5zSn+nywhKpcjWLTNpV0n3HY0QcsUX1Zz86SWpnC0MHbQlxxpilKTXOJubJlZY6mfWCS1Rhs9q
F7zywxI2KBd8lDLbS1ZArWsQdaMXPynIaM2Ed3JSxwSNDWI1R7ft9iRJr+d/HDFlM2zOTZ1EuEva
JMK9DlxsILiz/LJb+t0m/vFw0j3wCcNqgmcyFe66JITNr+BsqbkmBkKUVN43VzH9tqjLQplLjX02
QstkkVOalEsqHqRFBjERxA89vWJr/bYxsmrqq/w6tzl6pY4baFTQ18QRV7A0yW779brbLjCgl+Ez
ulmqd3oAARjmpOEj8Hvll42HF+iPWooEReBAv6ji1L98fS42pTDQcWCM7g9P3GKNykqOScbolBbY
ayoVgTC2MunVRuW9cSI35szRGgxUkRCJ7r8H2bgYguSdTv4ccDnqQ8obpRIW9MOQSLaqdLcfAgvz
+ioo8wS8wxBPCeeMaHVVNRlDTK9t0N2ee9VFxCF0PbC5/x1TutBexp584a60TzDG8COO2kx3Vbj7
5IhcSzKjKoEOkZE+nmNeD/Nm8KlfoTnSHSUstQIsXom8uElcGT7DzyHhB2Dz2+3JTcgCH/FRkMaV
Bih+uvd+gWCNVx3Hu1pPqBE1IqWUd3oT1skZ7P3LUbTfvY/t9grNWZITBE631M4td15it1NzRaNv
aP4vCiD7yGKMr9q8qbjicQI85Usllf7vVcW0izPQ7vkQpt7sfdg4uuuCm5GwFXV48FszlH4itfDS
PDn1rjkCvfPGvgavJjqTwjjemf88VYWTgMNfVfqd1X0T0IGbX5t3O1KB/3YjMAfVMwXh98ycYMIM
yka9K2OtiiZzYvK5jMY1M4hp0PPwIwp/RTkLXiMdDT0WioggsD2wNvdX7Kl6tDSiZXAdiHlmkjA3
zqPzgfftWXaohh0GKJhRp08Hu9PvH+cnaPOrDZVqrhZqiGT/e9Z+LtVwSFOqWmkhsV6kyciyyQJI
79p6uKiEYO+ZiZ/zcu5wnc4NIlvlwUXQIqNXh8hWsFbBw78Mb041zE9oOucP0NnhCu34BWBIOXBa
lsqG+FPSkmTtmvIBkFLhC6TQ8WWbUfAVyF3GaseOzhX6aYZtbUvOYdWY0gVyP9nIzX/3xp1fyJQ5
3RmM+P95RKtMVY+iIVW5Hv7P7V1faEojJ9EpOkKtHg3Ejl7ZRB/NvOyoRTITAjh7NXVi48WWGMWk
VFVdpD725iSnSpOyMBhiMTg0ONGRD4L6SQ1q4VdbnWCoVnp8vOXQpL0u57vZwoY/mPb+hrmwP4js
ovNaL7bI1DLYDVilA5Mi3lnnHS6Uo0gtNYGaFR3n0PJgcgEz2MOMyTQH/Vl40CpOlul0kB00gxSs
cayrpXdq1REF+d3HM7FpKEakYuBLr2+yFlj1zthUaeBgfugNyF/xCed0NCdDDUuAE1XWnnW5cUcz
3T8iGXGrBllBBv6LvrGgku2tkU2+k5uUyIpxOu2juM6h8+m7Z1ZfwT43TpzsD7A2Cb7E7QGJ0uXT
yyd4630+pIuCGXjrzQW/m5KmNT6qrFUISP5xAUwCwHU7fzGD6QCAwKqdysQyY5jQUxt3a7GxUxbu
Vkp2kqPBBHe8t7GhZKEC8vcMMfFp6G7KDNIHGQt5olX5DXOwVRgvhLUTIHsd29sg1WquPMNhr2dg
4E7/a3eKICJPvJRr8Yu+oRMeon1XETYMj/b5IzEue68HglYRgKdLpUOeNTJkLaJk55m+PnqM6ycs
UZ2q06arzoFNhSWaBPVsOvq5lequwPr9cvNzcU2HyCrkCJrEkLCNgekk1ij1Uqnj1n4R6UY5bwXJ
9iaxtsk28x32EY6WQYqq5tTq8F6h0zBXYZb0FXhlreuJqTMxl86xtNDwdn9zuljWmefV2zcTjAnV
sWmSSLfm2rna6UOxMVHxAO9LwiJlb9/bkFLQPnfU+nI+VN3Ev4OotDXxzHn4+CybO+BG4tbax8KL
Bda9xuegPuJ2kWOodoslEjz5TQadn96811PXYjXbYPpHxFfiZSYE77UOs7dbRniL6cddTYUdryJY
CbQSwwCl7yDDFVFkdQC4ptDS2va6WKdk8UrsoArfqW8Xg8p2GCIIUbp2PVzLHCLAMSlPJbvCq0Wb
L39BcuVfv5nHRD49geVlmOuiV3MMSVx2GFhX9lRdiP+2Hp4VQ/pGGYvFNRsWnb4AmiSsoCQYZ7ZF
uerlEBF0JeuIK7elmGyb4fAUle0Kha/vvWHBQmAkoKmySx/PHBwtFTJDgceXx908/w6WEh1nkPBB
FovF/eaxf0qTL2ELDaPqjyUnxHc4pjCejJjVQ49+PsXDahy6mBl5rmQhxAiJgCJAdpKzdlUWtRkH
M7TqCBXmfFG3HdX20PElQEC6N0Pwz0TLpi7OpBrTKqicM6HInew+7usPTnCLiAgurTGBp1FFQhyW
h9BdS/wTJ5g7FvVx5uBCxDrQhgqlvkBCVT2EjChinS9eRZY7f6OAbKS2NiZUoxw45hAmAgYVeuVy
rK263+mpzpmwR5R2OCFYvWmyKsriLVWNrDYVXb98baB4We6Gm5gdwyuQH+FXwG4BAGR2V9ZTTk+L
rYPG4HhSEUL8trUo1V5vfrEyzvnAolKrWuYD2by7mSQmMvjza9MyEAxywgRG0cvxkpta7fVBjV6S
uU3B349D7sXA1PM0nbfPJr0BL3914+C+rlVxeI+I7sJi//fQHn2ksHIxcby6r7Y3fzpPBLU2XWBW
5DD3Eq/V29N4Z4DtYTATSKYTfAwOwK7lin2QX1DitEHCHeEfZusJPT3MNrtF06RBAmjAcYE+oRjJ
rE+EJ/ZFWzzSGGiathh6pbB+SYz6OJ1iH0HxlqX1bjd6zr/1LDSI6gqzLlIOkCZciA3JzLbYn8hq
gaCzIXxFBQjAOGVZbwg2yum76LM63+Bqq9gqS0dxpKYQ8gTOOtWsd+QIdJtp1vuOwJ8olpTyYK34
fTuXKY8/jWxromiDrbOSxau0VND5QxYD/nFVpdpsW6hVcLdaYDUo3hANFD915XiOiIhHmU11e24g
Ds0witHLqQKTk1u3c7NRTZLH+1+I3L6GGC/v2s5KvMEHR1V6oIl5fmvURRJ9W69vbaTwmrCohFoS
GOFB6ZffHl2D9t4f6hTLKJZqrzsdizmkcq0AMsconse3+z8QMeK3llEbnWzrzcVYurdAT6sgGDaS
GitI8nYSGEEDqjlPF1446OIje0MkOjKn0mMozXGXKKyhqGfFBs39xS/irdXOw1Hw37MWrr76MGQU
v6CTMW4RQPW8f2YDQbtGsOpBXlLIYZ55VlMcPmoQzE9GmUSTkE8/cmlz9DmFgak7WiXWVT3jGMPG
REZ13c0IBTq1q8mqAmq586ot7iFGxg2P18tCOae9hcY7xb38XFf9lSCsoftMvOQ2LshUArGfKzWN
tDLuuLtIpLS1eezvnTxvhJdGrb+IlUqYP4AjwDWp1Ni7usRN+bDvp9+lP44J7Wz5Yo0me9Mip7PS
1G1eRDhaMMhFJJRp6kPq8qY3AoN5ljM+1PH3KSYjTtkRaMBvr8PwaTAXLVSZFMQWI5uId0/famLS
nRAdN+Vst8GGmF84qH2g/b/YlcbMknTkFlPRNRZqdo2+Q1oanMcGquC1MAMAsGGmInlu0u3IMuDI
gbkfZ7S5pBj/mG2aNkeHmsQ1oQIA86Y9k2xS1ezrKAJH9/CADTluafCr8fzJbE9RhjCjjqH4PohA
/VIpO3aVllNnKw4lHNMKdKCRYUqmkCsM5G3la2EXhNEmTU+r634jQHvNHIjNK5EB2kn8SwobPgE7
Xhsyhn8Ki4SLOmFchQKnjHujczk4XqhvT6J27iRwPqwKlhxuGUBYvHSM4FeHA15+6k9hI6emm4CP
d40tY5LJ2L4F80rKAqapnQVhCCFcDOVAChBFSqVpPMqnqNLeNGiyBW/QIJod189w2P0WUO0YyhAo
vfPRTQJQgxH5rnqBPgHEIzH24+k191z2eSGKzs9azMPiZngMJUXwNz+uacUSTUxpFZhg5H5f3F8E
LY61VD+wditQ0HbSzlruu8+dYGuOTt/vtDL5mysjOohNRFj5S4iZB66JCNGCdEuDvoJO08VdwaF6
tVIYjgBDRBR3diCN2u9eUyZqB0NUZ7+SSy9715aXXdYAHdG75DIvLlWleM3vjxY0ZRSHKBA+8X4H
W5JRp3/hOoH1TBImEif3riKhx7yYy1aRyouKr4vMy6anXJmKT0ULXKCzFwADFZO1lVzJayKB9wkm
dPPuiwbBzs6TMe1BtHwF3dDX3WWbGObm85w3Tllo1kaSv7Fa2RY8VoiNBXmIQITnljkr7vpqZyZ7
ed59YC6rSkeefsI1sdCfj8VCRDdU+2nOsPngAvULZvUINxgPtuIlPMqDNUOlPB+SSHNo++2UlbVM
BI+pqCYNz4Uth/2UBu6Dulb6F0RjtsGLiOD+0I0jACkpFttl4e3L/rhtvwd2kyCYeLkLsh+1mXGA
ZE0FTSLX/ZJTl+lYq0aEtSLsQa47SaF3LR/03RoLuCuNO5EgVJPmnYkSI0VEAERwR0sYPfugaQte
19Gbvs4tWPDUZvZGhepln2TzswF/qkHBOXLUp2W35SszOpcQVaSyazEi7BMGN5HI/OgfWfkZOIF6
wfMVQJs0lqp2WuJCAWQyUtJWW03z8DUoEjI2FNO+MoFSYuk4yrP8NEZLiLv0016d/qkxQoZfvRqG
3vJAjexovhCf05GzJAuP+/wqqFG4Ew76hnDaH1axnTm/wDTBMaUMwGy1li//TJZzTcnHQrtxR5QE
ltxh4Fl2lGKrStf03aEBvMBdxRIQQYENO4/6PnoYHa2HkgFN0imQU4zhESCMZOpoDteqLwHBi4sG
oGphjl7tgnm40OXZ31MCvvHznSH10qLDVOZC8AsPtehM4QkLqMACYrRJ7cWjy9s5jC3iGz+fFk3E
Q4DMbnwlClXxWjItAeadnO+yOYlxhCfEXOOV58P5T5efEEDWUJbaklQYzQRoGWJRrPODuYLtliIV
TQixCDk28rkwNhxHxYyhuUTyyx5llSTK6kHtpywXg3S8wsucBywULIOBejsHx7uf/63q2dJ2PVAa
65KPaD7Y0dR0ouIqNVxLN6/fHblSiUB3EajkoSltvL9pTNQPFL61/Z7uoBPNbo/xXoetX0I22Sd7
8/e+UfbfnLwrnAUfZ9Et7QSOhKNH/dIVe3+aN4IUl/Xl8HLGm4+NdO48cvDcLvoK/iWB+1VoxPcM
2xW9CyPR5bZE1gj8aI0FCpx7g4hLO/PtLZn6crCth/yx0LLRvWL1qZYADQfgPiZVg+ppCxHx7Kj+
7NAspDvKMjMZuZYNRTnF6gh7XDW33NRvZg+zqvas2Jo8UPEUOlcEK0wQquV/9LOPoy4j0bL+Dam4
yhHAfw95f/i1F2J5MBckcLJkPZQQ73vU9QVYCsDg7jLAi7KhwFLLygg4hNhdNKKFuvFMNqO+5b5v
v1YmfGcDu8oJZNLPyU6PEZuq5U4HGC6IbfBs7JCyge92l92rqebDe60XXphktPOWigAsjMv6KEie
kPzYriOn/HU7xpfseJSpSQatOh1K4blI2Zp1jPEL4ENjogBx3nMxxpeKcOcB6ubyBBMAliILetKz
e1kA6LVW8jxBb0S6BZYA9RO02F5IcpzlxtblC0WThoT3BtmfrgovNDUIV7ZtbKBC/C/UmBGxCtUk
JUxVQS89tjDlGf9mMQUzIDXGuBRnW92OB+rWRD1Q8fZdaXzffshY7Sj2pg0Mg1bjGZ5rAF+6eOgf
bia9ceU9Shh3OAdOl8tKDJr6RePC1ndKoHemYzXLloQQk1m0h+dvVjGbJllgxtYswza/CL+eSeen
X7dk6oV9vHcS2lcUgj4mF46xFZFGlt7fKwBV5aFKCNxwm6xz0S4Y6cgf+2hLoZDgngupegmN1IVS
iy0rH/dxVeujHaOalC0JF7rhKusNntMmc4yyqQdXRzk9a3zAPYgKgeeH022Fwlks/tdYhRnxmx1r
er9cJJAZa8q0yj0uc7uNuNzY827xnY6BcfiLMnrA/6jI3JaRpukE4In9m3n5kegBfu3OoSK634YU
wYiGU2YuhYbD3XvF61vK0FLR6LYjZV5riFi/XKDXPaXtgkDzyGIKtcXctJ5npv6nNuoUUOp6et2i
O6dq0xHnimo+5jFywTgeAFIPUNPdB73R22MRwd4sE5fZ8F5sBYYBWSb+lJFITzSpjlxT/Q/1e4AH
LpU3dKXuF3Fr7ZAcgD8sbVgnPezXklpEoH2t+38eYzL8dSJfINPfjuhAB804agYva60T234fgeUi
8DAV2fWjGEIsoIKk7fn/aXN05EU97ScMMhzHv2xO9RexKKShQ3elVYce10Uae9UHDHzfst76IczR
+n/uD4lUlz12/+T555nxMdzAfFfMlI1Jkg/ZI6EsKqawBHVlU68aKYlxcwgIFEexyPJqC5jV14Pv
HQepSxKFv2sXfLizY0d163j5kB03Fiuzx+04oTiFEP6DTJjYilnErg7kQmwSiS2zSv+4rV+J37Zk
zymu0isNE2LvTpsJwa0fl3i+zgsYeFUOa36oZ/lJkXQsmLwORJfuRAjeSCaWFzR8LRi0yFbmSnl/
Br9JvViJa3OGP9+ck79wJc68LXSx6o+YCH3Pg19Z7z0ULUh39TWwARBe61Svpqnvc7L/YzCNAuUH
MaLbuMNJXX9x/jobyGu/OSDU+RgqXr/9hHVeOe6znWJ9sJfaIiY1cE2BGfFCisV0qhMi7kFppIQJ
sX1XF6tydg/Qw8jIcJMjU/e0BY02NHM3eGA9LDUQS3Bha673dm1Lio1VFaDlA1fsF/Pw79tTwhFp
gSo/kkiWF4DfKY4C3YIJlqtOKijaG6Hsxo690qlA6HRq5vnRoSeYVqIJfusxDEjAkf4EqDkKB7pl
tKcHkmhGd8Ss/67x/KXWop7sN3l2Kw/6IQD9QkhmzyUClCMMaWFzUfirN7GrcgHODeTgk9XYPVD2
VnTVbpAFmcEBM8588wqSoXKOvqXbJOhlHvJ6nV56WZ8qJqO1Y6KjICILiCNxdN7eedoLkA4vAHPV
StwU6c3V4uyvwHrsbU4d+krgW7RLIhbptp0b3cO898NgY99Y+iap97UHJFSO3fwg48oIOwHViEnd
o7zvOktc7ytlBLqz5dzd69HDJk3duFD/yEr3sMvIZUNNYJjZLHlSzUrFNBRonuvC1gaTVU0spWnq
uHvlpMIW5fzYU26d+PpXAxvJK+deEW7J888OP+lX7/Nhl+1qa8ZkU6HUoERS5KjI0zCIi42vDPfG
FcwoXGmIZ8JoU/v4uMuzSxvlbkCma70h4MWgKS6scUJGak/u3xLRySdoQkrnudVcvzTeK7xoXakB
NNp+zXrsY56jvVcgBSvC3swZTXhc77JZhkoyS6LQHD6LyEwz+35+XB/QsOk7Thu+x1Zym6fVsBDn
GrIwOwdpNZTBw8pKciAIiA/76jKkMsQkKE1Gi3R0xrGNiVBtir5tg5nDBPu53+IwfzbwumbBqtQR
cCk1ShqOjyV04g1tWwh/KI+EjJ9LsSGAmNbtTVHKv6WUvX+tBXKTVB2srNxu5Q3voegngCCwDE31
yNcNrfSaqiD4P3YU1RuQpkeEUjs9XhKLA5qqIKujPn6FgSitRT/iDA2hAAt+CzwQLznSlqVVEHRg
5fP+jjj0ZTZWaJ7JIQc0dhmMpWCnQuzF09Y/tGDsar7CUSJ3inooqZah1WkXOr0O73AlBvIuPQX9
8SH9XB76qi1HMRzNBPFNXhpaeozh/zWKv3oAQFnX61EPsaVfsyyuZQiIS25Dz0sZf343hNjBlfqF
36ZzYQTchgEOJgD+BZIWx+wQUjg9yEKxPSUCK4iYeFOnT3xKPGc/odKYAlEBvTux/Grh0x28GQwU
9XT8O8rZYCyPQ7lLAnrLEi5QmS5Y42mPfs1R+saMvzdkgV0Wi/F5E3Vuhgf1MduLAIacUuPK5ZH4
bT/kuaH8sM5zbN+kouhwmT4FTAKYlwu15uFwgoZHVUo+uIbDBYvp3cKgHHGAR2CwHCSd0+VkugRO
Yw6R59RHhYgtxwiUEo8OCmWRINCa6JEekYiHKsypmYLd2KRi1JBwU8oLxqmwa5D+k7FF32qHeYkH
qeZLThkI0kNpIkxtm4qTXMpgbaBHdXz7zY/s7SvL/1tuOK8nnRVToi6FaaClth+Y1Ymggy8Yztds
O1NE1n5UEIWs4K83Gh1hy3xkmJ/cXJh34FkF1LgKr7HEKHzsIZjETU+X6rPBmfSd+mzByipr0Kl9
jARQpgexxlbcGt5tUF27ebyf9wXF6GTZjD/g3zfkYQ/ekXVKrt3fAK2GIIe9IOwzNMytFytAgzpl
ckNQyh9BchstkPUIvOyhutdT2ScT+liCnZRyB5wnYWdmjmZlDkLhuKTJFioedrq/NmMLxPRSS24s
MYHLRpNoAraj/lj998jmni+yBLtMQ8BlVKk1/rYYqdVhhnycreP0jtpr/4RT4QCEFAsqSpNVUSi/
udtzjOw0+8cmv/2HnQaQod1s2ry8zysJhhJrspHf1IARVlEQ7H4UGY2rMARVjrbdzI1IJVV4cnxV
f4/jf0tNqoiClzimPYcZH6oA6uU3GSDlsx/wkGrSP8bD15BkA5s/lf3Y8oLqEAzfpmSs22AVffUc
HvKIud8Divh58ro7/I3BqU+Mo6tzPSGCcb0DVkOxq319eLIyGXTf+eZa5HBHZiDIIECl57YXb9he
JNzlc4NNkYtNMpeyehVmmOxRnNRvVpF/SRkcOSBzGKspWYcyGyjd0U9cZQjUH0b5ZzU4bVczbULa
VD760MA/NpHWVtob5w84ywF+u6wqmByMpx4fo4v4ne/dDq2V3tiP7plX7lvoUT7lkPAMRmuOimTN
MNaxOBEVlQqsikyIPKEX79IP7N/79FnIuelhU7oi/jHFfknUfemQE1DUdIrPmK5YYPiuZpn2AYTo
zuGptRNdJNkzv+80u98MwZ1YO68rS6EnplpGhZqJwjb0k+0lHJoF+EhEvKa840pRxg3UtXE/7WxL
5mpaXoLAemBTX91LTtvBMJxCd+VO0+Qsh0BdolKeuQ9NCivCAEVslbajirEv0WAqXse353s6vJl6
H43oSc9Y8X4TWBw/WKDi5ye1m6+wknu1Nc5JsJLP2C8ag3ar41bXR/+PYSYCIYe33x6nHxi/ZcBz
R4lqWMAVTkK36sbtLz4W9Du5WmKmfbpB6PB4psO0YomE0awv3eWrHY0XlJrLaJbvbnIhiry3Ei0X
U+1uaduLpEEd76q3d+StJcTIMtMoPVJfMsZ8Uw03/Jpfuf9E4YjiVMUktSPE4oWVT8M2NnB+yi7E
633OqVvALkvEpLE2kyib0S5XBm+uLeSg7/gS1atXcUnmgUR3M56uyg7LmJGwYJcLMrmCEAYtgWuT
VOwdlLEvN/79BprhI83tbBA8QxWXJH2MM4QLaYz2dy2Jd6AWTLY61epsSNfrgMtT4RAa+SN/B/zL
g1M5RHXSqJ0gtKSF/Ae8pNfRone6d+6a+jFs0lmDS0kgLoOzGwAJdxlJLmGq6hvEZVanucYmTKnp
eawJqewlkU136o0QP3J/KJoEzWIGFwIHXWvLBeGWqzCQ3WJw0ALD/icbS5VHl2rDXqjHs2cNmH+F
NRD3uFT9+fFPZvgruOmhp751DTXToR1r9Xud9qzpnnEo4LDicc2lX5TUzPi7WSXm/Z/gJPIwvhBe
rcV19q9VnoaiV+xsOLSPKT8JNtV/K3B/UuKOC54g9Mm6Egv+BVm6eaTXg8ZMrElJZmuNoFRjxN4s
zxNYgsq5FTdmtmlBVqIBa+EGp+3frb7AiVTeeHm9YldzvsuYUAPd9kgVBz6V2yk4wL9gj62nVNHh
FqtTsCCk+1OzvY1A7lBvaoSxkojIRwKAIIhlUswNuE0ZrRyT65WJj8ULzrHRFJtsARN73hYpUbUI
eZfjzRALE8H1h/6/Zl46c7nuupTi8n19HGtpYOM0qsJeiCd01kSpaAlbD4xQ2J0n0abkpgXT1OTC
y54cBvQbc06HFzW2qv/VvzVlkANvCqf1tZ02BpVGcS4U+9ow3gPWyvgFtYB5gQ4uygAKuMjSy8Tp
zOSXYRIXGvoi4JfJopnlTkT9BIZ0fONpDM44NsonMPBhVyCuzTP6rbWfwqBkczZG3l2cNdKNaC6h
ZuZLXomFQ9e8RWjDwVf54zBSEhVTZBX0IolDAbobiQ8yM5CPUcruj6eOa0ZThsIaNGJvUeeXIY2f
wYOxcTH6W3uzJlDMr4DxbDI51bFlhpjuc/bdHy4OOYEmw5/tra1PWOJ3epLLIk6pPht/RAdAVyQf
OIeQ3TEhx0jqkaL3xgS+0qfXqTroYpgEsvPphfAGap8hQ/ksXAejtw2kMAAD7vrqSrtaqQYr568b
zUzplgczrQIkVxHc/Z3BWem3xtJdLBewoDnlEaKCMnwGRfHnFgfi/+RVB2eC1W8s9m+KhuP05YVO
0aJIr1DxOyzR1QrwFQMG7e2adTfGZ81mMgw+ymESvFtW6nffJNMI48oVLEpXyKQXGBfbQ4L5MvDp
wJ9wXiILmWYAc8rYR7zP002myC1jEA6talvoKiPhT4ldDlalF/M+6/r+ix8fTrmg7uexbGiyov5n
sLzyD+5ViQ0ztXlDHB8YCQ+ALLT9EkaMgvlwMA33fRxHUjxUZ3mQggPLz3uQR0q/ExgMUuwJESIP
A/v85YxEVVCvu8N/XOYsAZcmx93kuDzcaf5mnQcmaz/SC7LJvKvSLh3Th2KcA3GKARjlpzZkRlq8
PMcM68tS5DuEi2lSCagaMQpwfUzSj4yFjcoLmq6BtEKMSLBOBrc82eQIgD4lGjTYMT4pD+XuEPf7
UxufRhYhytIf2fVaAqW0+edI/eeEd0AVSRv9i1sfhYPmav8w+Q0HykD3WwdecGRln3728n/nwm8O
ibQqkCrUVSR75c9hkndrNq3FOFMC2uEutKHLJS4U0ngsUSiU1SyvWuk3ViLTad0FQQFPaXdeJ1s6
0jmT8xGrEYER6GNN+y0rPmZEfR3S9l6HD9rYBBYN2I0pQVGREW0ldByZw0oZH4BXubBCWivHXyqw
2cdF9XNBRKiarTdjkEWWOdTV7sE43WZze3iBtX9vY6NrfVdv6W8Gq66rd0KrnmNkqH4D02CVrLj7
K2tvQ+Sc3NBvFqddgNmkOKtcDkfrSMvyRGN99LL1HPgZPr6NfDZL/VAuzA09WbFywTQ16CwUHwGX
8JAlPpR4vxVn5XTLKmqNe94OzKfFakAGAPgOBCro1DOHbC5gNJ1eXczu5LzOtChPfhIyFhsTZ1yn
Og7fpWLGi4GCwH5tvgRS1Pe1beNLz6dbDs/LcpMEEqK3axjkbKv844jWVVc1mAromQeryEfbiizu
Aa9fWTkSwqnQF1k9PrKmuLX3r/iYc6GcaRPIX3jViH90cjF4t0UZjoM1q2i8LgJk2j0g2entfNJM
4viwKCmnqOU1848tfVI7hQemApEeP+bZfIHpk3T7bj/eDlCihG2tT+rZ5LOT9+/8UFR7VouKIbtF
5MlwZaapZA8tcSAp/sopiKWZ9jPc+Cz8Auo5rN5V/VsxSX88mKFEBZltLuaG29ClNVuTJ16+K3iM
m6EPCNqjOWsK1eMdHD1+Kb1mXhk4JsxRA50nG42m8u6cxWDDBVWYqC5udvnwJyzPKDUkQNMmCXte
vFO48MmsidG6huaza/KUMzlIOdTDGNLwa2uePsbjbAMFLG6FmmQvBiDnXHNuLGMtZ1+TKOo+Kuy5
zrmCIwwavEsfUlXa1fjIKMThdMjmj61Ow/X/R5tB0QXFKanaRojjJyVWMVyWIm4qOg27O11HTI0S
GQDDNGBiSa2iXDwjhWbiFZyprnXnIBFal8hdFG4DmD1mHo/6ejMuMjEGvK5aM5tKpl21A506Lein
yEYSiHhQGS/h9442T6+miIAcB9Rz9d35JNo8ZRIBIhkkwXGP2yL2FIcgKfVTOwRXD33mJTjkMs/B
P2fb7BRPX+481Ixn+wFnH12womj0hpfmCEK2WwJ0IJsw+2UzEiE2jnnFd+SUS4ZBGTf6+wCPebhq
bWrQGQfH8QAw+sHQTfyZNiPhNPBCgEa//10VfvlbB18F2a/IzFXjWFxcQYj96UqrLBPfH9Fjhfjd
+KoznUE/LrqBGJkIKExkFVpfD5/BiyXDOCTzCOeo1jXtjw8IeAJ3UWDTrWaVTPFel3XlszrQFsQ0
Ou9msmNBMjMAnJ6pkzipc41kLo5V1Sl6xP5Er5BexVaWJZvwBrjWIrHLf6u8PcsgDD1P/7fJ9pB9
g5GZIKmS1/jRJvO1q8LQXUaZV04BWRLkyoX/kKcAI9gJTRCFgOBfgqBJ5w2mnXZXBJgdVlGaM8n2
cMTJgby0wZ1ZVZaEajLZzJ3F+h9+I2dIPqU0vkS2OhxgDP2xJaSPPyyow81ldfva21MlUsjOngEe
UX6389lNAeFR+9bqd8jpvGbMlj6qmSfyFfISt4vWPmtOKFv6vZWTc2LWTk4eGlQk1Hi1MB9aq3uu
L785SYiiSGR0zrlIAIVKCk22dhP67A6rBcRFOGjW5GOkR+PB+OOpigX92Mai+pzulxyA/2pSpzX7
tfOZ7MSp0G7Vp32fLcmoeuZnwyfqHRZWdLOC/89EoJ0tHtszQvqxfbEbykJPFOQHXs46xOgJgobH
UN8uaSuv/mjV/Kau/KiloW6z0RnPRYTXV4rIeIzULZr20ghoeeAn8Ge2v8mLYkWIs2n9fXUrviVR
UiAWjjB25+mpKRoAOrHLDR6MLFuw6hLiaMSun7hcK1FzDfwVj3mG41eOZKf7EzeqDa2WWP/jOK62
WmmBZX4mw7FfK9gHl2zfx4JrU4UK2T+hSjFbf2qoQyPpt7gYCDAQZvKaf92bhVMYNOYQXTvdTFy1
A41emDGITsoWUlRK9U6EEFFhGUWhZliAT58x9t6es9ZpxWnRz46zHsA8NOEbAxRXyHLtlaSYRvvJ
5JvhB+FBMB1VRntplF7GpqqC9lTHJI1bN10q9qESld9ccq3eo8q38Jx5ehh/noL8HO2y4jmCnh0W
/2SIjRIue8WC9ACVlJq/VyzMBk9UTIh86NnsNKGF5hNcRM8rRSBG5a0ZnoGYCB4KSgohptMEz00u
Snk52hYhXShO0WM4/H5oXCLFVZgaVjsAcUBAmPMV8LyaPRGhMbZ+T+bX5VVZYUGcjJ/+iJGUAChk
28fvRVqDqQuEhySmNEWHG3lWgT6CgovC7L6L87rMAlOdxfoANU4wsOu43tEX+/gRuNFqtNNJcCIA
KubjtFdw9aKt9NeDC0D6NtKJ0WlXvH8Efsg0sPL59zC+jNRHb+t0gpTgVARt7SMJbqo1fLvpxsin
GSSQCIsOmi3vutsMKxvmukXK6W+s7ZBUnmTOzX/ILWbseXe4UteFSRtnDlLEsk7UigZV9kfFN6uM
BN9iA+jc6aq1GS8DXHjT1bfEFS/VRsu1AW3Dk1PXjuUbObp8pU9euphatFamuUFmqy7efv0PwjyD
f81NiaXQh5fxHMtAL78xEI/vCj0hTEcs8uXmXgaxf/cQQ7EjnbYYrix7hBY24OUzCtjZ6aQ6vG35
Hc/BQnebPxhtWgEN63kaaZyN65+VcoK0CIAURZO4fXqN9oUJ5YOfXI98YEUYQjMXkqAWxe039uGg
+TWXEpdK8zwrCLD/VudOEpcMrc3qsL87p3ZkRnj0UKU53piFu6XgHIqoncbfIKY8e6t8Vop2O40X
w4Wxt2oRau6svYbiqGVtLJjJUdDJdHPrCVfaLmJMKTzAWGE0YQixJGltXvlIte+5Lsjc05JXlntC
wqRuzSVqWMehZMtqXjQ6lgwXzko4fsqLNGFupbBtZRd7cnC7iZhYGMxHK/aFUfM/bU8io+9XY5pQ
MHQnMz2KH7fA/0UEYtYuwVUsjGwkGBvoiHbwDEhf50G366fy/t+aZRyg9suIr33bdgUrD00VZrUG
LUgwIVbhyhcArVF6maLd2r0ay+kHn/tzrqTDCxYy8HNzZTQTQUdRVER1TVPGkX6XCq2hJx5NeQqR
vBnpv2SjVaj3k8y6P/GAcydJOKeLdm8OHqO3zhqtKa46OktawGn2ICApX7sAE6JnAY+PynXt5w4i
X6p6j4lCDfkqEXVnvc51HANy3PQpbm5IIn5LehB4+UahIxcVeUTjr+oGNaFzraxGhol8ZOcvtvtm
j/1yDeiGNKJ/elM/jhea0mU+QxDc2ZtE80flP0GfDGPNk4POPHp9bH3VryBosvowWW0jzujRsOSs
aKC99Z+2JW/txXLZHF9CAyxm9Is4KOgNzS+h6B9tqr7lm63giMWQuwoVeEha8jzlvo7SlgQtRMJE
SIC3DIoSkYt05t967+L96/ODlfYFJ/MgRU1j1H5/PGJ01/pSLK+lX/jaww6Jst6cQUYZ0+chd21r
5Oj28U+U5llaTcZLeqoCkDkFE84HSuYFG+Wy4y+OBwhbCh/+wglq5BKEWzcxcHgGo8xRoZEwXNWv
4mszNtDcAffg1AB7gA4XsdiCNdo1FznkkunFPSzclqX67D1g9tVRiYxOwWVIPj0LNtAyV4cl6TWr
aGbz6T2kehxt2fFrJQ/BoWl0+npiRnZ55XbSCabPfaqepRJdGvT8F4TfhI8AdLR6M2PowkhZ3YKU
5kumylvfNQnPFsB3bkZXgV3vYzEVmSfvlTN6OH3yWswJshfv02qev2rMOT9Q6wLpy/DrAAufkHoV
oS2G1jNxYm7kw0SqJXRPkmsKGGlGN8sLwCokn+TNins9X9Z3lzcS3P0Iapno45QuUwKdLJYF1jw5
BIaMA7Kq3qFB+VvAriJqAFP4cf4wdQmGRMK9Wvqu3G4TfbRuxNZ6CaXV5ffk9ivxdhty5k5M2xSH
qESQYg7Hp3onqdC1eKJy96fcQai10Y3vZ8c34d82lTWzFFFJRx/LOKIT5sUmDlBlJBzC5QiNAXA+
K29Mzi6ErcWk8gfF4kLxwLnis3cTKEMVRcD5bKqcO70n6kPxaTDTblAhbVmK9E68ooffkcwnBdzI
1mPV806fRh8LHZoURWmWDORj+E7/l55kO+NFH/kf6J3qAi51cNcgMK2+b8pWISCxBgsCx3amcBHQ
pfSFl+fsCbnd6z2FwbXyBFdboGLqQ0MAjmRU+DMsF/AHgf2UzmKu/ISt2cySFu+6iOmNF0U0taxB
gxPybaI9m57HpOUDbAIrscCBFukcUlIMEGUh+q1JlIo9vkaa6ElvL2dJVYf1pMtb1PjKwpaumbF1
UHfJbEkvYyhr9XH+LDytw57QQB3A+VK8mzsYoX7qAhuWwJeT+DTkLn7sbn9r+VQXU5sYioBwtGer
Y6JsTNv+OZ8h2nCE/7HecgYu3yxLcgFKhhMXD6wjfUPBzbSlwrQro4YncR/Wbcmo0hoKs9zSnXUz
ClelyXDzAgrIxSdhTtpOnf/O+gp82nLxe2XJoMjLx62wLA/j0o0dtpgprUTTSvkczJS0CToCDGUy
DPATo8Xtx7hlRellzT//FbizxjZJxBskbTC7bT9oku0iZxkHjtEU6emGta+BIiL6Of9C+LSNt9ye
zWURKVm2+2TY+GEk0AxGtoL0Y5Xxs/0Vm0lHkEBfV7lM4KLyX931ThpGO1VzSpjTqUFyXI6H7Rkr
6mxx5+IRWb7HLBnYFy+oyDt+56ap4vv6giAQe2sf6UD+Llw0J4/S1lFvDA+MZ1mCNYGEUCtZbIwT
0TkAHxSJuJk7B8S2odtozJJPHFypbDWgfk21872W58ae4AnktESowwOu8UhaLJ2qMuhCf/4qiGcn
8tCmK2YfXA4TJJTOQsXLyUfv5iKBQuc0klt5AMv/e/6RAYoSDOBDVbJ0m52fSWHqSGD3TRwbZdYW
51ob2wjGbPlwNNskrvsXedqFPydsHQSus/WlaCQek4Eg7DBv6Xp9H7uU48mkrvEUxU0/2bDR7MUN
HfZ+GMQUaBd2V5NXtvbqDpL83Xi63ipIv5ke3COgqoaRR0BnXgNW9VtGDLVrZOE5WMgsBI1RiUjc
4IO39M4MxKqv7iQAEmZOfbGwoQOpkwIV/qmQD0CEuUu9w1EsrX65CyBL0kTIVlqCIIe1a26l4i+H
h5s+61q/RJcpG3CodczBKNfAKrt4eiBA6RoKV52jAVjaeKspRqKu4Uvp564gkwbl/FKJaFl2I7hu
idtUehRqopIlQ3YE7fPbJRTh+qHxelth4JmKOhHIR0uEzzuMB5Y+vK1wbF+EDShX8WqGsTFesNRz
vTRSuo9K7fahMDHfnG+xyoHs5TL5GnTYTs8QkTMeTxPtM1/rePY3OJw1HoqxCeMBmPyHNh+RaVUz
o5Wx+2hVTeX6NX+8q187V8wtfVb7bu7km/s3XvmdAEqHDix2XSrtlz5cjBXa+ERw4WOScBWZ33Am
soDH5dgcWLP1U8/JVjAf31bUlzBvPNaoAKyRjuaEFb5q5pMATgCHplhPOyj77w/AvwAyS55EpEoO
MOHlOVuId5+QUbTK5hGo3qasyBM66TFmh0jz7GW3CQ7p7Lth8qC656hT5UfGll41s8h74Ucw0Xhn
p1ffILyqYXD0JqU2aVeNGib/jirXE8HOAVIKQ79//bNCELAU5fKuiySg0UVMeuS+VHK9O1nXWXCv
JbcTkJg160tA6gYC64BwFCSz5sfb7Kz5zs2aCe7WxOzUSErbkMYzGIgDJ+7Jl1xmqY/ziY9lCGVE
z9PlX1uDdIxdfUQRgkZMYlbeoFnIFdnxhCq2I46il5gbVyvsJkPjOrjMZumg2LflvAP0YN/TiBGT
5DWAa52/mSy/TFf29HDQQhL3QGJgV9mSEQUfLr9j59qXqVhLm5aZrjPKMVG9mqX90MUL5WWFDZ76
1Zppvm3XQ6QSsUgvgxiLSns5beHQdm4YwjbSXjWqY62jTdCmWtggh0irbEEdlru4V6A1lqIGq8N7
WmCw9p4+NBJmpgsm/G4UNgFM87YAr9AL7EWex9zmCw33sW7lJgK2i6xfnHVmEna8EcVx+foxze5i
8nq9pGRPsCpLl4zHs2kS/wBMR8Yl9+qpWGB28w2zQ/OHunVcUMkdxIEeKDsHxuEy3SJHTKiiOaQa
rBPZT4ZoNY/82S1PM1UET5sa7njCttKMqON5cDsNHJSaoudfxixahCogpwagk2ug6A+BO7kIb1bV
lZOXvorckjNks/AbTr9FCjzFQCZ4V9rde6pzag5Ebq7gXRRt1Bq1SIDYdJuZavkcLUo5f+aCHz4D
ScgUS55sBwTG4SBG4Ciw06C07rqg56MCu9fr1t/8J5dvVjgj7hWz3YZ+QSc8lehHnO696E6T21ut
1t3TxCMdQAE1n3q00/+TA/9vckSksVRqan/YbJnJ+FZ4Y0cjtaxVtO84OfNMfpem3m9UMEQtIXqp
NOxM+nXsXid4EFQ1nT367txFAkQKFeNBDrQhj480uzPM76hC+SCo4uiIqDYldq3VZyNcVBwRWXtm
tndbAjM5gDPEG6Lo7M9q2p1VkSvTpTyCbPdHelLjZdHqCCHLhBfZpPX12wCmJLHDH5EXcTTX5kEY
NkXR+3+hNQWLfDBFQDFnb6zm1VXYpSiSaYsSJEbJj7SW9muBcUQwuEKZuLkUtLKE8wEQCpQuhKxe
6Vt0kSnIE5aoxUE7XTR84qn8EmEeE6vJTRooKG1/eDpPwBNTClcr9cqxfuXvsnSwMuJir3MkDFG6
p65QS16z531V64f+WRszkiiNj8n9VJ+yaFvWmwkzFSYG37inZpTd6Pf3bNH1vmAtTn7Vdf8eUnUu
IBrG5YR0HfY0Bs7zRbpblCPHio34kKjkSGpY+WQ86v/HZ10oeCu66uGJNOYVKwOOhKB2v9Vfczyc
1MZV2dI/wF6Bzm0zA5C+LnNWN0BSudUxIY1DxP/Y6mXj/UKSW8yxUF1YC6wR8O5OnM62d3TO6e7F
kfi+6dk47CZcWE5Yy1nm55B7swiOK8GP3o/v+eVAoKJWjRRFVv39K30HYmvfg+7nufumVK+xQo+5
3Wupex/z2XH7qbLtZ8H3nkDH7pU5CfOCFqJDdEEg3cxTgeQr9WUKrSSs4Waj6RCpuNyPdKsHz8p7
xkvw7fkiPnQIs99f/2MX//2fhfgQN7lj97rRv3P2Jj35T8tkNSuup9XZOOfohPTjL3NEVHQlP7wF
OtdjVmwAy4ZGGwgUXDldSvovOmDBJlNFhhwDxIhYlUf55lKdSZ7xlyQWuhn/cNlH3nIGyg8ghxrG
Zm2ryIOQQum1+CxG5S9800A5m/Kag4pp4ou4JtIruwmLaeHxt2V+Q4jaK466yF7wn00yMvw21Qmz
AVkAJ3BUJEzw9RMEW1r25uRpDrxhpvMUa4+B7it5hm27jmtVP9lcO+QTqCLtkcUKu9jHh0cCMtTN
PDmvt80uW6QCbokFrXF+dc1TpC1pthlBwfaoAYywjlFHO5xckxtcVqZiylBERykQf73MlBRbVTOd
AtuL5db5RX9OtLcLSvjm0mKFniCJeDoTnJmEAo7FYzYCMxPXidT0YBE5Bk+PpZSYfgJCgqvsPYZ7
ljcXoROBsuSGzlJ3NgQoR+IHBTD+i9QGGHQyax+VuWZqc+L9t4rosp07ladzZAvVFx3XPmyaT+2s
B3lrE1Acq/izbR7vwDNJvlR2G+FEADtzrpbIEeJ1xE3/8D/srHgpd1kxigMLhL0lrPKKM0wqcfCl
L+5zowVPYvWYklCqb4mx6MymvqLl6fa/++UGbuDrJ+RYYdfehGLqb+A4TtdHJ2k9CYzUciMMFS3j
wt1XqXLoIrjQGeyR2j7ENxm2ne5oK9LGo8+twrNSIWDmJupm8A/WK6XTtEPIoLuehUcVzmkFzNqM
F5wgoPskWMFMifq18Ppv02IipgJ/foOJ4hiv5mlG8ynhjTfgCBbyVe5WDwbsyKjaQY1fnqo4y8OB
SVtB5z/HkYJqztgDT9a+ZnNWGxstX/8G1Ltckf2hh7Rt4/sSKAl2BFAfi3pSzoz/28N2crkYTIQB
Qyb4ccnj8sYsFLkQ5iiuye+iFOHb9TuDqJhvN09GuNlE5FcUMq/rtKkcQxwG9CHuH+yxUvPuWJDM
jotBq9QqfnJ3p0mAlaysuewG5+4ettPrXx1ysYvcYaXXxY1fXm2GPTzHfg51RGk512bA5posSZJz
iJIKJzNpHzw/eWrBQl265xohCpHH/QMLXWUhTB+vS2UX4cbvhc6/a3FKzj/NQC2qX1XG4xmDwXWf
3i57uxWf+59iMLXjU72RoYAIdqlaOK/6bgvac6Xf5c++HgDClCecvs5Rz4aACoZQIo8oNz9nYF+6
lnlFXkUf76ez17zQy7aZakmOKhpSnA1cx0u3fxR3362mQhFZu/kb7dI+a+bVlPfAjjrzcUzyAaJe
LN6uW/zlR0rRTNtGw7987rpJj5QeLBBlqbSrNF9f+WlMDe61QzzswXXnnl/vVFU8WiNyr6oIuGms
ne+SMk9eMqMiHpQ9myX78KGaAzXjoUxfTzniUvwIEjF+zCfyXUVqCvxcacMOzdN+XYOSnSTexJc+
yfYCeA0o/+K/InShs4NkzEOKXjXIGUo1FtPGbhpmK8VEaLJeJ8FtpDrkqb7DiF1/zLXLmHo8qIMs
IolbskvbTDFiKtTB2S2IH2xofaya1rroHuRGYK4Lk8wK9uTlXgF1sSxs5rVgqheLbaoiBxbDlll7
7sJoV9UuzDks4TKaG1OgyGjDU/3JU4gr9IzEEQGqrb4SKw4Y4xEi2ptLNAnWLi4aOS3Lc8vvYiXY
Ek/3utNwi0Zldp5/mEkI+Ew65jjyeOAcVx//wMugLEGMAW9PaMr3GnH8RpSQYwKE4Y1xhhV5mGq8
vFqfBwFOks8K5K8YPQP8aoSdZQYndotbJVTprdyruukRTy7XA2B0It+w/NcNwdw02ajwtQtjBpTY
zJ0NZPc5TQJy5nwyoL6vZRJzXrbAVkJU17QHZAf0vJ6abAxK9CVDu+aYbl3MZi4UN7KCz65rDnwe
a2vpG187yHCedHbZXrKRlOm6+OUkG4onOM+Y/ZWuPEXw4bnQdVPefOao8GrOYhh3yOVmRrMoAqjT
M5C11oF7OCMmPjrx6/6ndz1oUd0guOFyjLZj5rYHVtdAEcRFiFdaQK4FzlGRN5sEIfJv8stxRdxo
JzDNgUxC0l1nmJp2/6//dbBj+D51s0sU30YKAWB5sv9+A0lAj4v3W1Gm85/4ZwJlPPjp39vz0djr
GLc2UiTq9FBhP2JbMxYXXAz2zBsjBjuAZc26WSFFd7bOtS9rbTwg97uyS6+Mm4j8i658NihY3n89
C7/xOoT54mTT3GRKcvr8oVgH3Og8hO8Dmzxxcyu42uzxX34SJTwk7yMCHunbuf3JIMN8mK7RpQMq
+V/DqVEkEJH0BcCiPXlJC5kMzOpttPbdc4BZ9o+YjUw/z7RlifmfdkwTVUhMhLxPDrKku/4hkcD1
vUg/UQ7HD/IEWKc8LlSggn93MQv2SQhf93vl5R9x3DMxyqWj5s/MgtxzJDIkr+3Pa6qzyoHL+WLm
0CMqQs/hS4PbX5qJIqza/T8NOdq0lz/qaASUs0uSXJ95T6h4WJTayz/MHOh1QfvVTFDZ+NjQq3T7
vGww4N4TG1qMgJK9XZcjZhLAZ5Ri9jdEncrJMBFGycu9GOqHQ0Qmj4p18rBXFnVSmkRag7EMjVgl
g/a9agGUhDGNA9MlzufayYxCCtT4aINWdu4ejpb8NqpycRkNQPuo4MZDwSnafoCpM3zGKvlBTS3f
FFLXCmFCdpAiPvMxHBjEh6nEK2RiOGVosB0ggmInzh/oSYDiK6BnG/TNTZ2qTAlbvay1LZBnNHxL
n+nxNNF0xittT/D15oaNhw8TG/BDFcUXn4bJWmJZEgyQdE5RDq1xntNXycsWgWuM1v40kxp58sAW
FekBVcEZ/CAfCqhc1YYRR3QxgH3NHL2wAksarxqmHf9rcPYmRFtBJuy89ks6juB0ygoQ8yApXY34
lkKCTheLZuvM3GD6JmZ0BDwtF95LUX2ycWpQhCoyRnXFRK+b7M/mr+goKriEg6Ktz3UQF2RmjcZk
phX5WEHwygvs1nOtsTM4zw0egGKjKCJdgzdvNiaXaeR1B04DE1kEIse1k8UQbRfXddZc6eWgjltg
8N39s5YhnkKT6DWlOJ40pP7kSbY1Bpek38m1BB6PTV/nyqVUwP3/NOqDDMoUFM81iVRYC9rHJnh4
MKwGq6BcQnVlIb4zIW9+Rn0Ni3aBHuHFPe5IAjkr5p8F8mOnwNoHsrc1EFNnpmTc3C1eFjoCfmDs
J0UlCJsA4hT2WQfGQhNCJ7jT8HtYMCUwY00BqDlmGpiibJv5XDOHmkKzfF5FYOke2DYtusexjPDt
xzKKnXl5dfx0CX72/RVpFZPJ90JNvgZIWs+oL1PvdrDD0XIm+xlaOhHv/GwRjmt190+1v37JxdBj
J4kJvXKj+Ec8+rqEAhtXsZiPYu7RrDgBO+bUuXF2WzPyQgVuW8qo6jug34OuOXoBqBEWJWM6ZVzl
SmA7PjlpTGlN7ewywJhaY9P+Kgz2GS42pjrN+7i4QhTCfbf40l+elZE3CSquXFY1FDGgfbU7n2VY
pU5F/TVIC2GeOZRSv//Fej1gvnTMDW07GC6/Hk8WLxOFG8dcnsVrzv9wWLgPIqzjDKdRD0uNaU4Y
syhbMu2Q2ImCtOtJT/pfAgInwMWiK59ebV1JtENUpvT/s84Jxm/SirOvn/X7INnKxv9GaTGf+69D
qECU94JHuUaVs7mzIyqrX8HTh7kTOis7Ux7YlLieBbAW++PL9YWMy99TieCUnQ1h8AqZjuFqzByR
5NxgBkjoa65jz/SoDHrJRQ8R248mgETDgaK6bB86o37zhR4UiEC7YiO6mQ6qj97zqGvYa8vuakG7
igjQ9UXYDdXUivqMYuH+qSEbpGHFqZnl++LSJYw6C+uu+4EkA5lFFjVZ+GSGVqARWtLHkTBmqzkq
tnRhq7noFpGTEYGFegPfiqzgFOTrFIdjkbrQeVAer8biyp9rriJ+OW0Kq0dObcd9yLDKzJC/5RQM
pwCdnDPTH/VJd1Q698t6XqYoa7+9ZOQpZf6RPp1Zi55fvO3SGy748kvXJ5r2owSVpTsbS/1lyGA5
n3Fi3vPjFpx1pPC/rJwM8l+GMG1drstbvisJSbrHyPR1/JpCEzt5nitewRJPdIpSUidvUCMX3f0K
HdFUwQlYrSy6nGeN++L3DNe8AsQS1Z4Vri0DC+2QT3oJpt4A/MbhSjhvl4E5Ld9LOmRyD7M2JcHC
G5bwBtTHaeRtl4hjs9GcTybvJgbJFMqxhHIbYc8ZJgDKq/QDeUNAG9zU55V6yDQAxQwyL2MOprny
6CYEZZggMg85+7Z+E3ew2SC1IVcbOCc08huaxdieSxG8M1b1IjKynfdTihibK1Cz2tMgy60NcnVJ
833zA1pXVGzmtEZCopFX5hdgD+ZJ51NjQWqBB5JM5R4on/49MmUOoOMRtScOH1TMyWCxmBd1saZ8
+fEvXST/mypb/4no20vZtuEG06xTKfcMUfF48scX1kjqZnZATevc9aK9oX3LvVA5SX69LreX4Eua
hgIWQxdXRRxrOo7/sFbjzvLigwm/LFix9UCg9tj/OPHfUCdBSaQokidoTErykPyObqBiOX0dTQTU
1k+PbqdVDOF2UMjBmM71x4ahoDEnHWys8EAfrOjNPV93GlTj6Jtbsp/ExrEu69/tQYIWbu5imzBT
LWkX4tBNuD7bZlbmMiqIWdt39JpirQof8ZIOpFbosQXEMbMSL+yGcRU9HCC1QmcOj6mFxhajSjdR
P3Y21HfclSQHro9RT1Io8C8I3inZeFqQpp13dNggd0INN/1ToLBw+MoH9d+nLNefYBzhM+WWWRaJ
agM2LB42aoei6dIebUCifntqSDKHAXSQd5CmliwI9tFrd+JOGMqNIeGxhBvEkCf+mo47zBrUdFbT
QpOcFDGHYZjsplIEFGBs9MKRKolJQ/FF0WmIlh+0rlsREqxICXuHccqhxZDmaL2snplSDAm/qD+y
w8sMaUYtJb9VS1IRed9q2x4zal8nHlEr13gRhsoBWBWhSGnihcJX+u7HaW5Il9DLqtnkKXiZN1um
e44aJm8vidVq+Xk/rc9MO1vTVUKfnndL8f4YZKp8llJG2CmBC0RYNw0HEBL25XHJzekoW4/Ci5/g
DmHakNQD/CXLp0JQ2saXlowvo4bbvOkzO9WO9uDzBLPUXI/sSlpo7sqMhQ7QqlmnJq1mXmJH1HcG
VM+MxWKkdGNe9Nw3brmeH3zC8m9E18rETMHnHvSsGWes5xGgwDHtEVNDocezDHAAqKWqY/m4EC0b
rR6go7M8bxspkSrzfHvHpj37Ieco0YTYbEuR18/1KfjxkWaotZyCrcWUAZcQ4Uqdwk2FIw3cFog+
DTUE3Eo8t5N2Ydo5S559YeI/IPQ41VV0sWqzxQpd/I7T7i6Sn/TQ1QEgiEjcEKI52R5b1/25GPHi
sJP99Idf3JWTreptd1Nh/lP3reqvRSuzbE7c8EAWxjUJoq4EeeY/L0cvESYjhQNydIdDC0xos9+1
xK9jtySlOl/p/LXMU10m21agefWMw9M4gBE7u9BHVr0sl5AXoDuTIgNfuBD/ajN0bGYrOGF7Ravm
pAJsoxe6yUld77eR4qX4aviSKm70D3hwSenJRIuKNor0xwm9dAsDrt9tfehrrBhfGsqBPgRChMKt
WpAH8ObQNf0j1op8MTQmXuQfWyFaB5JO/ryU57bsDiEd4niwE8doLxeELVDr3I4erhrCPHARkWJy
SBILsE6NoDWXBp2fFR8q4jMitGIEUzKj5XJEzlH9zwu4L+yoY22ZTG/9OWBEUV/E+ONgXA3+oA9N
MRf2jr4pcFpIl974JOTUqEkDf/e9Vhr7Zap7wJCrUvLX6YK2EsDUm1hMTAgZE4tyAmhlAZsXf8w1
bKA1i19pJEv8zW3UaEqlrhbmT5zneyj5tlpWKWYtg7yBGqNHUIVypoaCOp6vc5V4lVYSncCQZZyv
Akt9FKRm3o1NPXa4yIA6D1RNuXS6PiwzcHZzaBwpLEfWgoEjEuEru+d98bDkyGJP/uIoZom3rhVK
fWlYHKa2L+FV+MsnqYshXnzNnkdTQtZUrf5JTsd+PrPndZEpsiFLUHDbxxkSIDPVXhxAg3/ndiiX
VGHKAbN0UC6AMCIGBqkQ0vqzzQlHhzg4Ao76vRqls3Ti/YI8YIdQ51TwMC7RyltLDeRVky+eip99
u15GyGrJKRQOCfFuXHA7fpfFuMHiRUEkY8qMjtNbQ16lRbMMOClJi9oaqzcgOTvZ3A/xJ6j8SIbt
RLWL/fu1raFDRTLPxEnH2rBXe8ey73VgziHhLItrad8cqi6ZAe5fUBgzCndtis80cumXpBDTeEzS
Wp1TSgMn/vRv4kLigffSZImbvwwTlNgJmE5eCGH8KxPIR1qmY+XXCfpcWxUgyHK75tdKhy+0ICqn
K591RQE8p2OqI40BEjyDplsY1rMwW4arRFQqYGWPkRBaIRxWt0nOYLPCczeAFYl2SgGywDW80eTY
Q1JEnE9QEoR6wM64WFAhRjJ66xqnXDSW+VVv5XHQYlYSJNTrm4LKtKrZlRiVIUzOPqeCopfnXjRp
Jjg9/vEEPTbNR2sd4SRPQJ64nIS6AmCcItniLSTpw82m/fU05ihlGKD511U/Cd/a8Tj1fS7S1kSm
OLfu5wehp4Ka8VISBv4/LQhNl60d6t5sh+HFIEdRcPm1kD7qr0tlWtimhlO7UytVr44BORHNwyG2
Ig1ZM0X7X17bFNjsSdWJ6jwSNqtkaDV9dLBkOnH4FOxzJJWYlvNLK33Sbz4Oqn9/+uYivbBItu+1
HPNeAqbcDjEvOgroFLR14I/wR9r+q4xpQET4xU+/lic7YvIJeyWRa2XV63JI7Ui0c+MkCx3PDk7L
JXSIAaWsEYEdAnIcJJtcQMyHocN7lopM8+130fAEea40h74nOnrcpnPQk1cdHNXvpZrHlkxkELns
6/TfQYQL+vWvJe0h77JZJyRL3q3KLM+A5oBOWhHu9irwEDuaguunjFbyB2LOjWNZ9x87hXieYnRQ
iWzPrk5CFwYnMps3+QtTQZqr5p9O+AFalj4qBEPJ4XEN4qb05WzJmeLjC+shu3YKJedYiTyjrBqu
9x2tCcDXMHbatro7b9P6xV+9efH8Eu2F1WAWBdhKrxlth6QAOJ+X8akd7AA9LNO+lKP3Yv7whn6O
GoZrkdh7T9IMiFO0KhlvPGyPNmE5erSxOpkOXZBk4Hkxp2+saj5kUWXINYkRPwmXFW/kRiGMaIIj
9cslJHeW4gXtIjMfvWNaDtEgQqM0NaPKU7hM4EFIWBJc7MJlKwggbIHD6lLu4+OqAOPKncAVotSs
VPm5AEUtmTmn2hjSl8GEdkP4eXV7ekD+WLIWZsHwPfLo28RSkwvWGFtHt6WkOr8AWPjKmB+Z9O84
QgpZ9o+H1nzFDL2t7rfFKcJ7+ntCUiBkglEntNlhyf62oQQqtjeaXT+yGEMBCs+1YaXlfsl4i4Zj
l5x21oACGxL4REFQOZ1++NjZud0IYfUSjasMTKX3NtuHxv0YMArS5nkyD4KtlLzShtP6TpVJYQtR
rbaG6ZqhkLUvpnUeQW1F6PF5I+kpmNE3LxTeJmtKuumrIBvPXEfGNmCbQqgWNuW4z2UhH6fjnZiu
AZc5HABn4QKmX9XKeDa9ZMkDKX/M8pXIO6Id+K0uD9r3vRx9J2KfZti8HqIQICZCxJCeQbOWyb7v
hz9HnRpqPAohs6zEDzpN+xpXb27bLLKB4lbSpGTmCIiJKIwURSJ2mErGvpRRgBubNNTpXRJ8aUw7
jihIxEBEJIilttiklUMGKZ8doFIq6Xlk0fGuCByWjHlLnTI2CDKzIeXV37PShWrfS6J9dcS7mV+p
GpmgDTvYpUXWPsSy5m/kLsp8wPprpbCQzgOsVgeRwbeETHAvU9UxuM3fKTZQnOxuP/2iN1dMuDdL
y0Zk1SQSYdlsGagw597AOi8BvTZbU2VILq139AdLePbHl42nn2kLGF6Ab8ZwCuNBHgtI40C/0ZZK
iu+iDCx3O96NDs5G2cefOrO/qeQjmxFSzw29xxzAq2KCAn4iGanl0MipQPlKyZ9gwhsIgPdKdJtB
QD/fOGWsE2glw+tkfY2NvEsFU1rgLireUi0AiUqzTx8xuYDUKqGQCTZ3MVJj8k9RuMPGp9oCqqOp
l/+Wfjmj38crOxjegeA6aUTBerCD1F/83joG3TmwGggHIpMiVENg2HV+nXM2KKpPmLW47oSk6sfe
39VsvO2G6X7nAYWZFJA2ukLRw9ixrqMeW3VpfYNa1fNai2gmpk/E96D4DvPWtwstSF41xg6RGFmv
gtZWnjJbYuUba+y++i5E7Ie/oLBGK5UTrL46yviV0xygKjQM7IwNMFUcl10M4ABsZdcwPaDBfNcS
X5ox51+7S+K0cSOiaI23R05NY6grA1WYIfJzjz0KYyxp7eFeYQc4KenCwe4pFCMIpNJEqJMrYOL5
TwODu/yxxKR5BYPQtxmrDqHcu62zJL49L3Rb7ZcSE6hyIKrR+/KUg6E3ENJSLqBcXpZsxC55vhBD
BUEhoogvclHjQj6l2RA5CYUv1/AVsFpFyjj+kiWLJYc97wSdrdNIPwr/Nu6ncCTFE7t9fchKWcV5
O61WkHI54wkid1QbcuUJHZhmID8RJuBTNIGKm4aFrsU4sRGbjqlALSDmLJz01SXBLjMj8NZRF3MD
J7fxu1f+KXsLYB8szXduaHdbzzODUu8gM+86MoTV8AdiSEYDS+R4W9nbpdIZXlIrVSYfENLnrggr
F8UBxKlIcRUhll1OltR5q+fcYAGM9zivln69L+1PMmwwXU/NGfOUfU/Gbjl+bv/E3h61E2oGErut
PClE8e1RTbciKGDZ0uWqQtEoTZ0lTt2TJmnl8tFnnQwigLtpg29GURfx5gDpetVfV7k2OE9AaKOr
Ha7ESXV5XaK4NJfIMpAFm/m4U3kVxUcdjEjvj6fdWT1s/S4WmmnNcMRfqpnykd6cPACJtvrcYfla
/3QSER+XpOXVFKqcDubp5UNjLN7GdUzX0vAH+fz6YthAa0rQksSnBveDvF44YhmPXelDw3gfg0qZ
rGUEpdaTfKPkN9sRFEusevLTwiQRDX7ip8l1IUcnruEqB86KSOKsHWwL172jW9/E9epOiGG25Ux3
W9JE/8B6aBrExpqnxRo6hJ7kGQTwWBKQWI6iWQvuPZOuoVyXKgAOn4dAmX7S625fR+alkpQkuBiY
goX7XDRYIcwpCBfzNGSF0MTWtdTprhOmF9EOQP3EB/1HQIGW+cCRcDKtZDIDrafJEFSXuJI461JG
yzYkVJGUlwDgxYSP6nCqx/2ijNQRM82SZ8/0U66/+Dg33HvgJD6VMT5Y3ooehIi4Pq1vxsGJvPJr
+JjkQgNPTJpAarMQeiq73VzHqPTOxDUD70JaJJDK2n45kcCfxVzkpIc0P4cHtTJEuBVObT6tuVAv
RNenxgNjYFcYr18g2TDSNW1+uH9HcG2cliGPfxog6pINw1h2ZOgaICIMKWVpe2fM9m0uciIt5hwL
YzlbSQbrU2WC4FfhU+dTlgDOaRrIhyjbsWJY0jeCyprX0gAexKOUmPBrE2NISX3JN1sCMMQI/4Ub
4V7UIm8exrBNXcDwgv8FV0jndSDc7jTuhgHqymNKD+Sc3m5sSgtT1yoRxeLZGoM/7Tfgokohega8
hXYereWbC3vFQWjQtvKCHjFYlA9CmWRPROVpM/JVHqFCiEE0Fg/OGnSGn06goy1Kym0npsjbSJvM
zAwzQpX7VTOe0PPqfeawyagRGIWAFAWLzVQTAhAPMlsSN7UEnXoo6p1vasMXm+p9duTRu1hEpMmn
APySt0cHYj5A8qiEOW3TGwrjJD4xF1Sjv2ziB/7wbo2Al7Nsjk52fk9twLpGJ3V/LqHfPygTQaVS
6eKfcDGED5z19vjA9hR9u161WCM8elEDF+hVPKcFRhL8wNVtDGDyJbURfcxzSlfwURT7yDvDjzy+
oAH7jZiSK+7HM19xzqocuC3qlEyTgGZ4o8rVdDX0PoTkmtGps5sXMdI59UxirOvFfJTUtZwXb1uf
AUkXVH/80lj3apCzcCuSIwIQbMth+ckJGo6peP6IE9yzV+RAsOfahYxen5J7tK6apb34U0Y3Hs11
UqwQ44pMwcuiq46E1XpsvMZb39L7jYq5+h1Njdp5bm/Q0wDf8UucihP/qETukIGfKvlkRDGe6sYP
8sAAx22u53/EkCKHNezw4fqpiM06ZMGez514r8zaNOc3nub+zIs633At6TRcWJSWjy6yRy5LNB/u
Zd4xyNa25AlrjSkQIJowsgIzLhlsezmCUHwpvCKOMqV4g8wtYHIt0Z818GsDDbayLu4sBHt7hNDL
jonQaq7ggnmyDrTEnvqnd9mcAvV1GsWE2aHN02DXGio+CjhlzSZBqCU0I12wrVeeA1HRj5x8bNth
xxO2g6D40zjw7KuP91zWwZGRqxE8q0pCJJcHAsSzKrkzUr0GfF6KttUq83KYfNbjaI1RekuAOR3x
1pUksGsprdcr3v3DYbEa1veRBXlBiZamw3yb4l07XQw1zXPK9vPdkiok3RG+PUQ05E3EtibVxWXk
AElTM2o4dPfIcK3PGlC5S1lC/Nsdh9cQPXYyuybPM8a03sfZ3y6erZuNmv6MqphYFGPD23hYv95/
gRTWK89pc03HycJJysj9xU2eThGX+pp4Z3kwBa2zlMQ1y7FmWq+dj5BsBEuQ83cPJedTQqwefdmD
syWa97vbkUiFkF8Z6N3pyPoKVlIZlqwKH8vhcKN14K2lLdEPTD31+qdV8hzep3Er9u0m3AWrYLmX
LCDWq4oudhm5eLa72ZAeYWUCl3HvBPBImz7kT+GTSgkO3Ztm3S6l3r/0aEjY6QbE+nUeMHZe5ucD
e40Fk6A04s+oDo9KcNLaSbJSccBbTbp1c6uQThwPbBRitFtsuXsx6BXYPrx+QMt4LuxTGZMbtvXz
Kgzn11oi9Faa0nKTQdnAgERc2ycKaDihycpOx33F+oX7JGLMP0WJbvGBygPyfZm6iYYAMXb9E3VE
DgqXZYHl7zrhh2M4pMGIrkhr30nHhKzCNFwMGoYyx8rcXMhr+8ku/rWDNW76YM2p9foIDRuckQoh
Wg44K/Z06THnhWLmEaKcqJ9xPhPA0X2A1QvyeMDIz2fNWys1qWnh6agGer4WQQHEGJI2yFHXewYA
IW1Y7EAu1W6lEZLw/Px0hiKJpnd3TVKg6x0TnXRoltBlwHTBTgewSA2A5EZD4p30fg1638p+B/pK
61Lz6sSoiHYdFfi7Y7y59BFDwBXT39v/jNc4z7u89mqodFGuIp/FJ4JmSOxzSf6hZNc3Bb3m6D42
iu/rVer0k2/ViMY8IiH1T9jjsOt8SYex15qkX+qbBgCHK934WdWCW/kpAmHSNLkxzfwHCki7ok3N
O5HmpA+e5+JeLk2kLYgoKnwV5P41Bj1o/BC2v+RLhGuv2GiZipwuVv2s3Y7Ou3RYBMD3NwNokF3/
DZ8sTUZ2qX0wxDst1cneBKczMmUe9l/mW0TSdRTDAlanst5m/TlIK+B1WvcrBnQuvr5Izksu26BD
5V5Tm2hfva/JxTLi8G8+GJMCNxOV5TsUls5J0Z8NIMuZy1zc6pWyVBxOaf6TMWuyZEQxiPtylGMF
UBSyyzy/KWTkkMYKRZxfWeOH5ldeFPDpX1YKYa+/2EbUYzdLLw9wfhGrudv5Ufwa6sZOi22ZUxEU
egYIVl+WH6w7YvADblbPv09soYzkz+ZWnsrJV1Yhd3qqR3CN6k+HEfhXHwzeGiHTgEbY4tX+aa1F
NXZbgGAVgyTvsPEFfVevIOiWeBkk2ljtRwq6HJziec0hAqK30/X3lU5Zc39Q7u8LyJaXaYRQ8V5M
dc7iQ/q6lmm2KmT7OoFJTQOqQHwQE47pjZVtCYry7yes/5qWWHhVPF/Dg9BKwYuvmy195sTHgk1O
6OdJMFPOqUwr9VyPmsBirLgoTJZrs2XcPrMEOxP66OKl1KOdTEFOSsLKRgOqu/uQjycZ0yDCHu+w
1uepSUqHg8XFmWxi8KkyMGenfnLS92jbwQKNiarb+RPiZP3NysBh9iyWQlT+0VtwbBJMsLlCXb7l
JgYAxHD17XYvC/RUwIDcb5cNAH6J6vOn8svGgWsLXhoIb56vgcFLuLxMnajx4mXgR+h00AqJ1uPc
lwmFNSlggPG3i2dKcaLdsW7GqpexENzupA7cR2WyWEcsaEtFIgH5PJCaMQxYvGNvASg0g2HjA2eQ
gZkbli0GkN8vkMzHelmKnb5/oYOzf/2VDwRC32zR0f0Fh6Wf/M11VqbceEOFBT5uvQ5bLJiHRb9M
a/hK9M8iK8kXggZfwWYL0dZPqZoAhqvyjieZHuCAfwfumJ9J0O4zteqwa9336IAE9h4c+jVSQAZK
jx1cg3HlXlXwp+mStFWaPr5SOerzmOz3CPN5jWp/bDt5Lfd/t1wdFy6uYwws+BOWjMuXreQ9I1Bx
Quy+iHf0Vz1wAVQePOcXlWxCfgCEx6cZqcoiSpaFv8/nbdBX9fPs/e6jRJvfeBGoQ3sOaV9Ua6aP
wzg4hZ7FOHWse0Ze/Xt0EVLwVHa609YB1UHdbcJKEsdaStFcFGy8YJSTYd+ACsU25JQonn4eZkAP
FxwUf/ZD61IDf3JNSbDXEXp/afV/Gv7d2MDvWhxfvDcRZop6dv0Gq9FlzwPQhD6Gj3gwhAohI1/F
obEC+lp/+bpwS9BLNdKjA8TOJz1MiB+GjqXxQrosrUypBYUpWj+dAwkwSLrMLuQYmm7h/x3VjuM9
iQixgmhpbmCdwpiHqhFfYasc3tEQIVrfMP1Jrz5ZHaJ3VqnxT4RbLqgWh21m1QwcwPil1YlpaiXV
eM458Ybn1RatKgRnxPeVI4HCHxtP0RwrhvcANnuMPqHHCodA9CN75J5ytXBQZi38GFmpcDJzPqVX
dulPEUKPynV7K4/hkgrbgzVsxPEf0Rw1ep495TD7kQSnNdnWlbTYrebeIQ3GHsBnWf3ZWAddfF5Q
fQfUxoomoXDDv//nb4L/rD6pSnnSHzYZ75aPFTf5OUArSWLwEmTNIuYzcibuFMdTXxOdCBPlFndY
nHfhRv7RrbCNl+8SXtKwwCR2B0Svt8lNUsNXR3AumGdQzViTkWunw67lCgYzHtSFuUGUMF0j0k9t
BaqRv5aNCVr711p/GqS5/koGBqLxh0X3lMyXUecrFZDfvPiGNP72coeVtA5zsa/rFlBBUwa5qYg0
s1LxaDQALzvoVyC1cELS+qJX59CNm2Yj6+j5TItDnYBbOJXP3Lw/mghnW2x3OBKDk0FUFw6CxzKh
2dWjVHzObzHLlHr20nkxOgHtDIT95je5n3jUTYjgtZh/Mk9zZctyahajsGKIKC4yMACfW2K6knzM
kovTIrTD3D2c10mMWs8L+fU7x86yeUzPC/cIqJV3POA8Vxc+nu5S6mEIBHOXMBXXUYumXfBDhm7S
QhTNybl7y8Wze5DqdCveQ7JegqoSozaa/GLqb+7GpBamQ3oCKlZMtMTy6HOC1iCL40MfMAaIxUP/
IjOHEhnAV9uT1f8hnoloerNKPazpzGzS3KKkuI0oKZYYlp5AG37xY8yCuH5R3b+/zcnV2bsMfRyD
pEJj3iBmrq+qWPRRIKKel2nju/K2WN12VsGgtqpUk+vLgkrbqBjxWcrWx2NO/hrnQZGD2tX8WR1I
VE4Uahx4m/MPsRbErNWo5kF77SZgTIMRbnBnHxaaX08t2f+LV6ogS2/xuG3DOrepQ/dTNqhCDEE+
5nOL7kB3cc3jK/OGdJW3/irtOEdenUB8PqDp/HWX/m+L1XsWPzp38p/DkSmN1WlOV7O5p/s7qOYa
Nd6vq4TdV+TwrRP9r47Tkw2YABu2VLHKrE+UkYBpLtrix7rFyE6+0CbkfU0LN34ITx/CIBLOhzwZ
WCGvKkC8e9BD15NQp6CTn2HqDYCYFOmZwXIgX9bZ2r0hyXHI8wEBi2zfwLe1ssjievNjr0T0b8UG
C9f2lm9oQ1LJOFEaZzbMlRBpZz/Y31wBdcrqYNtgLLiz/MYNnXXOP6U8Lfn6PV642bmVfPe1mqI2
1GUwCb7l56TLha7VRW5kBu3xrSxqW48EHRXSZCHjcZmQWE9E8IZEn5f/Bt1VHwmzTpSBbKXrKt+Z
YuOpSAZIRdc+2f0U1CySuciqMwZRkWz4A++OFbZ33frYl0yMFZbUHtnPslt4BMgzmEtHXX2wV51J
T3Ha6If3v3RrEX8wOWchYWIUg9mWF5HOq9ohSAKSqDRAkr+gRKFFEJP35I0v3SM3m9+Qw2j6i0L8
om/gRkDlgdLmbfTqQgbRCODaD9Xfv5pl2a7pLI7WJj6s6fl+OxHbo/CB+FLFett70QtsuiYlrSxB
Kp3oD2cmHq4Y33Dpu4+O12tQO850rXOKWQheIY8CPsJTiKrdQT0yPebqwojpsDVFRi8p05RRzHa1
uSk2tdrXuvDWAim+vUEIHQ96Kq/52tld3HoJ9pA5eNjTcuNMcIGiSJeykf35oCNUC6CE4c+vPYvP
uzINU2ZpdAtxrVe25r+T/zIl7h0c6Xn06dVcCA52A8xkPN87+FVpBTm7YNeeYgSUe3wV937GAPYM
a5oce7cMX/TZJflk5mCP7n6oAmqKjhy5lGpm+iWQ0lNPhM4iJB1k7Qh8GpoGl3qSz5+2u+/60GWL
itlugxgXRrwiCWgRFVrntRfK2d9wwDR+FMSSnQUOVuroAVv3GS66/HbuofVBVlCN5b8BkH0haOy7
CNUWxwL+U6qRZUkW0ecSe8yQGO0PGIevnO8LgRAk7viTlS2GID3+1norC+D3r6bWsEliDSWwhsEA
ceFJGyQGlVJQAyZ9s1IxF6Pwhhf4L6aRkd6SsCTP9YonTyFgbkoHWhsYv9VUfvp/aYDVqCEMXG+G
51XMnjjqWcQcjZhg9kVgnOXYh3xkY5BaAzJlT766uBrK9IQz5+c1DvIi4sYCig5uZbBmlkIDq5jp
yN+1kd6PUqcAuwXdEWtQH18fz4qIRzaYhNnhUgtSmqOzW1U6wrD9GVd3tCOBvViy0yrGYYA3uNZg
ZVbqIwcZ1crhOQbV4Nii83s9YZ8BUOaxkGsFpMcSUjQ14WKHfGTqrNWGg/lsKefzS9MbI0qzXSow
qKpCDjubedISyggGRXhhqjrsVCQdNWvjV/lDTBXjh5QYcRB5hvgkf+v6Pi2bDeLq1GcUpb/9Tzv+
AEWBlsnwYabxMZiUnFaF68U340AsJsixoCpft0HVjTOkZ6IozINjfGslbLdPcgGxk7zRc9Ci0ZQF
yH8yycgp3tqtaKSTjcD9xZ+Q9Zcs86jLR86tZm9/Sbuhj4LTNR4VlaUKivYQ0qcio9PjUP1Suwv4
O9uXXMIR4e/w1RCOFsxzkrGuvDWDuWx4mujwEguwWQrmM48zQKy/RAY7XzEtOjRuJbliPRZM2Xqx
XiMhOWToaomzCMnF0i2utPUusBh+7VC0ZWxqW0Opdw3+LT5h04AK4FZCFITktwwbDimdxNk+S4ic
r3Ev8DZOm1QfNfjdkaHCXvSgF9A7mpw2P8npD0HMqcbfDLikUaLOQLyb+dgLADgc9TngOQJMTKCD
iI9sDTS+Okt9a6Mi3wCB2VxI6rzGHPSiJgFy+oj7DLQig3HEqjCYegupqKSHvFLRlLidLuk+WC5B
rvpglg1HTfgGAcp5cP2sDmpN9MKDKlj2jxenz4WIkdhyDQ7MLkYiWIq5mckNHjHamsIdKtGMQqO/
sdFop6PtAc8SpktsRiu1M0v+OIzqt8Q8GufdkNVNl++SSGm3JxwRkc4mgeFGcb6MozZh/qGdsXR6
fSheKjUCjmW9BFyHvJfovNo3+Bl6VdDB0cIqI/yBfcBFXzBAcFT4kS51AEf8BOCALAMwif9XyakZ
dsQ7eh4WXOsLfagg9z4hYI/qFI85Pr8XpQvU2gjXtJRQK9XYRJ1VEufJuBF7Zdflah66pQPfBbLM
20QPxCaCJmJRhv2fzO9RgXuq5uJRiomqEFqoAOUb8lBAKtQsFu5scR2rvf1+vdSnaRz8mlUd8YD1
1ZGvidMpp3mBqC4rq60nDm7VX3nS8Nc5e6un7RKA7aRwQ10o52j9C8wIS+8uUS+f/S8RAbQ5vc9w
7MYU8Xj8nTW1eFw5LvDFY8Z7WpvfB6kyCSyON5IZEzuoHsVw0DaiYOYhe0LcmH+ib47aV4B75c6s
gyKtmCR3pKt9l2YC/xWxFGxQbc2Wt0g8IQYi5r3KOEVMmf0Sq+Yfd+t//Z8PMNZ1zjuX6DDVy8nt
G/KvFmqiLX6XWQ9wY9P/SiaM38f6U+qFiSehrEBSbnVaFTbWsmc2yhZqMvKFcLGBBLuNRj7A9l+M
GuYeCMP/4m5RILUbVLYVlpH5EJb2YvynRHp3G6SUZf5xblRenmE0brWN6jrid10twTnTxgx3mPQX
Wk95o9WG+HNxIfbfFozaEkcsE4HxPxxfR/9iA6aKjW1/gTZSHbrtpSzd4+DZEaanx5B8FQdLhYcn
5ZOapTTGiut/3sUvvy/o/0mvraggYDgWWOLZALOLjhRFZrTfxY0WeR+DbMydVyX5F0AtOnPjmVIG
v72bBTEukToziBvTSlud8VsYoOpRnPea86QHFRTvGwLwNmdmNP5UaClljCnro94L3+AJY3zZOqbg
SK0kNpa0h5zVncjBOyLI7atvBvb7pNNXiM3d0uEIQ+sbytoVxl7K2J11+yn5Zu9I9smBtg2hgBk7
Hp/yyqnP/R2Z7lebN/rKI1QBgpijvyR5i89VBB3futCM5f8nXF2hHC059y0NqsrlA60CYALlmKSp
KoIVMPtZqYjD0prim/i5GnqFEzPAknsQ/MJIkhxRx2v7uRqgs3JypZqLNOza7tsWscjV5I9hGM5A
pZQ4j0Uvxt9yuBMW4PrZIVusWuiqE3jhmuu4+910h9eR2BiXLuA4P7qkEvJqzN0UG2AFZvgcKEz1
wbEFOAj171GS0NAod3V2TLQeqcDMdaZEse+RWABfwIxxWP89tKdoklOkcyCN0GVqEd506I0sqCY4
+wenzWgKzVvuBWlUA8ZBYhYkwEAMBSDjlxOVpbmFaa0VBfVW4mGEebnL1LbmCNK3Eu+lZsCZZsOU
nuDrTUX2cTVv3QgkOtqFdvHwSGSezqKdj1zEvk3U3NncYwNFEdBMwnWvXUiwAO0oPS/66yaeZ1lo
rPIH/Sl7nJt2rJC4R0CRijCil6/pb9/lHaEvv/KDVyVDeqf1iTm2yyxKny5tKU/Yq+l+UcuGIymU
jFGzAEb3NXDwCKC+1MaD+mOXpMXcFRWVJhXHeahNxzv5oSwpaO8GJoOj1xp+/VHMj7y7oplzqKf7
7wNL0AnkprTBjoGKbX+6DnCTtMcpX29W8ct/uDlle9UNpPYguMHW19IdEstlDanziBBuQjZju/Kj
yF90bTOxLgHAqrzbFTjuBuacf5CjredMGNYwtCSH9pY3ToRXkJv0+22Q8x42sItiq+sR3U5vEx7S
pf9c/p0MkBOn5hmCzBGuWZYO29JxX7Tvv7xdd+IPLmwI/sPCaB8ygTUELM+1nqBtDeXbJvsxtQwA
L6rAgy7G/c2o/cACKKAE2gzPRAwvcKIPBubGm4sUeA/9GCvSbp98LbiyHli0MySwble74nnlPON+
fYGt9GjjomYpnl67M5njmkb211K5ZDPI7HXEfJ60h52qL2V4DE0tZD6BD9qkPkWGQMgmkMQQlN1G
nP5G6YkYKGfCnq0BT9tCYj0uUVLmMwWTRTopmuqnXpDGUBdKoPrsgivLJxPVRscPm1a9anRF1EUQ
EcJNmlFt0TkvL9jTc2nq8r1P4x22VRb+1+5dlQmreh9JgRjiHqzxJmOYYRm3l2zudiSo6opT2N0N
Skn32St39T30U4po2wp+h2j1Pcqd4N1w6UJa46cDvPqByfHvtoiQheYlizkw4L8NAGdkYQ4VsZpl
1atC/obO7TS7gnKT7/qqW1BfFRbjIIbZmsmrxwdQmRo5XvF6qB+1JFInooxNvk8GM45ngK3i8OAk
him5ca/WnFt1XFp/TAYxPrEeO6C4xL9kDL8fjudcoIcAhFK27/v5QLuBZEp8ZaA4ALlkWR0Pv6Aj
jU99BFA6WWPWpewRmY9EDqvfRJlAeJzLoEf+OURjojyW0bdFzmxNBlMVnAQ9BcAVpGQU5QA5wyVy
VVdsHKNeKUO+ISn6/fMJ8ofzfe5hbrItTPvzrL14+CctHyg3tBOEYFgZsexS1Z1b3ObrsCxImAW+
JT70/ViTBnw/ZjrYSjn3lJu1asZYA35j6RUcpxbEYPdakKrcvgOErcRbHfqQdgSMOStcALwLsfIP
vWMU7Ff1sflG00byn6LrgxvV62ri78oI1caoVnB16ZkVj4vemuC8gDtykYPRhr8xKuXRlG5J+uoJ
9hoEmdgzZaModhwv9Q1wiRoshGXEVf5/jrTpk93fhgsNqrRU0CM36Lsf2qQ489v44+qGRe61LvvJ
5MXU2MVwPRClr/fxuYbxek7Fjc/3TPi1956aCbKBj+GhNtFwz1yJVOsya3OMvf0SFxpoayn2sueH
qaji7Q07nvShKvi0SlaQjcJBGZWSdCq8FOplDz/OH2GuMU9suKFkAQBPdYI9Vk/1OaEJoKjXu8A3
v9iIu8PSNvFnHWrH5UZCiVXiCjYRdIFGSIikBQXvBfm5mxHWsgqpJ+ulTr1oQ8wjlEKoxG0CmiBv
5S4NmF5u/ejLvmSevKXvgKhWzqTGIP4+COG9zi7Msqy+kTAtOqaZq1Kj+96YrcFMkoQ4NPgGNyLJ
qsfXgRxuyPWtIrty8GvRPE2IgQKAefvriubhWeTSQQ9orhfgAkZtqj7sYiDrLXa2fj6F0kqjjvlw
+RAWg27OQ2Aya3nBOWM/5Oh/6xR5ghuKaR1NIB8vHkiDKaeFxhqk0q9yWkZ36RDNMNDbg9Ljah5C
ZgaraPBjXY9eFh7eW0q+Mj7LjCnHCObWfngIUH/nwVakHCGBTu7FwlpxNS1R3qrk+sWOUdKT0T4w
5xKd3UR+GJ2JkoqFIC5gEP7/gC6kQRI7v3g/eItayBEuJ0kTwgnkA9J204Nx7jmW1ErmBO9ic0aF
/QauHP/j/1B7yrdKd7M2czjM/+0pbFUCOy5IgUU3yo8raefqQd3Jd0dklNc/+525/J0cGJLDNuPp
ZDqd2Muhrwy4EmIka8RguiFAk/WVzhl1KSCsfNwMgF4c7p/zIh9PPR489yTg63juP3t/XSv14jHJ
y7z7fj3LuHch+zrcSJulwu/Wj/LN+rVxOyAR4Lo1VGK6kRf25+nSTPIn34+wiDGmBxAP0RvijCT0
Z1qP8rUAweWX2fASkkLJzfM0lBfRfrlR38phmSHRHmN0Sv0UsS8wpwY7VSwwHPoI1zNfXixkVict
/k1pcgMHa/AbSDmia4cOndqwplHGX4Dk0TS/JVAE4+urn4MiGsJwg6D+1ohkQ6JMTWYzKtl+KHXH
Cd06zCQSq2HuN3gtT9B2GLsmPRRp1NIMujL3RJtOY+/kBLkDniA1Ubjxm21ELc2j56gn32YwBg+g
3gDDZ5kZt7ZBk4itP11y5UA4hSrmVkSiDAmg6TgnyPau0bm//rhP5n/EbAR0vcqatb89LT4C+bq2
8bmGLnfyZofMMlbuWLTm+fEBSquVC23FiLkHRHP1+DjKjv+E0JhqRC/ZbaKB3dkPlulrMNW6oc8d
vXqJz2l5J5zC6ZARBNGkKjl31Dhw5ufFLLbn26ZB2sYtvVaVlZwlTmhK4rx175wUtSeAs2CiYD6S
D306AJrK+FGEG99oQMiG4qjJLlpI3oyHBQcbUGiPKTJvLpYIVdtoaDFMDAV16kSO2/LUqQ/I8cFl
Ht4PD6IcpVrOViv/F0GHRF8etzc4/vox9WSc6Y2L+OBX6DpwwdvxZFrH7g78kd1W+5BiE1si8bW6
t3TknJIdnx9dR2TjvBlRS28kMgnIwE4ZvIsUTsoDTdP9Zw86nNf/goCWHpWOGgmrSXpOZugjN/Wp
SvBwafVls4f5ieB6dXJtYSCXdRVvK3oB6U3UpOkrHbQamOBREkOItru7p6nlk1sctaB17EGiutzl
L3NX+cTEyuJIvdXsPTVVc9BprUT1Al1loPTCrJOqxzDqTNDPFIH9vL9yYj5syVtrmqUbJVutWwEX
gRhSYVMp0VhMe6lTh5JvV3kQ6S/GmvMLYPWdM6PZO8d9afs9WhB1DYpz6G4y6k0VKjZqyxx4dmu6
Ubt3Q6GFIW4f6RsLEvhAJm5w7SLw14MU6FdCAvd5vEiSCc9jMs2wmheIAEl6aOjTIURo0xUeCO3K
X5A0YBoz+qirLSz8/HpoPBkljKfai5sGYA+ABxFLekmj5WUUx6ePsDUi6pTfzIxNsmU/ASDD7vMH
TAxo4QhFLaozwW5kHiHozOlW0l56roTwtFGFKEWsgfCGxIl82B03A9NQx+X6YFjOC3k2qduYKgRZ
YaPepc4uf5uRQXGXLLGJwuaBc99ey8saGRjx58HryDHscAhRPfWY7ldk+3uSM7g5+875HWTeh7wq
8D0WxXsvVxiOMVya0YCBc1jfUw+OvC/loDTpmM6l2MCOmQ+W4tVfkMN7gHV7hFnWOwhJ1is28R/r
fwbrUKafRrwmUa639hBqgdYe8cl1kOVidkpFbOVUtU6qU3j3JVq8LqTzr04spO+1KrQYf1CeTrp1
HUOdf5BNOEo0O5Sq7plXiOVcs4LJzameXTX1wkKLxiQVlH2XSwp8XnX6h6nRhY8rbsoZ3gNE9zvX
38uRTjjnytFY3iqyr8ednnhE8tlmrt/1WehXFwyV8zjlpVzvqHY7sQqURyVCgPsY3NwUliq0xzrd
j8fcbG/kCLGn+jvqxZeSKKJA124gegQynCmsScdYzxYh75emofQx18Hlv2Ps+ZF17yB2LUzoABzK
NCvLrlTBexaU80mr9t1qFqGVG33iWPtF3m9VKNXb4cNfIUvyTvxdFLjoblYd4hFuBCoWnfYaFKwL
yIzZucRvlngo9XflyZC7ZrxqhO80exkXsZHxgQNNE2NT0NQ6EF0Zau1S9EDMY8q+kaLyTbGpSS1t
rOq7gK1GkBXuIChaZx9vECBi325P8eB0DS8JoNsBWe7+8Dhh7zIgWB3CCmU1warx3/8o8C9FlpDL
Q+/n+njnmt61X32VBERQCx4c97fIeRBu/3F74Pb05ltzFVWelTLJ9IH2zQqT+kNqNNDlpAKHXs9Q
g/JrlOt5CoIktUAvT+o27uELTL0yw8wduUPwZ2B4lB3+eM/or1UMhMqxZPyxZPhLe+OTz+m11pp8
kWx7Nmh9m1Lhq67qdjuCynacZ61J6hC5Agxl+MaycAzwK++S3Ia3E2LNQDMx8AqHRUSfv+cRvq8L
1l8VMYAumqxKrExDTOTLjvNp7kIVPyswRdGFOlnTWXHAfFp2rRjJ/bTMF4R8ZgcDj3Ca028uWVtP
GuLTnvgHik+hgRnvSJXy871UiWP+6kVeP8qjs099zdx5vzHlelRD2OjbSeVj1iSsxdP71tgM9j8+
VbTgTqZ74wTjBsCn9bq7dAZKsSYnrPPcd2f8hW2qSBd8eMiKjRJgwF/1fvwIdWxYRCh2nAJPtmiW
IaDYPuz4CGKQgHrXeSaZCykLgZ7mOWPQXcu5497gDORNxhpjlBVZsrMtEENaiefsAdr9H94bVJ5R
eBB/q2u4BbQUqMS+SsKAmk6uvip2gCxf29esZPej35MwE2h12Z2ZN7j2Q8ZWu+30R3zoPlkkrn4p
Tfk/Dw/CNXnbn1a3dAzxZlL8TAlzV8mp07bpeIAeKeK1mvSev8xrkp3+idyRjqsaKGcodVDSR8G5
zaQUXb5Dvo+eR5KwrGbs4SiXjarCDN4O3NAOA1+JpYnc4iaScAo5iN3/HxG1B0GQvezAEmDK7Y94
AdNVh/K9qOI9xVjKF/97hAZKODKjX4GHviaOrgI1Xy9wpqb7Bb+XPM4OjoZM47ZZbYKCnhPoudUu
TQ9JzXaJe4Fokja8QA4fLXRJWyV59oioLIEmcnOZNxAGP1B0qE17daeBybZ8rjMpV4zp91SKZYAG
E5bxdzNCEvKLN5YBCK5rhK1z9evZ1CRQw/Rd7wa1nd4+xVFfkKJs7cJwkgIWdDmUovMyAdPEtVG4
8SX4R/yGb5ozyKQ82p7QeoSkf3VR+oDvthMO1E617w9O3fJt/B74Jus1k7Ill5ZgfaLCVOeAdzxs
W43RxPIjSPPKua6ITwmqV9zMnFL0BxdhsiOn58WMwTTRhiWoHgKbGIO03CbAKyYTnNy0fZ3in1a4
GlOuarxk1GQbMDwZjlhhhpEz41cNg+7EbWMS3Kf1ZSWYgWppI9c=
`pragma protect end_protected
