// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Umc9GvJbMA2V1NMA1Ws4SQYmLSUlKKg4qZcDbYk1TW+2qveQLSzR2dhIJMPouQReW+G9EXt02/Bo
TkDwLZ1dNmtfacM92jFqr5EmoHYqNJhd/tH3diQTb3mZG5dt+/iqapLzExH5hNdG3HmfqJe7Prta
Tkb1/XpnooFIQvV2UFtQYyVFDNsoboF8RN6EYs6jYeDVGGyQPwSybTN8rGYi0SUvR+1D7xg4M8g5
bpLSDccna82sKdMFX6c2s+b7y/pkDZFq8v8Fxn1pg9GlObIdXeIcaWVoHbaQ/nw5Nybj0+VEtnma
WnORRd4dQtv2nn/kYioTFeupfz75TZdlwqTG5Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8176)
6SxT7TGrEr/gtNncC8cA5q+UhS1tGffau7aUAQrev6l9sCXvcyrsP9Zp656c5je5vsW2rmYaKF8O
iAfIflfPFczZ3dIERDPqVdJAdVV1dU4CamEeStgXqz7oyRoIwyGEhMwn3Ufbwjj/j0qVo6QlRFAc
4+vs/7Wx0wW6kCx9sVBJnTh0XpHvsE0BdeBFpC/m1agGdDcG9Du3T7Sdr163dbZUyVKj/hxCe6c0
b3YxQdcn1iBnaapS3OJ/4m+xW+xDLKwU2MtKoLW86ppvZI82DzyTsSs+Eo01Q3vz5uIWOh/xHOBt
wIkHGsXrCcfee+e0vdqTSFWmbeopmbhk7ppXUxpGely9TYFIP5f3WN1qLWeusfDGXjpH+48t1zwY
rx/MIgc3LLXROjCZgKluwf1gKL5SnHEKXPkyxN6LbcAVjqr8nLImDiDns/jhPHOyWT8jmiKHC3iC
bptpAG76MHaVrR+ucSi9k3ecsu0WsF8ZCThtsJ9Hxip5To1LJI+ftp9Ap6WjkVeU6i59hLptFU9j
Wk03yGW2ldABY1FwnpTHz8snEM9TgH8/xi0dv9sjhmIz5WK0tOG3OUBx+z2xkeud5johPQV3SR3Y
/LhPFp6LNTsbAefoCQkZYMHQAjKcqOrxAq+31zwqtzDIJhutrjcaz6WNUt9NklhMMSt+J8h+b+D7
Rpu3tC9Xl+/MmDSk4mT+ZStquGxZUfc5uQgS2JSdV/plPv6h1UZJWZ5P5pjVMaP4VutxRcIOV1l2
toiW5ubmxI7Y84sEXxPLbbZgzTkJURmLkeNdFGndwPhCkgA1O7sbbhpLDFJikvm7R+Pj/SkNWwSE
PTaJDsKopkLFrQ5QyBGHn9FBzJtSx8rL8+ybDqcIoy1TyT9wXff5OiOqrjxJR4hwj7mp3fRhmKht
dUiZAv3KDQ7JeNqdtCHVvApzvyfBtEUolvN5my1+QONqNSC0JiQaoyvkYOVZSRHsNeS3l2cRq2sc
XkVOM+pK1E41mUKzA21wRkN/XzC73Pan9TfT6RyWtdefi/D5vUwInOwNcqncFJhusoo4qax7ESVc
6QQjzFstgpeSMdwH06YlgpoyOrpsTBWZaleEkVoQPhnvgkD7U/uIIpwKB8qicPc5gWoOQav6E2HH
RUj+7IZDjIXlynKI2Zqr0y9InPhVC0UwCggxG9+rgwF4z7N2D0K7JGNMGFsKWgC7Lp+1OnQEiSiF
2uKiz9Jq3ktkGlSZJAjfuKJUb149a21+2N6kSyDVDsRm+gxcRjakrhbtJUZI8CF8EmbUjyQ2cju0
yEPz/LZORL6vrIf0OrNzryEOXJxUgJT8CH3XeU9pUzAMX3sBFQvAbsyayyrqE3WvOLevXSsTVJBO
gYYpDP3PZVpsm3H1UDJhQTWbCi+6GcJWcwFPX/3sn1s4TFAi+KDoowj2uctjfwJQb1pNldNQL1mz
ZP0Dn586gHymo2TCFymqWWO2OSNZEEtVRqVDOzo9162asHVVJa78zVfdj5wMokT3JguQMrxR67b1
pkwf2s2VD67G0KPuyrPd61pehJ9ggKl2wFAHCvQNgV2Tk0ldZAS+T8J/xudWuLUrkC97tV1sO37C
Quplvc9jmxyQrDLjZ1RJY6XCZzDs9wdd3kenFtrMPjp0dl2J6Rkggd223SE7UfPzU4bzsdJL28Gx
Ko+4NNhMrVCvk9mFM+oRH7dlxeEXtfQEN1gAGEcUiYRYPHXHABFrwsh5nSqOKznlUT9zLgf0P7GC
4lYelUWTBF2wfOYov22afXmrnM6TgS/WLc2JLJALZg19FTg9VWX8N8PZNysAQtAxVfoVaZNII2Cl
S/tR+GasoGijILFKidPk1kVuEXjxKmZ5nj+TTVAQAtDEcrQBkiBrIGgPj+AFheeJ1pYVUXe5FB9c
0oAiMJj13IAlph49MzoIAOIY9ur2GmI4gF9hjpTAalWe/jyrSCCKhs5vQc5ov8D4tPFLOXjI/Q9Y
Pm68TGS21eC0OHvJ3/uub9HgXkShybb9kKTo4B13WZqSN35PJs4wBIbc3IKNl0EhdqGMvspa4hoj
MutvZl6Zt7+HuUrDPj8A20sQCGlfL+icmlDaP0Px8Zi6D8W/TL9ucsK9zqZDYw/TlYWpKX91wE1T
AO3L94E/ZUyGRyj0BarXfV0B9s/TdNMFuk4n81P+ZNwxrEx2o1uv9FojnHkL8UMevqtkphwf1yG0
rHwh2oiSPKMItfhSrGU2Pt60GjMmFOScHRnB2FXlJlAusRbs422GuPuAloNtKGvRIQ2x8qDaMLLh
FAz/aT7X03HdA/L2SDLNyM25DQgw1Oi0MfDpFCpllx2g9BO4kdummCA4wSpN1kyR4F5/+ckpgTSb
GpBeXtbpbxfnBA9Nd1ZkoASD87cFGolfFl99x3aWyEcCpEKuIblFEJJSFQM+Qh8nboUxYbC0YvCB
A621GqsZlOYS2wcs+s7IhMC9/JbubhKrpd6W0+F69s1fY+SrLSHZzsAK4Ci6NgpL4rvMg3JnutmR
OFOKhXWNRyPUuI/m1NXEeriZ7Nqjerf3J7G1cGxIJR/cXuOD3IvxB+OEaPt2KqndH0epm+j9dxbz
35ewlqgnuYZUOWzaCTn7i4dy0aQgKovPG4HMefc7vTQWnQnPeEqwfiWgNQ4n+kVsEzODv6bdEF2Y
V4+hGKBotNO+vb3Xa9ErdDLPMN8L69g75SBWLm622eNqZLT0yaimxyZpJh1MNnBVgdniLoT9TVRp
UN6YFAqc9uLwnJDR8Vh0xIDP4YJBS/QoIVaRRCheGC1E+vYnb0Ntq4b+YozUYwI2V++9hG2CJni9
rNmlLiDgLhHPVNGeI4d8mP1opXsqWGTV0x+42rnYU1czKrlyHrqomKTvSEiWWMD9OTGIhb9Hux+j
xplW6qXjryT+vfZ+i+/QbQyXMwMBiQBv07XOzcpO39yn0W0Q/G2at4v+YcR7/rsixoawflO6HTgR
+HlQqmp2xKQ1peVXAO1D+8B1jRrIhrXzVvbx4dxU6h8X3kibzyj897LgXSvsQAfTPU93nEy1TEw7
FIJQim9XQ7b48ZLkfgq/wh3MCszaryW8wfdqT1/j2LOKFQzUtv8WMch/Cq37mjAOgG0/l12slG5X
vJbwtgP9gBRea6oelxrzbYHLEHVZxkIbxJL99JPYP5E8sBR9T3+Xx5ZkAfSDabIJN5ySJYM6Tl3l
eym8eFnNjP/HtS89Kq/DeMYWcaNcJUcG+Co6kodBv0QXXHenghtao6PUMXCVZzq6vfEcqmGGvYsT
7b1WVpRi/v0t61kKBDQkUZluVrrDfSbi2Q2a3WyAdiUgo+iefeCEYAjJKWsXcd9qhsLZIerbjcF2
wn9vEZbiQtOS852QNOzaVPSRBQvqv2zrVXpSpd+wJRg8YEcCcrUFPCMh2b/OJ5POiNFA6qTZkvS0
pnGLSEWVN9sKyhp2DvWGzK6GsXMs08FKKP3TvMfdyFv1sfbZE0tkF92oD82/Cuu+qWdFFFe3SNwm
gN7UQTHBE0FOPr/lr26DKHsf6SkaG88v1rHg6UXxthZEbel4G60nd3M+C6V3TVdm8wNhDF6O7+bd
R6so0XutXEFz8GrxgmMt6S61+dBUdtzDv25MBG9eyijwwGn/Ht9EqVi+CPH9slEHsAzX2JUVfThM
MAVSK6XlEZ7DGnwwblXq9oYUSEu5cWwd4IqH5LAAkGDquhyi6STEIbgBY34pZTQ+EOCqT86k5jvO
IWscqLt6XQ7nrK79zoxqiHd+Z6ouGp1f7//7qSuXK030RX2/NyYtaGKJQ/FmdIq3VCwdq6p/fvCX
CsIPb8PpnlwsHLAu0Uqubj43vDv4YgIZ1KHx19UyXe7cfeEmzxDWkXnFkw6Hg2dYlvYuMqAu+ENR
ni4bHbSTrxxhmzdVviTmMGsOIx/SZ0riNraBWOXhSQDhfxagF/KcT36KrdDQeBJtdg4Me132oKc/
VUmI+yR5DHJ6vLtKqiSCB7J8OkzNsxzMw/HJeKyKON3Ezoz3OlGLhKDj7jKbluVXrjiqRy27aPLb
ixlBhjEX/97Royp990DQrU/GZ+a/fftiiFSKwSlJXQRR7Em28F54L8mPUNgIMf4YE1ACJZiSw8e4
eActxRqShAs2SSLBCn48sXrdSH8x9BI7AqFhJzz+QsRoGDb+mR19Nqan8iw9XUwGWzth/Ole9dSM
a5EaNsI4p2cgtXYAM1vp4SPgzKJ7q3hkL26zcPyQMdDbq6CrRZDAkwUa4BZXrArkXWvuMvBkjMKS
0iqXHrgxRti5uokD/mAQ90UXFl62UkuFUUszo5UedzU5iqk+P0wtm67l0r86/S0wd3201LLQQQvI
gISUrgN4Z4h8IXzuQDKXZdZeIw7awtqsj6V35yRzU8z1Rmzevm3GICZsG//k2neRgLhh+kd+L19+
kt3/+velKjTsF0n5dxHuyJFVJsqI3VJPXEnFrP0ASsxQi/FS2iCANkpE8BLUxAuQ+3AIQQhTZCmd
794qT9c/MIVmjFFZf0nFAc7DTLy82RZ1ASfEI+K+J1ie01fIe6gK/SNXFEvshmSJaswl+I6ku6ob
hLcpBBV94uRZckY64xooLJzA7Oxa8PAzvhlasuSimIeO+6kxYNunbQH5rEB7pcBKekV9dvQkRuBg
PvT2fslRpL/q1+XIcOMJYY9FHyLy9u8d7b9A+w29oix4bimDlyS3uYQelvb8Q9eNpz2RdFmvdqi4
A6CNLxjSB8N3Fb3FuWnmIaG/vfnD3d+fPJz+LXC1au58ol5swxktbXJ0AsH7d5dryT2VlZ6hYwGH
wD0a5MSuDGJbqBXp1IN64AgY17AQOlSKnqfcZH9jD+9j3ybd0bOEpiJWtOXY6119RxbJX+atOgsC
MT/R7mJrgJZuSiDyYn/4EjFBtEeVYQnJ2RytT4AYmW31FMCD49g+9nfGpYnvu9fokBC0P61+/ucL
YoGwvokStaOhTfup1GkZqsb7Jki3bxpZCynN/5tcWZZKicBIWJw+Trr2HdBpg6fEYaLHjb7ZZVsx
HG7PcbqiwSMMBbwT75gxeqE2lP2EICuUH+kZQlfhp0sWgL9gQoa2tXLoSkHrxAYJjxOXeG0ulZil
127eh+UH8eVjwHn1pIZQxMt7i3mLNs1H4P2AYX13C5lAzLF8VsvZStxZnVQbWAfPWQCJ5kebr5QK
QCkcOWoz7MrQGm7G/lSq+e6+Mk53NKCvbQPHekIRqIpaABeS4sRGzmybEuc7jX+oQVOmoHBP6t9w
RtGrlLaRY4s7zq140Fn9kktmRDW2QqjT0u21dUcDp2Qu1Oacll43lQjk3PxX+ST3aTt3pxGM6rnY
FUQsKjUdHa0CMPzgWcqmJfZVnoRd5YnUjTWr//I8xKaCSNCv15uzqQ2RgXKEJQmWKy0T+w+3NJOE
KDZSq1KPhmjwbiUl0Pd2osPQvC0zud+h4+lqrTvRYS0C6kEIaoa/aLJAn7JVG7vNdwedVjNvPmZK
2XBa4hGEZTw7oW5eS7jgt8DjeykgcsU5PrRnYN6GvO+tfS/wOzKsE0PmwaSTqSxvT6vV3TPQ7mvy
c7urWzuQYWEBzaTwDz+a9s0KOjuFOSbywwIy2+MKYn9a6ksvAJbN/9TXE5nG+cnPFu1LuKSnbwbG
Z5pXG6u+nUoW0pkwFjSvNofZvlkTHGMzVBrkrDaWUOGmQpvB0FcoX6WION2Kiz9tClV/FyIUSqVj
6UKlxU4A7PB8EcYRZUaofF8Otz1jadNyJQ+oAGXpZJzPaoSsaV90LY//NFGtrzdDrS9DstYr/OAQ
hKf7xaxo8DxHN0A/r0Nq9wYuISgqMbyPjCzskuDfkDMcUqkyIroE/xwpek/XtAOmQ42jSZzWPZgc
R4UGNCRDPBUOuRolsX/cWSdi+lGLS3e+PFEjsKd/ZGG2J1kf7EYmkJTfqSEMOHwR8eD57c8XTvOq
ged/vSGx4IKawkxDddvPBMaRLGs7DSKG10Bw3WS6n/CYoCfhhlp6hlz3KlcI/ClSJMCZ0Pbdn2rU
kpnsMoUa30JKbKHwtpVr+ocn9Q+RxYI00hlSMP/g2JR6OVwfpPYKaWuytizfg9Yd8ddYDOtCqnBu
g6PpNb8MOsdbrhBbNO5j+cHye6JLKtcrhssybBYwg+R/EWptADf8v6XhRPH6aFBKQO+IvG0LK3Lu
Igvv2LqP0aBk1bCkLHC5ShHR2/RJRfEBHluYBO6cex1WYtMqon1DwqgOIYWdhA/4Pqfv5e4rXEVb
qxNDwc1zcfwwKxyP5keaQbs2eHPqIWBo1J7AG19ggR0UgXJnzYkRB8HatIRgJGbbO+dI1tp1pgVF
Uv0wjpwae1YJi+/g0VVDWMG82zT3IQjASu9vAnT4pA3DU53aBQlpsyIeFz8gFyvITWc3v1pwj5es
SBSHJqfSGzUEjAHNRSXEXcME7aj3G/3CuVxIly53uNDB/+dqlKAJ+WEwpBE+gVi+u5wKV1XRpYvs
jl5pm+1wRMaYauGG9ejp6FVyIGow6s/jZxZosYoyaUEAo0bgd40+I7QCJyq6QeIhjRn3yDbUZUiX
O0aYW9frMsxW8eMXw7T9C/CIoNOS0uXIvFvHHx0jZ1iVTX2l/2IpTQ+fNoNEZgc+LwCokhkO8DTF
S9RwzVdvtK717i8mjLMe5TZOsa8FJSJ9yzShVodo8bDd2hl+PBkQzP0KwDCM32WXaN43JMV0dgbB
f0XrkXXgvCRU139Bx0ISI3uTEbdmkAQfrQRuCqIaUb3cLQuCYzrXetCwJsczVlzvU2DEtHokNrzj
Uq4eF+YfycxhT6s35+BMqFZ956N8ZZQc35BGju5LzPweBahPt9oZC3bI/8xXGstGdnKULpykLQSm
kqyvieTuMeSdBzhLR00uPEl7LzmI01/QZ/NG6ym1lskS7NZblC0jI4oR3gkTWf4OtPJZ5l+p0MDe
3NZUe0nNuR+mid+tB/cC+0tYQPXNEmsdSkcrsStdYJsIyTuAbbWqQam1crfkKg4YXfajfibrpKKA
QyMF3WQQ7QgSkh658Yddm1ZMt6NsDmslEwdFbit9Hptzsgd93LabGn7iGQnJ5pq7axU22SGpp7cu
pK1tnfRWaqJ9AeU969qNwofGci9knex5VzGaQSbOArHY3+a1w1ExA3tjLCRfP01eAhhogIiJULzS
33lhUmXbC8ZgSiGQPJeq0ddo8k42iSpheJcLl7iuHriA6BOPCe0eqLJore3moSqgJjeHYBBqmt55
pnL4fTC3bSr1MCKzVxORrt/am9B99vXA5+rfXZP+0MqKO70qyK/HTOSMeslu00SSE+cBYXuRBC4/
hupMJGxYiwn77GYZPop7eN6ipgt+7gW+UDkKnPfvC61TuZiaNeq0esSod6G3AjFFmY7n+KvtqGZK
JdpN+rtPJM/D1wu1PQ3kxaspBLHYaYUKnbKQPPu8SvAhMCAP07EKxttggK5/ye7sczpAbJXzXtsV
fqr22fixpn2KVkdx75CbZOUG2cs5zh986zX4mDENZQ57kIoZ/RDWuqFVUTeF3UIx7GLpg9GrViJ2
TanM4Baq9ZA/lNlcMMW4zCOLsihB+lQ9x/ckSsSC3dKX6aIM2Vv57CZE43EWpxAKmOfIPXIKvP/T
5xS0ajuJxSJGAs63qDcHlo+w0hI9NdaJhnsAU5qh4gtwBj1kwb3zHxWmx8+Sfizw/YyEMEG88q0P
WZcpuvondU8GrfExHFVkjkotVBjGVQucuiGcVFSUGo2YVlqwOfaamtOo9dIjeRg+t+C6KofRLNXb
5S8i5hMZFZvwrgvKpO1Eb5tmW0VUZ9aWfJwhPhEimRZzq6MPAjLEEYPdT/mGvM6+abHAwfWJfjYn
O2LRhjQ3IwHJptBy5T0d/7mBpI4kBCKb2LK24kid7vT+R2/Z23FRLgdTfraSkpAyCECO0kgO7N1G
6mH2Z4equGFome8sGq+L7yEnmcKFH+wPE0XqhF/JxfH3GcaIdkFUN7saeldsQNEt4x9jhXDsVBOS
mtD+/EoVQXk5n8KbBYupYn2f5+uXdMfTm8cMoLjef8+Z3hWpEDcI7tYiXfwL++mfFYTOu0iZzS9C
WRnCPCkgdEOgS9Roys1lkhDaGC93oVg2FmOHu4btQNQ9oP14i/R0o/Alzwum5L71W8q/I6QMOoce
PZGJwBa1y8fxXDJ9KVjWFzVGeLMIA478tYWFvCVGouN+IagfwVWJEZ4R8PabjOTBNphFdBG/1ZDI
8/tD16NrWr33WudTeB5D/HMMVMtSqfU7JeffZJkisd538DwQMJW5c7A4DPoUe7D3YoAMPVxcCLnw
n+P6X/h0tYFMmYw8E3I79v5tpOOpu4+lUQ3k4J3DXf0laZQLmsFKzPWsyjH2a1ID4273xrJ0yM3P
o45lyxRqHOQpOLgZi6cYzs1rp4RQgP69A8fuPTSjgBa+lfyGeXvOHLpLcfQmSLlyT4PWnVSsDj7H
UX7Nbsoxwh+QCTElTXgQU2K6GqCTyDlxreneu1hbBD1YjjRugxcN8pgqXmSASt+Gp5j8UI9TZXlu
aL/4kIyvRfXQPmGzv4R9Ih4gbg+qHIplRY4QaH6OWQ8LsLDYV5bspjcwAskQ4Bd34k2uc2GXKRju
e4sg7/VghvtE3FV4tg/UjWBeun0gmwshFfDyuNcbxE0CXzjBJBHHPSsR3cGp5lgombGfizwybyvJ
PTkv+a+7k52CDu5UMHtg3n8wIQvjt/hLxVxKNUwSe+OI5/MqXq5ayI9lsWEBoEWzJBBtkvVFbF4L
VKV/c9O130ORTqe8jNPmcznForc2NoJ3hBvOx+wdsj5UF9apTMXYqJv3WrOJWeqMe+3ENIrtFPWY
AuYLUljKeDudEfOB80yfufZ8DU5GsuC7McTFtbFuOt1NneYkAwpq0IDs5rnN2GLzz1alzpPZZzRH
HhQKmsDJ9vtDZdhc051CZrUCtyYMmf19FqlyPyrdWkXFHNWSAvxS+OOnTMnTYohotqHSnFnAClBl
AYwIdT4khX6puF/MpWlfhksPPZqWxPxiQkuiBMoYjN3OkRuj4jC2jHXWK5iAuM204+wjbYRhgEQF
c/OEZs+HDmhx93HKw+m+wOlVNJi2Z6JH51+NJUpWBHvaeUdrH5rFDz7GbgfIw8d+i9IPaLsmJ0xW
hlTxuOLQdooPxbmdSlfBAdZgKA7laxW7gcjMSOaxiPcojqdv3M0tmqq5cxa1SN0eQg+AlRIzUEcc
/yw/Yhtbty/qOvCnyGFvS+pQVguHVd+/G49JXNInHoOxbL6JzBaI2xZtghYrwbUgcnUmPA6j2mQV
9kLRJIanHul7NgA6W5kOkaR3tSoezhiD9ljhm0O68k6gzOL6zwhudDb5qp9rJL+Os8fSOZrORJRr
a3EYpnLMDgTeKr7ITuuu5NWFUjg+xkzW0K6uerO3E1HiQwqSSSNiQ8KLMZcVVmZZfASJDyk1H8DF
bfA0tHGyMb4aSmwlpYnP5UjUSxoRYJfZvk7VtbFl6dC4GfTb9Jft0WNILsTU1t6h/quNXDP6Zz4+
jKJx/igUnPiYBLqr5V8lbkKkOHTKOPLrfg0OGmAEKNxBtbWn1xMeOroAcg5+GVA5IaHOjvtS/PVQ
5PdIwtozRO4yOjAw/d8Q8gO+KQCPYtcYQo95VICzL9HdoajOHd1G7HlX207aC9ZbZrL+W9Oah17G
DyFreDa11xLP5jGo4DD4pT9Pu8KNWJSaDc5PLvpFhigMgHQOluPCcZL/spGlGyiYiKPQuPiQhZ2t
/wb3PDdo3L6yJLA+H8QJzggwyhtaCQldpKwCt3COd9SJu1INzsMky67ZUmDyPWqXpP0A9N2ovwNJ
JgY5GRnRjMV5IQrCzyJnZBQZY81taVLbKSU1+oTx9wBzxv2ruJ4Q5fNOmwS3xRA1kpWSzO6crON6
iDT4bZF3/Rcwzi+B+7F8t6jEga5wgiQ+dPGUBd2q/aJwywcJX7et+V6q99FvBEOAvSw1j0UjV7yr
o8/XqqQFSR+FpW4FSnz1zXV6D+/BxhmQDJkOYXELbrZ7idGr7aMUxLj7e5DUCZeWpm7D3Jt34EMQ
DXIA3+aaTHIXRj2+ik5nbxSCW/9hjDpYLVAL2zMYiAAGUnEVvxQH3SUs3kH5WV/U0x24m2fv6aH/
OQWCBmMQOzcZR7opiWC4mZBxAV+Co9GtaXIHN/eQgfMDlyn+oAuN/8W/xh8pT63EHwAF9qRCl7kF
0Wqh7TLRy3MqS+5epR2nRTbukGBiDvNGWZkdXWcuZDzm1uYJ1pNYWzSaUh4+7FqP2MeTh3ThYHzs
bGqUaAUTVdaOZf2WcjoJAMavcEVFE33dFkLugHcEcyuh2oqV2TBK/SRz1dklx1nhr9LjAfzd0S91
6vj1zuxVOEUFuFcGPm7stmlxAbS6HfllhXC4S+TddDgjFQBXbkNgPIuDXt7KafvrOSMn25Tv0jyb
lvOkcqLwCg68wP5q7Sm3WUKco/ho/JCGAzy3koBHJB2Z3mVW6i+zElD3zTk/Kw+Y1S4o19OkKQy4
nFICSK/wCp3yy9GcA+ADuM0mOIwahnEKOTGVEIrktdFXxoMomd0ERYMq1OU96W9iOIkBrhTIk9bg
xWzX0mUnTFxFRKjdL6rQagHmXFuGCHjBaNiiJd65C7RRsfzqR+wTgxe7D5n2ziuPKYlvTpy9P2bA
BN+CDpTAvGZy/sQhaWOClCuhIDcKIRQsr+zlSym46kOTEoSuBBK/oabo7fpXSzIrDs9asskCYGiP
8huf4s0+VPVJvRhgR+M3EDghvI94yWdvgIQzFSHx36sCq/t/Gpl4hwB8RKclN9ooKeWZ6y7EDe+D
Y9K+sb/uQPNwx9fzF21U4py2K1j9ic8wzHoC9tCg9IaCIaJZDSaOJu67oAlxHyFnsfFA1duaPk4O
KxuSGNCbRTsnqWO5J3jQF4E1OL2zh+MAQQ==
`pragma protect end_protected
