// system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_clk,       //     clk.clk
		input  wire        reset_reset_n, //   reset.reset_n
		output wire [12:0] sdram_addr,    //   sdram.addr
		output wire [1:0]  sdram_ba,      //        .ba
		output wire        sdram_cas_n,   //        .cas_n
		output wire        sdram_cke,     //        .cke
		output wire        sdram_cs_n,    //        .cs_n
		inout  wire [15:0] sdram_dq,      //        .dq
		output wire [1:0]  sdram_dqm,     //        .dqm
		output wire        sdram_ras_n,   //        .ras_n
		output wire        sdram_we_n,    //        .we_n
		output wire        sdram_1_clk    // sdram_1.clk
	);

	wire         altpll_0_c0_clk;                                                     // altpll_0:c0 -> [irq_mapper:clk, manager:clk, manager_jtag_uart:clk, mm_interconnect_0:altpll_0_c0_clk, performance_counter_0:clk, rst_controller_001:clk, rst_controller_002:clk, sdram:clk, shared_ocm:clk, worker_0:clk_clk]
	wire  [31:0] manager_data_master_readdata;                                        // mm_interconnect_0:manager_data_master_readdata -> manager:d_readdata
	wire         manager_data_master_waitrequest;                                     // mm_interconnect_0:manager_data_master_waitrequest -> manager:d_waitrequest
	wire         manager_data_master_debugaccess;                                     // manager:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:manager_data_master_debugaccess
	wire  [27:0] manager_data_master_address;                                         // manager:d_address -> mm_interconnect_0:manager_data_master_address
	wire   [3:0] manager_data_master_byteenable;                                      // manager:d_byteenable -> mm_interconnect_0:manager_data_master_byteenable
	wire         manager_data_master_read;                                            // manager:d_read -> mm_interconnect_0:manager_data_master_read
	wire         manager_data_master_readdatavalid;                                   // mm_interconnect_0:manager_data_master_readdatavalid -> manager:d_readdatavalid
	wire         manager_data_master_write;                                           // manager:d_write -> mm_interconnect_0:manager_data_master_write
	wire  [31:0] manager_data_master_writedata;                                       // manager:d_writedata -> mm_interconnect_0:manager_data_master_writedata
	wire  [31:0] manager_instruction_master_readdata;                                 // mm_interconnect_0:manager_instruction_master_readdata -> manager:i_readdata
	wire         manager_instruction_master_waitrequest;                              // mm_interconnect_0:manager_instruction_master_waitrequest -> manager:i_waitrequest
	wire  [27:0] manager_instruction_master_address;                                  // manager:i_address -> mm_interconnect_0:manager_instruction_master_address
	wire         manager_instruction_master_read;                                     // manager:i_read -> mm_interconnect_0:manager_instruction_master_read
	wire         manager_instruction_master_readdatavalid;                            // mm_interconnect_0:manager_instruction_master_readdatavalid -> manager:i_readdatavalid
	wire         worker_0_worker_out_waitrequest;                                     // mm_interconnect_0:worker_0_worker_out_waitrequest -> worker_0:worker_out_waitrequest
	wire  [31:0] worker_0_worker_out_readdata;                                        // mm_interconnect_0:worker_0_worker_out_readdata -> worker_0:worker_out_readdata
	wire         worker_0_worker_out_debugaccess;                                     // worker_0:worker_out_debugaccess -> mm_interconnect_0:worker_0_worker_out_debugaccess
	wire  [27:0] worker_0_worker_out_address;                                         // worker_0:worker_out_address -> mm_interconnect_0:worker_0_worker_out_address
	wire         worker_0_worker_out_read;                                            // worker_0:worker_out_read -> mm_interconnect_0:worker_0_worker_out_read
	wire   [3:0] worker_0_worker_out_byteenable;                                      // worker_0:worker_out_byteenable -> mm_interconnect_0:worker_0_worker_out_byteenable
	wire         worker_0_worker_out_readdatavalid;                                   // mm_interconnect_0:worker_0_worker_out_readdatavalid -> worker_0:worker_out_readdatavalid
	wire  [31:0] worker_0_worker_out_writedata;                                       // worker_0:worker_out_writedata -> mm_interconnect_0:worker_0_worker_out_writedata
	wire         worker_0_worker_out_write;                                           // worker_0:worker_out_write -> mm_interconnect_0:worker_0_worker_out_write
	wire   [0:0] worker_0_worker_out_burstcount;                                      // worker_0:worker_out_burstcount -> mm_interconnect_0:worker_0_worker_out_burstcount
	wire         mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_chipselect;    // mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_chipselect -> manager_jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_readdata;      // manager_jtag_uart:av_readdata -> mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_waitrequest;   // manager_jtag_uart:av_waitrequest -> mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_address;       // mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_address -> manager_jtag_uart:av_address
	wire         mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read;          // mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_read -> manager_jtag_uart:av_read_n
	wire         mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write;         // mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_write -> manager_jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_writedata;     // mm_interconnect_0:manager_jtag_uart_avalon_jtag_slave_writedata -> manager_jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_readdata;      // performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	wire   [4:0] mm_interconnect_0_performance_counter_0_control_slave_address;       // mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	wire         mm_interconnect_0_performance_counter_0_control_slave_begintransfer; // mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	wire         mm_interconnect_0_performance_counter_0_control_slave_write;         // mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_writedata;     // mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	wire  [31:0] mm_interconnect_0_manager_debug_mem_slave_readdata;                  // manager:debug_mem_slave_readdata -> mm_interconnect_0:manager_debug_mem_slave_readdata
	wire         mm_interconnect_0_manager_debug_mem_slave_waitrequest;               // manager:debug_mem_slave_waitrequest -> mm_interconnect_0:manager_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_manager_debug_mem_slave_debugaccess;               // mm_interconnect_0:manager_debug_mem_slave_debugaccess -> manager:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_manager_debug_mem_slave_address;                   // mm_interconnect_0:manager_debug_mem_slave_address -> manager:debug_mem_slave_address
	wire         mm_interconnect_0_manager_debug_mem_slave_read;                      // mm_interconnect_0:manager_debug_mem_slave_read -> manager:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_manager_debug_mem_slave_byteenable;                // mm_interconnect_0:manager_debug_mem_slave_byteenable -> manager:debug_mem_slave_byteenable
	wire         mm_interconnect_0_manager_debug_mem_slave_write;                     // mm_interconnect_0:manager_debug_mem_slave_write -> manager:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_manager_debug_mem_slave_writedata;                 // mm_interconnect_0:manager_debug_mem_slave_writedata -> manager:debug_mem_slave_writedata
	wire         mm_interconnect_0_shared_ocm_s1_chipselect;                          // mm_interconnect_0:shared_ocm_s1_chipselect -> shared_ocm:chipselect
	wire  [31:0] mm_interconnect_0_shared_ocm_s1_readdata;                            // shared_ocm:readdata -> mm_interconnect_0:shared_ocm_s1_readdata
	wire   [7:0] mm_interconnect_0_shared_ocm_s1_address;                             // mm_interconnect_0:shared_ocm_s1_address -> shared_ocm:address
	wire   [3:0] mm_interconnect_0_shared_ocm_s1_byteenable;                          // mm_interconnect_0:shared_ocm_s1_byteenable -> shared_ocm:byteenable
	wire         mm_interconnect_0_shared_ocm_s1_write;                               // mm_interconnect_0:shared_ocm_s1_write -> shared_ocm:write
	wire  [31:0] mm_interconnect_0_shared_ocm_s1_writedata;                           // mm_interconnect_0:shared_ocm_s1_writedata -> shared_ocm:writedata
	wire         mm_interconnect_0_shared_ocm_s1_clken;                               // mm_interconnect_0:shared_ocm_s1_clken -> shared_ocm:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                               // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                 // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                              // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                  // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                     // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                               // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                            // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                    // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         irq_mapper_receiver0_irq;                                            // manager_jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] manager_irq_irq;                                                     // irq_mapper:sender_irq -> manager:irq
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> altpll_0:reset
	wire         manager_debug_reset_request_reset;                                   // manager:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [irq_mapper:reset, manager:reset_n, manager_jtag_uart:rst_n, mm_interconnect_0:manager_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, shared_ocm:reset]
	wire         rst_controller_001_reset_out_reset_req;                              // rst_controller_001:reset_req -> [manager:reset_req, rst_translator:reset_req_in, shared_ocm:reset_req]
	wire         rst_controller_002_reset_out_reset;                                  // rst_controller_002:reset_out -> [mm_interconnect_0:performance_counter_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:worker_0_reset_reset_bridge_in_reset_reset, performance_counter_0:reset_n]

	system_altpll_0 altpll_0 (
		.clk                (clk_clk),                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (altpll_0_c0_clk),                //                    c0.clk
		.c1                 (sdram_1_clk),                    //                    c1.clk
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.areset             (1'b0),                           //           (terminated)
		.locked             (),                               //           (terminated)
		.phasedone          (),                               //           (terminated)
		.phasecounterselect (4'b0000),                        //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0)                            //           (terminated)
	);

	system_manager manager (
		.clk                                 (altpll_0_c0_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                //                          .reset_req
		.d_address                           (manager_data_master_address),                           //               data_master.address
		.d_byteenable                        (manager_data_master_byteenable),                        //                          .byteenable
		.d_read                              (manager_data_master_read),                              //                          .read
		.d_readdata                          (manager_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (manager_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (manager_data_master_write),                             //                          .write
		.d_writedata                         (manager_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (manager_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (manager_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (manager_instruction_master_address),                    //        instruction_master.address
		.i_read                              (manager_instruction_master_read),                       //                          .read
		.i_readdata                          (manager_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (manager_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (manager_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (manager_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (manager_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_manager_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_manager_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_manager_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_manager_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_manager_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_manager_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_manager_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_manager_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	system_manager_jtag_uart manager_jtag_uart (
		.clk            (altpll_0_c0_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                               //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                           //               irq.irq
	);

	system_performance_counter_0 performance_counter_0 (
		.clk           (altpll_0_c0_clk),                                                     //           clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                                 //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_0_control_slave_writedata)      //              .writedata
	);

	system_sdram sdram (
		.clk            (altpll_0_c0_clk),                          //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	system_shared_ocm shared_ocm (
		.address     (mm_interconnect_0_shared_ocm_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_shared_ocm_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_shared_ocm_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_shared_ocm_s1_write),      //       .write
		.readdata    (mm_interconnect_0_shared_ocm_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_shared_ocm_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_shared_ocm_s1_byteenable), //       .byteenable
		.address2    (),                                           //     s2.address
		.chipselect2 (),                                           //       .chipselect
		.clken2      (),                                           //       .clken
		.write2      (),                                           //       .write
		.readdata2   (),                                           //       .readdata
		.writedata2  (),                                           //       .writedata
		.byteenable2 (),                                           //       .byteenable
		.clk         (altpll_0_c0_clk),                            //   clk1.clk
		.reset       (rst_controller_001_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	system_worker_0 worker_0 (
		.clk_clk                  (altpll_0_c0_clk),                   //        clk.clk
		.reset_reset_n            (reset_reset_n),                     //      reset.reset_n
		.worker_out_waitrequest   (worker_0_worker_out_waitrequest),   // worker_out.waitrequest
		.worker_out_readdata      (worker_0_worker_out_readdata),      //           .readdata
		.worker_out_readdatavalid (worker_0_worker_out_readdatavalid), //           .readdatavalid
		.worker_out_burstcount    (worker_0_worker_out_burstcount),    //           .burstcount
		.worker_out_writedata     (worker_0_worker_out_writedata),     //           .writedata
		.worker_out_address       (worker_0_worker_out_address),       //           .address
		.worker_out_write         (worker_0_worker_out_write),         //           .write
		.worker_out_read          (worker_0_worker_out_read),          //           .read
		.worker_out_byteenable    (worker_0_worker_out_byteenable),    //           .byteenable
		.worker_out_debugaccess   (worker_0_worker_out_debugaccess)    //           .debugaccess
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                         (altpll_0_c0_clk),                                                     //                                       altpll_0_c0.clk
		.manager_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                                  //               manager_reset_reset_bridge_in_reset.reset
		.performance_counter_0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                  // performance_counter_0_reset_reset_bridge_in_reset.reset
		.worker_0_reset_reset_bridge_in_reset_reset              (rst_controller_002_reset_out_reset),                                  //              worker_0_reset_reset_bridge_in_reset.reset
		.manager_data_master_address                             (manager_data_master_address),                                         //                               manager_data_master.address
		.manager_data_master_waitrequest                         (manager_data_master_waitrequest),                                     //                                                  .waitrequest
		.manager_data_master_byteenable                          (manager_data_master_byteenable),                                      //                                                  .byteenable
		.manager_data_master_read                                (manager_data_master_read),                                            //                                                  .read
		.manager_data_master_readdata                            (manager_data_master_readdata),                                        //                                                  .readdata
		.manager_data_master_readdatavalid                       (manager_data_master_readdatavalid),                                   //                                                  .readdatavalid
		.manager_data_master_write                               (manager_data_master_write),                                           //                                                  .write
		.manager_data_master_writedata                           (manager_data_master_writedata),                                       //                                                  .writedata
		.manager_data_master_debugaccess                         (manager_data_master_debugaccess),                                     //                                                  .debugaccess
		.manager_instruction_master_address                      (manager_instruction_master_address),                                  //                        manager_instruction_master.address
		.manager_instruction_master_waitrequest                  (manager_instruction_master_waitrequest),                              //                                                  .waitrequest
		.manager_instruction_master_read                         (manager_instruction_master_read),                                     //                                                  .read
		.manager_instruction_master_readdata                     (manager_instruction_master_readdata),                                 //                                                  .readdata
		.manager_instruction_master_readdatavalid                (manager_instruction_master_readdatavalid),                            //                                                  .readdatavalid
		.worker_0_worker_out_address                             (worker_0_worker_out_address),                                         //                               worker_0_worker_out.address
		.worker_0_worker_out_waitrequest                         (worker_0_worker_out_waitrequest),                                     //                                                  .waitrequest
		.worker_0_worker_out_burstcount                          (worker_0_worker_out_burstcount),                                      //                                                  .burstcount
		.worker_0_worker_out_byteenable                          (worker_0_worker_out_byteenable),                                      //                                                  .byteenable
		.worker_0_worker_out_read                                (worker_0_worker_out_read),                                            //                                                  .read
		.worker_0_worker_out_readdata                            (worker_0_worker_out_readdata),                                        //                                                  .readdata
		.worker_0_worker_out_readdatavalid                       (worker_0_worker_out_readdatavalid),                                   //                                                  .readdatavalid
		.worker_0_worker_out_write                               (worker_0_worker_out_write),                                           //                                                  .write
		.worker_0_worker_out_writedata                           (worker_0_worker_out_writedata),                                       //                                                  .writedata
		.worker_0_worker_out_debugaccess                         (worker_0_worker_out_debugaccess),                                     //                                                  .debugaccess
		.manager_debug_mem_slave_address                         (mm_interconnect_0_manager_debug_mem_slave_address),                   //                           manager_debug_mem_slave.address
		.manager_debug_mem_slave_write                           (mm_interconnect_0_manager_debug_mem_slave_write),                     //                                                  .write
		.manager_debug_mem_slave_read                            (mm_interconnect_0_manager_debug_mem_slave_read),                      //                                                  .read
		.manager_debug_mem_slave_readdata                        (mm_interconnect_0_manager_debug_mem_slave_readdata),                  //                                                  .readdata
		.manager_debug_mem_slave_writedata                       (mm_interconnect_0_manager_debug_mem_slave_writedata),                 //                                                  .writedata
		.manager_debug_mem_slave_byteenable                      (mm_interconnect_0_manager_debug_mem_slave_byteenable),                //                                                  .byteenable
		.manager_debug_mem_slave_waitrequest                     (mm_interconnect_0_manager_debug_mem_slave_waitrequest),               //                                                  .waitrequest
		.manager_debug_mem_slave_debugaccess                     (mm_interconnect_0_manager_debug_mem_slave_debugaccess),               //                                                  .debugaccess
		.manager_jtag_uart_avalon_jtag_slave_address             (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_address),       //               manager_jtag_uart_avalon_jtag_slave.address
		.manager_jtag_uart_avalon_jtag_slave_write               (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_write),         //                                                  .write
		.manager_jtag_uart_avalon_jtag_slave_read                (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_read),          //                                                  .read
		.manager_jtag_uart_avalon_jtag_slave_readdata            (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_readdata),      //                                                  .readdata
		.manager_jtag_uart_avalon_jtag_slave_writedata           (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_writedata),     //                                                  .writedata
		.manager_jtag_uart_avalon_jtag_slave_waitrequest         (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_waitrequest),   //                                                  .waitrequest
		.manager_jtag_uart_avalon_jtag_slave_chipselect          (mm_interconnect_0_manager_jtag_uart_avalon_jtag_slave_chipselect),    //                                                  .chipselect
		.performance_counter_0_control_slave_address             (mm_interconnect_0_performance_counter_0_control_slave_address),       //               performance_counter_0_control_slave.address
		.performance_counter_0_control_slave_write               (mm_interconnect_0_performance_counter_0_control_slave_write),         //                                                  .write
		.performance_counter_0_control_slave_readdata            (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //                                                  .readdata
		.performance_counter_0_control_slave_writedata           (mm_interconnect_0_performance_counter_0_control_slave_writedata),     //                                                  .writedata
		.performance_counter_0_control_slave_begintransfer       (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //                                                  .begintransfer
		.sdram_s1_address                                        (mm_interconnect_0_sdram_s1_address),                                  //                                          sdram_s1.address
		.sdram_s1_write                                          (mm_interconnect_0_sdram_s1_write),                                    //                                                  .write
		.sdram_s1_read                                           (mm_interconnect_0_sdram_s1_read),                                     //                                                  .read
		.sdram_s1_readdata                                       (mm_interconnect_0_sdram_s1_readdata),                                 //                                                  .readdata
		.sdram_s1_writedata                                      (mm_interconnect_0_sdram_s1_writedata),                                //                                                  .writedata
		.sdram_s1_byteenable                                     (mm_interconnect_0_sdram_s1_byteenable),                               //                                                  .byteenable
		.sdram_s1_readdatavalid                                  (mm_interconnect_0_sdram_s1_readdatavalid),                            //                                                  .readdatavalid
		.sdram_s1_waitrequest                                    (mm_interconnect_0_sdram_s1_waitrequest),                              //                                                  .waitrequest
		.sdram_s1_chipselect                                     (mm_interconnect_0_sdram_s1_chipselect),                               //                                                  .chipselect
		.shared_ocm_s1_address                                   (mm_interconnect_0_shared_ocm_s1_address),                             //                                     shared_ocm_s1.address
		.shared_ocm_s1_write                                     (mm_interconnect_0_shared_ocm_s1_write),                               //                                                  .write
		.shared_ocm_s1_readdata                                  (mm_interconnect_0_shared_ocm_s1_readdata),                            //                                                  .readdata
		.shared_ocm_s1_writedata                                 (mm_interconnect_0_shared_ocm_s1_writedata),                           //                                                  .writedata
		.shared_ocm_s1_byteenable                                (mm_interconnect_0_shared_ocm_s1_byteenable),                          //                                                  .byteenable
		.shared_ocm_s1_chipselect                                (mm_interconnect_0_shared_ocm_s1_chipselect),                          //                                                  .chipselect
		.shared_ocm_s1_clken                                     (mm_interconnect_0_shared_ocm_s1_clken)                                //                                                  .clken
	);

	system_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (manager_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                    // reset_in0.reset
		.reset_in1      (manager_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                           //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (manager_debug_reset_request_reset),      // reset_in1.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_0_c0_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
