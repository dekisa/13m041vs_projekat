��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh�QN��f��ID�k{��`Q�
=�O�I���*��9��K��H
g���B$8�������#IG��u�������.���9,�J*L������h��g�dLCm�}q�����I�j�A=g��(c�w�~?����q�Ρɽ���hE��gAN�kD�g�r�	07�L�MfA�?���<f�'6�Wܞt���Բ�`��d�lcDHZ��xv՝�LE:�f�C�W9 a�
? ������p�?yR�|}W�n���'���k��7#6Q$�F]�}e�Td�>�X���qS�����.�����Щ�%,�D��|U��C;�r����A䝁��7'H��j�k�gs9�"�x=�A]+ܸ�։|VI�ن�/�mo��v�z�c��.�@�y)I�7 ��_q���Ċ�P;����o�TI������=5�rJ�:���5+N�����>�d���jڛPaaj|�{��i�
�\�nr�Vu�^;4YUX��X��*�+k���n�+�X?c+��J!��4p��4I|#�%<�P����eky��Lz��qs_�JJ�W꿼��mY
g^}IYG�����i �je�M� �Ql�{f �;�kU�� �)��UT�~�#����`�NDA{[� )}�y�7�A�f���l�;ړx(LO1d�i$��P���ܛn!��rj� ҽ������y��b�-溼Z�V����O�uб����J7$��8hX�"�b�qs�t  𥳐�=�O�~.��w�*�-�6m�)Lm�'��_�']�ϕA�u�lC;��J�AK|��YP�s�������q���sl4�s���ת�r\�ݺ�BJ	�O?�M��-vc�4�I��A��,;�l�2���0�
|���m?����jk
[���j*{i�]�vY��Q+v���Eo���ǐph���j�@�:;C�u�s�UU�����4y��2�v��C���F����csL���ɮGo}п�������*Y�q,�;�a'P*��ݵ�'>l��n̓��J��4�򌈹���eӣp+�'�4#��D�HBx��L�<n��ng^���me�ͅU
�k'�e4�a�v]�Lw0�>��XuiZ˃A���)$C����Y,R1ې8P8����9����[�|�Z�{g=���*�9�Q
�޽W��F���P�'�;zyZqcfof)�.rC�
�B��S$ey`�C��~�˚$�'�L�K�#�E���t�����q�a
@5�#ƚJ@0ʄ�-!��i8�g�k�QZ�BM�#�2?��4��y�9n�&�{y*��j��ƥ�V�L}a˧㒆b[`P��:�tV���F���i9����,S'È_Xd������;��V��A'���c�( ��.���I�g���ۂ!�(���<�C�<-2��	�+��u���%�cX��]�j��'T�R��7ȱ���yU�!+6�
���׬��,ӫ�j�F��b��9֎�ZWd�/QW'���-j6.vϿ�iQ ���i�y
��&0>q3
D@9�[���f��ن���ʟ��l�96�]��q��&#|驍*uӛ���}qR���7���G.F�Z�l�&��9w������;�SM�aI�����H��6)����f*L0t�Y�Y
��F�((|�c�ѕ�(�N���i���s��c&����6U�Lo=o�#��7?|�w{�4��c5�����De*;����z0�#b���K��gj�o((b�����{?hl�Ѕ�C�-{(�f�,�e �D�C�+8��Gg���<��!��+JT��������fS\to�O6߾G�������Rf�zh(��=|�im�EjF���&%��F�[S��!H6�D�<£yLd�G�5N쀺�}���J�?vM��C�Ci7�[KB_Q�9��W��;�f8��1�̿e�:���Ȼ5N��K���ء�(���,��_�NX��th߁�BR�?)�fv�L�]H���Y�	c��b�	�X�*Wҏ*���U[�Վ��O�����
�H��Q� KG��k���F�5s�3�A�S��x$v�eN��f$���W�vEZ�r��.�5P�f�����9i�`r�����ׅ�d�zJ��1�~;@��[m�O�+?���JR��{�{^��%�����rQw��Z�[	���_�Ǳ=�h�%&O3a�*����!��]Rf�	�ϔ𗿑g��d�'���Lh�<��K�!xd�k5`u�cT&�*�mg�'��YU�&	�z$��x�1i�o�@�/&��dNyx�v�ݖU�)J�  �C�&-qMg�8s�<�rp�yʹ�RuϝM�����Ur�C��b_�y[k�����K~0iyL�Z��	����*D�?��l��p:�L"~v�� a�w��4�?I�;/2A������5�K"	�QV-��N���7�1ӾO�� ���0����b���e��^�$�39ll���ρ�j�R*�t�]+~G���Y��*(��e��	�K��`S
I�Q�CX��b����@vmDg�ȯ�+�D�X��"�wM*�n�1�i-�%�sݮ�S��mVMP�tW�d{ne����l������O}T >T�D3�2����U��7�ُ�B����]ϓl�EI�	%��/iG��J���Q�>]B�cd�$��K#f��IR����8����C"|��R��=�9�}�Z.���s�w��s��d?��5b"��K!6l�?�6���������V;����s�"�]#�8NGDU*��֭�yp��4�A��6�r랛�5�o!��MƝ'el���-��;{*�R�t��{�]���6�Rm�D��$+zݎT>.����Z�0�$k)K�Xs�-vp|�d��f�ï�
 ��8_���p�F����P����р��b���e��Z(�V^�)v+�^�{_(姅�|��H�����9� f&��vMI��9����iJ�����C����Z�-��a��E\(]}j�ڼ#,\�]ay�v�?^�Z�������03�@�Z�#ɋj$��=p�f�X{�F3�H>��6�j�M3jt�A��("9���2�+��@�g� |�����D��s<�SH�:B$�ħ�X�b�:�\�MbUv3���k��D�Vo'��m*Ƈ�_.'^X!	�#�.@��d�x���yl=^^E����MV]\�-�Ly��3<�耫�'���������a��Y!��p ʹ��AR)�u�p��J}�2���K�s&2ۘj����T�êN�����fA� ��o�N7t���V�����̱�#�(�*���ԛ�U��M1�rf��{����ƱLR;zGkt�����1����C���@/�K~krЎ0��vG�[d�GB_��ˌ�+�a"�m[��~3] ���d�SJ�"N�qd�jj�e�=��:�(@\ì�o��1�V�l^.�W��8��sL�%nrK�	��UK�1��-7BӑVݭ���z96�(�d��K�]��i��f���=�c�aSӈB�~j�<�/�o�v@hQ+Z\�h��^�}�B{m���:"�P�5,M�6Hދ���v!��-�IÌ�E�n�)��WR�s�)ߜ���h��"����M����4Qy>Q��F�	�0�z�0]T]M��s��!6����
������a��9����/�5-�+/hW��%��|3��/ՙ���ދeZ�+5gV�2A?��Y!��`�`��<�'�,�jۚ��p�v{8�B���$��;ب�1��Z`yĕ�X�b.9���t+>������� ��T��/ҎTy!Q����6�&wO��C1U��E�נ泶7�-�A7�4)r�=9�!���>���9[��k��m����α��� ��׾xb��ǒ���_/x}ߔ��3V���J�s�6:��$��ӓg� ��o�	8e��+��RW�p��'vtuA���Uk[A�|��Lѡ\U��e'�Y¬�V��+��0���_\����Z�AY?qO\�x�� ����Ԗq�%l�o)Pkw������L�5c>	�p��\v|���>#�'%�����a��g�R����q<aד�D�:��_��N[�ȼ��z]����mo���ܪן�6jHz-�v�U�!4��"���e������cd�{�^��
���:or���K�o_cIh�[�&�񫆔Mh����e=�ꟕ����(���!,�K�l��7�1�`�� H˚:�ӛ�{���z!KChFl�U���|��;�gr��g�'�Ԝ\Z^Y�d�(����G�nOi�!;�0���$�M&�<�a�f��=?��;�n���z�2��W���2Cv��SU��	a�Y�SE���;T�ʯ{��ۀ�Ä�m�~�O��F� �IA�q�K��x<d�u�;�̿�/�9��tz���W�N�G���p�����0��Otcv�
6��֜�1DV��ϕ5���b�˪Sf��t_���Qm��G,A�7���K��p΍���]f	š溉��/��W�y�`�.�UUD�E��Ғ��{���Z�Hۗ�BSS|��g��#6�j�ly���F�FVw��St�����MG�����Sd2����G��*3t�&�0�<�>����h�M�i��"w 䣜���o%rš�����m?�����0,�S�z5V����x'��˾�@�`H�14�b����t�k42�T93BP숧���K� y��yt\?�hE��S���#�g3#�S"'.Z��UAH�H80�3p�� ���fT��)��>ioo4u(m��KŅ�tאF�^��؂bɧ\Vq#�o�??5ø�H2�<OިT��΃�h�1��ke��
1ۦ+��2�R���O�9����=1 ��D��DK�M��߈�ϓQF�������",�{�s���"�	l��[�a����	+�>e,e�}�=ؤ�}�K١�C7w�(�C���A���~�k�2��3ʝ]8*�,}�m�2w��H�8�3�����������L?cԫ����#7�'�r]�gy�D�L,5��<��*���N�xRk��^�.��� �T�����C�S�*��W�V�&Kr����:Kx9��
��4����~QR�#�8��������ܫ�>�*��*�	��<z%=���yI�S��+��`�?�+��� ��`��b����:Wcc����0M%���f'Ӑb��sAb5�#N�jn�ovTc���vac��֦1��s�P�ӭ��9�N
"��~?�W
���m�	��Wa̬����w����A;esk&��j�d.�;�����
 ��#��o�=�O����g�����2�+�"G��, �3��='P��WX���Qx��/t�O�y�� ��Hn��3ǭ哧��3�Lg�ߨ��q����[��K*�j�[�Qx�,���*�H)�M���-H��k�lߠ����}��|���k���(7����͹O�9���9�p*Mi���&�Q����)l���|�iu$a�����0���
Q��Qɚ}V��dTx.���h�z���R�!��R�\�ѡDc�WUNmX��9�	��	�ћ�$�v!�ZX�:	���-���V�JTz;�dni��1�ȑ^��}�l_Ux5��;ð�q?�AѪ��?���.�Ty�ф}����R8I�V�s@!�YC�w0�#�#������5|v���.�1�Ԃ�#XϞ�F�o��V��l��g1>�a�1��o�I�3!S�z@`�'au��b_�]�i`[2Z���$�%M��b����΍=/��4�n6���/r�^tۑ�A�Kȸd����&����
#g}�#g��N���$LZ�QX���/ ��&����5�n�!}�2����};We�AEdo�N!�Â�r���u��p,?Bd,?\��ƺ�Ju���D�ф��9�.*7\���&oaXJ "l�K�٪r�=�߶����
6���{���ɚpW���K �y�5�gkp&0��c$��\�z�\
L-�V��I?���7��&'$��ٷz��'B#t�mk!]L%��Eơ
H|��(k���/h���� m.SB{�h/(����:&HoK�q�j��^H��>�s/66�?���K6��-?��x�#y��,B�׬��!�i��)d�{��Z)/qy���Nͪh����"�l�	�Q����5����
�c3>-���x�}��bZ�ݒ�� X� ۂ&���h�"��؋�)ڭ�[����3l���b�r�u7)X~q��.��o�9������ �uq��ވ�	ND7?�����ݩ �2Lr��x_�ՠ���9[�@����.�6�-�ӹ\|�(��j���Ax/W�v�	m��]�	8Ph�B;]j)��>�e=�8��׍�S�M�Q�'�X��ć\�(Yn��\�\㰑��B��:�W���{n�H�n*�ʯ�Z�T�8䬂�i�Y�]�S/�W M��A�?jit=½O�aS��|<�̶�3I�:����*N�X���J�h��Cf��$-1ɴ���3T�=>�ja�b �Ζ�i̅���'-Ze7�=t�>	!c���Q��_aN> �rb�NЖYe�h4y3���j���v� !zʣ��w`D���F�醷4Ԅ��:5(���1Or I��VR������P��`��f�#�(�R�t��èm�i+�́�=��Z�!m�ZzԤ9t��J���ͪ����2��6U���L���wv٠0T΢77���� m[?�D�s�� ��nIGƴ5���jt�agX��Eg��q���G��SQ���Tr�4+5� �@G-|K�0�GI!
Nf?��#�B�(<���9�$�jVH��y�����O��w�)� ,�9w)1s$�4�\�Z�$���;ya�;!hcdnH�[�.$$���g|���b8���ţ���[��/,�:�H��C
2��%|qL�8yVv܋ K^�9�u�%���W�SN�$�:���hg^���EX��_>j�8&��[�V�5����