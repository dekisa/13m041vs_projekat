��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�@�w�4s%�mH䖩�ᐌ��)ޢ���U^�����Kk%�}2�4�ZS�v��k�=����?�,��%̀%Q�Q�=�~�ےOz:77��rY͒�ܭ@�����5G�fw�![��-�l�4�;�W��9�d -:��5<�`7��=����4�Y���qŮ���T=~� J�h�0�df��G�+���,�2��b���>���촓8H��l.�.�l�v(0�P񲳮B�Cc�Sy�tֱ�{u�^�x�k2
#�_ҮE}�Mz���W`x�HFcY�ԍ0�N���ŠZ�L�c��MH;~��Ưo�<��t<�H�Q5���C��br9Ǯ������/���Z,_���F�Z�O"䵲'��h�i�Xb)f��d���L��<>v1��Ld����^Öx��R�c.g��r"��jm0��$��u�\�n �H5J%f}I+q�]��Z:��9�6�a��K*��Ȓ�bG�+>tͦ9���<-�JDP�˥	݆���E���媓����M��ˮo�g����3	�nܚ9���L�Ƹ.Vc�ҽi^�H�$����i��J9�#_2cO��О�����Ȃ��4=����^p��BQ�_b"�+ܮ�N�	2��
�XWJK0���^($��W�Jӝ?�������ZE0c�!���nO�Upj��t��7Dq��ݴ�n�<�%�P���ŕ�]����/�B�g G/�F!n�P�'�gtM�V3-���_d�?eǭ0YE|?�":_J���e����]�����Oܕ�Rv��.(����lh��L���!�>�^Q����;��'7˗U��+�>��ll�_&�Ȝ��?�ˬ�B�\��e�4\+p`
y��c���X�&�g�N�3�(`6F; �(`��1�)��%��&S�Ԕ��~�2��MH�f���� �I�T-i�Zɿ�}7��,�,�Ź����j!��݌j�s�!�QG6�~���I�o��ɵ�����!�*�@���m�g�������X��BRK"�&��2�a~�~��)�\sUx\�Dp�� E��~#�Ʋ�k��0k�_o!v��l
��!����C0~*���[�I
x��K�xx�_=������d�W�`�rD뉏N*q}Y�@2@�O"���쭛+b���b��q��4H���,�1�h\��.�SF��{v�w���{!C�i$ $�Sz��m���P���MZ�Y�`|�Ŧ(��Q����&�J�zQ��ENW�~��a`T%�4��1�aySl�&�f �
�;z�Y��)�n��%)?�:n+�Wn���.�p�</��^�!)8T�׍�tȶ=�͊I'D�b��m�ү���R��������b[@v)�U���ִԦ��r�'��F(ٰ.V���cp�.9\����w+s��E���m�~�y�SȆ���xј���2'I�B�I4�W��=;Ҁ(������) �-J�
���e蟩�K���h�t+�G�m��aM��x�����B��Y���z��"Ip��D�����,Vtܴ*�2���;z�[_���9�YV�ލ�L����ja�Z�_�>D����E/H"&QW��m�77��;3��z��j���I�5r��ғY���&!�SN��=nM�����
�X�� �S[�-�P�l�RisP�����a�>�!�s�	=ep��,(����l���*��y`U��Iȥ��x��&�߅��Cs��3$��~_/(�����+"���S=�j���-H�a*'u4Q��|A��=���eX#
!�} \�X�ɚ���ֶ֊�y�?t�9a6�~�E����N׌��ZW�e)egE�P���W:�(MM^�	�H�~��~-<l�ѩC�JQ�~�쫟S^K����NE1C����u�Us��rhi-�ϚFF�@̡��(�lV�z�P ��eG-~�Y��R��z�q�%�&�:���g�9vO�*�pFfR:z{�����o=�7~y%�!�t�r�2�W���?IP��P^�o��"S�/�����z�����~ٿ"����Q��}��'o��2D��������`��n��Ei�����Ͼq�"����\;�j�i�An�k�wrg"W�},&��5i����8�M$-(�Ib1��{��k�ء}���&��FlL�b#��Z��{����.�R#=�ki�0�Q�4�ys9-��0c=�$���MN�`�P,��XW��d��r�4��X�E����/����0���>�������Uj�n�'�\*-N��L<�#v�	��*��VJ���8�����Md��������P��O�:Tj���J���7 �V�<&�c�V���芤b���.C<��Ҽ��&���#E&9B�6��/�6% +jLc'g�%iHa k�1�''wf\�֫e��h6�ϐlZ�L^������b� ����ڲ�*��11h7�������O��!n;H�|F�D��;�$�,�,�0N��̹��Ʊ�u�uya�_�Q�&U�v;Ao��yk���O騍ю��4����$�f�5J&֚�!Ҝ��rF*��+�٣�>���4f�0��|�W+W�������nKz��;��yiEA��Ū���6���D����~�) +gc�R'�V���h�t&�������W��Z~~�A���	�VOr:8��X�y��bo���4��@m�d)V���
tk_�okܐ���<��κ��f�Ynǳ-K�I��I�0=).���p���],��@Bj��R�#���D�D�C�)�i�=c�O�w�a��*,繸FYc��N��+T��ޮ��-�N���}��+J�)���J���f��[�n�K Jr�����B��cIPa�t�/H��d&��<��~�Y
�C��ɤ	�6�;t��/i� گ�Ԏ��0��=��K����W����F�jX*0��^Ϧ*���|�^s����zoG�8�/��AJ)!g���(�,lR�?:�~���$:�"-��T�[-K�|L����Zǃ���'<:�>���%�:���z{����;q9�0
QiA����Mh;q\/l��a�lPO�J�b`���zw	�8����̇x(Wr��3){`N	��v�a����qe�y�,��&o<D�H���F^�{됏����5Hh��!�����%V5f����`��\�C�q�|�1��	�$(�-���i ՆA�xw����z�61�sQ%� �N���|h�����w4�G����V}?����ś��i��J�����9k��0�>��������p� PJ�7�;�bD@�J�a0Y*��s����YF�m��!��2��f�c�Rh�Mz/�Ĳ;5:���D�C�N���ޠhj2]v� D)�^3ݺ�kT	���nJ-��?������7M��!�=��m(j��fh��/��ԧ%��Ǿ�.2�VL�v@�o�ȷ1�����X�J˜Y5<�c7�� �\Vo��ܺl��yS�� �I�d`��&�9�HΡ���\P���$u['2�ǃj��̓G�X<f�XUcG���7U�"�X�`��P(�Ę�E�w�zt�G+]� ����(r��F��x[� �����n��*�]J����!�-%�D�Z�	�r�H��:�[�'f<ii�l��ZP�E2*q�!�ik��_�Y�_XS~V��A�NU$&�6�]{�g7�2	�c?����
���,f�D��F8�\��t)���[�,���(~h���:h����g��	A���{q��,�E�p�0hf�����>ܠj���G�ء2;�D���3�TrMtazzv��D;��y�P��D�@T�p��f�B�`�W*�i�Q����d��� �c��Y�N�S�a��A2;��,F���<��M� /�p�&:k�X
��iGU����OT���T�_�m�� �m�~�<�*�x���	h�z���U�{�Qsw�fc�~+�ug�hQ۰1�e�&����/s�����ǲ�Jߚ�)�bko�y3��P��G׷	���tٛ�V˰5��^��^�n-K
ǧ�oEؘX�j���<ى���q�v���+�d-\��AC�׳B_������������Xfu������_��6���[�D�f��R��W*Jwݒ�b�<f�1� ����^85%/�r,Z�"J��3��+
>��g��o�)��Vb����J1��K��N*/��]PK(��dH�5�޼��Acp�	�Vh��sL��g���OS��*�-���
`Qnj���k���?6��ؚ��������S�,��k�iϿ���6��)�s:�-ڧh���yXt��*�c����`����'
)���/R�� {_���R����:����F%�{��󄆸z�<�.�t�a�h3h58�T�4�!U�k���A@i-�sX��]���I?��U�����mk��88T���t=S�ɋ�gQo����4��D��@��l��l\G@�&���8��m|*t�Hh42i	�۞h�t(�pb���@�OJ)���'/�A���x��Y4٘�Թ��U��/��1'���4�y��?��AO�Ir�>�ؾ�pg���hJ��W�C89�����Q*�\4rm}]Vf�ȑ�[8<��t��~Ϧ}�_-5U��I����QEm.J�~٣o��� $M��k��{�$d�e�r����<J��.��pf�7��(W�VY�O��t�I��Z�V��$�jMNG ~�����?�:�&=����G]�#6$AW���e�?N���	�ٲ����Z�o�>�!��g��0G�'Ks&�������9�	]��"���=�!��~����u|l/\1���6���!�^G��J��c\o��f��'L���W_]���{����e<�8���	>���v��z�	�l�S��E���嵅�������7�m�]��'��w�<�Ea0�ڎ��X]���D���F���M8|ZҸ,���)�?xV�#G,F��d�m��@ǂs̈́q莂��/�層T���{m�Yl��.9����5
�*w��,�7kT��fp��:�VH��Z*z��<����}�@'c���#�����hn�"����ij|��ʷ	Ƅ�S�� N�}��� :��m�:�,����l��ܕt��� ��=+��j�^+����z���~�y�}� p;b>~��+/��1���R����z�'�o��x��J&�+!N�d�`���d�$�?Zߜl��ƃ1@&��z[/c��B�
�DMf�s��� ��{/�i&�'O�)e9�w˄��A�w��66G�����n:��w��(ɾ�j���(pA)}���;}0�:�,�]��Gͫ�VH�&ާ��A	�6��RE�X%��6�n3"ڲ�	n�����}����G��}�ߢ��� ,��'�����g��2���	Y^rR�J��X��=��;G��~GD\.����H�|����-께�kJv~h?[�q{6݅Ɓ]�.���Y��s���5s�j��.'�F��xi�mf���[����>ʚIܢ��G��6^��T��Goh����,Q�����ޱx��.A*ԇ�P���`;��ݫ�4����
fT_4퉰Z܇��ʰ���=}r�G�Ry�kU(���j���7��Ї"VI�P�������Ua�� �e�-�P����M���E�^6�	��֬��6NY֗�ڿ+,iAdX��FF��\��,N*��@q�1��n����6�yg�גZ�Z��ј��亲?$Y1-
җ�&~�J�q�.��3-.S^�%����lKŕ�\�B����@��ͺ��G��kTg)�l�/��F��Ś �4Zװ�n�yN��*������	��Q��_�A��뺪^�%l�Zo  ڇ'E�T/��i�7�?W�(�|�+V>ajpT'xC	��Y�q��7����.�.���&���ρғr��;v��4�c��_�쪏[/(���@>���\��ÀV�,aQ��p%������8�ѓ��3���L�2�0@�,y�:.ɶmc\#���A����D�[���v�p���5�>ѴS��I�G=�aS�ypq��LB��<��в��QW���GM�*;3k�`o���u����tI��?��{Uo�����+�/��y������5QK���~)Zx3��-ե��?�X�K���=���a����]��M�7�6�V�;��+5�f�神Vl�IX��	�뱀pH�>U⟨R����sQԴ�B�t��[uX�yQwzXh>:|�`%0��6�
5��C�Y�9e�ߦCC���hG������R�U,64{O5wq��T�c�6}�r�ozQk�����֠^|n�I���_��^_�/sgb��^�ǏM������������.�/�ve�`0�<~W�dqf��Y�Km��9���[[K�QJ�ʨ;1pq|�׷�?��Th��`_E㱊��϶���w͏�'M;����P��
c�L3�!żL�w;��5�"G?)��2nʰP)�������#x��&�M�����3��.g��x-�!�,JzF�Vpa�\�2��lc�Q �5}�h!�3��;eAT�=<2��Ż�8�C��Zb��CO�^�a��p��Kˈ�^����X��ݢ� ��פ�f�Z�(��e�]�"��x`ȏFj}�� ��h9��9J&���aC=���1��5qQ�S�ʤ�F��:!�n_q|h/��c�mʂ�|w���������,cR%�@%Z/�G�*�]rh�2H�@E��� 5�>v��A�ŀib#sΛ���G�� ����������-��1�;�I�R!��4��L�qy�5��⃒���+��v�v�#(b+'�2��H6ώ>!A�6R��S��!����l����ֵTK$
�c�$��}��et�N���7�Y�	����,�gF>~y�-�p��f�c_�<��ln<����+��z7n:��Z25(�5R�Q�"K����4�t��s!�/+\���%B�c�v��{�le�B�p3v�$Ӗ&��M�q��k��UY<��K��D ����iX֢��#aѦDe}$:��iJ�*uTV-� ��e�L�(3��]Ci��&��sʊj�:��8p�w���2q���q�T�lUbF�����KkV-*��3�R�QL��Ϯ�������nQ.��x~ŮYXH�ef=&���=�x"X�'�4�§V)+J��w�FPJ,�]k�h��uw�}��թ�e]Ľ	�-�茂�e�)��fל���r����{dO�-��ˉ��0MO��0�`�V�}?�VӸ/�J���M��]�=FI�	QhbT����'r��*tێ��Ř�/�WdH�BFb���%�#����Jy�e!�^p��e�O�?��g�໴S�9�l!O0Jn�_��"�j �p�r���ja!BpU٠̓��٘��ƑJ�N��T1zH]�Q�E�h���G����!�ђY���e���nB���F)��%�$p��<�],���h�r�w���׀��Z���53qOi����X*�5�w@Xj�_R�R�5�cK�3���>�R���N�����4M�?��O�8ȧ��L`$�.�4���\B���i/%��)7u��"u������{G�!���k�HJ����B4+ŴP�����Qy��ia��&���B��E3wO�$v������Ȝ��*��ZiZ���N$k�r��Cy�|�Vi�ly�6:��d��������(f:k� �
C��ɟ]��~N���)��W�f�l�`'� a��J[�Q#���Q[�Y�˕ 5p�!�
�B���t[ �2��ej�,�5������yM�H�����[�m�0�Z��̖U��$����e�\�I_�0�J�H��!���Upܶ �Xv4���Þ�9���&B!���*.'��#)DF�* tQG@�Ea2e�v&��jC_)�u��F�<�RN�<�rp���V�#�z�Xdk�h����*�.�ľ�|yL�)���h0�ɇ5y��e�7�rԒ��_��޷5#+�P�HCs�*��֌d�*��:w�1g�r���=��R(d�KÙգx,�{L����R���`�dFʑ&n�BP����L{� x�9��p��ג�p���1�5��g�m� ,�v�s��)"�}��8��1�59c
��R)���i����J����{���p�Q�/��C�b�� ,�v�t�nQX�����d�d����
)��P�f���v#�A�r�RnJ�nַ}߰_(�
~��lOE��s��*f �J�o\�����

E�4$�k*�,7,3��W�*Tzq�$ ͏�D{ɞ4Yu�*h�Ǯ�P�� �<F�;���^5Y �%�w�hW����y7�Hg�EuU�ǈ���$e%�uc;�V��ʔ(�U�;�pn���hD��+ڭ�R��$j
���:����"�J���7%Y�� Ԋ-b �H
4�t��E�J[QF8-]lgw�w;�.�v�H��LM��t������`�E����i��^ҵu�A�^��s&�f������o:Z���� �7?H�%����sJ��?~�&gFM���!�myl��b4���N��w���C���������Db�L�"�,¬nfP����E(� �
Qt6���t�]'������	��p�����bS��bT.{�x��7v5$)a��N�é͵�@��I �
;ΫU��J,�_�~1�6s�#��I�;�K�X�x���4�%6f<H80l����o<�q�
�+tB�m��Gv*�Z��%F�5�m0{��jF^.@`��c,�%� ,)#��E�����|fH�-8�%:�*pY�
[Dt�]�^�U3�=�ʵ@jo9�b
��9�hZ��A
)�C�̰+�m1��Re�q(�飛8��eđ������b��َY���[��g�z�
��K�9�����JώuQ{��c��T�ji�����������?�W4Wr��X������� ?�X(�wH0�)��
��@|<5%+t�x�=�j$r;-�a-9�6���JM�4{��|f�w"��#���Lq��Qέs+��ec������x�#����b62���.�6�J�"ʼ{ʯ>��d����pQ��K�06i�
t>.�A�Y/�;ͬg��tX���`�$a|���]?iz��sClUf���T���hm�cL�׶3���40�8�@	�W_ƪ1�3�y_��b�k<*�$߿#�$(��c�$� p��N�l������6�����v(~�zX�}�=�^�~y�a���3���n�O��C�ևF�d��u���7[�78x0UEfR��s��&�]�c�p�$����r���*��`o#i��F���{s/8�SWc�� ^,d�@�,��&�����q:6�η��͒(�t,�~� ʕ���	�zfbP	0i���8Ֆ��$N�Eخwj�,lb�Ѝ3��b��re����>6n�#�?�TE+�Rv��jz��NY��ZH���Í�������K�ҠnJ&���Z]���x	K��y�T�Ov�{rV/�P�B:.��
�! <�{#��iZ�����P'��(7v�"M������������-1/�)ў�'�Qe{e^^r>�����a��η�y!�9zp[��qt�)��z�#��q�q�7��2��x��
��?gB?+�SW��⭖�O���<7�ՕӘN��r���;Gsf�+rSg�(��o���ϱ NB7f%���Q�9>&���
n�%��=�;��a�
;�P(��^�m��k0�nWOx*#$l�C}�6��JVS��<��� ��!T�~~EnI�B��ke�Ϟ�>?�h�'�}�El�c�����b�|�{%��U��������.B5�8o�&>��2cݯ��j�i/�P�HY{k�x���io�#������6r��������K<���o���J�\2���zԪ���~��"�P�%8l��hZ@@��	R�����G~��@��ɾ=)��!���#�i/��t�`�B��]�r�[�'�Z����Kl2��`s�)�;�R���\J���uz�����"���� Żj���08/N�:%xf��>�b��-����x'B���oż��W6�Ɋ����OǺo���*����W9z��Gu}���	�9&���g��28���h�T.8;�x����.ӂ��r�q,�����F:p��� ڬ4��8!�v�M���M�Ec�NS�V���!��"���?m� ���BN��6=A}����IL�K�+:���]����9� ��f%���7���T&>�ov�߷����v�rd_�6f(��M�(��.Gx�\���)78ڽNԛm�x��()�a?V�"�E��B�|Ֆ��N-D�\�#�e#.{ѢR(�$�ĕ���B�[5~�M%�hk��7q�j�J��GA��^�I�#%SI�~�z�Z��C<�)�/����(8WcP��,�����3{�P�dU۫�
���lY�Ōl���̬�����El�'�!�I��8@	C��¾���[	KA|���w��S��j����p���c�\�_��?��=��r#:B��۫����6*�ޘ��Tt�#1��E�r�L�k�S]��Z=ݡ�oq'o��
n���t����Ze��� <��>)�Ɍ8:�*�{����m5�"CHD������h�u��Xg�)��G����\׉������N�x��4P�f�OR�G���_zz�˔�Yj�j��zT�{ȑQ~ �_�(/�iC�~-1�N��[�����zX	?��;�M��>�+����;ed���*���ȥq�*�<�6�ܥ8f��"�$�DY��v|��}~&Xb&�(�)�o�`������޶�P�E&6�|T>Q�w�8 ��[ 8f���%,��	̀ͷX���H�\'�n��]���o��7P�D��SD�Q���r�V&]����GuT�s�~� 1 ��a�D��>\*��z��e�e�(J r��ܑ]o*|F�f[�S�{��F�t�X��eH����9ɦ��Z5Пے��KW�J�C�U湕ڬD�l���5ֹZG�Rq%5�%2]��1���qWQ�h�M�k�r�-�B>>�
�ƞc�􍼾�Y����6���8�5q��to��HC�x{Ǽ��Ti����/�I膚:��U�4��P�Ѕ��`Qg��hn�����{�N�Ahꦐ��L����@����'�_�(�8ҩ��V�Nu*�etl�v��l@;��3S6�:_�la�7����p�BF�B��ϥi�-���_c���4!k\�4F8n1�[Ќ�2����1z0�#*Z�B��eIK���H�#��-�.�-����1r��R{�d_,rC�����:S&˭��~�?D��f&���C������{�:�a�&N�t#�杒�/�Y�.J���P�d��Og�'�*:������m���C;uՠ������)C��5���3;ƧDi�����i@�*@�	%�n�.���l5��X�H�[�9R�k�R��K��]M=�	�ͨcU�)����Cy=R#$%U$M! 2��bX��W��dl���X��u���G �._�E� ����?��@'�&�  YV�kX��:	qPF�J�ִ���{����H��y�wa��L���)}�s�XX�!1/C%�M�?�c���8��V}�Hq)@T a���Y�h�@���U���ni7�����Zĭ^|����ۤV|4!r^ƃ��1wD@�<�ą�S'�t^�nzW���G�F��ȝ�#2�(/uBv�k0WB�p4˸�Z��C�ҀI�|�5^q�`p�7	�V��Z���#'�HΚF	�����W�6H� �s�q�Uv���_�n3�y\���*M�*%���d���Q���f��K�KJ����G}S�i�{�����iw�w���Qo$���{[���u(�5^4���ؚ٥�T�A�a����~��?+�`dg�m_J+>h�s�q��CSr�X�y`��F��5�ɵ�Zt.�u흖�rqpN@x�H�2o��N�A"kP�s���h��c�5Z������}�>�9'�z3p���%��/���!~��j��R�D�m�#x��a����H� gȈ1�.�S*UNXf�jnK ՜��kJD.��4~�B����?�U�^��}Ëd��R�+��~����N{ǽ��`5Ȼ���SߒY����M���Ư�|�P��a�c�J��8��P��j�"B���kz��]�_�XKZ֥P��?W��������	�\>}&. nY�#��e�'�Ի�(-�nJzw؋�9U ����C�b���ؐ?-B5O��D�g�	�qp2�>,�Pfڠrҧ��f��:vaYgu�'���cԛ�O�l��?�@��
��Y��Ě�e��G�&8��5p�c��?��l-�NK�P�]��ld�』����Іqp#���_�D�+���DOO���2]��Ÿu��͠�wY�g�)T�5W�M�V%r<��S�6?���1i���>W1� ����y��=�fȠ+�i�Hi��U�f ���H�}_��Nol�JX~b�t=̐��'����~`��ڊ��Ƌ-y`�Ȑ�ŌxB%�5m ��t��yx���]l�|޹9��ٟ�ĘE�,� ~����C��7��~a-;%{���oHP�2�qῆ�3�3r	Z��ˊ�����������<�����;�^?�0����i���5c��/�H���d�!B7X�yDzȎ_>�K/���'Yu8/���rR3}쟊���.q�r:�P��ZP�u��^,8!����@�Ќy+zR�S�@c�����c�b���
����La�WJ�T��b��~������E�R���r��![�~�2��kpmO�ܫ�S��q��/�m�J���쓲�*A&zac�{���?��FO��ŭ�6��M)2�=au�<���+3��Sa��Q�{#
g��	ގA�Jڠ������H�Xg�a�@�G#�Dx�l{�5�ZjLlɩA9�$+%N��?�L�MA[VP)1Hl���/(�W<��b��3DL��P�g���2����iӱ�Pp>G��hq���G����@S�$T����ю��OI5�_�0?8��bO��5���alՉ=��6`[B�<����������6��[��e�ˆ|�`�ѹ8O����~��H����{��ga�ɷ�}gj��i؃�GU����`	➳�~ѵ�A�$���!��PM7���im	i�
R�;#v*��a�{+k�x��=���f� ��Р�ī<d��'�ak���^���j���F*��s����_��s�">l_!���"��;�s(�\_�ƙ �~�	��,d��4���(���OI��ܞ��i��~5���]����+>j�ö�l���+{`q<��_��ƁAj��|?�j� ���P8W���!���5�G��F�'�����5G��_w[T�Ҩ�T���UF�>�&K`�̎o�n.�y����!@Fc�x�3��`ͺ�ὲ�<�H;Ń�
y�I@
L?����f��KO�!A`�~�� �a�b�f�c����J2��+0��%	Rr����zpVx�m��_P���
����;h9�G��W��c�"}�R�:����FMa+��0��sj�dXg�s���6o�m�)� ������jӛY�k���M�^l�@=���u����9IfWk�fUk���I�dңqvU�Iy�{��w��2[�1��_����zU\VGMCF/�Ƚ;����|I^|�OU�;�g���wm1|*#XoUj��5��i�GqHS�ЭeDmLx������y�||����q��1!�ܾ�tW,Mf&��D���ZWox��ſ9�?DE<Y(��l}*{�A��T1�?�+'Ծ�J�yq���^
S�O������;Cm
yՐ�u4����ٍp�����ȾH!��g��>i?'t�[�T�uJt�A
X�\N�h��云�6G�<��௴I|�>��F�Z��}x包
�����͊9��ϑd$j���t)l2n�$Y���2Xc<$�мZ9��q�z2�V�@6�\Y|<3IN�Yc��^,����w�IEx��q͹�ZPI���w'��tz��\������D�c���`TH�U4�3_�R^��Np�+:d&gťʦ��'V3���U�]Q���{��%�^|�ʻ�{b��q��6T֦�X���r'V�Ʒ����2X.}lF
����g_�|����hh��s��ݑ�ebt�фL&� ���샴kg���K��S�=*��?�JP�γk���^0)�����1�bScVa��t~I����$�l{D|���D5����b��mӌ�9���>� �K�&|�b���ҏ�;S&ӌ��3/�s
Vk�A���9dQ���J�o��?��K!���p�D����PV]\������?����de�$�O�����}_� $(w;[��2�V�ȁE��-�kca�)�&\�[���6���dE{�؅Ty$���X�.��@�Zդu��N��Q����Al��0�|��?ƝQ�S�8x�8�!��ü	������C2n4'��S��kF/�"�^`{�Z֯�=����o&=B�v��*����D��>X�_`�c�xB�-�OcD*@^v=ϴv�O/�#�sj���]����eH���`�@N��2�-8��o�'r4����f�Q4tl��nt=��p����|�\�h\��{|�����Ѣ�l��z��	�D�6�^X���Ķ!�� ��t�L�ĉ72�҈KbN�Jd�w&"kЈG��fy�ܤ�9���+��9e�Ճ26��Ƭ^w�A~Yj�)C�F�gWx����Ӕ�s�s>?�?:m��a�zZ��]�2Nk��򟲫��a�P�l�v2��Jkã� �u�)��cjj�85.�a
��U� �Ǔ��|9��6��u��E�z�*�|�����!Ev��,�0�������9�yg��`�ce0���w��"y���h��RZ��䖎�N�caO�
���6ӵ�q�K-��9��Ko#�YK7���Qv�������C?EJ����l�S��-�k�
Aj�U�F �wn��$;���K���PS,��g%M��vu��G��U�uD�=@�uHHitPo�_
E$���L��s<>�v�K��X>���v3��z���C�=���������h��P�	��<R�����  k�YdG}���楆���i����eY����Ao�܈����z�;����n��k;흌P�Sȿ����ds���Ӈ��n��R���3wE�����)��*��vV�tU��(��	�mn��CG�!���sJ%��#�E�ȳ@A��H'Q'�����'QP)��I'Fj�E>g�s�E��%W���>�d��*>�)`y�Ю.����8#h�����[3$Շ�X�/��d���%�h8����ɻ2�dS.dT��� ��Y��xQ\L-�7k�������=�]*-q�yZ���o-�����I�YDn9Q���T*�Rܿ��[ͥ��gF�h'�R	�����r���kKZ?Dr}}��h� %�쳬��k,�v�iFMN���\� ���"���?�	5P����r�߾ڞwDPI��hei28��E�|FǮw=??n�⛞g$�2	>��B�>݂^�N6��Z�8�m��6�}�f� �Eb��	��(|>��&��)��r�9ѿ�������Z�����̈́�*.�˗	����'o=��Z)G[;��ͮ�{C9^��k�/��;�tQ�F���a4��+@[��R0���z�-��?`�5����+O�q2��ihZ�A����~_*� ��l1�p����x��	�����Շ�J
�ti�����ڊ@|B�:��k.�\ݱ/P��-��<��i�;����9�=&�����Y��$��FDgsBZ��3�j�������z�yL/��k��%G0�l�
��@��K��D̱ŪBM	X)F��J�$��	W�Aa@��(4��Bځ��;�S5��2���v�W2X���̞�b�i�{�8��L )}VФ�r��?��7��V	�{��E*G.�ŀ�m���o��5R(��x�0��g[4$���V�4�s!����OA"���t��."/��TU���o��g�k$�*�c��v EZW�,V�W��"����M�y~�uL���[9�މ������(�٫8`��]�W�R'_�\�w���뉚	byc��7��B����E��u�t[E}.�Nu�q��Z@�.�ζf4Hg�hަW�OlJ�2�/��U|(mqN�?�9u��z����C:�k��a��6!-&�����A�h��VRp?��P)�%��avs\�,	�?k'��}����ѽ�BB�Q7:�r#���� ۰����|sԤ9[�n� �ϴ�Z�DIw���w�x ��}b��lʞ�8�:�X+��2_�?�Ρ�{_�ZN\.j�F��2 uh�&JI�1�K��}�����m� 0M�����5��|��u��)(�&�������?ؗ�|�7�D��5�Ȏ�������ߴS�a�\�.�s ����C�9�>�P1��j?@u'���ChR����3`��ƸgH�w�eb6���S٨��_ ]'����O7Ӿ���w�k?��3[���6���-%�XZ{�|�����8R$�VO\�B�C*=�: )��ɚ@F�����UhD;��+W�&s��[M&z�CX�1�q��
�9�؏��vI�~���z�N��eu�������Q0�^����Ʉz��t��mzp��uuo�@V��2Ő.c�\_�����!}��+����?����Cr��]�z���Y_��z���=�ڶ;��)!g*�V�����/�+�(�'k��~��I2�qY�.�K��N����f������M��O�G����Mz��/��	o�����d2�+g�ہ�֌��Ř�A�c���*Υnf_��đS'�&�<Ȫ=S�!47��k����,�K9P�v�+��l�b-xr5��~�N$1j@��&T[J�z��-�^ԍ�H��hξZPS�&I��H3���2Ģ��g�����:�Z�٥v��{������X���E]��5�
�S��6̾��+t���[�E-�nta �K�wd��N�,���s���Q�:�3)�b�*�37��dS�V��W�L�F41
�\PaJ���p����w�t���(Q%�P��׸"Tk�A5(�Z(���ǜ6�%�>e��7��Ws�|��Œh�s�P�%�4'�q$R�D�za��Fr�nEҗr����m�l��YHeӐ@�Cg�8!��a��6�j�#�ǭ�|~"O�R����p�$��h�_
Ғ��()�> �b�-ċ��� �#< ��r�/hT��	B}� �$�g�1Y��,���6�V���`�R�\��H�V/(���ǚj�pb�f[��zح"��g$-�j�5Ξi���Tu�/rZ��2�i�@��;t���.*<S�v�)��o
����ڎi��c�̙�W8���	�����O���f>S���wj3�G]")�^2ڢ�}�Jz�7�f?Ŋ��?�%l�5º�Gg�ѭ[��� v�3to�ƙ
���QcO����A����o�>�����RzB?EA��S�t���ԓ��A�s*���Q ���H��u��D��L���)���s�^a=>^o�{�~���Y8�aӏ���)i=!`�}���I��-CM��L%��b���i���t� ~�$�̊]�� 1���$��e�۸����@ :j�b`�_GQ��h��h���kR��wqjAA��Zm���ڶ�.=��4������G$3���I�����C�Z�z�6*'�HB[D��ۃ���%1TY6�u����\B+b����ǿ��O�+��:mH�0�a-����k?��j1B��
��g�������X��ɓ^��ή2��V��/5gU�L>�,�,���_�t�� �}o�*���%�2f}4�2��$Ӄ�����iI�ە���;I�J���F+s����-5� �E������v�sV�L��N�q���m	�_�B@�1`_{GT�ퟣ��W��N�i�Y�R�z�U�mA<|�z����]�+\98�:����j`�	�-�%�h+2Ri6Zw���#Sq"%���W���������h]9��5��M�́�
>r�4�U�(�b��gP'�f�du�5��E����K,?�}��J����Gc0R�Y����A>���JY��~��c�����G����GBjk��cl��3]ȸ	�kg�oƕ
qA�K������	�42��e(^�]���/8�u�(HN6˪��'�����#ڌ��4Q�Th��&'s����W�hE��Bn�"!��'��~�rӶ*F,������[��<�"��rZ�Hu��֪��N��b\��i��奯	E��D6��?F�ŝ� ���qG��+p��?}6Х�$N�Bp�o�9��C��� ���~/ƅ�Ole�#���L#��Y�ұ�IUK}��A���s�U�M�ϵ�&?wy8�ؿ(�='�I^�V�����uo�Y'�u����ޔ�7񷻏[n�������s�(�II�s'�C�1�����`k��>�����kڵI���fe��߀Wd���
��ӆ�=J�?YaPiָ�N:o��/�S�g��W>��<�#�`i᷒��ۓ��Np?�kkޞ�|�H\�����U}Îv��\����[Y�{���I���4x�6iܣ�7m��[�9<|��߶��l��B��B������Ւ����I�)���	�?+��c��z�TX���2��g��� �%���T9��5��qՓ������>�#��)F	r�^ר(Bɩj�	��GD*��Ky���ϡn�`�ɫ��Zs�o����� 1:�֨��C罸���<�k�C��D�=�9���aݴA5���T��Z��������5�jx~a�_��1��Mc�V�?��1�a˪��F�-;YǶ� ��E�[���Ú��BG�����W��a�����0
��(��0?j�h�<�8�ſ�(\�d�F��2͵Zv�-��d�sЖ�/y�3 E�Z��4�u1*uj^Z���Lj#����w�8�f��9x�v2�]�Ln9���I�����Carb�]�E /�'�=h��\x���7hm#W�G�u��3T���Y�ώ�O9.:])� �~�RJ,��龈�q����8_���v����@Ю*W��g�a@�D��%��~n�����>%�9�]�8�%�^K�󗦠�-M��HǥhH7zS�-G�L����X���ǵ����Nyv�V+�܁���5o������"���G���#�+{��+9��W�X_MT�� 70��k��$�ҵŪ�E!^���r��k5���HȺ�y�H�xA^�K����;6��$-�@��E� "9dC��v�¥`�|�ua:nT!��S�IΗ���<\�0BV[�"a΃��i�����[��#��V�:��V�,�l@��%�;g�'`�w,�5��q#�̒���ω��E�ǳ;%���Q�C	��/��t�S�]b- ���)n��s Ce@w_2�����lȹ�_�%:z��qY�2H=�$�#� ��A��|�d�T���|�ptN�" �#f���O�A,%���d_OS�V���y�㢵L��ن�Tf�r��`�Åw%Z�����l�,aI�ލ��N�:M�1��`�#�F�@���[N�q�p��d�R�N>��[>�H��޸C���K$��4��:�.��?%�"o��?�昸	v�eոV�\��E��%1�j��Y�Np~vT�6 �_\w�e
޷�i�@��Ǚ�H�v_�]��ö�O>��y��T�:!�^�y��7�j��h�߈�K�J��d֡a�س��N/E�
��h�-��ދ�p�����/eV�vn�iGǊ�OK�����5�_s���Ȣ�	|{(��$xlO#u&z�p�	��y�d�o^7��!gO�ߒ��.�e������.�OQ��e��&���i��N-]Yl�Aޅ����X���E�:��u�0ub�߂%����v:�Z:d���i�j�l��'�#S�������?*4���Q��.����E`Br:Y+?:^j�k� '���O)�X���{FD��"Yp�����}������]
�nT�	��@��}���5*����(2���R����U���V!��g7UT9�n���V��9`�(5����%x������/B��%�1�^�w���oc�E쳣��X�g�Wc��m �ş�He^��5�r�[�����
��&�C�[���#�\��H�5�߲]�t�Lw�V꘧�mjG��_�M)>����h�ZD�b�l��.`��ᇺ��}K=|�c��{3iy�~�MZ��"�d>�zoN[D˔rޓ$�U�M:t�sF���6�~��?���A¾���� )��*�8w[�|=<��T��f�Y��bXڽ��Պ ߴ��`"o�g�z ��W,}�P��y=S�s@��S�g��Tf�]N�3�T����c�����K���7����f���R
�'�&ğ����9�T+q�2���.�練}�ʭ(.���+�����d󻝲��E���P���lCZ���u�YI*\�:И����Ԋҧ	�r[z=�S7(>���Okp�T��SQm���p*��>C��*�T�	����\�;���,y:
:�0� O,$nHr�_�)�c��e��.mp%h���I-�%��Rf����W�x��o�ld��
t�F$�|=���+� ˢ)][v85<|b�ήaizHS��g���[FWX��F��K����kDkY�G@�!�(�p,�ҨL[��x+ǶY�=���m���|��9��=a�Ĝ�]{.��I�>�b$XD�"�A���Ϳ�D���צs1Ҹ�m��!�i7�Tv����W`@p��e�M��n�&	�A^���̎��"��m�G���΁|"G�*cx��wy��"�|��/�#Ǣ����O�����8x���Mt^i�*vTݿ�ҭ���+z��<&+8]ȋ<����1�����2rU}Z�Q�(�HRf�&E= &��-��^{��.\^��4:��tj)i^����?7�^Z�_�i�JjX���tmzS�Q}\n�	Q����|�������)z�y�T�vW.p���:|����%�y�}ò����s�F�3�=���@�p��e�~KN\�Rx�+A��d/����蓮M�=���X�P(DZD��Ԩ�Ȏ��R�����
�����a�?�r�^��.�Y��5�%b��Zk�:b
�� W,gtjD�ŊuIǐђy8K�2tH���I���2�jk���]���5�`��:e2�q��-M�
P���ֶ�V��-�TC�S���0�3�2].����M�]��7}��)��� e?R/����h�(}Fk��g����zM�l%~s�{�F��O������l§�ʸ��2bR��cn��Hm�\a�aO~�h��b?��|aLT0�.d�Qk6�O�3!�i
�f�ZW�"۝_4x��i}i��!�5nw���[�AXg�M,Jԉ�^�>�� �����c������e�eoc�O�eL�wb�Y�P��ͬ��\�R`��Ӂ�@n�J���#��z�n�&�H��?c�S�������]�����N��_dC:#Ǔ/��TaK'I��&nu^�� ��3�U�+�0$��V�1qբ����b�#����F�~Z�>m10��7�U�<�v��9��R�d�>����W�6����+g	�X����U�կR���~��N9>����}`;o�[($"i#�6?�9v{�٭�"ޗ���X��=��.}��pd&�(�v�l��an���b�}��tO�MG�z�Z�_�F&��<��dj��FV0^Q`J�im�q:�C���Gܣ\��l]bMxm�i)tx�Q��Pj�y�R1ϒ���hm(�#M��d�1-6�7h����_&�y�7y�ngz�U[���r��[Eϒ�LҚ���#��[ �O���"B+0҅#�MU>���,�	S�����v< �@�3h�jsHC࠶Ů�硑�w��z�$b�<��\I׏z���;�2��{T��r��8$�`I�d�%���ۀ��'x���]�/E�=m�K.'���ck_<ҫ(���2��dh'���j	g��lZ̔�^�=��B 8�'lxچ�O�J~=�`t���g�<�*��[��i1.�Vg�����hF+�׍�[���ܶ%u��1N����8h�����>���ڋz�?pOqF�݋�|�B ���5N�Xb�G� -��*��5]���������_�+R��0!�ӆ��bTz�+�KG��@E���!�I<��-��pã��0]�S1�*�f�0�'v@�!7�H��o;h$�ԩ�ƌ2�qf3v�o��1�� �@�܂��k�������G�?[@�B��,Td�,:�`U����-��Ժ4\Ycg��a�!ŝ��ʡ@VK��9m�ra	��<�
�N8��:��d5*��(o �E8�}zT�O��]��h��%b~ޟq��^f3�*Y�{AX�eN�"Ȧ�6�2m�R�� ����aQ��ץ9c�>q�������z�@X,V��P�P'"�Y����u�idM�ap��Y����p��_��FQ�D�7�m&};aξp6��m���ts��5������ܟJ��z=�)� d�~Sț�)'9������VN/�����t�*��]��l�����V3�/!�.~�|�g9����kA<���
O~2�͒��'��s֘8�oz��m����7,���#�ETJ����>e�az(�E~�%��j�W�s]v`�JE�pJ^b_ϲ�?�4M|����
���1�k���	�4ŝ!�z�g�Y�#x��F��)�A�8;�M�~<V��D�غmj��:k$��V*�z����48Ƿ�dS�y
� 滯�n�6�m�n �Z�(�;:������M�Cy��0q-@�#o��ො��9=
g�V�r5G�Ls��?^"<���Uq���σJ���b< ��<��N��\.�t'�cZ�����f=���)�y��pS�҇������].���۫s��_J�eQq���M��0h��U���>J��ZG�@`x7������A�D�9O�>C3�9��y<S��Gb�־��In�J]�H"����_0O�FX�����{]t�� O�_�{Wu:�v�7�7=��n�jsi�v�@