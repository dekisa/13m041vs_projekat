��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����Ղ6dJ5c��~�Z���ͳ�����t�Ay�~7�3��;�G��_��+{�S=�$ vJՋ= ?����DQ�Lv~�hvp�!Mrzy?ڔf��E a��b	7��s�&չb/��Z�F�bb�%U�A+3�k��<�m+�uG��u�zVG&���j,��D�2�@P������EjZ��%,�p�28N6����EZY��pç-�֢���@���#���wʯ�6,q�'#,[�vH��A!f��}�Q��0��:���ba�r�Oۚϣ�V9��P;�Hjԃa��ֽ�>Ym	.�����q)�YPv,g�%5��L^2���q����&���d�OtP�Υ4�=���Oқ�
[0�A��`���Wį�!u�(��r�B�y.0�nvZ��+�B�v��Sln�7�|�$^`��${�ڴ��$�fm��EH01x2�8d��O2IdQ��!����vJM>���8�T�t���rd� ��0[Ѩ��`*�%�y�S�YuO�Z$��R��R���!�t�\��R-����=��t�'��ȶId��.�7ė:�p�Qwꃥ������GVpl�\�Fm�@n���k�G����F��ӓ��V����Q�Rr�b\���@�5¥�C���.�/�T6�Z 3>�O�2�Gk�C5l�bJ�Iu�x��� 3��b~�,����T�]E�4�_Xuzf�/�"�%����+�|��*�:DľQ��T:���p����H��P���$/��0\\"Hb�c�8�z2��F��$��=�5ְj@=Iz�B*�� (��[���[zn���ɖ2{��P�[�Y3T�7t�c�ѹ�k����0|mq��_�?G!=�%�%jd���@��(�B �O����E:d��VVKJ0�"��65z���I���TZ%a��k�H �G@W�ôȪ̙�hA����)��S[h=Q;������=ssb��)l�eo��s�2Q`�ا<��x��v2�?�{����Vv������/r��H�C�l���uX(U�u��ܶ��y�۴���� ��Ș��W��XԅҴ����b8WI����)���ӣ����
���]�[�N�7�3��+�;wIw�qd_�A%�T����P�*Gz��Q-�j�f�y�;6��AP�D��aCp�!����2��������ZOp>��푈/�檓ñUI�ϖ���𰺸X�O�`]�H�n����-�CU�^��Y���ë��хН�bR9�[�E���,c3}+�sw�c<g#(fb)u�74�p�$7>e�~�=�*is>)?�J2:]��GI���K���H
���1�8���1w_�؞������\"a+~(�!cvY|��\ʏ���M^��v�8�%b(rXX���w�x�.t��M��[�T���e����$�2B��t��iI��0��ɻ�-V�)t;y�+j�V�$i$c�=̍�N���bE�;w@xMͺO ��Ear�-�u���N�e�K`�-�my\�d%2'��IN�ާ�}OQ[�9 ��z���������M��us3��`T��)��\��y��cQԼ�o� 0��S>N/�>�V��P�Bk��iw�����Zy�8�DNEҎ�`	�ѻ�ztCe� ���~ڕ[G(���}R6�����P@�0���KRB�5���ۢ���`��`-�T5�!c0�`���RđlD���>��8\��,���+x��~<մ�`P��Œ��K��i�����fj��Aj�������њ�5$ne�q�o$���픵�v�ݑ/k�h��4,�HM����m��a�~���@{�Ŷ��3�:�x�V���P�:A
�Wg/�`,������J��5�M���zuC&�?�)�3��_JH���*f۷<o��ug ^7���Is����oB�?������~;�/����`��2ڏ>������X�Hqq�w���p��G�&]�9�K�\����:q��]�z���l�E�wIA�CJ)y{`�O]�����h)���>��Dt0_�]Q���9aK�ǈQ�(TT�J	�ӎ�N�s���a��ӳ���c�q�U9��=l�V_]�6=���l>C�w�>��Z�;�i��i��e�t�>�����:�Y�M�&m>��֒��R����X���t����y��+~JkE7V���ؔ��6b�J���e��e�6�����h'��,D�f�1BH�&�T��d K�mO�239!�l�>Ɵ���>L�[G��y�7�I�4G��92g��K�q_��NH�x)vaeS��hZ���#2�ȋ<���
ϟ"ۇ���Q�&������B�����&~@�\od,�`QT�?�~p��H����U$�V_�Kz�S;��w>Z�
/��E��]��3�\;X������.zM� ����5ə-!��-���A����/�R$i~����p�߷yŖ���95���1.Z5���|9vʊ8��:�=Ձ� r��z���G~T�w�	E�>wq��h�Pn��ӿqɹ�G܀p�َY�N2�H��3ЕJ�⚊:�:��t�-h+2T�жX{ps�Q� �Jm��}����W�[��˱Ra�GzP�K˷1�ȣժA��&�OUd	O*��f��l�2~:��*��R�k��|m��|�	$a7�����H�g�#,���%a��2r��mn7�p����%)���PyP7����� ��a�����h��>�4i����>]�(�1�?�V���.�럴I��EOH�c�?`wk�F`S��G�u/��$To���\u�t�ψ��	�ɽA"e��avo7o��K�-���W �c�S����u���ֺg��)�A�T��q���w����k�������'2����*E�m�4K.���ٟ�"mVD���EhK9�*�s6�CFSf��F"rҶ�+]1�ߘV�����_P��$s�|�	�����h����-5��:�1XD�b��#��f���%��,�=K��V�GBReE"pw�2+��KcՅuM��������A�Af9���[%х��h\,E��V��4���9nE־j�����+۫� �j�f����S6��tB���?Bz������f����¤|��
�����
e�Ɋ��X�kE��¢�k4�(�c�NX��_���U_%�?N�=9�ԭb*�< !C)�J �������"tSB�hN�q������0w(b�:�z�a�z��J�������z����E�o�v�f"�|�_R�?�Ə��Ba� �0"@���nV��_�S��H]�}˼��]���n!hLH����~,�I�j�]��zDҍ$E)\� �6�l�D�W�*2��fT~�BPB
����_>:2,��E��{Q��x�q�uM��Ν鶓%f�+����ì���Y`6J(�cw(���2����t�g�L�i��iӘ��������L��F�'R6�$CZ;�9A~9n-)�� �N�gz��+��X���s�.f�p������z^�r�6���� $�	Y>�?�o��ʐ�8(	~ַ&lV��(�v�
:2��Q�MNRp���9��H�,��T���Z������<�1� �>]��V^�#ĕM4���B)��m~g���_���D/�0���݄��,�Q�{9���^��vtb�%�� �d˚��SS������2U����C;[C����6X����� �c6YǢI5�,� �ju�H'�+g\!{�>�U!HZ�E�C���OAD��������$p�&mt}�#&��4�)[��Ẉ���&h̉�s�iq��)mEU���}d�.��角a���Ĉ+jQ�AWJ�vZ�e`Ⱕ^g#o�K力*�v�:jNk�a���fRC�F]�Q�{b`�d���_��R�Óm��;օ���]ɰ���KeBg�Suc1Q�^`4)X	�v/cآ�T�E��s�
ܭL��0���捸��.�^΄�D�0wY��F���?;#��r4��A���^<�0�ؐ4fL���P��p�0�^��N�Ջ�����!𿖴�.�����K����ƉKB�1�ռ�e�!V��O��⏤�z��J&H3�Fm�*B�֦�T�݂�!��z��"5��-�;G�cm���R��0�G�������ZLI����֢5|V�KJfz�(�hr�#y\�=)0��C�S+�y
{��ȝ� ��8�7B�b^F���B�`	귆���]�Z�17&y۰97�9��+5��86G@�5$ٌ���|�1b����+��zvxb^�Y�B�I��6:Ý(X�׃D�uj��B�U7�v�|6f|�ᡸWM�~l����J��թ2ǎ����(��ʼ��3��	O�4�s ��^�	�@�VjN����k^�g��$�Qe��`R-3-YPV���(�PLo�P�w�е��e��=`�$m=�H�a|�6�Z;�Ø]�����'�|ú5?�r��*r��P�)��̃`1pk<�Ab��m��H�TcT��!���R��.^�.��7e�F����U���[w=��ه�K��>��e��c�V�\íxq�y����Vãօ[����i~��
���l��H�<*���_g�|X��Q���F��֙�P���V�-	��q��
��On��6�e�C� �ɖoM�$�&�i��ȕcb����g9��.����e�r�!JZh��Y�/QE�mb2�7�-���	0_�
`_ŝ�,�]�N;�5�?Q~J�]+ѧ���~z��o)'�W��u�
�K� 
���(DTS��[�$â�`(O�q �Y(�y$6���r�U�^W�W�c�j�l� �/������)7��#.b�-�R_�8<G��i"�T��j��W�ޙ:�����d���a� �@��ȸ�*ܭ�Jr�t����n� ��Pڼ3�f�xeU�n��@(B��%(�h�1n��Ɂk�lL�3�W�P0��_���[|���D�Ha�E+�?��cC1S>��ӽ���@�+ �W�l�%�]�5AI  Gx�%]������� f%8�΀��Vh�ܱ�e��g���eo}��&��~h|#6��Hϻ�%Q������c�=v�Ke��$ώ.tI�}l������8�{�28߿|��ծń`$K�<�
Do�PH�%��(�n��.�{'�_e]�R��*�A)��Q�B��}�#��1;���V�����Iz�� �&����>��=�gZ��~���A��E�&I�#	e�(E�L�����p!i�����(:AH���B��N������÷?�S�}��ґ����H���:!��#�D�ѐ�;"(�qt�ҫ���{�3��,�	��8���'�VF�	��D���|�ĤWn��/�?��KdFR���(`��8Z�d�+��;KZ�U��O
�(8��&f!r�����#��2�('�@�U�������<� T��|��,aD��͉`� ���^=	l�Fh̄*��+J��آ��y3���~��Ʋ�Kɨ\�,�I�|��HO��/��f��fR�NT�WNL���{�V������f�\�0���}DZ,��]���\9�	��L��E�t�����A�hXrص�g� |�@Ȏ�O����hE��a�y�^{�N���~��������$��V.���G0���Yn�@��iyr�dKa�"In8�gǝC�e;S��=�K4tj�Ù4�PDD��[��&�Y1�-{���~��UNo�l��6�?-S��_]m��n�N��vf(���G-$rҊ�W]=\V���ࠞI�ϓ�q��X^< �� �d��� u���ʊܶ����v ���;�nTW9Y�(�t]��\5��?�!G4��vK���Gs��"�)&݌��"�6-�^�n$iՖs�Uj��p��(1E?����;w��f�3���M՛�͔)��\*��\�yMLn���>���ݏ�Ŋ�����_7�����]D�ҽ�7(1ژ��Pdab�����`�d�~&�X�⢣�FX*Ig[�3Q��t���"�x/Bf���V`�j\��">��Lu��BfB����D�x�2w.���`ghy���qaH��s����pDP�?ā��D�	���'��VG�$j���$��:U�.¿!}��5�Rw�x�傖���!�8D޳���(�n����Ukdp��>�.�[ϴL����]�υ��{pD	V��ČD:��c,��OҭoY�ȝ�?��Jx;L��.E%~JNˮM'M0ޠ:.�D���H��̱�w�("�7 ��-C�4���
�4J���������|��&e[�{7���so�w-�c���i%>S&���;�T_�'~&��-}������9��__�s��$���yr��M��wo���fN�s�L)�۠���Y8�eK_�jL_�T��ӈпܩwxPK��ޔW�Y���WD�tu8m�L��wu�Θ�k���]��,Jk*[bTՄ}�w�~�m�.V,�O�vw11��_�|;��Uo{E0-��Re��Sko'���~#Č=}q}Y#�>�X���^Z�+�⹹��p)�;�����Y+)��g�'�:\���l�1�Z�S�v���Y��-�$F\���%�Y��L��`wˣ�z��˛��?]��@7��z���|l݊�ߒ�MF���.��N��hb�;�z�ރ�\lܞ�f�n��һ�[��^lP�S�A>�"�	�`�d*a,)���o�a��K�� ��0�3�ࠪl�d�5ԓ�Y�����V��]zβu�<��A�&y����D�<��8rha�U�Ԯ��b?�`�:�>�����9����J�.p�G�Gnz2L�r+(���#��xQș�d+�k�˚�+̀����k�_S>��V����F�G��4�w=�Ȫ/�Aݳ�
<����L��Ӊ��d��pQ�m����[��#&Mg$��	I�q%
�9DT�ɭ4W����ݚ����}�<���Q<��,��$�z�aM`�*���?FTơ�AK�5�'�D�^q������w��-*�֞cEQӨ�m�����v�@dIG̯����Nw��YڟK���2��<	j�T�b��̄��Xy5#ѽ�gФ�m�":�p�q����5�H�����߮v��9Nq�;89B�d^!I�O�;*��qŞ�����G��UEu_XCΏ.�x	�W�H$���l��n�����i��۽�8
���ڶۭ=1@�� �@�o�-�Oc��7PCa��~l�M8�	萺2[E���aY&���=�\�>�P�@.�PڢX]���[{=�fX	�V��2rW�ɾ|��ϳ��?�4t��>@��E���6�a����s :�C�Db�F�c����t�5����^�3
#c�#"��DvM�j�Cm����P �x�B�0�Iw$B	��HT�}:�GM���1������CP��8���#V�i̧(�b������EK�K����'�
���oB��M�
 ��ޘԷ��97�`�L1{2���*�l},���I�f5�5�D�ò1t���II����L �k�}����-S�M\�8�[��5]���͔a�cI�o9�ҹ�^U����h�f��-A��h|9�3W�o%W_�pд��d8�;p;ҝSɫ0p��܎�00
oa������R�4�6��B��$�ׄ����T�}`)�lھ�~�D�X�3�%��V�z�n?��sL.^!%����v	�K�$��c���T��dNq�oD��Go�������0ݭ���hϰ7�C|N�Q�ox�R�h�E(epZ�����_�ܭ�(�� �K�������\[�pVwb7��I�9���wfW���C���H��ѕ�����$�㷟�Ӊ��T��B�.e���:�`�8#�ay�h���wV����B}��j{H�Z�R��+5�/��,�r��G�h&P�Z��a�?jb��y6O���We�H>)�WD��%�A��������A]�xNI�@/��U%����E e$���Db8�l������>)����� Wa�M'����Hg"֯��$%a�q�eT1�K�r��	���S�o1�2���>+����Z� �����@��v�@$������׋]��tr�o��-�NA,�B�q�!�0r��+P{Z�R��#O�Q�:8�P��m��7���-ʬs<0�Ԛo�4ߩ��lw���g&����͈���''�Ws"��mmO)��n��2���8 XCb��G���O���0Z I,eA�&�8l׷�!0�Bq��(G�hd����襺)�膣�N��fF���U�cXxx�G��3���d�qo�l=䂝�;�7v�Ͱ��.��8y2����S48v^b����T7
�����R���n�ғT�m�["�R�R�c��!��}}���b��t:� Y)t��c���]�|/����fDw����RLW�-v����яT�(�����e=%D�����bX�y��8A� ����C3�����h��AS�-�!���cHK���3�0��b�,�N�hl��f{�ئ��Ğ���i���F�Oޅ)b���Bv�(Y�e����J����Hfi�8+`����[]����
p)�pi����8��k����]��+��g��"��8��Q�Py���J�R@�ϑq}�|UC�ϙ^>���
��m���M�.C��hz�#[] 35�4���a�����\M:�o�Ǹ^)P�����:U�$��?��A/�N���G�B�i��.�R.��n.���w��ۣp4��%ֿπ���'S/n����_A�aR�����m���:s��R׻��-N4�%k��d�%/Ѐ)�.1"�	@x�%�n44�Xq�j��Q��bJ:�EO���0\̫�[���_�O�p{�c�C�7������z���2�����M�	���F�������[�y�OF�m���=�D�c�׸WMC���K��~�!�PX��sڵ���(O���R��Lg͉�}�!1�k)w�iLL�k��2~���5���{}�-h�
�]].k�+�-b�<J,��ظ��KE�'?f�=�3yfWs8$�Ha�<>_k;e]_f�7�Μ�����\��d�O��}����F�8����$ΨП�8�m7B~WvTŁIUM�~�e�t��7�3;|@���x�c��v���d�>�x�,�{
%�Z�ؖ�i�fx�D3&�� \�
�:C�6��j�G�ٶޯ*1ة��ac܄�,�b|��qԲ�T�����<hWX{Q��ĝ��?'�>A:����9*�J��Mlչ $��aV;zD,�AVc����t��L��Ú6��-�0����\g��<���#E������hx�c�j� �cb"�Ds:�Q��5�T�Qk �#��Y���{��'y�M� y��xtg���O�Z�X��&��SH/� �@���zZA�mm����t�� ʋ�κ����U?L;R��K�[fĶ����e<��{�ɻ�t������SWAx�ս��/q�_Y�m�Y��As<&���v�˴�(%VD'�ܖ`s_f�ɹ���<���:��|�I5y���i�=�5��ȩ�#���eS_���xO�6ϝE�i�5�&���BR������aȲ�ۻ�kd@��ǩ�\�>D ͈p���<�N8��k����rb��Au�)�U\CF��N��Wf���e��5��<�cL%D���W�/�Ş�SIO)�x�˸��Z(h��#!L.p�M�pyמ�ړ��4vj/4,�F��l2��ː1�����Y��,�M����j��UqU%��j|R:S�Q�Dp��zK����ye.F
�+�S�Ea{�Vع)c�[b�F5f�J�tϭ���GJ=l՞<���U��1�!S�u�/���Pʵ.X��d���%��ێ�(#
1���WkxS�zxG�ӟ�=P�,$4�)M�u��e$(�ޯs��QR>̕�C����Ź�<��8�P��/�K ��v~;�kޔ�4P.��O��p?��!�#�J��wT����FB�ʆV���%U̐�s�U���P{�2��ɨ܋A~�{�T�5���[ǐI�K	��*� Vr��������Gr�kN+a= @���S���Ιt�T4�DN�~��
`2_||.����>#����	���j&*����- -�_VsgfH��tЅ�p9�Tΰ�!"�}W�-��H�}�7T��ɔ�GKgӕ,�}5|]��G�0,�Sf�����������$��l������n����V��<��?�A���VS��և �_��B��Js#�O�2��^:��$3����ԫ�� �4�!��a6����.ppH}k �{"�1����cP�C�yZ>�G�E�g1e�2�b���_�0���4�ܓl��|r�ZsX��wX+� �}U��L��.��B����-+���*��rP���1�BE��g�r2�hџ��cխ���s�v�'� ~81�V�:ZCz��$�f�4s��o�����O���{�wr�O�^