// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
udWEo6+GgHgMJB5EVOIV04XWJgHdUtCBMmdv9UYvTUormuxEmSRvBX7vj4qoNhNs+rm2xq3KKRCJ
Xphiju08HlYWJY+yj6+9iIreZBoaJEn1u/4I/Pojkf7+6t2Qd/KqSKTwpDlHTBfIDhbrmfDSlBN0
h6itwSu0YrOJwkTrqfdRzENDgiRTnLFmSGfqM6VobL4xEBH2obzwEkNF/SOWCRSjPeZHeytXqRya
JM3WQvtYRkpTpooSoin3b7Kui3145jrO5mhk7GofbdjASqx4j3s95QkUnkaYv6a2w1tMk1O06YpQ
+l5vh4pY+MRayk4onGj3OWRPQWKC3bwiCdeLqw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17904)
LWLmq/LCjxoSBy1gB1Vc/gNemJKMdfMxkL8wuqonFc9x5f+Y/3Typ6xthcVQBZvxHjTel+vjzIhm
xXRpyzdKZip3T4ULoIAPdMTfPEucEM9t8grtUGz23Ap5sZBReVCh79KVHRlAIfdwbp0qUfW2Dr6o
/1LxyjNpMTKczgS524mMxgCfIlheoebjqF7Wc55snNHnORpF+r8SwkYTGIRVuijNzaAE4Iuj/A2c
+sN1dKSUxV0Bk2VpSAuMzfiCgy6KP/vkNlyHEzJZ3UFBs0XbgiK1WSyjQnaQQFEp6I+BmBlveUdr
jSTw9hNAPR+AqYg5rZMQFPCDjGW5BUz1iezhCSzIfWsf8PVTTMvmmpLu5JTpG0KOTPpIjuOoW08c
nNqbRzD87xVh4E1Q1S4awlGfyTHufuYGygbb4yqp014/Sjf5DFCdVSk/LFBIEiJsWLOvq9QAQURZ
Y7dxhW0sLaTzqc4Gr5oUPVwMX913uQ9ThnkKoTnhdC+aYkIPg3ak9h7/D+ELA/W7vTV+izFEPQrb
eInLa6aeiOh4LCTnX+IbbB/ED2XEMRusXE4pMubGSIGuLDmTIgfrC3YxrKXxiNGozDcXC6Xf2+p0
yC2Zku54sest2QgEDZeH4zh3WGNTKwVdVWFDmEqO/D4FhooxaRe+nxUP3TnsGrj5uKXODazBNrvT
RbCZ467gS9jR5m82AujBF5vgNEUW50Cow2APOgGRlDNQTaAjWp6QJZscjD+yZSLqNANarSMBTIeQ
ezdyFNuduj6KeA/Pq5s3CRhMGq+8BPFG59+5za2Oht4qJPHSNuZZ/umG7/5rUbEBbmpQ+Efm1Jfy
6n6d8dUD9r6BencAS+pPbszJisrHrCoiHxcuT6kH7Own7Lhqah1ocKXFRhDikYgAtht1krwC3lDW
pgwVcB+Ttmx9SviJD7vOb+bKeYX8d55U8aKwi+G4qsUApGQc0fnkv3ezLmQDndNa/UD7qEfxsSxK
FqZ/m7vNSniQd5CL9H59GK2v14slC/x9QI1cOC3dSQ/nj/Ci1thTuyfOvHACy7ZucIFsNrOjqjiy
UIPjjcPVOMm/WquokfWCV+ngQnN3RvfgxTnX+bUWXUPtYzq6siy915YVHkhTbA3gCSokMfwUngR0
JsJNxYtCcQVuDeZx0uEgJSd+IdQUGBebH/Gu4Ip63GAXOyQ5DmYsAPT8Kzjy0V4JsmjQ5IcH48p/
sphqTC4pPIxkpQ8r9u5sjoCkwlPweYCrnRCGFqCjym8XDX63MSXzHWmHTha3rFLiCL9YaotfU93J
WkKc4mnDiOrmo4zF01CsIYAktW523FDUjRA8ek1Ba4cqBIiKA606Pbedgn5Ma8GNq7XgT0vJ3DXS
3grcIQCwi43b6/cnG+VCIXlU/AQ/1oO6uQEnRkar8cKusGHZEYK9QSvVYQXUIrqdaxiJYO2zW+bF
qb9/gckTUYZ8Tdxx+DiN3RwOmr/27+Cdj9qQaoS3VbpZyYrYAdlf3snQf6r7jBYYMU+MoTyZpVkt
nHzbULWH3MfYhCS+tS1n6bDlP5qhMtn+Qj/sd9+j4SY+wmWmRJYeSFy3WRgNkimIimhCa4n+/qQ8
BECc2k4aAaLMHgRi8hm0ORrPFiWYba/YNzhJ1l26L43igk4Mj+BX1XMN+sMjfAlex+qUjWFlJIGw
3yLbcegUwzI49zCwse/ysoXtOoT66d3LE/tQf0JedYSSK7nl2RPtZEb2CWwFOmTaL3sAHksFdWt1
kcoRXPpbcxjR+PvwK+pfGDjY5E0M9nrVc4It7xHu8xVQa5BZps4l58bUdYyttWb/AjF+D4jUf7gJ
FgDapMO2iISorF3UUinn+MBzvQkyfdi9TxvZtywZnOek1aVEtGC4mACT4TQUSVVQ256fDJ0dxYE+
McDe0b2/lpk+nHD+RfhdGux6d+0Yzne4kzSnC2/cILfHmLJs5po4x2nvdTyqFwOXCxKwChTDpamQ
LxifiY+dW9zBiEik/VLNpfRW3DyfIEaGBSgTGM7VPCLu9Fqx27+c4S0y6Md14Bo/5OZeEbZHENr5
vtCBRlc/04IwPoJWkPgTatKdcj/vRhUkZI1O5LzOFNsFSoOmyotI3dk6aspA7vYDa8bf7DNlw931
S4ryuyEjdJhABQnf9i/HWoz5UVX02rzYQ7pDa892yKELacvd4HvdNYw2CPCdcR8fLVWtBdCnp4x7
ebanU5DvbOpZParHX66DaMYJ5aOyNMeaE2PNK/gOjqvE7Q1arg9I/R5g0Xj0nLyoeJN7awiDpC5X
mFzFD6QeXpfz6g4rP3BJkS/AnfAq4M4lw6C40PLPnprwFhnnrOnEVUiLDapGsNkqYZRmlRUHMk7c
DPpNPdogCY/g0YX0R2PjLytqjwNhcgF8bkS3y97QeWY6BspGGrZwPewBsD2Uw2c00sZWV6WE5uwt
QZtf7LGHfgbbgK/lWfjb4CsxAYrZFcYbiKO1dNg3CRCeJ3UdGW3q2S5mTn01Rt2QweqCovOp1JQO
466OLV8Oq5ZPZIju8+aS9vslsk9NS4DdJ2T2X45ltLR4YzFj4ce/QTp1ZYuym0W9izDKUGPzoIUJ
fDL0kGJhhanvcrCGTQcKt/p/ttiwMqqSpF+4A4yEdiCOw3VBIvAA+8xxFn/CTUkYf0iwCRBNmDOW
/NTDx+UGnWjWIWJpetuuGM1f6KUZ/Q3/UXJzvfKfpbJcvtTBi/NSvOO5jh9cvsRRqdYXCH9R5xnI
PdmKeEjL4sdXNgbI76f+eIfI7zjrBYSpyommm64xj8KnKjvS4Zu5gTmki/QIQNsCBmOWCB4/+k61
gBJmDanAouEGgHx9hBJpvptOU8S4YxM9+W1NbhxmW/96dcj8XMcnS2DAD6ciM9mMLVZOyoi8zb9c
M0GT0nXSP1to6MI0k35nuVxIVXWTdZH4kHI8l8XdwTeRKm1FBNk4FNA/+n6PoJZCaP+Qa5+1UK81
8d5LKYfrH70q/ilPqOFKxYhX4Eb+1mgmoBicuPtrciFHeGgq+tdX0PKppeNnjxzwbEAazDes/wYi
5ccyAPNJKIQxJ+6nNOdRQF63N0etLJhDuHknQCIre+WY1TZmAUXegY6GLghpRzfHbFGaS6ldbg+F
2aR2H8Q7nLJPy0BUFY+5f2SGMNnnBBdCmcISD+bnimGpI/oBr7Hs06tzOXJXlJltgryfiCPmVre6
LI7xyv3MrwcM66N/jLuhcPpgYqQqUsUqXgod1To+az0zpiaKVYpGGqniPF/CzL5DNopvDy3THBm1
we0mfKU9M0q1sy+n9Y1flqNARocWVQaBJGBrDJrJ7l4mYjF5Q5qExzJyaH07BiDH6pwwtWPk88ht
3v1LETpY94mBbeSqp+IOTPydpEqGkKM1gRrKmvZCOdmQZYyOoMWb7DybFllqROlqFxQUehCYazxK
gyDXNKeJ9YbxzROCfdRrBjeeovDLGgNiENTZlrLErUfxkgX8A7uewD6UB4rQQQss4Y5a8WP+ImfW
rH+M97BbToxua9nCsddIKeEz4KenYT7VaJqptYyZog+gcFdkW3CnLY+raJPdm0Q+/hrY+pptBnKj
Yk6rRybPtNR1zGfB35d0l++ZBHBipAwZ1Mv5wAOAGQbK7Tf5QnBUZuAkiYsafMGeN4OInFMCimsk
uM37+KlxP2f8n4hhR/2zoTHtW1H0623SG44JEvVkwtrJ+6KiWJNJigs4Zquoxz2mpKvTMDPrpexS
M4EytiA0KoaqOJPFpMlQt5WpzQr52GqLRrAuQzF2G8KR1cnNigydKkE5IBCX81d08hLj/179p0lr
PqexfuQm6F+2fy9CkPzWPI20TU7KrJo8LFMlzp+JQ41d8MQSAZT6ZAFgdkNG2UlBPpfCPbPzGzMU
gCILttn5XNDYPT18ggdULT1/78OJRjW3UL3GZB6XRGV7dYs1U4WcRiBF0749sLKfe7j2V1mWquv2
VUaeeCXu70rPRbPK8gwwjxHrJPNrFI4qpaVuCNC/n+gQzxm2gRj8+xPBMaCRznh5a0qZ2A3iPHgt
JX1tvsNXiORNldlI4R7r6KoQXQZtORLtPmcxk+mhKzgq7Z17AWxj2nBsZpHTfKAAfnwb0T1fBkFo
wDubpVHIewFHtKByy6kZMKOuvfhhaoIHGuDtSxQYrK2QW2llA+rcbQkMRI2K7tWaSrohbM5zI4aJ
Y1pXV7v2i4sxq3lUzkaytM+OtE+v+GKzbE6TtizmM3x0VKHh0oUHjUHbkMhmGpQO8krPYHYjK2wT
+wBIRdPXbwJ1DRV1GNzgnB5kzf+TRNYNjZgRB1xW/MrEEdHqak/tdLVaEAa1NpF8zDDZtJb+HFKU
uF4PlUy4DvW17hbPP9/n19qBgVQ/aa7/Xfw1V+qyLwGxhH9E82cIttwEYnoEijFufp1cBbKWjlDh
YwuGNFzSDTSQ7qChb5saIl6jQC/y4ZBiwEhrUOR6vhB0SNU/GNezB8qXno+GkVHs/WAYknNRt4Of
m6ffBXfVAwZ5/yxqPPlW9DjJhf3yCjmjqPk8JmjAm4wcUuczuJojzlZ8dAYI1yNz+nV+AV3bmtcj
ESJCXNIsejfYNb1b3b4d/Rmj6Mu7BI5WAtK/FFsCUKai3Y18uOx5BeGvHaYve/3ypeI/+gNv8IYq
2QvI71YOd2JPbx9yjZ/Fbz6uk5uFqnq/NHl4k9GOJNiU06i/IKRAUp1Hy4DwngqBSvMD0Q/rlOnn
pZTfuFQi90PrTbw/ZSxEjZphEEPAjVUsQy2qJfZj1m81BfaknPKHqqN2/32KLb8/nL9Byskhhs70
twQt9N/2Xp/6T2xwenLQ4NS30pphZT4q1K5mZ27xwIBJryXiy/U/tsH4JSdWrAWQrGwZxctZ6ewh
pNHVdwW1YXrcgaOlVsn8biEAVWYx2eE/S110tmRXuBL2RHUJfDlQGUKEl7OGwigUm/hHlYI3tsWf
GtFnxU+0IcLE9R64AClxa9AjuIFNjzryk63R2awMdSqx28AFDp7d+5Xc0zcgt6OHgS/NV1SjMV5b
Froa9NDcDrqwDBfDvQOeieiJJFpLpjyS9zlUTmZrrfBySKJEk8//7XwZzx4E6JsecebxTcgaTxvK
/nZXwlJQXTwXTmaq2of9Pc+bu+cZut+avvYEE6SKEY7LoYC3/BCjouxNJoog+3b/GBbs5jWjWqYg
Usix7o80+H8DTdMFpYOlZOZrtwnPzH+FUOX5tMgjZ8VfEN57wpDkKRadsBV5P0gpXpiPACnkx+8i
PHGUpJ/wmv6hyNRJEZSZebhfFyU5lXtAi55myhI6fWLrdJ0aYUcaalHwNgkdyFm9zcOXPlOLyaxz
0zFttJA+8EtD43PyF0UU2ns649nEGAr94Mm2ATBtL3zsOQiuh+fk/kXcPzUo6wi7sb6MOcEJvW4a
+yYWxv9iYEEw+9NolwCo7zMwnJbR9FiuvOoRPRsLrmn4+8wW/BbJ1wC4yviPxFaePpcMrHlos3ik
dlo4WxgRzz2N+Rk8afcvdDyOVFJbpUOSRGrkCX03VqVvmncxNtCdNv0mViV0fuFHBOFKDmoMMQ/A
zPahGPhg1K/wxnKVjYYikZYsOHUpmgR+9I55hl2YV3uI1k28enMmwONTcMzASy7hqjj2dzbF0TSg
xH5VLVWdarnDGgZ39VY2YjPueDGDhnWl+r2HSfQT9BLkIFIW/vAXtcUCT7wf388o+pKgYC+NvGoB
KdDcLsQs9YImQVwSARkdVhmmS+RCTKp3qk/ZSOfViRBKD+qUTYCRpyR8KsyNnuUzG9jKOf1V96pW
/CzIHdTndEJnWHjUfUkXNYUoufzWHGqK1ZBqJupnYbLiiFTO7OQH/l33xN4uZTSZClxJ5rNPUY+p
Pwqvw+rOq2X8Lgxq6+ATBKHvt05sg2qkrMojnHlqS7jTazcHSSnH2JSY/wfLzRtzgsHPwpwW0WM8
N7QhWvJG9AvI4brWUxbLZGEHJsOqs+5uRdRMCnsyE8IatnpxuNgiCCXjpCX3rnYBTrcQMwCLddQt
WgWQR1oaI/oxC0TErpaM01MYl3Z3VOAhGCLhrJRcI3Xi+Dln2L/54rnZfsOmSPhqZEhdG4wd7RE+
TKfxjbA8xjXtA0PPfsys4xn7c2GcKQMZXrEGTIbbaRrhKQtnHzl3k4VNKvvsCQgrI98bFobyDT1V
9y8N3JadO50FshhFkxJgWElLe188J9yqyjuPEsghKjMF2ULiCyl0JnCxmydNAp8hzQ40bxbYGwEp
jxBX3ewV2rTuUe0BlXeQ1BmPocDemTFdzelGZvOnxSiV+vaFSSDM9zR6n6cwetC2gx2HDQOQzW+l
m1zg9IcktdL9hhdAPXfQDuHsN1CuKmaEJFMNziFMVvsbsRZDT3BSq4yEOTE3T2hGKw6YU9XNnU5r
5bXIBvrO4TaDor+h3uwq1qcQTyi7Rl4IHlNZNfN8Ko3HlBlQeDR+IrvRmsiEpNTwzTt+L148M8GL
VBKpMTH4VyMdf+2eJSN17GRsyO1Dz28AP4vrmy0ntHQTbvbt2hx1uf+YArfq95zWUMliVszrVVgu
ARBS7wCGPxmG8glaIXwV+A/3KAjH3SV/w5AkNFhYn3rcS7SNduOiwgYqO+Xb1/NSS62jG1CEN9zf
ZV7aAxYqaNeWL/vVczsGaegdWujTuOnNg39pmue9zufoXnwrePMraG3NeYkBpzVmPcXBL2N9Tr0p
04C51yEFh1Bo3TOuOfY/ZNOsEOpa4lu2qzZLDD2JpYUdhUup6Hs64K4THPWXmJisZZ4ixQ6KnoNu
ZeerwFCIURehvh8gLgtU7L96nuzCBbB71lxJgfH1lcdCqu5kkkPYCZtSH4EAgv1YGoyebtafnLbU
wmME+8QH7u3NMP8FPTD3J6SxhaC1pP/xjajbn625M+qbGfLNf+Pru0Bq+vV4eCjLc5vb9N0Toeng
OE4ZCaXg7jQ0KmqKGTiy+ffl9TeU9B357+ewL53PovEPxiFxnE05gsHSe5YWegBrkQ/lBnBu/CCJ
Y3mru6lbG9aPDkceA7f+ZNaFmWOT0ov5kx9ABNihMizO6a2VxLmQKc2G5p11JsLbYSojZuGg+E89
gpjsgh1UUzuiG3gqEp6lW4Gs6QjdstO9qo9f1GW/fBKG1zhUz7mcwOvWf28DpWpWC+CFxyBXaWp5
GjjVIxgoza+//IqHi2jyllY6Zu+3vmRWmRUBvIeqvrrKbVs9mg77YaE/NZHrHAXGr6meLnfDeAls
2xuf9Y+tp82sApUpohMpvp+eiefBOH252EsdzMlgq0QIAEy9jN+vYKa+AFE9t1anu5GkArnf9unZ
9CtGl5t59F9ODhHggWRm8zikgSp0MWuvOvQbQ05iDk8HhwDGpsB6IGR7JV+q55a7HpMlZdn6VJDi
lCg9RNH9l+FdUfaeuBnH8ZLBbYdlE8xRTlyWNXpUzpPIPPRrD2by7zwGHB1cauhS7AvLTqho93Sr
dlx2NY+SyclomxJNsiIr2BRsa+Cz7X5jH9sL21ZpHq8sq6YULhCuY7WwX47OlCw81Zt2RMcqZ35T
cqtE4bz5wT7qq387+jg8qAfLS3a+RxH4DZjakVMaFbFJZd7sCzTuczeG43xm6aWirULoxyxUx26w
cRK1t1gsMLhT/B56Q5DtbsiJWj0ukfHxu/0UxXJNhTW4TaHviO/2vpomCRCPS15uznEyGqSF0jB0
6xD5h2m0EnamI36mI7z8Af25/rAJAgtJ2yncpVPEUYzSwojrkcHbYUSly/n3tN8jkfNsSmuWZuE8
Hm7B6zZjaYEWy1jRB2EQ9JUxib9IrBVH2S9nTw1wcLT9YLOk9Qio58G/Vbn15GstELipsUE4q97Z
z7S7zAA39vgC6gAixTQQL0fxIHV1fUqD4fkvj7O+c7mtMi6y9WwCKqBtS5k2ncS1v7HtoLnroP5p
P+vMdDlxWpo6GHJwYdL+sbkow3ktIr239liECngnFfI8JXzP1e+LvscDG0wqV7DvIwr+0+mlPEIg
1CgVv43HClxzD4cnUJgvZ+NnFc+czYwXvZjqcadGi+7izoMTlbpyzbL4BXoN/o1/8/24INcDNHvC
AHkwgasjvIQgaPS+cF4uIT4aw/HAL3aYVrcbShz6JoU+zJJNRiF98XR6R3iiHRl6Cr6Pv6aW4YyO
PBaTTGbGS2/BECHRTTjGHT8NsYjeF1sChH8h+YRHH4fMxyBLECPw5ExGI7Vusss40QfoDczcU2Tn
+5aeko89yVzt+834t5PS967RQZsWJIvhjvYyFJUMfYeGQqIAUtmdAJD7o95XZvMkCWaKSUiJlczb
qOA0rZo/IcHEtUklvIeTyYAzdroneBxpf4tlguL/9fZnXmLonztUJCODr7f42BWNAlqt0gPivl8d
c8LdjbGlHxyvik6xFArQ055XTMVKfLCADcvNxAfs7LsOJX5FSH2MBDuxq9kC6Mcu14LduAhiQEx0
x66LuUxZCHydzqZbJ3REq+RxGXjeYgDg3Wuhr37oicAqArcIAeWk5VGQdsMhRz8Y7VTDlbMWFIgl
GAX7WALfwn3lvUFnTio6jVL3ERIlMJG4W4LIjrJPEe1iC5/X9n4lJW9CavVFFjZhoQTvMTpY3vhf
K7DWW2NJqSoV/xSLukGoFFRQJk6FQg9m9ppa2s7Po+7mKe2/iKV/UmuR0es24nOfLqX5SRrKLQnr
R6WDC1Aa7haHu/fgi6yM+pxlfV8vM8z/OGuLUw/CydoRv9coE10/uhsl7tRCR4L9MnRT2jNrIfJP
EtF+VOdM4Zrz81UUltdhIpfEpAeEf4Y1r2AmBJQH8D2cmdvipoRrBR1boHrZhuhxxvtmoz9OFOim
amyW6GqUV0cfHp6b/ksCyDv3e2Oru9H6mk8YpZqjkMj2O1VikiqK3ZhpDqLo+NyefvaUmh89d7hV
pJArXOmWXOQqxpD3w7m7ukr1sogVTSaHpYXnE5nwRxe3Ve0i2SjDbAbmpVTo+TlD2F44sOud4XYP
l+2GGvfy+tC2ws8hVMcNFQ/l/M0NM25siWZ/Owjs53GEwpMekPEuG0JqJs06bmFiJp2Du7bz9n47
lOUClw8rZFS/ejX1Oe5M8M0dDAqrKM2zzUgF+FifRcfJ1NADd4RgiGwU8KJFpnM1rFnobNPa/2ll
HLN1pJ1aeQrWNcI8c0HjGP4wPa0YmgzDPC7CAwPhCjaWmJ3BHMqPLFvUBTkNQRg+llOG7Smb4ZKH
Ohym8HvGxZbrgLMy0Si/Je0TJ/W8IM/fnsT8YOoDhRCa+Zc0Em/iFVxHcFg4ULWYLwHb2L3wb1Qv
YC73M5ux48DyO3PHNehRHP4SWDm9gEhdoW5qr9cME32YEHtINb3I91C+VAjESq4hmsM9WanQvOAu
eAri7WrfG4pWYdxzyyPT+tEZSKfUESn8F6xTnNoy7SDNs1YGiJcPAeQXcTAG7pucrbJnOJW8ZUIn
EypixG6KJYopAnrmhYynpkQ7IGUOEGmjFFX+B+3ss/nid3LC52BCqa4tP97jsDfNXLwnlCWvan5y
npxH3ZgHY7AzbqGkNx8XdIzA+gVrKBr/4TSzdSrt+0u7qmc1xKCCJofpJRU3Rf6asRnto/vzcPm0
vwQpXuTkMx9xdgO5n1z0794NYe2sdGPmNTMmpXQE7309RVts/xhDwGObzuk1tv7Y5gh6Uzft/2dc
hqE4OLMeEbe8Cd879CJD1/5gZZePHEWnYxGOoNX57atzwxFYf1ZJRjSLahBfgVEIsFng4ElupOrb
3YthJ1Tf0G+TyC5CGtmgA556EE7j0lENDZUFQ3nayxgoTQYTE2VatBewP0DKWq+ApR/dyrbGawv5
rWXjBqMP3IwMM2bSwRaMVQntFz5FoQHtf1SCOVB/HQCPAENaZ0w8mkLdtVm/7oh6vKFiqrH4SIce
bgGvQFXlET3tFsuQbj+45Vr1jdHI/ADoAuwzcpsxxU0lu1wfx8JbEY6UktDAUZSgw+r4hyg1jwVF
dEaw4gqnpq1WYI0G+uHGfBZ8ykAWBWF2YU66VDiqorONx6wfn2TYqIfBCBQsnJC5LJVTGHswkQIF
TTAHCDLgZcMoSed0moJ5pDlf+3cMrSSc9NeLDFnKzXKPqN/Gy4HNLNqR5EAlGeVbj2OTys0/8Hm3
NRnOPqRGMREZFNu1LWoPnAO6yp3T1bCdU8LDj9j+x8zJxC7tgtvupjnjHcZxOekfs3uykhN26Zw9
82fPGMryUG6d5+of5N0vAiZWetazUJupS89kYYohNZ6b43cqu7OuuAKqXuOMk2ndLCxa3+on47Gn
qd7IhdUSgnH1CjKP6s+1YMC0Un//NEyAa2GWM0hr3mQVFg7sAwU/kemyCoAW57ItU3H/SobpqXa+
QAhedDrV/mlua0vTpi+p1caVfWpRO9uwmhvixkH8Q/bD22LJ2qvM/Z3QRH324SAleRD5NYHzZXTp
scHgdehp+dG40jTtw/ZhMPDzGiNEUqs7msWDsavN78/LO4nG7bGatCRVNfBC+DTxihWzmkF/5Mde
q0+scTK6t6UpVr9xmvZt8XNTWrGYuMlAeU0kpNpELZ10aCkBO5+D/LmDUvVCPlCj42dilDtcOnjj
aRDUsscaf95Yq/n0NkPZJJvFkK+mdq7QpSu0mYwElB5R8MXAtfyy3ZqyJkMNfOM/FGfzSa9zS1ji
hCGXvQnLx731ON0duGvL3bfhOGs3B9/1vHI+Vbx7R7dPcQl5sg02HzuqgPEV5h1ift4lVMwZeNAa
GDwMVou8LVS2sMAqJb4VI+NujrhJJDAIhcLyoaMlrKDGH2YSIZ7SYbgfSAirIKNsFWgdw3Dr3RSB
fu8uJFWNQj0x/sdvWRus8NzaUiQBzkMnboTPFyYlkrKBCep4dhFWYeQ38F/Wc2q4SmoccmYvrKeL
RPoGXisma9fA+z9eBT+J1zrErDRj7zbZI6+RI1nNqB5lKUYpdC6af+KrgBes2kPq4lSolmvOBoox
3t+zcTBkNk6dPyO3TGdGPNGue4qhaVTONXFRjLMO7E8ykORAAdl2V8IObAxlEP7kD3jatCduVYS5
i7q1+kUIzlOlarucjrqeVTym/L+MrnCKylEoM1O5KKBoSiUO91sGHE9Qv/SUOrj/YnIAW7aPNPbn
W3oXKql7Fks7EDBreEJQZ4feKdAUK3KfJRucUxmZoqPvJsIAelYMgrpJkTYLRqwAwKyb6HR8r1WN
U0278x2Vru6ldQQq/Tt1Y/0dzEa6rc2dVVjaHcSJfs40hi7QKiWMWAXNjTRgbwV2vy6H4cv421v3
bLEnxkhG5RVhRXffGkTc0ND5P2vpGbu1GTib/UXMmLz085BSo4UBaJ5VP0MvhEyWNj0wpQp+0U6L
6YZeCbHVdnUsPxN/cxOKxBiNlzcgT6015owstJMVZ8KXzTSDXfwblx03v3Knx/ne4FQ2sHFdEHpT
J5Hs9jIp1fe2GM8RuGa8MpFB/mqX3bN21Dg1mkYaSLOaT0e63iwUfH43NB31AEF44w63aNmbVDis
hdKbPC8+Yjd7/rfVAEA0hAU0D3NkhQB3B/0VQXNoauaJQ6X+g7jp7JZWJC9A6Vby82ixbDgUiuIf
jrMF5lhXscekfdCkfmzcLSD2qWQ9Ubj2ckV0oOIDaVbry/ZCQBsP1X9E5lEqRVt6PfKUwi5lETpk
MGL2sn7S/PyJpI1nIzzI1qNCr564Waqtjw0zvhujAAoWmSZsHSbrX3UFmOmv181CbjYj6r8H7V71
TmPOTUNCHpZSdyGDU3Ai5KkXfSYpQpes3RqakBZDWP8UvlCy3SCMPjjWo3JsY7YbmXT2dLhuwM8s
bn5FcL3q6DoqoZ1uQsPZPmFioiQ/2o1Ef88pRWUdr+e1AFQHmgH82PnLkvcBBdU8ieZrBtXdH6sB
zXOM4DhBQt3M/toA/7prbjCEputPvvJyXvbhcEF5ygDkX1RcMpziv8rWUC3wfXm4Td6/jB6jr/J4
roPFQk0NonVJ8fqcyr8VzXAV2Pve+561Th02FdCrU0ZMxGJqXMncRT95H+x5mkxAzzPC5zznOhSX
ufjIGhd74ztMnqxG0aKuAdocjBjnEzB/U7oKOL19RWCMtxu4JjsHctC103cXQrvmcq0JHVYscpjw
jrN/CKJPHpSJmcKSHY3KUCr/3jNoTCMVRiwvhS79QsT8F9MquCYdGL78BqLlRZpTtN/Nq5QMcjIq
zWO/yL9/aFXzV+8l5Bo2vz9p5sdHgcNO6zu32C5tKXWbgtflpRajx2cCK5ka2WTfkSP8FJ5OTgGx
VUxsBRpyjARZlffUH5E9UYbU6QdUG/c6YvolEKXLWhTGIH7327kkYXr0Std+v7+bC2sP16FXoOHW
3HmsNQWt297AFIW/kSinYlUnMd3srP738unh2nx/qg/8+lzQxB/JMDiPNn/GYdXGSQrXZAwUvwJA
HTZrvX0wtqEMi8QzS7s1I5jefezrWs6xkvipNzH0hkQkfq3RQfl1Xs5L9KlOz8KtV90O94RM4WHJ
aIjOP/qtV62QufzgIkrCymzKy3zxErpHSxjD4NMoCHxzhc5BHiJKa1TCG9zjPg+Iq44Zo2mHCX/v
Nmjb+5LUpZXXS8+eibLBHfB4vFsGHxpruPp8mkMRdfW5h2A6qdyi1rKpfPf9YeQRlp+OHWnFb5mj
SF4SlJl+9a08XyD9uCsyxSLPPHQFCorsNmkUDkfcG6h+jFgnbjtjRMKIip50CKGXF9mK+oHYU1yq
UUhZ+B8PxwK2nQZT6Pb2K7HTjQ9k4BH3uitO84NiC+s6DAc1ZuSnFhDVpkjMJNKblotI3K542haL
1ZeIMalDUrs7SZ95OouJjv1Z+fnODuBVW49FvXxfsMN+6ivnzgZjmlsRw+38Dh7DfxveXkH2Hajz
Mtla4D87N6Zd2LRevfiETkviSfmp+I9RY8sLezDoEoulUj5v/TzOSq2/+j3VHAXtBFwM3Wp73iU+
LCN5vbwL9vemEwBCC3Zza4Kylhbzf69TQ0PJOVeTW//Ib7Acnh3he6t7HJ7IsiWgrlhfHHW4AHLc
6ItcYo1UTR2MvDgqq3Cwj0EgoNrtrxZXrwCH7zviJpHX3O/bBruUNKF9iU5b3ZEf12eYZycJoScG
a+QjKZfDCx9vLAcrcTr95rd0MeqwRJ+STh6DHTgYSDn5u1nNWpHrjGp+lC/uSyB2+L5SgraM209A
5u7QqMOvzDII3WeNtmLUPEmulQRZs2PoEO1GEA2JTqIsHSPXJbJLBpSu/8UPMkwoiLnBAC8RApN3
jD9e7uq0njc4dntdWjyRoNrmpNeE1PmAPRgRejVHZ5VCmv5JSJUproZ1t/uvXMC0AiZ1rAnb9OFP
kG4ah7iXK82j1gaeHho9ylMGrOaYKecvkMJ6kSxOVO8GUJFJzyRX6BMBrdC8iLYlHE27hUUta31i
2Kbff690DRDhAb2jdYkVhfDGiMrPQ1VQ+P2emYsUp47l3FsvFmoPdshmz8l1L9D/BccKBCvPFzHN
/qPGV9CR5zjnZNwhuNqyGz1w9uWtKYqt15fTqH3JwLPE9OPPyNbqtjV6l36FTqgvFLKrrmNA2VeJ
1RXOvQD2qyo1PpH0n+jAzsi0Rt51yxejiPAN1wpczwUqXQcOfYMo1RwMDhTm8UlOakGVdA9Au9ai
+10MPocNb6qQnjkRVHm5RDVyzOahPttUF75OxLPU+s/wPUVoliJ2+oK2b9l77QlRk3Ng1Sj9qGwz
+pr9aT9QiONq2F23JDfpE55jBoJrH81D9mQ1BqUQqc/7NeJl9ZNQDAtXfPXQswOyweerSmkAvPMp
8fY7kY+SThw/9ghRx1lBaTvx1yd+WNn/+srbBf1WG0zK4dILy4jz4BuHUw963pbC1PhIQGwLLu0j
iyHrXRn54KtJjfPxxJyaalQA4yNorOM+/xFJw6DeMCGo2PSbfKMvmKYPelBSBBpxKC2BrpUiFAdX
Qk884IBFT+56sdtRSzb01WpDwwzsfwQ+kk9WGYJnG41BlC/PiQkd3iJi5LXufo44HPddytBmCR05
z4Qg1tLzFsMBkMewysjip2W6i3UjSlR/PD0Pe4kNpBWHuplp/7cL9TDRu2KuJ1qB4px3fjrrxqSl
mXQwmT30Wds8svB4yIa2NFSwg4hxe7hPQWK1HgHVeLLLior0sFnGVytaPS8qyFuIcSWb10YE2Tsk
9QggHFHGCyOJhFVy1ALbfZ42M69dJ9Q5Oad1BP2hpKqXtLLuTaJu/Q22m7gfSpmv6dRP/9ndYFWV
SKQRH2OOV0ZHdOq5H9ZfohikZjKNn67yOC46wiKW126Oxk9NFc8XMccfbuBw1bM3yTK/cjimLRo3
zJWwEz12bVPzqtu68jYjegqRRz/2ZYciFPFCu6iUGiUDkDM1K3RasjlSlJbaBFqy5hR6ZomgepPR
ru/A8cPnY4tga6pGLOWaOxLiy3QsD0972TOp3rM5fGqAXrpUPzz7RbsSyeYDv6fPAd7UGP4D9pCO
4u9I3v2AYR9PMAzBgfyPi3OVU3ha/tOcNE5/IkWpb5V8AQHBbgGKYKQDCVkutNXbywybaICS+ArA
XYLSZpEUcB+dw0QOafQXlnrheg0L6S7+FcRmPVfhcpXs/349jx4sPVCoD4xhLAEK56LRFRM1z6t/
0wpih2Cid/20fIIjziNhCrjmd9UX51ugBAW+4AIqXUo84B/gL//m8Vqj4+cfoCSizaHBxkn871Wv
crXAE5ocSyMCALuNP7vqNO9N4+BSIQnV1D6euazM8pMd+QGza76WPBs3RLvssx77acS3rwLZfVEm
R1ZZYj87FReD2bt+JLLKarA/7jmJyOVK5mZegJ/1mUmwwMMVjfsD6zZeF2Zs5Xg7/3nOSnsKj4Dr
2N+aTT8sUnRaFMr8mJzzsvGNhfCaWgJT9p4hD/uh0RsWu8+zfHF2gEbY8cAR6E/5VEx+14KC3Ztc
KlU/e0PNmWazu16RmpyUt5lca7ihWzL/M0NgwAqWzJpTcgLUSkUhPYI+YG64jGwG9ES48aJUPZ4A
9cMC0voGLEcupI8vDCYqZ5efDNO2Y/BomxlNhfBfEvr2XyT25gr/plk9eNm+kbyTX8YerJX7xaQO
63mM+eWURn4pV7y/GdaymKGl/oKimn3raqNBObjWDgPsEWvkIT/tGETnxTI9XTpn9gpsLOUav0/a
Yrsq8oVXDrrPsh5flCmHnI0XfnHOoGC3omzh8IZF8Yulf95jdWN7HynpPBjJzOp7oloM41du1zm5
OoXuURsNn5YdSJfLaRcUVaHFrljBSsyojaJHGxv8MqlgnQbbN48EiuQ7acPpN6wLExSFR60nWgM2
YQU5NwfXmE7LNOkodJemf6qM88zkCm9AtL/HG0beOqOldqgLkYIQtGhBK//ioexMRjiRlGG+ewkD
qUHIIq0VQpb52/r8u+LYIoZshNmPitIUws64OfYPA41h+sc2s8lBrAXHcLnacSLDh6vWjSFc1ivP
IDAdJTuNQh7CI0vqSK1kP196S1cD2A/YiSIPeeZCLAKfTRGv/qxxZc6gxGWMYy75whxelHPsbj6h
eUxxF9ahr+K1dvigrj/hENoLKZT8FyxgcaYqLO51oJu0TcUPqugxsYpqNSW/TSdxM4PlwCltQKae
5lE3iIBNvpCI7cCkrkNp8eGCEbJxl6skXiY/7OROgYOOy2ZUNHmtbjF6PeacSfa2b6DbfPKYoDHy
zw5uVqa5UYONRDeyaE747kYn2Doof1u2AoUStsVYEEOkqTw5Q4LSlq4ERjvja9IuTxwKh59+qd31
SFDlNrkOVu6gBInn1S7vJXIg1Z+PX36dS+3/8R5hHQZTYyeHGU8S27/n0At2XZT/OhG3/cITiAnj
JKjLP0y+lWyYbYB+gZZZXzw9vpq5ugf2m005lBKoQD+fuHm47IuLpR8S0UZK5OfcZ5DKFtmNEo6c
NbgoMbaajCP/sgE2jVo47+67BtN7s422gYBjVwvE6nPMHxYvjrCDzuBSR6dWHKLOddE7/vb3wwur
x3i3fXAlOSriVyvf2rdFeAVxKpJ/bmF0MkvTRYgenVO/DVKDpinytQ1NpW+2NAjqs8GgWcsLPdIj
j7Lp2B7X7fhFtKgwk6hddtfXf3ahpG+HL6bZ66o8iAWZYjHiNOBX+NcGf5amm5fI/TnEk9U+QbHg
yV77piL8w1RTpRA6tbq4gvq8QOfLWdf7wkHTOLdf+FzmOV9flzczAx1Lp6iTrnHijAuT0o8YaC34
TbAOyHWkrTNEecO8fszIyeg3EOTB2+Ie9+K6bV9FdySDmno+EElqWoiuM9sXirvBbvLUw1qKUbvN
tZfBhv623cWbjCfKjdCKsk64DzAg3Q+v/tWS96LuUPnZR79hlzMs27rYXpXf9DsrXZdfYSXvraeZ
3V8k+hXOatRD2v+mVPhpsLhJ4sck+WENrTQzBTKWgivULk/oHX1+6vvmKxITi655bCAoNK517yal
nwU8wt0zlvfWBXSeoamFB4jgPjMYsR3Dt3rO+z9Tai09hDB92yuAZFk1LAqP78yqwn+ntIes9Ul0
sutFNn4JCJFrxKAqYJGOuO2vg76s4+O4omsYK2XP34HaMeS27xDr9SQPyFEvGnk/yjJC9SclpWfc
m5x61y3a2y7WcOnJrOZ8eVyeNLVtH9gI/CdszjO+O8TiOrN/PRu2Mh/BpYAZtuahWpE1wgvUPpbj
MrU9gypWXH3lCB815yi+nCDr15ABdtf5ALK65Uh/6+8DO4ZVKnnxUcFVLFJik3OPvcLZvnNiX0V9
C41U9PBQmzopDgDULkjzW3UpRTHqxNUiyUwnpcWhE3TnLhlKmP5RuqKabE5RNdosucuC8fraNzQM
Y7om9yfjfqgd4wxz3NquHVWEfbE6YijH6YN0Bq1907lL7wgCYNCltgiZRKQe0a7TSvCzv6mhKEuW
xbjKg9XMMYurUdceoMj4ABkBHlJIdsyDH4WqDctSDUpcOWNAsd4bpCtXGLTTb6/cnLLJTUbz1pI2
dN58Lc7+z7GtoZ0jn1Nq/wOoyuA85BLxn6KfCU6h1foIYS+mDmLx48+ra9Eo0dK909u9rDMVfDI9
USTX9mxgXzfj+03pvoebr+oi2Vi3WX8RDg3iez7RNG9qh0kJeAquE8vQN71DTneFhj1tdFlM/Gmy
eG+Z9bhL0AFbFxfaSJB0onKMOi6OML7Pw7U9oMpY5YR9tsYamj+nlMrANR5b6/cmZUS/tXlGbftd
1rGa3Cpm9AxkmvG4PVBn0+iQIH6aFTfXOSQm7U9//xwUBzRSmCz+CKSZMayuT2tK/Lyiuu63ZWpP
dEfn+Ddb/qvLKvf7NyzKejqGhlxQ1didaHxYtHmwBPcZPVqYMG7rwTUY5QbcIIqQ+dLi+/PQ12QI
73sXhCgqroJO42Y/7HNAopij85/eSCfWGRWoarc5oeLEMBQoIxXJQ/o649Wywu+1LfN1ktJcCUxx
k+2jyfqYwt30JlTo+qAFciIfMmnAHhS8lXnaCnRLsEtdVUILWbdr/14ctqFiSm629vFYG61DBRle
TAmhKdC4ZmmG3vOeO+DMhAaLlCA8yJZrxMb+gGDuj1iXqWV++pNxJqkgmRSVNs9sCC1jxvjtF/Wa
SmbCTiOaj2Hfjw9SMi0H1ag6GIcJW6cEjyHnbjANSE1JPssfB0XP6uwmECHTITUqULOH66BQhWWV
RDPHIhNL5ttFmr/q5nguI9EPpIHP0KMaU5mKSoZ7Na3ZsYA4WXqMnctM7JKu2VOA7yHjEPkune2p
1NuP11jABIdh2uQ5+OQUzNqHxL2O6TTP64KjKHN7dgnKo4akZBLVU9T0cni4rx77lo0xfD16oW2N
4MY870W56q99x32dgBNnOAHTP/cWEgSlEwvQBTqaSqb6+q5xqXI5S+VGf33WjzKbrndI3HsPl+wK
GcSxelQbTTHhVUvlXXZwtHcyyIkGERgxa27KcKsSJZzAbkp+RQaq4z3qq1CAfKVdII3sSH1Bv8U3
TiM7gWKBig7yd4HYUwQmxDWD8kQuWnqPpFcX0T8skB5GZpyS/q0wPHkU3B5Y8dESr2GbmYh3Unqq
mn4FZe5lLfPVdwX1dR8m2C3l/h6s0+ypGOqyFeJIJSrkwP1n0wUlBDlmR3T16XQ+P+0GXlb9wfi4
tGbKzacLrgvm/cnG4ePkYSauiB0Z0HPybIe5LlYDt+lNMbrDQRI5Vw/cj+UWAGC3AmkYdtIOi/0c
GyrAjJs3+chXUu05P5rZVTegjhoQs+1NyBz1V7MVIcAmLWAlALUMnOPpIWZ8vvcWygIUka5WpkXU
XU9G5W1WWAk2w6ncXW+Dma+Df8r0cJ62eH5KbzJ5BP6yQDqQf/93usU0CDvucQVuAN6fkhOSlwmF
3qCG/iBPNNBxGlOJ3ABYCb9EpbnAVON+VjFutgiObXTpg+/AAoDIK4Wbrx7xj0hgUdb0tbyVGrRl
LW+ovbmCJojxpmsRvVOaUVZqV6RyTszMgUud5oK182IOYLNbu9c5gLhQVvwWfVPsTVCof7WIF33h
PCXP1eiUIdjp1arZ3APuqxh1ZHIZEeERmTOScwMNATLOfRAQr24jKX8aFa/h/aGz5YzN//EjEgZm
G75kTJ91TjdxyeaRXRpd/DDBYYmNPtpmaFF5fKEPNd3tNFmOaF2R67A+xREUG5F6BHXMZ+pVHZwn
BJWtdfDFEafUjYSZUgep65Qqh6y0V8P7g9UpfTMDtBE2C10yG6QJaoK07sb2ByvSUEKsMdNMah0P
SFRwx1uOcOC8zvt0JShmodAJqnK8BtX2+nDf4Cu4G0RPzpqZv1WDDhcJQPcAIIGlbTy+KwOH2kJf
TK1gU2Me40bWy6Mlq5H0RTAHp5X0aVwt+StzVEf3alP30WoiXUixsRomw/I1zgWxtF8FlhOyz+I1
p+vR39UyP/gqKZgqZKaNbnNodvPkWVh0X34SPGZl7zjx4/R2W5D2jgRkMEXvdF7z2iPjTZZ6hhqS
+k+nWX3VaJTlIfXjUHUrMqqtWo3m9xfFeLWWJtNtxO/en4IPi/SV6Xdon8Ukm/e7xtCbdFztkv3+
B6VFTZdA4HV9pURfIrfT7exQ0KO76dcnq2aJ930mRFK91SJv1j4Cye4cIjMuFsVF6xang7K2DmgS
iUVeKpZ6JPfoBjnsbIu90Ur9rTxvArDvxkPuNAw5YFokhgl+hdtciwiiTeOEXt3ysYWHBjG0e4fO
w06+oEfHrawGWR4meZcMhUsbbmxgkowTaj5CqDltt2zn9U/oybLAPr24CX7+T+3Hbau2XBl1tDz0
jySKoKcuT8CpP7FF2MfEt3SxszES4r+9ZrtQby79ep278gSNiNzDHYCI585A1gocmIMmAEQ2hSuI
lHyWYYTYaFXCrOX+I6GLro71NNh6GgzqtlMTllZbkk7URUQUPi6Gi97b2dCejV3r9JoQvD2KKWa/
96gI0ab21S2FXzmjTDffJb1EdeRrFqPdmQ3DQBytOlo6Glx2hYWsp8clmcHx3vVXrdPMvOk8HCN3
HYKz6/6xCOf7cIICV9G1siven2/ThvcWJntayTwtIk3AqFi/PT2ZPwl1WDLYwuTrWuc0N7wDxXDR
ZiUxTaygj38OGiI/GSeNcXsW9nwL6v0QQOdUt/9qO4jvbZhsSo/Cp1NNccCKrBf4X0BAOWXfnhgL
jxgBu3dfhuZhCCtqQFuhdXMUqU7es1SOeLl1KZrgSCYhgagGjn3aC28MAbn8jXVv+rcNkAASe2kV
CD/4T0x8VcYTtE/xmd4t7U16qda16f6c4MsTXNHT2Dv2hKRPFz6abOTTAoebBp5uTpIve4CgyoPb
5XEQDNNSZ6bJQw1cewaR8vNaKtCpsuUdpsLjhaGhHKhnB0B9Wb7rHkv9nG68ymCBIwd2pOwpqCFS
tdzvJpnXDbslodNOAULH5+N2/zDfpyCpm704Ty34Tbnv46P14C92o3AMS1RT0k30XzxktDEwIuCl
Kqmp4HPoT9AJ536cW0uk5GfZwgiyrHmVKZt/uq3+7bHCA6TaCVce990wfUaooBDYUNublfOlF0up
gYL8zshsj3+A0441ttvjo84R7vn0cDCGTA0G/3ZS7R9MOEsAxbCtA68qL46T0bOmTVbsvi9SYd1S
1KW54QSjQMLkcot3lKy6bNeT1ButTr82jAjE89ady3JZXGmaMkQmzc84TX9Hlu240MPOUW2oBKpB
BMqZZoOB5NthY/YNc3RAR6AjhAllKlq+PSL3a+yz/x7VHzc4473BjjMbEwnDjPQe25T3duFL6+JZ
L6o/KOntelgodeyV7d4789BzGeLRfWjaN/O9cQooAurx1TAPZZvRuKJlBB3bggo8DdiZYCvNFCDc
cYJx0/zIpyAmR3GmAHeFdLgY1BpmXqz9Lg0+loQAmrizeB1WdkigyLq6yYyRco/vWxgA+T6Zf54D
PMg6u9WxbpZpRJ0nBjVj6YNB8pZn9z4SWgnXJmU3yv10t8Uk0JssZOGIlfCpoB3T5MD2taYbcx8U
tBl21ry1yl0odfof74+Zv2ZPdIkDg9pF54DmdOhWOmOn4dMqI5y/N57cP4gCB8fHhhvWbGBuKriN
HBdWxDHfk//jtgfjEwcB73VwCmZE4upu1ja05CYqYBElLZnVK2U0/D5P6TLCq4gBEYusGZZREUj0
22BdUyfVE46YZIKQu7gI0bZoj7qMWA6DxG054ETqn1imz9MVNHDH3pdSI2aEDaNILcpsvtI1P1fm
xe6FP48b0p1EJyceW4UE/Y0CTaWgOvGtyajDjhopKtf9xK0al1kIlVSLaufqBPbrOOrYrvWidU1S
bQ7bUsqTzHR9gUTMsA2sPApc5bdGYXiRAsPSzgZMhRXd1WQbPuMa4XAbrTKrJO7Qw+IGLDniam1K
viRWohbJWEdt0fl7+0L/+V9mPikrGKYuAppIjHK5bm3g81FfREMVojAWJkXbFRedc7kv8se/fy3i
wUi9dcHrqnvJgEXYUFJHt3O8RpONdRXw6qb7U9gW5TwiFa7G2KpIFfbfswbku9Sd42j2PM3s9HYm
foTjvFWpOp5IvgvnP4LyAKhNsRYjJWvpEqdNv0VqTfwUA0C4/qi/7QYlrgFnDN1Uq8/N8n4D0VmQ
ppp0+JEKlRSazIAzFBncYyQHs7TLoLSmZ2m1xlSo+pEkKsjaT7GwQ7PSiLdyJUpCp0ZBA0bi+3I6
gTQB3Mg+S9qTHc6VTvK9x5YM0DEE0nLV3DRr2Jb8v5ReTj36GA3uGkoyfTECjfpQpIpnSYfgpQtH
6A56oWq8FWyiAj9tgM/Zvfx7Z+62SQTaMd1U1pdfpREC/tuYQagD9EuDqhTBpZKFQN7PItpROkCz
o3YhcznjBA8dW3gKeracSS6W15gy5cZNdKWlZoUZRlLQUsCPwnZtXL59H2cFv6eZliFUuJJD89GS
LLBRml3Um0EYTU0CBWH8wq3B+YsbGrCPLnph2xgsMr5BYWH3YYYNZsHO7Ct/mNHUIEDqxllzeHQ7
QHb+/PHDLu6WTa/kIVK10gz++0mWC2YFgcKAkyiw0nKEOZY4FLxNjJ5h1vncEUcMBgxns9kELjLP
PWVcN9eIEmPLiDPUprPD2YC4ji3b0AlPvZK38XjEybwSYtbnxwSXMcMOTZOsPqkUxm6dJvjlCRnL
FNBMyljujtp/twugpOubxh3lnGJqQSgmCSnyj4+nXuqMSuYxnjrnsKZRDWgje8x9ga/c+HtDxreR
nXAqxoW/1wzjrw1QX8X9Nor+VqiqubRyDLm4CFaeAGwn5uMwFYkmRZBvmAsMqqq+JFo9ET8Epa5f
s9bfsAMj1d+Zfg5jwnELh9dbotBWVhYFNsuBhGkYSJPKu3+9LxtK24pV/qEyCEHrablxLg2mKgmm
prlsiDVYfj0iRjd1o9OGNKdOPi3gqaA6yo3Auc11FVU3nizQB+fEgqCBy1uoNdiBHbN71SsFmWb0
71TItlTq4zdGhz9zBf3nYrlk4IkX0hTur2Es2H0I+XmFYRu2XfXtwKWIJZL1HBUAgoEgFVkKibXU
YuVgim0v0dH/AmY37AM7HMKxvYwDN6jtm4g5PVkRpyBZb87FMHEF0pGDVpYEyrAZAIzwtbSFPy8l
jwA8+ZYrLvYfRYrYx6WucLHv5blt51/XqtAd/LYW4aNYfTdYaE2Z1ztg43QhAT+QTXrLwzBUS0nV
lsxqCeG+w2AJfPYLZcoPQ2g/LAoSTp7dYMpMISN4KPg4PzMr4ndvARiYOjh2z2FApXaKja0lUW6N
jatOYDdeoDfCYHvVyC52/x+PjQ93T8fON/RV3mJMWXlntccSpPhuXpe2OBfC7th6bqaluIvJudxa
zuHtdQQuBa59BYA0YWr9hk2cb7B98R22yFGufBCImBg/bukjtPwUND2zLhpPzlgm/zwMboZyHarG
RSyuRaxbosAQkLM4VVilLng8mEJ8s/xcKO0jp0LM/r9fwklkKKQLL7nLS0B+sc0lSwREAPJl8SLN
w2QIY/C0bpEfNYivM7vBeFSvszn/dthplF9pw/BUsNFboQbwd4MostsX0r86CMdHNnSq45g/HbCT
Vg93IeMplMTYmtyPc5Yx4V8a59H2/7BUYRvvJHTxq1/td5JGAMXYttVcXkLQDRBHjb9dYdA53zNe
aDsty5D15Jhson3Di1EH7FTMMphrgjb3AaQYkP4Ifb3ZEEFWWq67z7sXHmZGM6H4iJfITM0MW4Xi
2DqdhHLfKb4zuP9wQsPcBWs/4AwVfBNbR5BVQpEeeC1vg/9uQBH596v7suo26qUBSpOuHsIyOpMP
bBU6CIweLTyIEe+h/WLynbU+9b+OeNniZYmMEoaSyBiPUfLaP+m/URRvseZlRTSnAY9NPBrtmOEv
ySvu1wVSiaVmvJecRnQbC2kqTIplGOKqYcj9jNrEMe4R4VqSQIjS6B2QH2n7lCiKpkKqtjlcwHcY
RoVloi0bx8ZPLHVyOpFgVf+PHXarZujQOzpBP4XRi4NoWrKlP3kRcufaVayWUZGBIkA/zshvbgKR
uvcepQjvVBEM88EuK+/D76r+akBh33H9l98IHv2v9nU0Ilf74my6yg0LZrNOQT0BYRspEow22QSA
v8AmFvnBnFnKsn6UhMPD+U4ka3g3Pk0JmqCqoiT0vBl52bEqLdH37reteDgMbo6LOvxmsocA11jq
iEIhBAf1wj+whWGX5I/ACDseDSxkRq5MgwhftMNZUYqans9TkeMbwUZam1OgE1UpK+hL89wlTOsn
wF7+S4YvFAYmWVSm1+mflc5rlPxRBJwQFCXWx92wUETWucjworRbVvmJ4dGIHOetARo7o8xXbQM9
e/qC0EvKlrInF5KwwHxinvEZrc8wKTOIOTUlQ4v8o1sm1kHKjHS0QWQWqluy9CFI6wTPhLITnTma
Le5AYrQ4wfw+Tm8up3foulSQSsEiuf65Fws5cD7uuBYWRdnjy3u5KbXBkz+tT+s+p0+W739DMo2s
bvMBjltTXvrtaPuvhc5N02/2b8KwD730pSXt7YFl0iR6t0CWxbA8SENSn+CW+w6wal7i90fSucpk
ILhO2fG2tCGn+tj9fOB7Usd1xvtLy7PDD+j3VkcVMWhRaX3JcDLY9liQWoJmAfZyWAM7hLpfIUCC
vJy2bnVMgEFRzXh90VOJTj6Lg6ABFm+E9iVhTA1kg9Iq/WoYnniX+N90sqCQBU4RmqDsAAri5o6a
TMAkfLro7o+DecdpwpK6OpnXLyJT9qk6iBNtJXKSfKSHMQsTFyFrfPxc3aQUOj3dBAb9sori/qLU
zujCF2ebcXvn7C93j+Zo7P5TZdSLMEllLjiegGHa8l7rWVG9UMCrTHmikQf4YPp/LLci3cAbRjgG
ECffrJKk+nhxTNdDNT2zwd/MGtc2zKJgyn5v+m/9mWQ1gnntrTQUfOSOCtwsr4M6zioChYAK4JYC
SM6NxnKQ
`pragma protect end_protected
