// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:27 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ul0hM/S8MZsr4pgBYjiMuPHzR5WcVR/c2p/8PtFFYYm8j2iMP5beQekHRffudPrP
h4bZGNjtkLIJSChYpvZ9OQciEEow6iFXdoKugSlYYG4eypGCbcM221DbdeuPn5vA
p6Zf/svCTQAqHn6NMA4AlzQ1NO4G1jnH5oKX08ATAHQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28608)
b4TwpehN2Z23VTMJtI5qvIotS4+LeDCMVv5n8Zx5FuHb4Wdvmo+9MgJ3A59wznHh
H63BZpx0LifVDidsO+nIGcb7QfYaqatlGGj2khztBIm1TDUqZ8rrft6G5aoQVboQ
nYPxMrejWmFUx5+WCkUvQsWKPDm+OrIKvs4xrbjFY51CSWm+mYC60i8Tpzddz5u7
rgqi4XY6A4zv4IEPFTSBzVklz/1Bp+Re8VYUi+ifLVza4oD82YF7rdob50vgCf3u
J+A2c/KQKhkIIcNmgDch/rix84xrmoblJDEk1GtAigl9HEaFw6EKcd6z0ztM1q7W
U/u+wCcu2qd5ALoTSWo2F7/mGGIDa/NUHyfA48v4S9S87d5dd+cIYGp6CBBI3BWw
XPh7+8go7ZY2YLY1Soqrln8GP93miAeLz4/eCF81pZ89J6rV0qxST2H1tFRBneNT
LameiJ3Rihp2NiY7zVrn0sCwhiXZIR4+eJvsPEa/FZ1GGRn3rXhDUcXdkxH4DRbU
hi+/Xs4XhTaIlQxS3QH50HlNoN2CX3oBqONT4DRQ1waR06vEbNTblLHBiV6rTuYQ
T7m8YiCzRsaLFgHeW+6ar5dhbwsJIH/wf5WKJfQ+Um0Dd3Lcdimfgn1D09WN/Gtd
2JgLgdu0UC/EGTBfZJe4tCOJBH1Qbb95V3NFAtyYEMl8jvi7PsrxHOb/7zAjNJb6
SCT8xoHWhpXG0QyUsHPlZTJx7feSFizXYVlUZenPQZ7B/SfsS6rGTqmP/PTvuW/J
JbveDuvtC1633diEm1yL9fm6ixy3yTU+Ba0cuFc8QduLPoVlCWJpYk1TvNFvtFuC
V8y2kvW9mvKzMzEW9dJSRBlBOnTPQPKL1SUr6MZtgxdH4xi0eZLkYw3qobOQQLuT
Pj35BNPZwdsvCSqa324mjTfQOKWjNvYVf3/oj3jZNbMMK7WCH+NnTrPw/dt59FDc
kcvrZjK+c1d8u/IXfq5Sw2AosXxDvsnCf2mEnnyL8Laq2Y2XHnvyfk+cSxEbtNQR
XEpcKHkh/dz19h5yARwDyShKhyUS97ijrpL9tc09fLIrYc7yHfcSVc2qZg7d0a1R
dPqNG7F3Jj/YavCy7ifTxC4Zykw9LC+nGyq9ULsl0phax11emFxTJYJRC2GfbKaN
qlCMY2KIk0UBPf8VzEbm/tF66Vy5OUk5ykPavvT7XnWbgO6z8GdzjlfSzH7vtI1f
iHLirbKf+OQ8dJDCF1FHlOVTXaOMz+VQp3Pcl4XZiUMUv/DN3DoZI4UGSGlEWFwR
OCHq0lXSKFCaRCq+yOSJ5DsAosZOJpaa5uk1/c0sD+tG0jtbDK75hxPqKiC9SYV4
gOBuMx1hy1vtxC2pfj9C8iTqa2cKBhnapOQwjeRNBR6L5yP+CIlfpFyzTlOcO4tr
FuCdueSTaYdT/SP0SdHRqLRP1aVvV2+Rtm9/QH42lN6zdTBpz0e0Op+vTSEqv32E
glNK00o1PdQAPZuuAfyvt5vAmYYzgPc8Vc0Z89jCLS+MTmCRvf0s22CZsP6aPwj5
OIuK4e+v4liNxSjMiYdBwWERzsUVKZQqZIUrhzqMR0k/LForpExBNqcT9CrQmeq/
0zGNwDiL5ubdlisWZQV0I5E2xV9B84lXV/684QRsV04fVUhZk4csRF9kBJ4SGYaQ
g1VbjH1t55HNH0Exdc59rtcgWBaV3pAFZSFooUVpAZbidndd5R81wxWwLfkloEPO
UEfyaNV8uoD3WFlTVM+8qdWg39KCf7wmRZw0VFllHey0Wo4Z1RZt1Uj4TLaD7zYs
5xs5TYDE14/V/3CYZ2ZidoYji3YiiSiargHEs2XHdeRRcExQL+5DLRqBtW+tI9oc
gZXKjyLpxtj2NsPxi+N/quaEX9gSHwBj/vyEAnXWZFfJyFJ4gcCI+sPIbNwowioh
3KYTqOFMLUp3BptpXPdYt6wG1/c/Q4rVIr9FvzB8RR0ZlX1JNDjUD2B8RebAWhH3
RTwEqe6tG14OL30djIilUc9raiMuGYoI6S1ZeW7UpFztobWNNyUqfj9tGdDhayo9
ZL37HMT4O1KDmO0IrgKr8IJ5qwshl3xoE/ICXe1eelD3Q1Q4hkXoDUZHuFQCphXb
MnIglEI8XabII3HrZrDQmCtHo2RHz44NbYCKWM7/D+502HmT3YVUfZTdP1HnQ3lr
rkoHSJuHywGsL599VPhhu9Cd68Zk2cjKuxoIE+UZMPxvhallPjurpTMtZt9gB1BZ
3Qe+9LUyLIxkEAgGqOIi3Y7ED2krWaD6GtRmnUXF3T71koO9RZThUHRx+jnuk7DQ
PD2E6YmVDMDnxNvvujwHG1GWi7wZ67X4grGwK6Vir7I+08HweFQZ37gJln0lddZr
DBquLsktYyQFk0N7Phnx0X0G2lY8K68O8aMijDKJdIeYfE1cp95/Yk95K1Uwj4mC
iUES2G2TIL1prxH0fo4ygknxNjbwX2AuuZW054/xzGZebd83+SJdzn9MvdXp4cuA
9xR4cBWnsnH/p+UdDyusjyaB/rfqscxtUfrAhYBud9ZdXhx4kh6T5JX1ZA5h36Zp
7j3KfKJwTzUkzDbrE4bFAya1Dg2zmuU6fZL9Iw/ermfKbxuon4+wPQJKNWv3vwp/
yWfFI3pVt4ZDACrb+h/m+mT7JNHubSQ06NxIBtNOZVe6mjDMvh3xKsLegAckFUGm
Ik7+FgwGJLS7R1LM/TkJqVkOm/rbaVsCSpqyCPg+hjJ+SuZWt7cFQgD3A6T6/7bJ
pQKXaGb3fhmyTCQ7V4q6qwO19WiJn6NNCiOEVQqMnMnrIuOZYDMqfIB/qpx94s/H
D2hvcEm9/4dWCCiVtTadcW8RMBqHquk2dGhyYdXcuHD44giRhem6mri4jDjD4Oao
CZdnXImnt/g86oR1ycRAutIO4r5TNQjtuDWa1HVPhsbmKOvEw1RPCq/knafGXcoX
pOLVd0jwzljYcy7wwgFz4WWJwaxZzShAyCJM7GkyuA+6L2pC4N6uHpSH9ms09SXs
MdVUK9iBJz+v162vT7beL04w3E4yL5AuD6t1W8/jq6rS/Q3YEyVwdDPNIUI5mubQ
AIuweK9YYOyhBPHzYGi7kpguJTaSs3y2ddLlT3mS5suvL1VjIkhJ4tiu2Z6qm1Rw
/Pd7wcqPj2c7UU4o5UHUzuIv5joewtuCJJjr8fB3cUNf3NJXHKGklMFuI14LOZ9Z
kznADpgFuMfakn8dOU8mPMh3R1YhubxTMvp9SfUQpZ67+X6KFI6Yvo1sKbJpJ40h
IrfLvU3EB2gs7Bue5p++pTogXoOwjwYuJ2YL6jJ5VcYiaAi93HsLjDKM48TkN2KC
jPIuPMVFbQBS/3HgElZTckYT5RLHCdIN1tErs0BjSO1G+fYm4kB2bBl+doZIipbN
lKGyzRMIC3ZQF0YhtHz+doLwO+upNt6OfdnNYqjCAdy2AJaO7oMQtAiDu7WvPl3L
Bxln9ZR0KzS4WLE/SFMlV53YCsjll+5KX8v5PGJKOuvAroGNznwH70Cft79vRUlG
gZ40htEfmB1jUu5/q7kZmlINS/0CnUA7xwoc8HCJSLOheaBKuraenSFDhuIZESn6
7AwL1B1ycYKFBTVUcyiPA+MRiV6XrBSkvwEHNeUBHhVuc8Lqia0ZhJrXwfpTzyaI
jY5JPTSxAvohAcCtStCZCrqLZKzR6GDsp1s5DAoQMldJ8DiAK+uWFbr/DDrrSR5v
uLBpBaq00V4D0c5NZfWhpKX65Q4XvlQLPdfjcTZMAoJ3aiYQ2nLxOvx2jPZxTves
g9s85vEdb/U0JD+DbkCUCbpfmQae6snFhrIPel3xsfBNk4IUgjpSf+oghdN4tws5
vz6ZB3fMwA/PgCqNxZ8uE/gE+gchciSBFkllVdRgk+V9VRjBH3/IPRJXRbBJLRME
aQW2eUQuxfUEehXduMnB/HAZ7rESK9uMPz5FB9ZbauPre62zXMtOORb67QEnE2jD
pGk4w5lZXWmIYBxrwUC1XiSyHi1lKuRAtFnV+1Gav5OxPzM397AVex0Y+CnDoVmm
pQuecF99YcFFs/I0NTtWBkJq+p8ycpd7ldvFVZWeHQS7YorMqfmWxfw+VmSgZuqH
1PTH+lBliFhKP6BLVQKu9GQJ1G2TEyYh3SiDbwNHOgm4N/afiVuezyUVJeqVFzqd
3cnplMqePRSDrBWs5ayHAgunvLoTtKiCvzv3oH7lx5mTfj//b6cgxMt8KdNgRuro
4jXIvPfHHBSONeiCmuOcvleVyRFsP/XGo9pm3DF3lVoUHevMoQhIrWTE3x7botVX
II6OAcaRJinz+hoAQEbG/9YxymBVDiIj3d/kSbSbKdQOukEAetdakYfJxde2XO+I
7uDq0BacvJQ8+4M3d/7QzmIBpb+SPNA+NBz/wd9Of6c6HKJl/sZdPCFpLRVqu/Yz
/6P8EaNzNefJpJwuxzT3tQ+csepp6c6704FT7889uuSH6y8KBM7DuU4oKy5o9fFH
VlosRbo9gzB2txk9q8ZSxCai5cAhMBsBfP+/I2eCLuBcKu1CnytjkCfC9zSFT99+
ngl7zsWhS4adnkKN8ziDfVS8qoaZawpmSzbUy8cPYpEgirUbzXI8Rs1L8akNQCik
NlLoPyHD509bwL0ILN7BiCe7IAL1lKVOlEXQ6uRWoyXtwHH70L/I0piZ+nim0GrJ
bG6bSF3ATRsEVCXPnKkBiG+eM6arWHM/4Bop7Y49SheOmbrIETLuJpsjbqwGrgvK
w1rOUv3wokbWw4MXptmDV9KRLYZR+VbFnMFJAFNvuBlM6nxfLcNIa5JLiHatbM5I
u9MIZ3t+fdaty4puetW6H0tsQTmO2/vBg7hgUixucLesEfGkJmmmc56ECZpZZkDf
nxgzPFVsNtQ0moN6EoxbCUJwYnw6QMVByEgvuectD/BFVzncuFB4g5u5hlDyihvY
Xgi/j34+gBFbbWkGe84fiYMYiRwloj4lK5q80IAqxkZwojTMmY7qmaJq/WLzZ48N
x1aZ4vbZ2VVxW5pd612/mXLH9l9VuVBQ3Oh8OKQvF+t6ovdBYMTllGUc3PnwRVq2
G13RUcWdr8Afccz+7Nfqe6DkjgO7PHY0aj7DYnFrV/15N10pK6ojC8yDtJXQIgk4
YiFCr/GLyBKUABa/ITKz87AqHMJgjzksjm9QlCMbyw5gxjLs/yGKBx99ndBadIvo
vweDFGSxPxGuz7IRmdW0HEXQjjVogLFFcXW/Xh2LmXp25cSbLRl2os73bgXzq3Ys
ddj0yRrSj8pitzBfIChqZIZaigYbPDQBIy4Rr05JqKVkp5H8S+8iGhuW/2MQkP+Z
VxTP8XXh3UHm4VgsI6h2aGb3IgqCm9kezyZUvghdPJH4tj/tBTilLt9jHmVRKFOf
iWqpc81O5WJkJb/BfyKs131zwdoM9r9o1nfZkrmipEq3rdU45LfJ6kTQLukDvrDf
RCvSRee0rPEzFi96NF75JBdNP5KR6whYOR6OpRddBSUToDy3gLNMmQPvQW6gN5GF
/yF3lLXpDiwCPyFnJw4u4ocWOumsNTUAGtAq2Trls18B2MdhOYcFunETozsC/2PD
kUfTuOOz9V+i/DNTYgB/RRLhSscQ+zFhcTZyJQxdiTJUAq3+cEMKfpL/uLH5WeZz
V0/kckCDjLXA0rQ7MMqBoAyodoyA/eT7C+VAuVWW5JCcRCm+toM1Ijq3PtM2+0Tv
RqD2JSPBfscH06ilt6KR0PxxuJiXyHCg1Bc9br8rpgzqOYty+L0Tr7mF0sE/8dYI
JnbfSYuvG5Ky0q/sb0JdpOAWPKeT2nW7ZViM/CHC12SBn4Ctq9cTnLFhCSE/XLxW
bV+7ZxAhYZs6eXBjpatFff9UGdgYX2aRWGuq7Zw6B1fO/qtWWFFBWApz76W1lCph
dc0r8CHJUPQgXDWaG1tEvLKKxBua7DwJ4BMWZVhT4iNPwAnA41QLOaE7PFlig1q4
+n5UCdTvfeBFIvYSIfo9X2GFvSIBl5MusN4FETMrdcKMi/UXNf3hdQZ29fFxtGKq
OZuX60McebPAZlf3PO1zzEKyb3tbFVJ6EH0V9Ay1yeoP5KD5c8i2E59dlLdhxjzs
0bV6guJQDdiRb//TMKgrQC1GmIj/NtfVVR6q1pgqzT6YKjJpznWQ9rHcSH+BguX1
16NH4/AI1fOI0y0B4yvKNsZqUXmzQfQe//vvpRplZ+tQkUZM8x0bbwX4emrSt6uf
sAeUnaDEI3VouzGB9EPM4pRDDshXuUdj0gficsRI6hRxHTP+pVl+P5rJSGst8Ytf
xu8Xo+G8YZdZyASi2M7/3KaAsO53AzB6JYjqH2TPF9FSOQfMWrrNctkw48dfMg3s
U1ChEJoqOS3R6zGJ98W34KsoTnUPVaxPOdT19to3zwKhl1Zbet9Q8Ty31tG1KJ06
O8Dp6oXsSEfyKR2DO/5UCFEgyEvPRcBZ+SysCsvU6q1VSeatoDJWCA5gO5YCKA3H
6ueuyouQDVcJXKb7ILP8Pc5DDyDILoGiClcI3r7NjQRr5P3jkDHfBFqOGjkauJ4m
fJZZGj86oHAQcKTT8OpvgMiP3jh1GDb0aXlgfDhlD0WPMO9RxN6OaRjHAfV394jm
MLuxGBjhUd4PJgpnYisiruHjjiJaAkhMS8aXXcWq079Vd0ix6yWGQnbuIPbAr8yf
OXeV9nrHEdIZlX1i4LPL6Kol3jeB5BPWhRYezC2Sko3Hzq8Rg0yGwbBSW19Tzzn5
C58ABiDBdipnKHlnzAj3gc7GhU3MQiaXBqqL9rLorm5ExWcVBSUyte9nio1WDdUq
HKhveP2UWFyeSs3RR3TSnaCdgaLCG5AqBdhBvedudI3H7haxBY5ZHp+EtXF0eXAA
ykAizeBD9nlFAaifoOkBtOFVOFYkRoInlR4h/hJFmTfGcacJmFbSr+pS8zJqaJZd
xvoTRWYQkhEUsxfVRscfxhPEwMxyeybveQNSUH5d4Lv7zoE6Qm8ug+TMtAYMIN7R
s/c7YImW4I5VVLNZRC6DTjs384Shz0Ogr+pahL/RYj692bzadexFIoO+PrlwqA0K
/FSzrY1dJSnNAlhqMy4vWr3PlgthUZVc/knqBmI07OLVevhNFysgOjkALAFY7IYS
UsykolCib3vtzrJQpf+je01tBUhyqpvnurHaPnPzPGQ3YrnRvcyHoZ9lo8tIK8Zn
imsAjh3Tzxb/F/S/Zx8p68NPfYsO24VbMiKxFkzrFoIAcmyC1zJM+k4u3CDMBs1u
31cEjUmir6bd8iZdYxbip2vrWkcDH2EhgumiUbHJUEA3ZbFg5rIArhvfY4RYlWH5
xBghsDeH5/R2fIy3sX3y73WEZLEDQAbQGQk0ADFj0w7hiGfvG6/zc3PH/JHXyodG
DTkIw8OSwAzJG+GZlLLbl3T7ibMT8jtMVDGVBEIGf0VG6x/z0KxosWs0Z7FphmRt
W4z3PhOygkCJXoAoh7kWTbXb9tYQ+2p9LdR57iELW1zWny++z5QV2Me32Q5i7MD4
pgCVPInW1B0skaiBuM1rRY96q02fn43u+UWFa7tlxt9GSmzmZFFbBm0kv76xj9wx
C8oJwcyibQpiwwFXU6lKPSEl0FzAXZ/HuONVdTsGJMQHHXWJehBKpM7uWLL2S5TP
8CxvgSNSc1yXIDt/OFRamZGNahFG8XpTSJ3i7zENzbik5DTbMPCZVEenfnIJnMFb
r6dyy0QoCNddzEhXVn38pX4WCmVFTRJ67FfFFckTX8ZyKIxhXRAXO/pxFnogjtWD
E5g28/vvJzEFHkezcl05CGJVSRIGtsGsRCL1AQ8vHKSaImhWjVSXH9UxnmZmbGn8
7AuDdXFxJpGRhTTwL6qx2jIeRLmBElRmSyhIp8JdYBDe/QOpEFEoKIGIa1oVrROy
sDQQlTmXis13YhV0zTyzJJIjGVA872PtLnFZ++W8gu//jzrpQwS3eWO/yjDpDxub
kc1kKxRq2OUSh0jU2Wq9WzInAyTM2f+i8QRvy1vUiLisbTeFu/LiNk+MPRmvjm5J
LX5QGO9pV7EPfTTNPt4R5o+FjBo4NKZxX7q9bjGQLMh3fvdP1v5RPGV00CtrqIhP
DT7/hRyuX59Ae55tC8rybTiFTJZpKteK15lC7MvidjoWn88x9x41TGNPbqjTQlH6
VAhDBLS2R3H3U8YKOzS9kcPFcyiOfTJx+m85I5dybSZIMdREJRXQDzX8Gyj8gLYV
YyOp/Ka2x2Boptgb1KH199Fmn3GiQtcERldcutoWjeTOAb69Ce0mmdFwjg0Q9iiV
SwvgOUj1UygCKgS+BHYzr6fi/9LxUXO6Uogp8oSonRrY7NS1LdtZ2fiW8x5QlHAY
m0n+q/6KxJFeX2RyMkXnd/XVKYsJxkstFuPfYEx0B6iNbaC0RTe9rsHOeZda53Jb
6w8OCgcj1Rq1OhowiR5kvry08psRs/RpK79LzTNVbKTBC+ftNf70dMkQaGakR0hH
VPbbS5h3u8fyp/yzIzrp50/Ld/xfdWS03btuHjKCEglC4OloQW/qcJzj28K4XMwE
3mefB0EYn0QehQU3HDuHvh2n1lprRQvCW5Ku2U3/4JGlbgNZENeapNHveV1SoF3a
uOIIJsJJWKUv8tsolGykSeKlzvAgkQCK9NwurZ9ZHbLiF72dLkqZrXSClO9r+14J
UWkHZSZnuzlwsJiJMAdHJaeMaSt6aPtdCrkO58cv+jLtwfvmo+QaNBwwk9PgULrS
d020S4j1TdHmsi4m6BkskNC4HqPBTYe/NmkNceO99rWUIVN0bJJB4/B4lMLwM0uo
zKsHYGPH8J4ne2DHdrSk4G+9tdKfKnerACJavM9tnS8ICdeQcQJUAIdl1GrDlN9J
6CVBKxTXvRxIdxZo51I/Up2Tiwd64zt1nhUbEvRpWwQsW18KiF8z5ld3aRHm0oHa
cfJcgc0sx/aTmo8lm/2HlgBnpxLVX8bOTbeGJZB5onaw4T5qqVCctwu5OMxVVqrw
sFcK4ASJgWZ4fQ8Y5/ARxbH5KKGVFjeiDHYuH5tLd4i+0DVkTiY5MrY8PH8J1Rj2
SDMa9SksjbtOpua+ONq1PPzwlR7+kXvKbFoaa/VlqNMDvfZPYEd0yg0fLLfG2YFl
NrLtheptd6bkpxrl9VVSzNDtA57uKiXKpjp8p9ZIWMs1nIBHTnbRHJ9nZxWPYUp6
IQsf8WtDy1DZ4VZakjnh8roVU9/zcaaKp/V64QEMo0qgA8oEU+Ht1p6qi0zPZLbn
ANIi/mKOndaHGGi8WnheE0WRPdkvoZedBJzFVvbcCuH0iWX06f0y/WyWf++CWpKU
mlYll6r/iH7YI5BoY1G8SkVjBF8+1/W57UWaSit2yjLkwpkDX+q2Deaq7+s0hsU0
hQX4EVtA7XfpxsWhcGEFdQ/z01/CwMyxkZ4k5FO+FNGp1Xl1+O+ZzXjKJiiRJsfu
Lz+VpvyztIHRw2H0lK0SAb+nNQ57yIuMubGcVvNgtklrVuUfTcV2vWUCrJsTpA+e
XoxbyPjvK5LlWTDtBZp2BFUJLBeZKRtEmhaIS6vxIC/rGc6dN7skH3MJF4kRFyGE
cs97/jbPOoV2S8bzpgq0XQctDRK7516mnb+NlJZEoiqqbJmmvqPu+jE/I15+SnaL
57STH5zxtRet8n59q4l7lYtEIn9cH48xQyfLf16tjPOn1L5Kkkog4j7aFaM/EGaM
uKvC9f89S6fI4D5HxfUytuYr9RgPKi9MYKwLsymt9ufjIuCWFkmojssV5xB+wfUv
PY4Wbrny/5u1bhe22KREIwC4ItIVs9CdXF9kqawdVWpYoQDvcqV5RkRNzdA1PR0E
frpwLifMYd7SALhRcjvlbi8iqby6u7EN6TAs98I01LmBeGEt1H5LzuvgYmqt+aTS
Db9pywOZrM8mIZejhLQnv/yxTGpJlT5yZ6MhW/cS6TOEA7+Lqx0/09ZvJlHKxoNW
Z4Zn0McrOqPpQFiquP37/jGnoZbRFGZGD43uZy3YgVGiAzTxVMUgCueHy5VYstvU
Bs/CrPqkQM24ZMWJZiYcL9qdwf77pNbnj8bOh3CTEPlExfCatC7kuY4pU8ZBuL2Y
z5Fi7b1Zlk7D8aVctjiQqz+pFWSGeHyWt8dKUWx0VGJ0icFx4Xj9GsAB8tA88DEK
7YsHTzkGvapo5FfudQr9AjHgN1OGiIe68PVoiy9J257jeZc2rskQAZBnrBQidhhb
0q5/BKjomveoF7hLbljazXb8fgZ8KbLhNvOij4qT7pQMLsxubh8dCnN6OqzLSAnu
MYSMrOFbsRahtmQyyVq04l9MUoCBLPg4JFDufO+c8ZxgtiQPhIIIpBcGqa6SIjgJ
D7FL/P6X26eUgM18MgPU/0YlmEM9PvjS1DgvOF0M4zfcQtBnxwjf9uCUcZNoX9Fi
XAICLPuMbdHqpD+J+IMhzsNSViT5RJYgnBxAhik1E/1BPLdE0vUEW3qxHsR9krDp
zB0UrzbImIX10tploVfLw6sxhOZ6t32LCYTjEtA3EhSpzZBF4tmYzdjOmH0/n6gW
9wMoxQvezRkJMCyLvxKHzdw8nli5oRhhj0KTqD+pUj+Una31hjG7dgLQaLBBqjNk
vFIFanh1BrXuXdLVPNLoGBBkx7Rv+wRmYKOjr3au5mCQZq54AHt3hHk4t1i06h9T
9wyCU96pymDA5ipP6qLOlpnBIxOAh4rw3AYXSjymS4XOyxuQPdonW06J/x83nzKg
wfVf/H/NsknTnGsNlnqnouOYvaIC0nQmQfm88MHIwLNhbuiqmuTDOcVxgOvCXybu
Sh1kFKOVTXbnkfpv5p1x4Csp5khww2VA+AloBbSmRd942poIrVAqDl4pPWjCirpd
VdczYvH/Z0EEVATruXeDJRSadpHQlbnSrjnNUsMXfXX9GsOwaS5wCicoSHwbiRhE
q2aN9d9JEzIh9WstgYfpr24lPU//aMbk1pBAOeXXgC4i9hJ1sWnXMTpxyEkhh/SN
znVuxpP+YljE/U/8Lrt0/B6zgJ4NLsr0+TKq1O3K042r/LBFyqVLdevEaOKGvIoV
/LPX+QiGKpaUQYZ0YW5tayu+oS5zGHy/Fs6Jz6IiLE79AjT+F4Cbmodzhg7HAFoI
1RpcoLd9oMCXsQbI8z5B6Q67m1RQYfdfoPS/Fvyfp5vKkCde69lZg+GYNTpFZ+4O
DFg+DvbgfLhzLwKGxDYgLn4pJya/8NrPpb0/6CwB5DD/Pd9d/x1jwj7TmzVSDK/p
mM+HPmc89W4g4XdsRF7K5nDbnnE5Y0P5J8BnKhP8vAv2uFiJ9qKApN80alJD67jH
8rjTaID01fUhn/tkiMCArkCZ1EVCaVIBFnHIbrj+Zy46HKe7dWr+3nkXnSF4k/3K
XFP7gFIEaH0zeD66F7p6ec9ZbrYYo5ua9qmY+o1eQBc8q19RqeXzirjz1PYBcff9
mZCoA2p1HXVzs8oVr58smptZNTZ6ZZfd2QP+v67+B6/Id5griCzF8j94K45cQ+Ot
RRu64vUSdM7Bh+h8O+irxEh/dZxwf+zexoDA77sQLvnYPrv08cYtAqXpn73L8+WX
K1ua6xHDhNZrxqECudQ0DuPZah0j29BcB+zudhfORPlfyeI9lmw9tAdivAVwhRah
3MhyEFEP/8LJzi1oMscjOnUItbTXZ6mF+Nq6Yrdf4UZt23cTvoSIZj3z16wWqyRd
HGLSL5FqsnGCiR6+56j2Z7PHeWprsD7jPBOka/6O8Ti2EgBPw3NjwSgtfuNRYpRv
PYQpZbiQ4qtcwJ0LtkemyB0v95WsU1nYVPvtldEVTb5IbeAMzqRo9ubZ/oNwG7qu
jEB3ecLqFXaUboXtZ2Wr7+wXA9N4CFJqvaBN9rQV+VZIzMqCQI+cg2RVh7MxfgPf
5iVRksotZZkpbavbtB2uC7qjQKgcWK5+/Y2WS6HjIutNWZ9ymTqR/7zg1uI+cwDe
qV9zf/+iXA0EtJdUd146jDngMHEC3Sp+m7fkgu9BcSk9XnnQXbuucI7YaMm5y27W
PPkbqMo7H/HA6XP5ztHSeREUrPI/z/Du1dClGmPXLDPnhgDWZj4q1GSoBjfafr7Y
FHH/6p9PxImF8jvzH0IdKjIB4/znd2IWsdblE7TKr7rskuy++w7SC3nrs4JU1OX6
cehGMuTgVKfIbZ99Dfv0eNa5js03C0GsHQLmixSD6OQeFwu019KVrKRgXlhxKGwT
KB7wnUHlMUzF98RclqGvYu5HXjKPQFLpsPpDLNGSfgHkW4MX9ySRln580/gUtBTO
LXnveSDNPHduh5s3eZaTFFXhIDlt5eKMo0zVrLMLNPBibmSMGdBrqw463CCQAaBl
7giiGm1q3u3rJEr3u8aWLy9NicsLhBh2CdOSbGyim1gxy2HlP449MYvGSFmLjhvk
/vFiBclrnT8a41K4tdZYq95N240aTl9fpNqH+9ag8Fg4IqAvV3H4o0kt+27nNjZ7
g55396aM/7atHMY6d0KAPS95QZVqA99kQpSL/9wpZ3FxEozv3p2tNj9S1cQce8NV
9B0Kdlqq9cWtGxOXMJUb3yWmIRMEgTUtjOqkYzWof+XpJtzXk11oI9S2yJ5N94W/
vXJxVtXGzkT/qhN/rmQ9UQqNA3qAOCUTp4XCWO8qC0rnHVXDVJsX1EkbE8k0CMEo
iK3G8blol2bALfloW5SkRx9t8aJJUqPGMbB0Zp37NfS9LQedf+jCzBq/8QTftq3g
pj1H7+69bb0MX7LJ9CkqQMRmROr64x7uneZqhbYlhavgcUUA5LcBgqk6J/LlyPuC
CkkRbkzH+6uO3Qd5WVuw/BawiZ9At0Vy+cTfuO8W+vL0P1CviXHZWXJSpYS6FOzZ
os26UUWynQCJevM2g1VLuEibbgzK9xqyOm8Bk30OZ2tCaDmGEDqYFbc+ipUGYiA4
vG0Dh72n5b/IByFH5FcR3ohc8nZjMTmZ2P/5ecHWGizwKcqRuohTmAz3wkskFxx/
WRujlkn/Z/59xi/QvQXdxsNMzvmWkDThWaFUEur2Ni9mfk6+cHbePJFLkV0ebEp6
r2WX5Wcg7oXwhKf0G2bJglD4ezOE7ZpZwPrGAh5XFSPDkYgeZnY3GSO7jof/tiLD
KSL5UZj+KKboBU/MzAMVDm7Ox2XHkTUyn71Gc33WoyYiB/eqrovD5R4e9LiE6sWq
giUxcdWP0GibG/1h4zRM44T2L1+7jIuecaAH2JR7qpZK0MD45Ss8nkowEO9fjp5m
GGpisURVU6yIeyAzqOj5fSTPHRPIkLLOqXAzlZEyXySK5ld3aSaY8dgNIs+4vp5w
b1PiZ9R0pQvi0CYhiaDgHDanf8nOhGrX8d+OJDxpkGytyIhQr93+IWwrZdaYwtD9
eLg+k/yuRndvL5zKAw3zW1XHW/DvvgB5B+INhDX9Qg7QMalKhG400ZwaK0TK145g
EXsR4grgrWDfnVtj88vY7N57yC7oKV5pt5DEL1Jk2DfCvqjUDX58d5MLRqQJ2jzS
k8rjx/LWgVGUIBm1FjE0cDxJZxEuW5Nt9a6F1ClhJ9hc050hnQaCLUbEwPyUyyHR
R+MYhLHAp26mu5numFpN5R1Sfyh4SSrUIg+e5oapVNKor/dbRmn7Ssi9HxZp5EVX
kqSB2G380HH2r5pfrec2L6sCu9DD7z5xX1eKMHGZBXmwk8/oQi+CM0uXC+eajC7N
Ai4UNcw424HKVWBnlAWvWPNZDI3UqmooO/IX6nRhuv8ZYap+NcF++AxL/Gr22sqq
x6usMIEB/Zwkq7qB+GjKFwFy8ZBGKzNCR4/YxGbqCc2Dd8JDA39mZymIUw7DKozl
tR5bn3Bm9m9n36qE6pWKmix+OneJckMa6dTAQkYc2qDqiQmrixrVp6cVFHKY1VE3
IDdV4LGYHPu5yk49E3TSp8GDmTx5mHAVnuPTZmSZxM0ha6CTBGQroVU1uxjZlUad
6CVa/PQD3QKVlf8fugQ3AoZ8zY9/PAPRvBu+bL+SJ+iHYESgl8PnqOJVRKcAP5rQ
uyhffFcqJCtKMYxFUVvipLezFs/guoRRrhzqDqDMdyAVfyiuHYpEI+dkdtCz6EZ6
64c9SywAzhbXE3pixPtQQYV5bYWLxPGCUnUwpzU8HyRW/BpwPN/aKGVTGAmtl7FH
lzTrUgH8hEeByHLn7yX0ixX4u+1pI2etRVSVHHlCuHO7nQTJ1NBqDehInLc7vd35
QpFR+qNxJYejL2zy6qt5m1xMvxHpMgcdValCi3sc/UJFoW3S75DeK0foP9ym8wJn
OIQ2tPLVVnoXz36diLySsZb1FXIpKBsKjan4BAnxAwQPLQ9kRxTV7wpFmLkvSm+u
Bq30tciNi9eKGDOt4Ejq04GoClDZXgR17ixOVljKmKdIwqL0QnZj+Dm0f6oLHSXM
Tg607JPTXyjkQdRqvCUN5GYhj6Xdm2MKh0ZQ7rulVdKKc134igtibvdvOVr1Zc8u
ZiKjza1APWCr3Gu2RoXee+NqFxZbdhaiNCqH7mbVTTMbg9luk8RGDGpzpyaODF+u
nzYaDn4KisHIT5K0RSYKnQg0W0cJ7ryMzsDpPnWj9qMG4SIBqC9bqEUJCnfkK/1X
02nUYlynsUl+Q+aIZkIzW2ImVa5aqBkLvBMnvBeZ/9iTVxBhOgSXso+dc2fmpKK+
j6O7OxQZU6TCsE7xkLAsW0e/i84ebEKpKANcdnFc1fBAVn0GmpOwMRG7ta2DxsJO
xfo6uwbdxeA0YQMQSI64alK9FuXSxR4kpzGgIVsZaBqisF9zS/HT2ZZO7Pp0UfIQ
tZGjvTQx47G/mqxdBvWdBFwEaqLLz9GKpfhZt/u2YvEqvFHqMCn2yrxqco/HxOJB
i2JAH7I0hROO2/4UhXahjaPtMhnqMwMtkMj4F+PiJDMc0qUwuihS+MSuOxAB5IRo
FAPJH2zM5HK3DWlOz9iSd3cZMpv6y+kDtFA0orqc/NSFseWeh8GoWnw4D1minjU0
qe0FiwI16QLyz/kXZiL11jfmeNGr/uzkNKbydwMZoiHPADB7m0CEsgdFONr0oJ1m
25CMerSECUFjTywT0GU7kOABPCLg7TwY2Pfvf1M2TTisGZIoa2f932jumgni3cUc
mfFMnhMwaIaMKUQkme2HQulxTfxfpwpzvlVMdPppYxUzMnuOX64JvNZ8wQwqcW6N
N+3LmqHYFosxXcNSyTAf9OFVBrfbV8gE8rrHJUHzksgdjThiIPCYadIgMIHB3Li1
sOD8ZLe0y7oXO5C/f5mDZz9QzDF5KuhetqyY6sDuQD2Bhp+Mo8//ukjTAhrWQSXl
Vxrh+uyGi8RHx/RCwzUaZrJ2kXCl7uoUg0SWQlktRNqVYTOBSLTWYvpMKsAicQ6S
UlBoOTl4hg1rCyM/voaeFK0/jzEJkDBbWuUtg6s6+9d887SdDIOatDs2wLtMjtxZ
P4xPjF+KNDIdPk3HDB0RUf1XyoRCK8CP0lFmjCsDiLHiFqaNoeKY7QfvL+btqEs5
oqHxdsm6A+HCWCmkgTCEB8H95zfb4Khi2OyWp3PEfcISdrJCtc25xAbGXU5g9iJx
Hdidm6GmrwJGUq24Qe1WJg0HV2cZdRsyK19Rm3sNEZ1BgEbGXlaTUOW1+GIyKFxQ
r+bAq29tGEckY6Z/SThac/VEMpY65kcxFQdfUfrC/4CI+8nJZABkdWPFCAjkLo/F
WXXovxfAHzw8GPCJIdSrdRnttWgyw3h6WhwfzuIIgO9FdRfvwLhltmtnCHCVWdJE
eVCs2H+z0cBeD0RYhLDd86zZyMnPjLoTs738Y9MlXWN7641oZTnGBjVSVKX2pnIV
91WhkuHSvxTcIuKVwdB0W/6ofKQs4eevSdVfXzWxFhTg/0NtS3Cfe5z+L51NVkHj
I0ECYDdzPzC8D7aGOJPsnRx15USl6KJcVl1UlHpOaZq4U3f15HppAM1Mrsu68Al7
S6Z+qeDP+xjGc0XEBNvVxqnv7v5ubzEL/PM6PRti8cxjRqNHB17LF3mQ5ZxRr7TY
geu3UikNdJDPsBTM66TZtgJkdjqEcOvs6xdkhMatr/+VUR+1rS7WmB1h2LKkUpZN
CUI6SyHtvjuwIpae2rxntAXNs9C7Fs5IuuPmgkKUQmoDgWEC99to2m9RNjrIgiQD
CZZ+sAeVz/dz6S3G8+6wVmaiPS1gKBWw7TOK9xaLczfn/J2RT03jiNzpz10oW+U0
gERFYuEqA5w9teHVkV6+cm+R+AmaRaLWVsb0OG5N2L8KQGS1PjglfrTzHfIuXrs2
bx0H7hFu1g443XDvoQ7Jk9XP0+TYOUmDGqS+0eyksjnUCAcDmvwfidspgVyLKnJ6
Gc0t9dKzOwSft0XzJ5KfwCMI9rnfwHY++rRdkMqasmk3JpDgppmYF0+bhrySiH/V
gJ6RCKXakytKcLztdRkKtlX9ZMEUqBPaWLH1Qw0+4RZVKQyyxBcU9oVmCnAg70jr
oi9VQdIdhHidKGTenx3zig+12bh4gI/WmaLI52RiVJ7u7eELqeOoPmshNQPGN+vo
6cSLMlTUooLVmyKmPq3dZ535h3ELEnYYGi7cupO7fJsHPjfxkOXgnZJfFGqTE36C
UwP1WfX1ZbkJLKGlVaBbVNlZ23Gf3Av81uyAO56zOxPLdYf3STOC7k4pKu9oGbQv
eXZZzGfLFFJV3h1IlpJWqY/8PjvV3D5+yvMq0MzEvlJdKM1xsrHGqFY03wHF2F+n
LFfazHQ0qPdeHEqNj0m+WGWtub9/+NaDC+QlF15ae3eDR1rA2Bxs0h3NlkVgHMOi
QLCq1/oZeEJAcp7Mud4thnYWzRAVLQm6o0zfwpjngGJYMxyO/6vculgiWo9LMkDM
u3bnW4y1aDvgDagzF+TZYHSrsI3pBadvVJ+omCpamqIyJll8JWnpFxv6zz5Qw57c
z/wxiSv68JtBbEKI9W1ErnP5cT6Tbv0r1NNJ+F3fJFKK/z4CPXfhRpdMcWNJ54Py
dBAeqq7H7eX4AjCDmF2F+Is/vEobSUzaZ90Rc4Tr1LniiugB6iWDn4BuqbEHVjtI
IacM0Vca69HxOHgr+M41wTt7l0c8ow5vUguorOWTjF371C6tGwcLXgn0+Omv6bpI
cFRJfuMf/fg1DJPaKNvKAME/+/FdcE2lpEum0HkfVU17Hh3AoXjXZKPpH8pHS8td
Lc3zhg/O6CjE7PeTx24e0BFomdy8e9UYYLvtRgqAyXTMb1zJhRWwn/D13WyU6o2K
hxQrGKj2A6GQGfHjqybGXbk5+ooIYzoPnQPbWBWLBPYmasdKa7gVVgWfZNZ+YnRS
Drqu/OdWrdsBZVDiUi9NW7zCXleQoZgi5BzzMGIhCpbdldi0hviFlsWBuJfO/ciR
lW/GTQIeeeeAkI9OmpDVjIe8fozPjFgd7sw2zoyimBZXeDuMtzTeCnnXbiGU2OMU
AK0ECJ78kuwW+D8vlKpKGT5hOhCCxzGFV9U352i3E7IsakYuC1MRcMcf+yngr9Dc
7MS/AYnZFJv79EXv0hx7ew/ih+4dNHiAOs8iuhcDWmsLSQbp1nUVwaa4mfAwYvj/
GXlEZM5lxcPeaI/oFI9vv7mwTXY0lL2FRVYehleAPuIcWjjJAsqwssJWwJdbvtfw
uIHKDAuHZl3S1rujcp9SSN5mZ4MpUNQ5p4llHwPM0mTUW0JB3fBB1xi5/ZIuDvcS
ePYYLlLjokp4yV5k45QQ0kz/jxyDPmsFv5dHVKj8YFSPIASn4zj2c/2FbS9w3a1H
MgorW/e9R7ApmYvXWrRnUlvC5vDw294jiHTDxlTOPGiLi9/4sideK4xe+JNhwKR3
VtZHkckHzOz8q1TmDI3VnST9QSH3YwKWTy10hZO2O+BcndDQdEIcUG9gVxGL6YyB
BcI7z8k8320QteREy38WwgwKdioEpqvuBUBPNbRVqHsCeQOgo+1WgA7I43L6HZo6
MGJgRSIMEeREIeCM4YHEgMDhJaAehDfhlugb16IRyEQuqbDfhp8xLJIb+gd+5r+B
7wxq2Ibq9XpD9NDHzjrHKxkqm/r18Izeg8NktvT0Z0Tjzt2gSzqHbUAS4L8telP+
Mw1a+Kx9P7dyaD7DTvQMjlP+FSEunrMRBZ4rW0VPP2VxLuO5F09oSpweXC4WqpzX
Zl5dgpjtWf/jgFS1mZV5nxPSbzIFb0uHHd7aZfQHL2iJIHyC3BpHuwFQIUQuHvjW
uR1mbRMP4wfd0XFQotAIcTCPiZrwxmm/vwinH/2XYBZ+o8dRp4v/ffsCm/kTeN98
VNAPNppUxCxS6ZvLbHG4li8U56exVVsXppDfB8dIjEtQgE5KFAqi5/+h3vSmkl4o
dkqmV/nq5iuG/JXCi4duUyI1KpfoAEgLV63xcMqWfWeeQ03o3J2G2B0TSkRVqSX5
N6OB8wMJm2uTjWYlOPhtkL+dlyN2ic82xtHxa5LMyDS5OTHDwUdmmb0XOoI/upU5
S5v63jd/18AscLt1SAoIXlRBxt4hOSnCEorjhLZUAe7HW4YL02eU4ArqKzJriFAd
OZhUJl1HcBKjciI/ExXEAsfQdVgrHRgCi/U4x8tVFJ/32qcUJ2Zutw6R/4UshlyR
ztKFB8rIAGW1fTAKNOLafz86faC49u3fvxUHh8IlIQXhtiXsFpxcvsIx6nNGWUgt
jcfCs8Vg3EQ3hK9Qxe1uSxOXUK0s1VGYV5HXbdGsjF5baXMUplPp6/eChFQH5xX/
hg/M5LP5/t3ogVXyCEnxpvb//EPgFu3/JhIJ96iv+D5wO65bel559mYySUEkAXRh
MmVCdmz5D13kzKtnz5XVgc/bc2PdEQcZgrPZCrC8K3mtefK7taoUegChFD79yHi/
LzkCnt7Ugqlg67+VXcnp4CFgyLaZtobKeeOkjt0dFM9t2XM2Pd5dnle0E8dheGfN
+A8goXUQzJwCVBMkygMMJULPwUwNhK0I8B8qBeGKPtaqhpty0d2RD7JJtx1S5wNh
gY+FpVXCe9B6yDEORGxNzxyuOMV6Eq0bLpWNtWSQkIAAHVlzRjlVTxEzssZAUiDa
b6PN1zzBsv65v8pZoHwSlsH3Udfj6k/r5TlgSH1me4TqInecVwTSPw7VXsGLTZKE
0YZCKJfRR4Ay4EkGVNU0HjD9a2xzBnt3Sb2qVF0TSCJlqD5hlCO/zCqueMW99e2g
aMNaq3yVZsW5S3I2u7tUvMQZO3IdvCXB9U3lYIHhWmsmSz8fWakJV0sMjV2z+HJZ
TLsOB2FZsART99UvRVV9Ur8VUVg+jqw41NPgUU2dS+HexBz1SeCWCQAzGzy4riKJ
hxWuwhsPKa/k4UhukAHiRT8ZmRaYEU975KsQ0/JhrdY4bj/LpK6GCJYNQlMQbxL+
6cjC5bsUPruPawcccbSVJTaIuOoIavgNQPxDlYxKp1DGVpv3XJhk+jWbu8pno2QZ
OWSO28fKBZsdjER/4z0infuyDBzrMUO1c4lAmrbUFb1x5Yhsks8w+BtFeBaO4E38
UTVaKhCO1iO3XZ1uKJdfKDAybvwJhWz4sMAKHOI/UiudyqipbwcXEXHiQGJ820cg
1zWfqbiBTh5fGVDczNZTUQ9ZKTo15FwziRjCa1A+wQdUK7+G4+TATntqt2dzlWUF
X89IGZwxU2ZPQ6bqX8xUaDcdk7eCW1r8t3F6gWT4Bi5TmVhRYn+Ey9mMZYucasmU
I908tbN0z0ZCfZXXXvlrGuurki21RKg6Ve7K8WyrCRiFmQce9Ip0JipXY9Akpn2L
41kwmVuXytXSlgzwQAyrkhjtE4J4GWpxzD6BuYlrHgdSfuNp4DflmadcLgiEugwM
qIzkpTlypH2VYX71qTcqdGtPvkzvupx0AwQBaWP8wOoIVlWVLAEaPICp5lJ8+wz2
Cf6ZMlrj59xmN9UQthkcuekLZK3uVNzJ5yptmfC42tZ8lKMClFO5ALj1WlMkEyaX
twW+XjtCogWAOdhiK20aB28rvbwtmxy6DHS2hjlAclNw76xPiTpgqqKMlC1ORi43
3Dvf6YoWqnHA4r3/LCnncJa+3HcMWat23x6+FwyHU7b/2VVjLe3N7dg+/unGYMIQ
CmlhcSibGGN41IfaozGlqKQtOaj7ZhBVqOUve2LWBrSgCetHDRBdLrRQSsFtfzkS
936Q6jumrMvV1zgvqv4SZmMw4kzqVmAJOLRb2n+615xO/Fk5EwGbvPPMe5CgLHiR
G9KkwddHWUsBGmdAKhF4dRbIYLZzdttLiqy5AR4By+W1Rwn8Z2CcXcPsZqLMej6u
1IwXQmPg/Pj2KD2w9eOabHhxdfkWVEMwEYeQvBkgurM8NOleowQTeTsDtbxe4Sur
UMgBtMSjGxv+jY/2TCSgnmthyaUXIXhawsAXTESt4mmtcsH3YenQt2JQw5lv0lSS
gayMCZexwEL5USLQCNUW9R5TdtKdfEmJeZNmaqYl2Sa2dOhLJjnK1MW5bRjtE7Ov
wo57LHQbvJkuueOJtLJHYaTkKYdoPfLRRS9qofT5uUfIsMl7g+SCtr3NU9QEFwc9
7wQ2F28nB7aUTly+L+zWg1g58DNHE4v0P/edPx/lsXPw/OBq5xq/beszj03I4F6B
dXcGVhI8ln2oHtdV4ecNddQD3W+J55lWoFz4dmuYuV3T1n7aR/sGblJ3/MvTdPOf
DnM+4HhzaC+KyYsJyQYQMSDtlAiVPs07ZH0Z4zx5iwH0aNJsvxiY3QfM2q0ToIN2
PCinfth6STFgJJKtS7X8jHNvuhZLW9ZS91EwzU4PPBRCGJpH98j3GfDnX6QcpQz4
DO1LZlZNMvP6l5Jcn3giALFv6vJn7szZW4kQ4e9iDefuPMj0OIncVVCPhLJJnE/N
xPQAt/9VeUt0yKou/qHZQi0BjosnLEUu5HUobgBNar827Kl37X2M0tC2v93DeSbD
VyvlFjnm93xgfMAgFRVZBUxYeWfPwrKGvdlXoHEkydvZnSk7mQRTwig8EcdgLRhd
ecrtIp91oq6r6aPl7MF7Y7+iSLnm4loATZBbWm1KLYdDsQ/Ct9PxE1qWEqN8UHHt
Mw3Yc3NOt85FbNamFK9L26VZtVk3pVZMtwdgUVJanf6igjKS0zOcNx3+tnNbkRtw
nhzaE8AYWe7d0j3zNyZper0kbgJi+rdstLMR0veit1EdndYB6fFSpIvTfjGc2py5
b5ZmmpvBq92h897dbITSRaHWvW3nGzXITYzWZ1N/s8k3sydLvkCpwKXsvYcObLrC
eOl352RBGqZUTUGAdRwTf76JF23s/i8fxwtLGS6DKcmerTSZnzOHPYwyfPA7TuOB
vlFKl9BFERasG90k58LICKrTcE32Y0mjNWjRq8D7nWrciRJAm9NTlmv4J1WsbVzB
hlXLrHgfJxjk5FmG+Itti57fl58wZJBRLu+/ywLANP3En2pOqQLwf/crip4us29M
wOMLFZ5gdxmdGRy7T4hrFD1QNCvxlSFYl5E6VlnLTthSFaCSS0fYew7m6jsyF+xp
JjSfUNA1+PECUBIJpwoOQ3r9yjmvE8aIANg8DHEKkhzD18YT3cpNBXafymPZQWrL
8yC/AUVslZrdf/RE0Jg/Ngi3j1H6CBQdKWPXUW5M372fTPtB0O9YMxdGOeBZkHQg
7/daSCIqpTHketOA1w21WFw/tkzRZH0UDpXnJm17BCkvRYNafmPi4/+dK3/h2jf5
pHuWlGAl/O2I//+vlP/NMqyq5JcwNq8MG8vEpcPwt24bjXPqNLRw4zESl2kbrwBO
DmN413NYdR3DviNZ6Q1vjMa7oPG4IZRaGHpa9Sm7t2VpwOQMjhxb8McvTA+pSYXH
hdvyjsyaqaGqSNAkje8Jk/GN6thWjl9Y3DPLYhSkQPt0v5vJDD5naBcPd4OHuDMI
mW5BYgKoT9Z+WhA+DViQm3yEI5SbVbZL7dE/w9M3d0BWotAbb4Eedv6qBvkk/hGe
N5GYNIlSVYQ0ZQDbzyZSbpMNHEbdMuE6AgQctsi/Ds+OkrW1kuFXr0v2upW/7Nsf
la0FxL7AzUzCLDvxHO+kpv4hfVa7VNSu9TiJLpltkGMz53mba6I01HRJKNQovyr/
BPvsOXteXNyEwp0ytHBMRuxZJjROt0RHFa+eOKFsM01EemCanj29dn5arFMlA6Fu
nkhmPZGLP+++l+T0pNPlCSS/i82SVe1fp/SDA90boCo64ml0b/fdYTUTWyMGK+OC
GTJEVU0Ug6XnsYD/rP8cNeAFna7Z637GscyJOMFFFWTMFzPmE5N8ihUClYa3/oj9
olDmEABmeJWSCddPt7CP42rcBiUXTltwP9t20sq8OmcKN5xklXMAlZ7qoF6HXpuW
nd5gb6HWK29WJTtgns3wc6tHd9rioH0PlKMzFEdyM3dz7j4J02utsxh6Z3kQtyRX
gBZvLionW9ZIuaKgpqIboftwfXheyuyrbVY5l0LGa0Del0Tj71zk+Tjp4jzZBwJh
LTD9YU1Bwrnnghc29yOFqMbWjV6bmvDsSVjz7JElgFQ1DNazaGhvTSrUEUqAVuwC
geDH7SoaeNYSlB9PQyDWoJmHplMCFN31MmQrIxuUCXJ0xyXKhx6h8TeMradnzBrV
fMuGy+5jTKcZJvXt/aLbDnjbsBBv4Fzk2WwY4yycRawjduiI4NsOVDc3nT47R13u
uQLtbaqIJc/PuiU68niZAIStsZ+MMfdOkoysyj2LOhBut+Blw+AG+19m1Pmf9mrQ
2get5Ln4wo/AGkoT6dyU5iwUIcztAdp0v4fFqjRtXzBU6gGvUgOJBiDk6ODyyAIk
yOpWjLpwYVF2UuECWKfl8rBqiom+5kXqA0RtgJF7/RPn2xx6kGO7tI0UI0nrosa6
rDqi2kwM/oERAJ8mNq1D8bi5e70Frxtw86PTXXfAoc1n318qvvThPSYA0S3izoX6
dcSTcm6yN32a4xc2dUACJxNbRUlGwLQ4hNNwO9ZSmUQVOaOEmamKQMMvkV2isBpB
kGEJ6NynBg5Pu0OrqVL0w2/Ke12uxEAsqC6F1TDz/dFSaKk98z8eMtZscofBjGsB
e1wX7wPpwqGf74rdVpybb5pgBB0rtBwbOntOGTD7u4WqFMtZs2lKrfEkahUqZaMq
q5FmMH4lE9xRt41tJKx+GP0ael4DhOAZQZ/qXM1kd1AjCFjetMo0RTEPj5RykqmY
fh9/CJrvR4LrsfIoFQr2NC6lc2SCRDHIshHwjBVmU16RVVic9fMkpYV4Lms0oEuH
U+Ac5oO2/u3aMzQpoXYfaIf4VQIY+r5ht3OjqSETkah/Ge1rjiCjNV2euRNgYbIR
IjkYuJIjbOYTneQ5zK7+YrZ8RfM74/Cq7NzA1/czOjMokaLfUrGonIaEfNn3o74x
J74U+1BwtQe9873GSDKpGYkRNo9M4Qka1Ahn2t7gYCB3XTU+RvnrC0jQC6O87nYV
061CufMjL9gqSxzhOMdbxEwfFqEeZDjfudZbkbGFqwluza2jSY0wZv4xFWVK7PyZ
fDnO7+WH+8zm7/U3Q/jj61Py6C+7+U55qnDvgYDU8rlE/XC8mRIByS7uAfzS5yat
8C0pMAE17wTQ2q7bBZbx48zL0jCCR3zamwQoUxrh7l1ZNvy6jz3k87A1DGApIi30
MDWbMUdoWVWmVjrxO81C+KXP9vqp3oNwHHqicwXPEOdjoRqL8ZTIrhFw9s81DZXG
tmy+//EZRuiWmveB5VZzwl03ubgTo+nkkCG52wa4XfPTD3ysSWS0o1CMkgKDyT1g
wnY50hIeOuWrlEKVcgvqkJez/Cy4M27JL2abN9uzKoeEMBmk4xwq2f1RibiyI07Q
PeiKwYuVCM3e2fgwkinaEvwzdQubhWLI99eW6a0LH6cJ8EHBmZYwxYQQctKFWHHs
D+6SjIW6TLrm699Z3V1ur6YujMCzpUoOtsSv6Xf7WBZPbhw3XuBqxShJx4XMzqPt
ulm2UtV10a4Rl/BnfxN6U8Jy+1dM1KlEK3ZrtCeCFK5NUXfXrvFpKKKqnsU5ku26
p36Gzn80dh7THN0bK2e2wkyerIdW12ahP69o1nRdr9hEi9AbJ2teZvQc9sbPlSvb
bYkOCnH4jpNrZ/qZmmTpMdty7O4e74Tlo+7nmuCjwnvCFCEoK0fJJvC1yiLVUo3G
ox/ZnCBE6HfSwFYE9i0QY9w6KsUUkJVC8rhI7hLQLiWPpwXCWyyaZMn2naZdrwl/
MTZp7t0fwn+z80aBwzmDzUjjLcbnQpuUhwK/J8hKOJRRYu88MhegCB1SJbcNAmqG
A6RwptrChaiR4BVNIkFp8m0PZqX8MOMwMUVwo/w9qEqvyMlwZ1LbqXXLGxuvgWFO
k/Ty1opZfWJve/w0oghJZ/OV4VhAdsV184caSN9EcVn4kZXbzoqntWfic2F5OQhd
ziYEq8SwH5CBm5cSJrvP8LwYLTMCH4z3jR0RIxcA58jDuQnxhoVWicZQAc1BBDWl
qgW6gQ/sHF4D9UVoxKTqYYMFLujUgtbcfbiH8064Xr5gKUaMilVCK9icmYFmieqX
q+ryA5d8Wj5I6cWUDS4W440R05XqsnGvnQ/XHsipJTtgzvFyHkYqaIr0C+Dkgxnn
TBGEmTdIx54ly0c5kGm60dfm+8gEvaAvgGJE6nMStogLKfdreWm9QnVbKWbzbsPw
23XmPl4FEM9AuBcigTOdw8GUzUHjlP+fV8CZ5x25o+RHsUcDxhWzFr7d1prNfSON
bVkSxgPZySuUQgOPw4XjcKnwI8SGrOFjJWydK+coSYDCrCto+hbpNVUHuI3s+sov
rFBbOA4gr50OjjrdknXLUF/y1bIA2Stb4MF0cUV2Z4G4qNLzTJPd66G+36JN3RTC
m4dFN+ej36TzJFGIKSATGM/0xNgvZxmMXLO/47bELE8KfXRoSik7nIBztJjkbEi9
B+/V1m300qG/UKRaGfkf5w/XXWQnH1ABkXGvjWqo3VpQydzPzyHyjy2geiAHet2P
lkukHPrWxbrOuJ7V8Qa+7utcfYnZwfwT6hpsjjywZQNjVo4123svy3G40vT1N6aE
u5CooiJ5URbGTRCBWeFZW3fcsWKvmC62pZMLGx3DOlh22izPFUMJ3bepA1lnEJ8N
y8Fei6yBE3AZccki6WqcsoJHTveBpeO1CpXBKVWZHVeAMqY9vuykxCWRr77DLpQX
TgUxVbdMEyVRBR4Y2eK65WdgRyCXz/BcHsvMdfvyPI/yOzB03ax4C7vY7xG6ZILo
YWoCzwfxl64nEMjserEWlTEuA8J0JKEicw+hqkuAep9mwcRWiYATwu3/pvXoarvH
zipuBTC+MAKk2h1iceEvf7TUt1ar2bWR7negRpufAashwc6d/PPhDPtF81S8oEAQ
C7UpVWBxaDy/tTKrlX7VRyhPEfjp4Dd09zTAWgCiLJsQmVhbJiLOp3JdCPj7Y9bm
6Ltv4skN1aQGIzVVMKEFx20fP3TZ2WrrY8nvQ6zntI9+WiRn4fj6Y9SIEuS0SSgJ
JhbWJtxDJN3jsguAj9Q7QurcEhHvqb/uF3rf4NAmjmbLr/WaB92W9fH4FuLR5mUR
BOdXhYSYmJcklCh5Qssvosi+riiMx3b1wSYaW58GJ6gj1mbHl70w61UzhnARFqJx
Hr7gueCwckTCJlgPuM+F7b7TTNty2iareu97Hrg9LXhmnH7maZWo8nIhKuYlMRui
cHe8AIiWR6OQaZjboxMTvgx1p5Q6jfUkyusm0ks6lRdRit3Z89NEknjnHNMqJc2u
TfDMPms8Ux3FbIFY8eckj/e3e0oqwn34htVcBmK5gQlMwdDFSe3NzFPblgQWCG6R
EDIlIJ6iKSn9Ia/liQyUdDqyo23vBcqJChhq1PkQXg/pEoWkjx19UTxjTRJdvia4
1y7yVckDqxJl1mbGWtMIDxdtZPsyq+geOfjBEzx9G1G4nX2Jj+mSWZYje0WXFG/N
I8cwZ8GZt9eh1ZKHFZAIWBhN9HCScIOCU5yG4fYFEHlBh5RbO3JIFMbbHqqVZKSL
9m7UR7dyn9QwEwlr0xdSnlK17ElBf//w0ft2AO87oj5n0zCDjonOHaCNVdId3I48
mJ2S/Wld5g40LlGlrewkUFoCDFX12kUWvRKv40ImUDjQXsRaMVt2d2x9vgPGPFmA
vSyzV/u0OodgS5TUupdvr+iumMKigta03bbLFF1AdWpJytWNC387EDhH2zRhsspF
Y0jFY/WEFcopScl2B30qU8CRoB5Rwq+G6vofFkJ7D6sGipRHxLEtpD90Lc7a/yEx
DDedLnERzSPIJt09OdWCUapxz2NnWCYVWw9lAbrhoxMOw2FEAbq+8NhIhHGEh1Du
ykrj4TwXS8caPLBzB+JzsOc1rzbSJ8A7PQWFbpqmCplCD282jFHPqLpab0P6AxBW
wc/9Cv3ZczMXHu5BIbcYdy13ik3/2TT1dLQtsBiUkiTRIaV0ZDEwxtfEoJ8rCYcK
+HOLzKvrB3zXm39JqTrZ4S/q1Odsruy8+tvwMk9zT0kEjaeNiasIm9EiHLEiSMcL
Bf2W3vJ4uOQ+txrITza0wQxE34TswbEAtPhfm75hVPfKwMMG3QzXOIjNN7eDdXKz
BrVtrjYZDA5arwMbQX88VjMZHukHNdu+nnfXwX6fG+dsHibwlItVQrca81afxhPx
LFZAlEXPMVVfoIDrrKLA9JBhbKtknR7Bzv11+ELYVIK5jk+2gJ1qu8FaW224UIqK
iFrNgHwprxOGNQVfhtg9GvW1xSmVcWvALEDIiYWDunNB9dzLMUVidQJvaKFLGoz/
2/pKqW79fC2ohA0SKx3OkWs5TxevRt8oCZtSILla+xTDG635ISsM0b/t5vYDgtdN
OWanNltWDGECRaJUl9iEpngwx2UzwdFqZtyguJrlXTiKY7TzADf4YyeN5KPEU5+Y
BWYzV4tCgzsy56916rM2k5bAjZF311yOPOR3eP+Uj80cFWOUk9ENT8bHnBhz+V1u
dWeXGD+299NjhPD2uMGdYMf+2kM6XGERyOpFmYc/0qD9shHKnb2CrA4ojZ4hbyab
W0V5jerxHvxTb+NRdA1ec7MyQ0PsvC9w5w46h53ZSDB6UMqeB8epcAG+dzeW9P3P
znQ8I+Trb1sLeOftsGibiLnnOGr5C13X030e/7+2z7GyMMmoSmwB584gz7axWbZW
DUD4gjZYsN2/k4UArVYEhbzfshu3VLnLJSwpOVFbMszhHqbWZMuxcYszK1X57OTm
zaRO8WXVCOxg9v+ZMM7BWsmQUa0Ijcnyswl/utmLx3iX0Ca+ZY4ymSqkmzguDDvf
1lKBdlDZBYNCsT8qbiACJZ7edBq3O5Glxe+ITUns1bDtyDizNMEoqlNavw8yWqU8
mgzL+TCBTG31opvNUNMJ9g8u+mOjWwlJM0M9anr+Q9HmIna95V2/6FgsJUeKS3rq
G1l4vb9QBRjl4nCL6yUskpF+3MWGRXOu3wD7EytLTe87iwqi9Ey442fDgbEHcx3W
i3pqVghzyIPl9SlrwJqmJGNmFKZ/BM4u3e3ouNYLgbR28bC6BzcAxM+iVDWldFwa
C8buZq2nJ9kTiDN+3a/v/i26OaQKF+cxzjohFMeOAtjHM0QVr2Pudmiqoh5GQMy+
dgf0Qxw2knsW/KGubZvHoo2ovTZJTfGjoGU5nm4jSi947qawGLyszGslu1/wRctH
58XJW0UTzFSLhQV94A+5dh9jf57d/oFw1rsCWXyKhICiAyS3mfpaqB9kTOg/xMZJ
8P0PN22vu10h1cisYHCTDeCLmjqplnR1Ss1GaeVC0ad9tbzpCpDNPVXroWMByWwe
sB/K/T7+IpI1NHTf9kQZSQqS9oZ22achjinxlv9Yg27+0pZ1ynH8mBwHkTBVuKr4
ZzBhgn5Iml4NJIf7YRwboLTgS1v/jZ5OqGE2IUz0x/P2ST0Jo4bpD4sKzF5w2UpB
Ctep1g/pU5N8anFqhSOYUEQDOCXsoUNTdcNmtjf9WVb+WyHjiKInLln1rN7mO6ck
kFM3TFPrnkzUdSu63El3BFFOztjn+/avyR8omlzV58wsypVup3Nt8dGgX2PalrFQ
nbikooEaqXeMbMX1u0p1PYQEi+u0oMPMmF0XDZbKFX0H4Q9IUcRCvzEGmZMdqnAw
UVPxbtwdQzdE8/po4T8RIdoZeNI0gWdx7sJzmAPsPYqi5G8Jeb8USIQ9HhtQsDAj
91A4sfb2KTXWp3pfUXeFxjXyMm6s4zhWViXJEB3sQA0e7Ym/tYxXU5AUDR3d4ILc
3X/5LiWiOgoOF0LBGaLhayoF9tdOYC5byGtaPJEj5iBE76d4I6EX/aZjW515vr92
UXFGWiBGMBOHgDxCJO+fyZMF6vkKGHJNrimUm6qci40+LdQG516Vjdpt4owSpDvf
MtDXFCYHeZtYPv3abStXczixJqU+HT8W7+3yp1P3AfYmXhQBu0TGH6IJHuYCzT6t
xqYMFKVIHreKRHj+SYcV3bK0xyK7hY6/CyfJnVAuFEaeK2VjnYFlc4Q7pZp+znbh
YJ0ZsyL5xZlmK7wwyukw0le+lc/T3vbNtCOOSZbdTMY08eVrG8OZozcFC8XoWu0s
9djQ2nDlkHZdDMLzNRxDW1zq5vGeCR5JwEPZsjVFb0xh+vtzgn2OGP4hkYJNVGph
51HioR5B+x54Lk9BvyifS4Y29SLLNIaOJazH567Z/pzdX5VnXANx/YiPpAaf2MPz
rUm50JgO+zbmqgO4ZQTIPNBME0lQnQVdeATGzW+1+ZahOKhi/fB4qPpoUYE6VELS
HEzc6zhxQqUqmYXLE1PTU2P1zGCA5GAVgqH7ycUVP9UkON2kA/JX54//qodIaGZ5
4wJO5LREOHBvPnlD88jg6bXtQXdE7fV4BghHxl8sEjb/YqSprY1qt4dr4oTdBmXq
EuiNHeIpuWDuPItrnMnBIAvgfy4Y+9NzZU08zzb7dpGbvUWnsK8wXgKcIqnKCys7
onOI7cYa8eoBwTEZpHcEZRXreKr6g3H9N+3V0KRtu6JsvuJqt9ccuugkdOxthqds
w9XQVTbaVdwz8jIYYwo2AWrBXr6lsdLehVElkPYk4VUo/DiyVXWxnVwYMq2LCZKV
ggdxkSCDB60ce0JChr6Rsp8jE6a+RCjoLSQI4SLmwSslvO/1mFo3WoGC8xjDFHw/
HMObr9WtdORTzqHaxhwfZsGfo7A2hG6OEqKuhXQ3tFBUPqMSj9Lw+jRp/hEg9q6G
+OFVv8ECRmCzQjz8E/Pq2MWrP87oa5ulQtib78WVx2Hu8lUqtyxHXOUBgp7eHzKy
AqOR2qeE7XGGCddaO4yI4bJsCP0Bp2/a1ED5g1E5bP4mJYztEqOSHUGTSeL2tghn
FsimT03B4M1PfD4CbdvYdRvrXvHpohLecvdJSwJjD9e7GI26XMsCjENp3PijDsz2
lGF6w+t4pdmQ7yzZJQ4VZLfI8Kc2uMokEjMgDuwjZyxVc7PgjSUiQWE6lp2COCKK
uJ/AK3pdogmiKVA/7DEa605Y5SIWBi2rTIv2KDNtQqNs886CEB5n93Cs5tH8S46J
HE3eWMsSyh9Yi3/uluX7bJO6o+1Ws+S+b97bca00Mja2LyN8pzuAXlfn7dEczA0o
Qo0Zvxqbph1RogK8C2hEkpZBb2qYO8d526GrvNmenHg0mie5/ht4/Xc2qFxWOwQq
eo6teELKQCHAO9csJ2mWY3zo8IpU37FEYbFBX3M486HjQoE9W5yU2GKVytirz0Yo
mP2wrWXEdtw7Og0dFPd3hSbWuZFSddEO/Gaf0fa7iJfGvgtbWGSTr1kgjpmV17N4
uGX1fPstf1EZ0HWPZ5pnTPpdOXajcy+2hELsXnI40PZMxrdG1+3/R/STNArB7omy
AF8mQM7OXIWFKvqzLRCQEudLkkkG7AXrgDlNXMltRtAL53ChWXYuVFQLipW02OrF
g84xztM9W+cIwh0UjHjiIe/2SmZDzg0avLAAGK0jsXJ/0zpb6cCf/WqEdmg4RWcA
YTfVycx54JAvYx/aHghJjCvK1gG4sNVsVP/teuhT6bwtRWNkzOz3lLK5iVhVWlRC
k1Xwm903Zrp/IJRHhuksN5H0PqqZmRoEYJQEm9xw35O/wcbTPOe5tg3u4SJsLpD/
10jxPfzxYSi/2VyKZs/MXFdLrbQAMQhZx2VfUFNgPoMA0G1+uzQF3cLss9Pv0XCf
2BUqbkYuzWNFpjYVXJ7BY7Ok/C7WNJ2Rh5VO1WKMIHveWUVuAsEQpVQ0jXsZf+dV
I5h1lS3yRK7oTUsKrP2uAO206/btAlR0oZ9tnLH+yFgNSA08QYlUjXIr50kQS0h0
4YI/d1HFBA61GYYylSd6zfen3m8k1a/VjMLZ3NlMTU82aj+aKhKpFCJzr+Nh3jvJ
2w8vygFmCEVDUPzg1QLDZOLqueohuAgNeKUQfD90QkCxLzev5Z9fXj/27qsNQboM
c+BomkemcytsyPHCTP3WEjRPta7vbCBAEyUJHgl+xW9D13PGEwkD9LfDSsUt4+Aw
OhreMCvKMRuWGYMAkrs7nHdIXfGWAjg8DV/Y4If43HF4gxUXrBrVI+tNQ4AuroHq
mIrBaFIIAbefUktCeS8ecgkBXfQTUVW9CfpMF7UWmnTyETL4UTfiTv+nOnEVW7kq
j7d10UpUKZVQVfZBILEtwCgxOfQTrVWvf470IelV/b2v/Lc9w4ifd307rnZGOeCL
t617GQHUrDii3wr7y4Ij6o4O0XMATt/rHifJ4T1k4CPFSgzI4yntj5OMQ9V2zyKc
SgUH9INc4z8hVKkbai6+7e6OLquhC3XQEXpUNBoDiicl/ka7dobCNy0G7aRXtxth
C0/Eb9Wg8dY6lmac9jxaQCvnmjRiGSpVwFrEKuHcwhHY5KUCGskGfEo6urLtQPiN
S3kpXTqfQXvL1HyQTo///epGzChjIckGikbVAKQXsgyUF06fTnys2DnOik8YT59M
l8T7lWKrOKPvfV+YjQOM1fOQtgLEeq/fk9os4Xnuksynqb9pz6Z1oI6W1wrKT8ul
AilllpmZ417NDR8MDcJIX+SmEf0jKPj+C2d/by/aNgQYsPbfYb5g58ZuC0J4vmdE
Ng/IxY88ydMwgfMyKC44Ga7mDa+Xln/rpVOJSYS6/ORKZFXxKAAmtGa808/YHNsV
DbblnmFvV29sDbNENqtXmi609HTr3SAuFkVGmq8QBCJhVo7LYwh/+SOk8Jf2t4sZ
9UPbgeQA1GjaBAAQP/3JQ0iJEwu3nDafIX3a1eISolDk899NgC+ZWlnssfD5aEG2
3GfNbEGzV7hud+YEUAbmqh4FOGRZJcNputTDgTNPjVF7zTmrM9Df4UMgLofHBHFE
m1el/lBPegT5pg9zKrUl4HedlAggF39Oh2ipisNdc2pNkAPTiGZjwsc+KmP3yPSl
ThN6KGqa9L5YNSB5plbuiuahsmyUQFTk3R1VKKmMaqt9o6dT1K+qDqjP9CxA0Gul
7I/fTIYX0wApJt7MeScUymYv2lXe6/5DcYuXZlYe5ZM8HAnzVcQ1DoTk/uOJNhFV
MokVZbf48YdRZZtfBcU+cOeGayXs7zWeelb4Qv5LmxTXQcXCReS59HvG8fTBPRje
afIhHJSUvB/JW8JDvgVD8JYfCR9PNBeHbCFS3zQCCfRjjzzfuel6dgb9FeUpXSDu
8OJ84aZt7pbBIWxD9DYF3qMGT+LCedFFLmPWGtrUgMh10cDL32nKV2Hx6nQnkSxw
WBISEwSEVoKRPC4IXh+NtNAJdKBtD3MWgWaKNWhOMyXLn/lFUJtYHqI2dD9gxviI
iV1ihhTlYIbr2rwydCnK2SpNJmgoqpaSHyiztf8rzs3lUBsL+2Gi6j8/q8hISWgc
b6MXOkV7HMfNswCh4tU5sfVzmqHaNxeZ4M1UHpZRKjtIXbIHVu8pAeR5TZptZGwh
eWh7Th32+PwNFgCThu8+XBfudZ0T/PkzfHYAQPgz7gwHYH5d6XJS7grH5Z3X6Gn1
TT3k5LEi+1VcL+qtYwQKPxP3QmQkkueoJUi0TuTXmASbQv/yU5rPua6Zfr7c2Pa1
53TbR8eTUYlXLkTnbkARBaIDjCzA8mnlv+QUjGraW/iLPPqbmbt3fX5LFH64NXLO
j7Cfy6u6sj2dongkmmxxXjlccmoRlSb02SeFV5P9XibZ1RR6EtS/l31ftQP7mFdM
sXvcB278Lb7GjLxa7N+7GR5siGd2pYXiy8Yb/x7bBGAggR4+IxX4yZKrk+EOOIZk
RWGTd39q5TRi7eaG0X0ntYL4heJlEysPruGw4sV+528OpRXSWoEk1RJbish/aeDJ
iMXUwdJvAePtjQi/vxcfyIGhvVIoZKMmapUTde6mBL20q+LDE//O3fyfmZUOZm5U
6XzPSFhWZt5/Ws4W1GD9V+lEWy2mEdoZikOBa0O49IAYJ9mSOBEqVhQwJ0kAB5cY
+gEvlkR4enKuCNbJl/elAkCnawl1c5ZpRmc7DB8s7CwwdTF78xUSPUolTUMzkaPs
aZrfkph6mMogvsfqNkGamXRPg+leHN2Sl/eJiso7mkYjDGWxefCEY26AocgM9xpE
Z65gjLsuAC6If6Y83/WxRM5thOdJ3Lq/RZq0nfOdz2F/3XNZ6Pl1bdJiUF+++tUH
J/2g9AhfBIEmIf+CW7NIueEPNaaG7I0nyib19pADfe+uvjdRC7QCUCapfy1GTQ5d
dBf8z5tA4O6DC16o9HPVJXstwGtD4yA/PaAy0+gmi8Y8EQWUkmuiuE6GyoNjGu+i
Z2MIHZCQ3SMdtTj1pjF0ZWmDw2SSIBs5t/U0hEOjoiK6oMjpCM2twV8Gv05Q6mrA
a3eJE7AZ5ezj/SQ5TqALmQj27r0uR5s5aPr3zbW9v2DROhzmQN0N4cg21QMo4cv+
cQvPFmpdA7oa928QS7gR7t0k6sJ64d/nzfGsPV6NI3Ux84OCABkgNa+KdrwIA/gB
yDgBaW1/QDORlhcW7eRovsOPHLafQmvjqePhkxFuM+W5C7M0RkfRTU9RWl+pNVKf
BTcjrWoUlQHnKNCzpV/WuJ09PDoGgqkTPPeDHRNhphN44mqlwGWneuocMKsHIt3N
BvsVJoCQtTI4WrsA+ZuYjT3dno03ntuTunRg0EHmaQsikMInK6EOx1Hz3LlR1wvy
aUZRlnx5KXZH2T45eD0nazi4ulmkCBheCDCjjk62mGBVxDQCfnjDjKfkOzu7/FLD
3x/WdtFP1pdthP5ZybpV6oqKmrB6SGlq0jgvYQ4ZVgzfnGi0wBbbS0XjpuKe5VjB
jiAVzdIMd9bafTLHvST4y0SJBPC/+RVbXMucwLVAmDFFepJREvBACcL2A5UpPIz2
Zwn9wRyfUf/VWqpEzz9qIlIq1yhOFunklMDrasRpNmwyGb75uhQuJwE78vkXSM4V
YjGISGJO6aluh7EvzMk2aMqwV9MSBVDWOwQe3lJmSIA6R4I96SMHiA+yMC9UTFk+
aV/ZgCLYfFe4wI2zQCwaMAHnrQe+HtqMOITZrIvRQRJjVz/0hh9RNX12dN5JeKnh
ZYSze1MWbk4WWnn8OIznnZfRGux0MCbRalMeZBmZkJYTqgf3Su5YY8d0+jRc8IpC
Qfp3j934bAy0l1PPTgwkSWnttTyx7RCLjLe3uV8QOGNtuhiSlhrhaMya6PerjEm2
awQ07C+sTbd44ONFzHUCwfx7GBuQ7tfGyyDU4m9aAQPd8QlVfApq1O+fK7fh70y2
wny4CEjyq+uQzIt4XLsutMW5o/GW6zLLC6F00su3Pj0bl33aGIB/jJIoabxH94CY
WIJ5zdcUhhWulxfcF55lV5c7PbLtWFDtjThrZPSSkYWpC1JFT9xfZpa0gP4j+uGX
G3VlXC1t3Hd9imSpjIS1Tq6B6gKmDGbJ6Iq9j62e8hYMcoAT86VYWWmjKLsnOCtj
ZnDUL1XxBLyiOIAnnX+HS2v5zZNepKSXW6fy5+jOolgRapa9fkMrRwnLGAFE3HWR
iZTRI2l1QvQbEBiEmXALH1XRK6e+CpUH4FTDOm7os2ggRqfZPIn7ODUA6Lu0zMq3
KZuK4Ovr3UkNFP+M/J7IN5f83HYa3OPnyWr5GvpdoAmqlld5RZHM7DhVdbYJgn+r
b87kJBx/dVbYUzkJGcQWrXX15mggfADn3AytKUJeZlyhc+6PnxqEBuC9JMHxFaqJ
R+PWotlRbHbTUSCnjK1CfbAXMnMpCVRYCHV5QNR2L9hcauM6RQGTA/Wa4n1RCbjY
gqYH8iK2klivxFNZGVo4qacHS9Kqy2lg7i4/iWql5cZEJ6qwE1MphIojnHMs75Th
5UFYfXsvwpL/GofD5cB6MmFdQg9gPuLymCI0AJdX1nPtZTwz8Y88aol0J1FMS5Dc
9jjMbV1ixxKFGfXYT7tIL1lf5l1HfRAoi38kGULf0NgRd8fEyCtS+nrdJ8X0h9Ew
QhLgCcxcXukTKej2xKeUWZkJnSo7F0NcgU1W4inNd926VjSaD69FuEnTRzjsslJH
kbwkE4Ku+hjdXi51WdKLSwbuNpJ2BcjkeXh4b0JnB3Fd9L5iMx0xaDJsubz9j5rE
/FsnFEw6wzYy9LIh0aLloVBMyCy9e2cLy3koy7r/nHOn/SVy/jqYSfFcDMMppXoR
e7loAENMGwlssjfi+lHqClKHM4v9FRlUuYqImBQsgXmSs77KdN4pMEmc3IH+KcKk
OkKxFifQJn2VyCmQ/+dTrCseIPfBdRuB72Uqsd3wtYybAKUA5oWLEvjqTrgIRhiL
b2K5Oylg1RaC/a7aKXQJZbPA9mACVb5UIDwRE6F1i8HPFMAICoIFtPVeeUlzVxoB
QQ6JZ933+6QJwf6uEodb3jKbxIXzgKhXq8HptZNbRx/er7SsmFaIGsUUpa3gNeuV
Wmgyy+IoP/66CofP7T/fqhj+Tm5TdBwsqyWz7w7Wdkbtd5GXj8tpWpmX/dvC0Jcu
pfUQppN26x1cHzllgIi4gq1CAa798ywLiV8mIe6+nyI8UNkSy17g9P2uxG7+jnrS
PBzN4CxrzVXkBGRvJrrc9aosxq/vau8Y2u8ClS0xVzoO/x9u/Ujjge5GPcB4jVIX
0+OMMX1d5ovPMYqBbNYnA4XqzmtfZWJuLlTrRKcam09eVt7DXT92oVzAxatr/BuK
tzQl6TiUj7hNaA3kso3K1MWFDRRS6B27QuixkIlAMlDlisn71GbtVK0KXcVOa7Gp
e+RjZp9HZN2CZVvtr0/MAQnJC/mIK1ZQpgelcQEGmWfWXBcmSQRnCvkuVhij1bOP
QusB8yRuHL18aHENPdIv+uYnxLhhS5N2JMMug8rNs5nLsJB7h9HN6PBsHZiWVIE+
dIDAPsNyzq35wz2ru8VykJCJ5racX/JvZIwuPIueA3AzHikjOjD7Yx6oggiAH74/
zxNO6t6UvfwpfbqgroCvWV6NuuEybISXW72r2QODLfLQXuIZHYyT1/c8g0tk/lVu
rw+4oqkseZJMpZWNqVfgwemPdas9plEl31AgJEvYkZBh3Rfp4Zme2DfI4Mbz4nDu
dop8FfEid6lGb6dsrqOHNBLLUrrvyW0fAfd2Qgr4LFp5aByf4SHMWWd2KNsdX8Tg
lzFFGybMcLSJRcWYdYsEGbU9yme6JxzJR5RB+/anBgiVFiEeKgGDnVIjv3BfkzuI
m/2YPqN9+ZWWLP84IkUMbiNuIPTbZ2a3wjt6piNWLqLmARr+MQnV5f6EZT6Fuxde
APcSJVUAqT95ubCFW3EuMByB4oSiW08mlWFn/uYHTTjzlGH5Z054+RffmgKYolOK
tJqbxzckHERakdjEyrxaBo0cK+6qVsa959dqzvO/F5ZdhFhukxsYyy82HpH2L1QH
GO5K7EeuxynzEWRvMY+LHevZQPa3KkJwSv4M1UuX2NyEjzrM/ABixIj9fQQB9eJ6
xXmiFYC/oQTC+os119R7KM1Kq6fgd7wxQ99UK3gJrCu9UWu3Ij0N07lK4hnq5tqO
+WXh00gYIHEzVojJJiVntXTVPgSp9fSwOXdktn4hl3nNVw1ufkrfbIbYgeHYer+3
UuEj089fWsZfh7jT9MgIz1ZHfuy033xHN3h6mD75A+FQ1L84zrsvrmMGmyqbkTg3
XVWri4ZHlnU8la7qcCFzLcSGuFmHgUhO99vA78zfcSma2ZGUufvo1Z196krZncVW
cAljG84R4qhmT5s+yl5ao2rUEo11474bHmLVwF/eHaAJ0wKCjl1tTlwb3NZYu9e/
bTJMtgUac0MUkRFsodpb5bFB23kJ2CpNzdqvRsaNkiH8SGnOohzPIecny2SzDaSI
N3O0UHZ1ylfar3iuI6Sh4oL0Cs8uhhBfIlVYjjd+nVl1jLZ34uNCRlqOdOdLMT1O
HQEf3PHDaEw7pcN9xtKDH46X9XgZhVh+8iN6GCmU/d5wjyqyvG9wOmTn4u4TzVLD
pz7tn+tXki8ffhf4jxlvQLpJnCCOZR+xVvNSxGHTsSORu7qdB173Zsezcvk7QaSt
ofRSuznZ9kCQbmYy8/2+SG7vnmOvvl2J3F0kysvG9YxsLiAsEfBB/HgKkDBnxjde
AruNO7cB+Dr7zfel2km3T38igs5w9Hom2CMbd4H3OAlS3gipr6K/kNygzaL+uKLd
euQNPOD3CQPJrC9sUw/5EVrcDuE5my8nHasldeb9JgtAKFvz4gAG6Z8VZfuR2Cam
k+n9vC3z/bN2jMPE+4vyKEKC+8zZ87EBeh+oC4NSGlUfZJrjHAUkm2xjuzXzfPSf
/43KDzEyBuEId1gX6sncK2TwkKR+rPhb5IuMr2MoyaJNbsO1qb8Kvq/BrBA2Ra7e
w8NzDTdTmr56w3HHsOesgoRwXg77+VPwXsfRA36cbUytFVhktjZA5XsXeBDccLkp
IKaqUCRTALY8eiH9JuxJSd0ZKt+lsFkoyV/BWOKSNdVzaijFib1dTa3MWH1p4jZ+
x7bsFwrtgD2XBZY0+sgokAz7M6uGCuWHonXog3UOvDXzlVQBPWeep31fr8crYgRb
prmQ76bLfDbEOg9Dt65kHtvqNZdt/PgFt5piGDoQbjDuHGQPp5WxfSqZA6RxZFRP
8w1JuDvHZBd30jFvod2BqTrB3saZSaSwfI+DMzq3mulxt6ktI6QeIM0UkZj54LI8
qKnubjcVuVohtFQ4fHpcym8tZ0vh0P2uD7F74p6jbRBEPIeIzoXJPXMGm3iy6VE7
koADmI6KdqnUE9Hq0iRGC0LFSuPXGMUnhaNjV+9ieUqcpdEzuQFxARxF75aSCMXJ
7spcxdyhmktVrqC+8pwmtXBR+hmATliVJJBypSYvQWinKseJw8PIFIzweg7V+ojM
A8AgGw6IoH2dJJEifDnWUsD+seouQAYATa7i6zjnfgIv2XDDwEKXpFFX+dkRZKlT
QLzLjuJphp7lqQsIeiufKQR6ily8qmwIRBAhP4PWIjcjnL6Tv9DDcli7D/TcSHVC
ySO5RBL8jwikMHYLyZVSSyYL7FaC0WTJ7SHRrSH3A50kEeEUDDbe0sHFLVW2UdTE
4hEvDqxrdiHTZHFUGCyHiyjzLNEtnTSEEXm+U3+n3nn3fu4pjaTHKVTqs5FTN+XB
0aewRECAmygvkVrZpKKi4dMrLySwDe033XaJTo7GBusz06IA7Z9WL0GjoxPH7J5s
OaHQbpxkVB3io9YLcIOuq5Emxt3c4Xvv86leVV3GuexroDbsLZwXi0664nOkWkC8
AmQ6MMGDutRKxxyBOc67ngQyn3DDBZtVhu76juRJCnsYZfOrRLn8Ck1IvhyZTYa9
z43hajwriDOz/6YP5kV3Ph7TfEImTDIUmoEMZPXSC0WDfo+78YoMtrp2kJLpQ2QT
oBC9e7m3ZCg8GTKrOqw3f/GEWuAASt45EEbQQDnFGHb2HYx2fBqhFhz/gLB7EbHY
H8SqK+ThFwNk8PFIogluoVfqXo1siNVmjc5KjG3k4s/Os4PGO1L6bKnmYDa6kIjE
+eobnndgHkcjVjQH+Hs8Bz+D/6ClN2f0UWcR1VWwPU9ORKa4Rbt4ctZYoq402qjf
AI0rs8tkMh/2X6rpmB7wnIF74WQ03D1NS/vKlfWI6eF6kP8DJmGQAsR8bed5JClb
cjS5yneVkG84SV3JumoLKh1pj4InNmNoIK5eeiUUuaRp0RlswqrYzys6bu5RBjbw
+Wc8AW6ch/pIQ/yOkr2psq9XKHotj+GgmPofzK/kGL1fUSLJCLzgKkCqhRI4OyYw
xVrewN50iGsLDUIHzpVwqhlzjTXLABQWY+XVr6euyN3ee/pHAf4LN4Qa3hnaihP9
gk23/3qDpYhPWBdkn96TFKHuyijr4LuonrwINLxNP+VRhI+McikJTD5jV94Oso/T
`pragma protect end_protected
