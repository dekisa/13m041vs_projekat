// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:23 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JWi5lF8G4zHlESMWwfl51k7zN6eBwQKQU6tMuYZJM36AidWvMKzaSPOUxBC+/ktZ
FBpRrErO104AqrPb6cJL/7k7agIgvv1nUERsXbKIwlLHA0+2nPxMqB61X3B579E6
libJE7nlnStPvdtpLcjAE+20GMz/I28KsIijZr/Sd0M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 39552)
iKnIYy3Fmiih9pUEpylOCjnNzTBbJT94UIQo/T7eUzq/rhWVOpYbGydEPLEemC0A
mi0HXaYd/KOTC8Np0JQSVSThD6AauMi2zGwJPLxkN2FwljfGjQ6Myhb/ff4kFnEl
9Q+iKFOYHH1H6yR+D836ggI6KSqFplyxeynZA9OjlOmo5w9qFTUOwEhw+i4x1TUi
o9juslulZQFkwc937OCyDdA+CbTcK6l03a8qyC5r+COXmxhN4F4OsiwXEU9HE6FA
y+CGtO6HxOOEDbrHaneackkgckY7iNTYq07+WQ25AmetQiZpqmj044lbiPdUZRrL
AJQUMcPH+tGszEfT3uXdj3fzNHBIQNOCSN8tW3E4o0nx5FMk3i3gDdfGTha5WZoC
rONZF1Ftv20IMkSVcRynEEZXVoFE52jHgp082lTNI5fw8we1FDU+Gd95fwjy7kJ8
X4gaBE6BTsGyFd1vvFqp4nKMNd+mcpCX+PiKuZ7fZ2b6uzCf4rLyvhVOD1oEnNiL
XpzSa6r7wF5sRfe0nRl7/B3A3oXfBgtFn1XMyGZlzp/6kHdxsOXppQJKfpC+KrWY
J09oVeIfSqjlgggfXnnoIlPSeHHILe9oP4Gp7eMD9BPNwgBevg+86KOg0flOvdGT
oYoErUgJHTHnn772Zosb9GyRfV+CWSvsKzFp9t5y62ndyMq/1XMuP9Wc3oLB5kFB
UOeXF12j9X8c0rl9Geo6Wut+Vk2XSx1hjOlimV/tHCv7VnH/r2pZUsd3gToCiW3x
fQ913gjY4t9cbUG5uhqjf+AYxb02pdlJqfyQHxnekw3sNjrm8iPQTUZXpgxJtkTs
yyb2em7BoIsYNd1Uz1XBI5D4vD5Ik3M+5OCguUhhj9z6p2vZfjmBJSdGCZzy18zd
xjkaGbr3eDEpRAO2zdwRMy7OccH+ajmLx2EZxHZ1VqcDRTlOIUO5jRIszMfn0yGV
sGkAx/PLZVUOqORkwM+dmUKO6iGQcaCxJcFlF/6Pk2ZEWuIqOEMK6joAuy7k7213
rFQjj+i8HJ8midLPWgBcdj9OpqEEpLUze0um0P9GxdH8mni9KGGhw5rR0Elw1q9V
CGRCdtEAc7hkwUprS7WHnwNy5kL/q/bEVJ2LVZqLQ6lNlObY0vx1pwsOWcnYchy8
ChWwVoM7ZBTOOXiR6bRsdhHXIgc7/jGPH2CdMDf+W4NkxHLQIuxWs0VGvUrFbhmR
W+Xz+YY/nd024uKlGgFCWQrhEtWHuSvxM3kJSV1YZ6+zBdGHtGOBu4rn+aSa/fKs
LXe4fZWZStjiAUWUj52Uc894Vzja2RahJpRHL/W0uwcHbcrAMexYSAQP2Ig1/jq3
NaUtI23sRHAoIpFBkTna+ALu3kFchcBana65yThxY2+3lhduKVmtN7vhNC2b3Vot
WhTsD/pmbhogxDFhs2qvFUGnmziQ9+xpMVhg/REGlhU0cS60uThM6YtJSawaXYxo
f+PeH+mu6sLDM3AKaV2yN4OmQeLwvS703HefcyP72ZxR1PjnnR9+6RWRJygF/N8K
fcxAg6tGJvHDSttNlcgmHLbmqsDBg6VOQdnE/6yzFnFxvryS8jSkeQZ5tkamXbvI
KZVOxS5xMc9dPt9I9fDCujztUtWNtyunp8csmtHvSnTQWIz5Gn+U8bc1c25PCFeF
X/ATzJUnCz/rJusZzvs93LIMUTzW9Tch9pP6Q19xdKrIqVsUwdq2r0K00P2b185I
J3fHslnvsZMm+16DW5Koufftm1TAVpptrd3Shy+Z0Z3DiNeAbwomx+GZBonuoFiI
qnKWH3hK9jjQmR8fdOmTWHscxK/zDRDM3+HHCWCLW3+h128g4dvicdReP05YXDSN
W9F0PuxixKlGjoiWBTDp95XkU7blsctCtukwHUWzHWtQRKTtzv+a8ddRHwvCXW+f
UNVdQrsSflEOF//+vXHMSW7JOg5Ck4HwsgncE+i/MVXXgjyEBpV/oqvWqJRsA//H
b99OTpBuy08Hr0TNjKJQjKjvC7zjpjsK4TKZMps+fkQM3VP1iHY4nzyXdhQ4S80p
TB0oqKLyGFY1JjqZP1hSyneqG83NUoWOxjypySqIZc2uCOcfL8fP9MCa1qIlezIE
6cVsH0g9YmhsW9gHBiAx4yNCX0l1khTjnVSY80s0wuF1uzpkV+aqUr1+APqKAdHN
e+OMD+9vEz8/OrWn/97uLseO4zGB0k1uiis/qy5NmogCEUDZc59lXtmKSULxWjQu
+m2j9qE6O8/Pec9PaBa1uZqg90aMubVyo5cE6CRJWoBIiz6aoTZux3bpNcndOEoQ
XKiUBNJ0tx+c5QW/8eeeeKEFmqA7gfshRqm/Pv7uS0HSeNh/61ufdPU1HXJLwaog
i+rC3wse6jhY8sM37IbitOMcl5Tc+AbRVIvd2NkZqzHTn5M3KcX1wm6ACsgtsSa8
EEqcAr2AeRqxKMnFUbvNskw3GXsUxTayIHeVt/Xb6K69br1gSMCII9kPfNnPqCWc
4Q6W7SWy1m/eyZg39sNiWtoqXjPL+6leoCVHq/ub1v5xAX510akSTA2IXi2xORj4
J2Gx7SS2w+jL3TnDsI1nXpbrBMeLvKeKawVhPJ+6gOaOQ9P+Zhpvqaed6qUFhA7A
5BPIFcyelq4krgwJjmQk/cIk+TcWB+gwpT5bH4xFuFzgwSaScGfAEXaRXHiIwt7j
Ts0u14ZvrFyxd4y3PVdj91h8+EuxDE8qEOVeGCboR9Mt3EUdO/0rH3TgJjTTOq7E
4Nxoj9lrK5aP6THp6RBmlAyooaRdhJu6Wymlrtj5rcKojJOXhXqwtfLApvHrKEO8
4XT5+Ab4QC/D7UOOie8zJFpJ2Dsuy0atyThJzBBeISbiMWOZVckiUEsYKC13/qwx
3ZJeq+0t7WH3vvy5T03cNfwiYA329bCVIHEFW4kTdmCfZ8bEqiCWLFZ569DXvWBB
9yeIgEXitYN2hk97bcE3YLo+6qAlO8TR0A/8/qQy81i4yLtzKm5+zK7z9bAmgURL
IbAS8ToLfBTo1SkshaC6QT6yu9/3/4hydEdRGXcOEDncFIewhxxmkrsB4ivuinDA
szpLMiIZNk2LNED/NfHkzy9bqn1fQYeBVYUHC6VW4z/8vB8huIRI2AYT49cUJOl0
otyI/+00tB7feluMnrLPQP2P8N21aBcgGlvdPPCae6HUnUj90zeGjlNq+Dywk2Ak
m/Z3c7rwGowZcQRRqpVuSquzKtihNqRF/a6++s7wOwwxWnala3PQiH+2iNYEyxHI
lnd9pyEyrq+Znab2h4bI+H3yz43zSlEvtZexki4yz55GAlUABLwF4Ig1U3/vVoTX
6aHU05tpe4IyWFyiZUm9zujgFVf4dT1/RcJywTHuCgydbaAEnWku708uCiSBe5w0
5hbgwlpn4B8TMH7y6oOQTBiAHGV0E7z6ijV0KZSnh6KgqSgr2wLlXZItKMtrCKTt
s3GWLOECxDyOcm4CwQC4N8pLPpWb32g5N4jeFv55REjpZxS9LcJU8GgZTSch927R
aTzkab6f+4zRO0d5vYNxa4+I0vCR+LcwLNnOMIlibYGbDAwdx71hGp6pGlQ/RBJW
0sbQoa1MMDzcQbJmSaGTXZqnQ8NiIx5F1aaeSRROjqyMqw19iuQZ+DAZAGwVMy8k
d21WvfOTW+MvZec2SAlVBtaphjUNohgmhK+H7YmkVofGhoU8hIaGzti8hvV/P4wv
rcyoQg4ohqSL/wG+fzdoQ9jqE60qYZMV1LFgXt7UxeA2Q8BerDM5XupZlSDIcG37
Q+rCzwvcBIJ7Nvue1pPM5ywPaPqZGks9RAHzXZnj16pzZNnkTsqlq+moki43PEl5
WAP0kAYFmi4fYrUTyU9BlDUZ7c64FSc6XozW+JfgKDVwsF/N4k325dLcdj8i4imY
ZZlYZv0bdC+yI/ubzjbpUrRhfWGooX4mZAUIqkZzcNncboFti4VtzQQS1F3cOZCn
f9Qw314JyXNkq2zeIYKKPrKH60Dp0wMidPlDbpxlwDva8W9BFta2gQyojopKJJuQ
ofYTaTI0X7OhiEXsVS/Zg1iJq9aEFEWuSBoJwITmoTYAcEsAuhHqF+gvBl3X1um4
a9njOu2cwJ3R3Cz2cThGgCWcUVNVLVTpBrDk2FLdFe3ir4issCTwuF8GpBGmd7sx
9UMZQ6UTRortIeE3mcoqIjcExJ1bGbpU9LSrZez7/TgeHhFfdf0Y6tZ2SCvpN80e
GY9yvJk7YgWzywWm1/C45k/JJ8kjN1FEGlnOdTls4KS7hzvZ9oTK86gtZl62Zi+5
73zIFwVuhVpT9ICn7TUsU90hDytlI16HWps5/oEgI6UAOceJb+Ct3WpAnisJ6ROe
iX5J+YPSzD/lnbLN2HEMp1aUkG6TZtYY5qqe9qXJNARvsRB8bHF+L2hbww/Xhf1x
/408RUqLCqEieNrYPb12lcsCCv0jtp+u12duTefXbyEqGhH2uhYe+lPRE4KuM+zC
6MabLAlrx+YOkS6i2toTCTKleto6+jbJgZkQw6Lzs8qvHUw59sLpDxDiZHweymaO
AX+xAiNNuBwETBDZVVT7URTUIaXOXtJAw6ZrTWzGOa8xl6KsArEazgDyBWCGFGxR
AAP2c56oHTyJKuR5ZYg7kOsxJpIkkY8N2QD5BllTKbiQeTzJ+44+ROYMt/OFZz1Z
3yddFlO094za2ZFzN18E9w5m0ML6PcbufbISjMNZoo8CjJEjpl6c2GO3GpaCwBSJ
BQMLQlpGjtUcm0EXvxCWnQjY+wI+AA6Z3oO3dagJZM82qZOcUiEO0g7JW/9PexqU
KZ5vz6ONTYn6C966yoH10tCmpc4UCH4J2GTM7yrmu8xs/DV0Iicbzo/6TW0Rjcz4
U199ktxw20dg8/x9XlzQMmSFG3kpEGJEfqYHDG/nbfRy0BIkIW+TmaWjyXVAF6Bc
DswU2+7lt0Hwd97/hy85Id7E+KiXwU9nSipJ7hc9c1EHtMn5zXCiNXyGvtLgygXv
ocZHvL+fU2NpKLP1b7W7u/Hsoxa+LBOuLBDxdZkPwAEVPie/Bi2D4CgEDQ7HdABy
/36BJDQrJaMYBh/LIXYaYcTMYiSmEyxP1S71UvG1CTuvlMp1/q4tMAMIBxotApgD
s3NE3eRngxaktIoUGSwSWcKIpN/QHnXZELHDYSuq/e3wfOsDdQCIGyVppjUSYsUz
jtqvVzVAXf4EKsN8akyIBPRDKKGfLe9M0a1E13Q9jxpMtv3zawnSqAqXJoTvTmjS
T9oNXxlRyxh+/JVMb4ObPUNFt9NtnRvmvhNjA0EjsyN7tIE0PMRwaE1i+pTuTCqY
7KBi/+gN1hfE/8oInhriKOZ/AhgU9r3wWcsCliwnfgq9RiiZxQJEgj/iFjXlMLq5
8U0BS2r1gFBS8cZK3pJNidfLDB9uIYBSlv9vsFl5En49xOPxT7BMCji0+oszKshS
s0qpbxwncihRwZBLx0vCEplifMMDIvxUGGwYULej554VTWBm7pjSdKX2Nmwk/MrP
C/QIf9k9K7du5HYyXVT+Qft/DEYEbXvParlDpotCiFWv9fkAZ5zvVc1xuiN254kF
HCynuUaKnYpVizRDybk4ZZUGvNwWBhg6Qr6EPRV2YJkNwRD2vJEl0ctUPWW7b88M
1a40HYULski3uW01ZGHND8W9j0RkCzQCwez9dYQTo40KHtzszgIqsbFmeMtDsPc8
8vqruuYWv3KxfBHQokIqEOjRJVwOpLkJxFUBdhrj82bdY78g1fE+bJA8JNm60rPt
8HqJtQiyA+16DHLP2LJLerJ/FgEQLsW9ER/u+lIkDxyk3wzYsxfmJz1N8fDrnyd/
e5E1PNp3dNowi0c3VlFk05XqOQh5Dggat3KltrQIccSRA43oh8QqsiAqQCd3tlz4
flWt3TbZCohKvFxmisNkyCev1eUgN6N31MGpAZgEE65vHuxTPkp7FCewgZjV0kxC
0eIGDNIUpEd17hHHJLmFIE/0x7SkcnjEgh+BrsWvmbNtZkfAie7+iy6e5xtANo7/
7YrlO0S0zbgmP684T+foxqXPBbi2qH4Wwv5w1d402jgOsHCI3TYB3KE1Su13Uovt
U1FM3Eh4AmCvCWyw4MUmlATzB6PBxJ0AVnCKMZsBmaqCEziRmW3ywKJzt8gmEpVg
zymOzCkN+OiFZBABd5vm1833Iq7z4GphcMGQbhnJyvYiZlrfp6CbS91LuBP4mRok
nAyVI6SHYKrQ6ZiApsfmsIXkbZxAkQkF75u9PDM9fADfWd4Dg/apsGwnImvPa64N
7hZXBjvzNsyA/lGxA8f74LFAzoUj0JIO3WnZn9LdpzOsl1UHE8PLA5J06upP7l8c
7+reC/7qZKVYe/zn/LvJBuzd8ZuOj1YtY0RGK2JBT9gE9HDfEKkXd1Yw8HKIp7iz
3166+9HmHwf5z0Wzd4yFTt6geqDcnOWuPSzoyrW+Y5d9s+E76WLzZ/eN4lBAwO0O
HKzw5M8czbao2MLxSE/Zc8D298VJGZw3WZc6gkJ6BtmKR+o/fnxCetxIHJ64qt7O
eSZXNxbn6z5ZWLLc2vLoChA4CAj2YdkEQgKySmdVtpl9q+b54lUY5O/1mBE7pLZ+
ljGbXnOLTVKNpq3QhotK0ZgfZ8IwGIw6mhNg19UzJsjwbrabK0r5GII7qqUYvOLT
rrEXSq4wrv5Xn/1t2kCcQf3uC+OzOlNa4z28N+seOOCbyPFVAGfcMLLwfi68X0qs
2OJ01FYBaROjN2QW8ZroREDFOmi5AXTi1rTksCzT8nOmP5jkwatctj1/r3Q9Dc+h
904huATU3frjFJ36voRuPVKhu1AbaHY1sBFRF8cvtrQmanZjroIvhRpLBsWYyVro
P85skY3Q3bBSa/CLHF7rDWMU00H7JgNpfBg/gP7Hv55bPrysKqKvm4WIhfSlePx7
INLOjBvaE4FAoniQbqirS9sotFwMovBs64nFeoieZvA/QUkP2DZoo74l7Egnnr34
OtSrWy/MIVF+jOWWB9bwZx2qETQBdPbI/iyxCB5sCUkx+7J0WTWTEVvisg6kULpg
1fqqpvZt01/2viyy2qJEhs1l3vIDedP8IP2PzB4bVEpeeFGTWerOKAWrgobq145w
48BsrM52BFVo9IyuBO6smX0T32s++MYQOP7cnehCrVKtYg5WJYjZe3ir3+B9AoW7
kfnFbN72QnnAzNVdMGOQihkhavVgMk7P715wbfGyRfQlcj/H/RHh4NqY6wC9xxTD
Q8f/BLWqEpDyGsV8ykosuSs1g0KCZqhUmoJpy1wdIQxQYWc2I7mISwZ5EbJruKMs
tkjPGuTJivissNeioFMSlaB9h46rjDhD0AamHYjSVypm0cKDnji8unl5wLlY+1i7
bxxTraVdm9ASifOJE7/TvRiGA0JqHJGr7MEquIU7ktm29u5SsMZVm4U90n7+j+TJ
VykkIZZiOtlObevjFcdufC5WPfoNNqfd2cmSXFfsMKjQDv4UGtI9JcgZd/RziQGX
X2Aa+BNcVHu4twjHjUR8iFd/BgTD/cwGDQuUuycGwIBDm/PqW5xUYmXovMTE8Lrh
0nszq/oe03w2GCay5v/e1vwlbGO3qUDRRPvgM/RTgU93vvRWU+Wlhf/CSYHjxpE7
rtxkzmqL1SpMl3nK28pnDIy4GOVdknaQ57ysllrIJ3oBfA/dOcoWvv4eSiAVNkeY
X/Rknnd/nJMw97Cc3jfttXh+r4m0BB34bHcX2f2lwXwkec1VjOWr2DS1tT6iLctj
1vM0baNY4vWGnuhwHG1gWyXyEMA/lF2kisadEdUw09QGzI22Gr3I5IR+wjutW5Ve
bDCc4JGiR2Fso6yoqN0DZB9AnLK3bBR3TkcDnRBCvbfxF8qCXJ6giUnzCQ2lZmXV
EkrmPsMfjkiA88KXWA3afsh/XH3LtO3w3O+3vMdViBOKBlX7FaoYV9/bl92IteBp
X2IYTCZnkBGfD1Uoszs5qVfUkVcKwHh9I8ZWE8fubCBUc207GOEoVINiGiJ6Mpz5
NeYT/0dEdJVDnl4g4fQjW2I/e+/QLigh2/R4J1nIJvpIvpSPvnKMRQbLZG7V35Iw
lm9xZd6I6YU2uUc8JgYsJyzLJLutM95ga8Znche0k2BEoM4/GUK4UPLOpiG9MywE
SeI4ulYMtPcrZlAXZVJ8ZvOUUhY3y+6DQkw2d9Ksy7otDcP8YuxWPK62Xeu4gF33
WLwYd2qx2/sSwjletAp3+QskJG3Ts+GHFqSp7uwQS4f6kyCJLjIHZVfc8axjob7X
y4ASQjWPx5HRu32cb54WqtNwN3kf3TGWDWWyS43u3TRegvH3MSJRKfGOT98HXxqk
cEoaQQ8WHIOCsaBOnPeV/BvtrnRQ4psr4A0L9tdMhaqtvpH38ENOX7CzyJascnbh
ZHGclFa7cNR5y99UsZ8a0DmDFXVQziLz3SyRqdEV1H+d9R4M/KPqY+sW13H9GFPc
zbBy3XCHuHTcTGc9IluyV8q/ls+QFfPHYLFTdEJ3EFRPC9z2n4L0QhmbbnGN0iCl
sCVcTUizq5Bp9MT6F5ENAZc8gCNbutNfrrrcikZTs0Cm0PmTYN9YPGGU4rhqlhAp
gaaSWJYshIicoyT8gLAs4tVAdWn2tiFFdcG4qF/5BW4bxQ7LyDnqmW6bWOJ7b+tl
z2akLxWtSsv0lJu2hyosM7ZU/D1FbQcfZTog2hR1C6sAH8b/LW/HL+cF6/66XrkN
KnuNLU/HwPFHnz5PESUyM22D6WZDKueQR75DEbKp6wuKnCE4bu0b7WaJWhCLqucD
IV8tgK149pkdZuRRNefrjiZ4hu2Pd50gd0YoxfHW9wj72pGWqF3wpPQFKQC/Y3t7
DJXzEn/cs8moZRgyERIMatWFTSTvpe65KiXtqozv/7FnXP+zABYFqgyx9tj68Lje
MLMW4Yy9G2gBOff8vUEieHH04V4VV5x6xrmLnsEew1YBXG88pvHXPk5vVkhQmtlN
cMUptEz/ZEyBYSCsz/niRIlHD+x2iD9itLwQ/B/3nCxMPHHCfox5S6tnHt52GhwM
pHnzZpi4kBTYxir+WjvKX+WvLCf5o/6hv70biotdIAngiCLZLp51P7AWghr6dRsk
m1Z1MpGqEoCtZZc6M8r4o5wRM480fM6+ULvL/7ZTvIWPW2qtu4+51/gOTsux9cmf
qZyS4PV3/ZKPO4+NF9ra1wICbrzK+801FZVVbIEXrKUsL7MipnI70/66DRdvp3vp
alsm5O1HCuhKdFPiYps8HDTXZRvxDacwe7RNmciamVSulVC8b9QTlh1f2Oo+3xhk
Rsf2o+IwacAt3zXlguk9dmNWNY6iY6AiOILweKAyvMrvtSuMBkX6DmKgUzm5s4vg
Rg3FXXONjNiOXrmzDwtj+spC9LzjoD4Y9AvKtsAGvo7OfRnK7eG7BHW8ujrd5qgY
xSHV3SC2FoNFJfFy4XEW9YSM5XUvwkNbFwlADbFO3H90F5FodN0WcVunCwz5x44F
nEw6oX/rjiqgqg8kgVHh+yuAjmQvtgWe6dXOEqhNX08nVXBbROVwifBT0CZr72G5
RpJe08lrDcMtuyDpZTU09A7dZ8PD3UejoUbIwserfZ3cWpatnRKwUMvPraA5jgx0
PTisR4FgdFcGaBUiiouir2ELYUl8e2M074vTrvE0ariYXsAA6L1y1X184jEXimGQ
MhI9Iy6NiEklkn5JvblFliQRi7ROaRz/E4sKoMhbiL2iXHkA+5AY2D6LEUKevpIN
ADCChbyHu5It669a6ytbh3v+gAqPyvSwcM66hcuLFh3PGg0CFYDGzU36k/X0M2Xr
Yl/K4P82c2xmVQa+subSpFui2bkvBoXOc3Ze1GvmT7heXL2/IerS0DH/do5Qjb/H
2oWGXySz1wOLH09f1O9ti5kl1XoS4yV5U91pfei90st/PfxlZtPW8lY5jRGimz6B
eKdyn4gbmm1IPwm1NyC7mP6WHa82AwVfV/cqj1us9HmZj1tGwM/nDsqITB9jRrCw
lonEXxkDwQAVK2di1PzLMl5M2VX4z8tP8CbN18QY20ri3tPmJOvoOtn5O7XLp+MS
TpLYW8fFLutwIxW/csoOHSfhRVVV5ZFDV+LDbeeXW7oqeT8xijrXVssgPXZUGBFn
+qBOFHCaDEwie3L4lmDpRsh9wC3lVYC7b9viduksDiIBkkjkU3ihuBBEyyBNowkY
AxFMR4QoDkhhmDC6lo+Clh+vL3WPEcvEsk0aiuXgtYYitbIeXiS4tAMee06q5mwV
gHJ+zKVlvdHNyd1bIhTVCzdM6l/N+VI6oYudxHkv4Bw55FvFY0WVxmItY7vs7ipo
3zampYZ8B69wKgoo+9VGE7HuTW93Rfm+ZB5XHVSWbitEq9GhzoSyUYQRHXANGq2K
6NubkQYHw42Te8t4UE6j0fQUvGXXYUP29tD1FEpkHjGqg3uPjOfQVrpkO74USnBr
dhOwwncXcrIG211lQUclVE1Ve7xQGOF9IHurGz5+1foP7nGI2vjuneW2ANYc+NC3
uYQ+B8fFnm0gbUZM1M3JCq2f57vN1g5L0hbOqfvyFId5/5YJRaHNKKo5OdoXxuIC
AdVlIEiy+LeedXFitrUhQeC3gKbFJu1AP+OzVa6CKZ/tv4gNvEX2f/h26w+RkwGb
4sMJ411lXaCjBoygDCaBaLGbSWvufEs8W8EjTVRU9FnCS+HB3bn9lqxTrILaPzfi
jJnAzUYNuwkFBlvr3MFH/h7zfH/ZMgiTse+zhxl8vrq0tkCCUvzEob3Bi3JBwXZ7
OWqNRxfoP/Htuq/byi0WtAolKJ6u/u4pnb26N2KhGrSwv3wt7UJqeyZgvtf/V7Ln
ymQiQbAg4GcSsE7MwgO4kdYo6PODS5k4U1L1gC4Fp/UfzkkkiWybFOy5YE1Unr9P
ghpvNnu9sQYtCHtnNUjCW2nPML8ZoujC4GvYHQdVm2gel/TkcITOwu+9yf7Ic02H
zuTUpalOgqZ6VyYgBIlNmOqhtZHk9TihcQj3Uh8A7nw5u+uK/nd/dCQr9jMKoFvJ
OmbL0QhQVN2Eu7wXqRDTR2VhfQa3muQXDaExYq6OjzMkOqfSN5NxTISKWrG0Syj8
lfz2o80TMNDB3zU1N8YGi7wOruCfH65JBcSXLPBiG5pzbQLlO3oello6D0Bm8X+C
5EYSNxQA5ZuStEtHdqY1QglP7LrUzPvG1BjJfSfRJ4DJdrATk9f3dvPFMJMffQFq
tOCfMJJutTh2lmhFDuaFsj+kcd4k2J67dZ/yXnNPNcO0A0WI3/IJ/+FazJx1nhde
tX8A2UsD3f6BW/yww5QzYNGz3Xz1mwfkXQ9frU5afHyZdJnf6GKS+Myq1Symxw5B
5qz+WdqRbdZaWThjk6NY+BQf3Q7aBI1sLFKABzjog3CxOQIjHzs9fTrdxb9Mnres
UTx1rl2bsnYKrXf17H7JEhaQcimbhJS82hMGlICZPMP62rcndkr9I7kipPY9/Oa9
KX2phE1k3i72ZJSkchIp88e/Mrad9otnmkGt7hngq/Karlxxboe3BVhJbWQJVW84
EVti1Mf21/7/SFRnbyh+nHIvQz3zJr6PkBfjwP3U2Ed5SQ+SaRKhXrl5Uf8zrdnO
qG/woFksBy2pQiroQPYxbvuOfekvZ/QXHT0kRjdVeF7lzHfSN/GhTG6PN8A3q27T
5NEoX+kGAWvEdQaobWhTB7WqGHIWMaHmc1uYTW7PlXRxksXrV902T+TZANKsDoM4
rHUCSWzGTEtpI1oejZS0/NZjC/JZM4IA5Os/KZTck8rIU/OMjuPY/FaV4lFHVl4j
rDTLlBZifGeMXVwDp/X9bn7667AjQT+xj/j916K8uwnVav5UgjZlLQwy1pezj75a
UrogfwdYwDL67eubTzcB8jREzPxGbpFc2kscFrVwI4LwMMMCSswyW6zO9/G5+iXk
DI1qxurUMwKyFiMp/r65vfAoWETi4q1HXaKgIYZkSLDg0PVnsEJgYDOku2uSGEPk
P7MwpH9/F1R60teugRRBq78/GXreC8dDbgIZXmViqm+k/9Ag+Q4mtHb0+vZU5vci
q3PVyFTG68wZP/hoNMqbshWMCIeC+1KN04sZSxXEmBedYN0mHEoyvM+t467Bm7CC
jppuQgwFyhG3VCU1vRQx42W701HUmC9DKLDc4tqbaQXa7fa2ene3xN7gKtJYCWPm
Mj9bYrmUA4EJ4PLIvL2BviLcsQsuSGyBqZs/4eO/18GfSsvO24lPJo9h4CVDpyKH
dSOfZlWGXOi6UbMZadlcYpE+5mkwsJahTt656H8OxwYKxyrEmC5gUFPHafacFEz5
CvPnzTcJN2NKgY4rwGuOyOd9mjkT8CLRWdwQNJ04ZwVWbiYe+x9Y3AOEeeAsPhbB
4ljcRkwJ6cUr+pXfILHBO5Z/XKsw8a1DZXOOmJqVYXhrUa3XNnKArQj4jeiDiGj2
/U27qFy8N8r95nA5ryLnnEaIOrMvSuDWJPGQjYHiq4wwEY0CfPFoeJJ9UXcBskQW
ehKKkwQ3XLPMQLH83LM2Ylsv6bPrEKSkoGVqNbnAebFhHCE3qsI2aWdRQuIc0L0x
TABlp8iwcBhp3CLIoU+imR8dD6sqaKyi8OuBjt38uj+Kgv6nFbLWfgnlKFLaluUr
i3btuupqovbNt8JgQx053VYLsVVtYyu3wr+/C5IYNG9XYuptLOznx4tBVsnb4yi8
uRDzJlk13M/9G8RObvF80M3QqzAuLE8tzhgJTstIq3xZJaFsb060UrZ3V4Ovvcih
1+x3LeZsIoQ+iVArkAnNxtLqQ0I/Rp4nCpNlZT/WT/EL6XzqLUdE5uKCSLM5cvxe
R2DmNzxslIUfCa6g0Cgk6Ob7rhS5LfAUXdH/x09ygDvVRDaTWUThWPxZbUUvLrNW
silpRuj0S9pfVKO38CMnLPOfYWNyEXeU/olLGmsLIfBOgFyAWhCEbmFYGyrNMWcT
q3NFMl/s1PqSKtRaCUijb55tkKaHLtWnH+sCttPJGXh3ug116Ix1aVzca6wEgmvG
EwW5g97fpd0HeoFIFhdgdsT4TSSJt+SsiIi3wN6/DmEymKeF9L5eCoV7oN1jzU0r
E0zytJJ2Cs8Xx5DUFl2MwSYLNwkn+g7MDvjgCwcZttCZdLP0aEaaJmWaZu5bmMyX
6dNIyw/2cAjgli7UFudT8Fp0TCw5mJgi55M0CaFkvc1hwPw4pqpuBsk5Dis/7Ri5
/b3voNYBnSHr/lVmIDnxQbw5SELQvbN+6uDrlg5AktmpvJr9bOaPviorKm7FFpBv
OcAntwCRfVzttmZTsZEtUNgbREGoQZBp2jLDeh/u88S3iQjMhc1eoPz40/+v3KtA
YiCUXuicF1QYE1QCfYQU/KL+Uh5g/IzIJa9r8TPIGIOfHSuCPXWAGwI5kE284o80
OVZTx0P0nP3WNkF8Q9Kp4yYJnuMfdt5UQ28hHhLKW0nVBX+gaMjuPGQr6Lit1zrm
oReFxwR9l4c4+OQIbPQBC/iFX2fJoZRXMg4cVRvgHroHdtBCQaNPtURXHoH0TZZp
HFW3u6+OiyQ8QlDIQ3pDKpZNPV7hngRV9N1EP/5MkBBSHEoMDS2MnEaAhYo+PdiX
rxjpw/3YurbTu76Ojo3FHTriB+1a8aLGNq2rLyLmy8jZXQLPLgkcJJKtYITxcGVC
D9fO659KYhVtbIbzelt1SVbqAPMn+ZhyFwCowN+0o5y9zHQGXjccdxCR6pKX4SiT
PaHE1GTaQjGirYG/++cipQmZKZXaAI9W5uexaDXnnJlTQtEGfyTE6dzjFC27Z5sU
NF56yzYhB5qI2snfaku2NTNfK2YBMTFs5zRQ0lwguu+JzUEfh1XuzIlori1/njfa
BBZpjtbhC0Rg5Cd4yNaNMqt/BohQNP7woZXcmv4PwO6ehDXqMxIggbaqPae5HzBM
OfgBIUgt3lr47a+Do7BBAvXoKuIWBS1VEXYpbF384fGf/fWSezyhJrMLkFwLl+jX
6MmTKXQA4GKVQbK7ARk3Zm8h2ROCCk1Gn8mqa65/ZtY6lSV5tkB6LvhduJWzQzV1
uJIXDdSxqAOk4ljs/p4G8KtObg4n1QLanlrEfPzJDkyVrMpM3HaErIziuL/5gjf4
22+sqLfv2c4+9cYHDVTXqvTJJlIKQdi3yGCaHUUDwTeeIZxL0eodAH4DgIWHy8ce
zVvRlsXB6t7S0CBkUlvSokWxocT+Phdr/bZC+V0Rb59L7ethyzDza9CrYyVfzJA8
mvU3WdJPKLnCnAxrwSKvoSRGAdWSh8QLOpsLJ24rzYxCCUphjKXd7oYsyJF+eJnS
Co4PNA+LlySqEMv8CxXhHh0QQ7Fbp//6JQer7NkvnD0oJXUx2uERr5riW2XQt5v4
c1fyQvbqUS20G7ukBizMP5L9J+YaoyQc0KoUdfBXpwhAS8tXqRViJZY+Oh5UF7pc
QSTYXxeaQHLJirX5sApdOhL/bdEbucUASqjC78cx6umRDTuLnamxUgKJuH+GpIHx
kcGPbMfR0mh4McqMmX9HAjUPFFIgY5M2wSQPggjSSSn33n3hqBhQppnvElII3FeR
do6bzscLJ1B0jHXCheNRb6UyMfaA3KbuRKGIxaPKS4YQ31/vnwlK226eKzLoZ966
uGOVKhMvix4CWoJWYu5WjTbUHY09z1/aM4KmdP0fvdKek5QSQdQOPX2X8mReY9zZ
TfQLLw2R35F7YcS9ryHtTZhUb6puXoKOtsMSEABcMEFAUCvhsdEbGkwjDzm7XdHM
qJJEuy9QTYCmg2Zcee6dl4By5dQYb/6VROFZO8kdgXyMfEv7owrQFasd5GdaAVKZ
jyuseVTVMQXGX8hFByybTKZxplijYMT67SGXOssJzuhU4w8K/3CWxnNJ2xMz9yUq
mJRRKsHWsoAKZmOSpLXChvdWlJspVzd03FoLZNIjN0b0TnZyc2hvKLRVtizA6BvY
BdQ2otpnLidlQiUQpOF4u0Z26CfL6tPQbfBXJyIqIGH1ZWeF3F5gY041sQrXbOgU
meh1Bt4KrA1skG00r9/BeZ+ndhMQVMlQfaKf5EChht2dNntXS6NcCeza2RZxNhCY
EFQuuGucMB+9b1yrQ5ujwlpdot4V0FU+aqSJz2Xo+NLwXyidjRDZientxC58reXs
0rRcKZPJcPRobraKO993SxPzyE3RK7+WENLWrr2OSE6ptOXihNyNZMqFsgNnktZc
l7Ov7r23GEkVU9Cmw8rzOw0cuNdyMbGW3E++6JGb1ZPrhf3n7xlzrc9sjV0lrkNA
Sg8ztEkRnYweDmacAxsoDUqVWdEyvR3Jmutpy0+Ymbx/HHAL500cwiJTk8Yl2PS6
KZ6evaF0XxVzI1s8UexukeTJ/qkzPFTGpSgmIsxYVfKDfNfT33scgHI23iP07Tde
0diYVIaznuBLVlz7qxDsAqujBU8dffizoeuOVwZZYB+FKrP/HdYlw77QQA8fBCcO
mE6YEw6NvCtVqUdzcExlxZSScAwOsnqYztL2HW/K3wJtm3m2WvV6Kyca57ziR9FK
HeKKVF2f062Ec38pDruUo75hhwWrvNTHLQagyJlrtrP6ufgqe1F0ZM5MotMU+Dwa
JxhRVJBZP/NJ1/1TsNDnQxmttev5Fg7rQ/rXARmY9bdq+5O+yICx6I7vZVdivAXR
0WvslgIgkD89WYfgcgT68cEeoYgrQK8pn+x2UBQ2SwVo+QpmmhTS8zwyYyJ57N/+
RASIKMao6UibyRCaPmXhaARn9kEL9TsqOAbLOL3QqOr9AwmbpXPFQZroNCEmR32J
5hO//8++FuYtSnuX8vfmLkx5eoUu+OhtQgKifNFG8PzEvdhQBpQcfPpFnIZel7QZ
EyT017jX48aecGecNcbVTJ7ApAbdmjgs97+eeRi42Ep4aC/IibcH25ndrBv6nIG1
6aZjf1fI1Rmw4phk2iQW9vcWonbvjYurv/bPDXIFORbM8jMmYreSxX9I45NsoYQD
2e0ict8VHnQcrKUjfjf2Lv31VPwwzJgCUOj1mVduIjjeiD+1gQWxWkq/Ej+hWZJg
dDQ1MDgOcCwIrE7B05gaAqcZSWyHsOV/2lj30rNLprS3rN40Ztyb5Tec/B0BXAHh
Lyd4vJzF1UKkFoNc/+pYuT2uGk3eQoK8Dub1O6CcWRRsRR1vkcfE8FPxLCNZRXkh
rH3nCwlkLF2aWwWbJs3WRgTBRDKgcTihnWUw+F9uI0NddkgXeYEbtflPQR2EXsNS
j/EIzsB0Ngjh44WB2NMYq1rddH/5FNwnpfjnjrHf7O5m8q4bOl7IWJapVbkU2/RS
6mQ7YOf6F3xvNWy64XgfsdJiqku2DHemjYxZdnvHBoticgbaeMFYm1wx+gIfCh11
CYtOxw4CcSSUCxhy0qIHXXOHGHKwqg8iPM74TCvAJ9X0PbcCcFROGnOMg2MRR68j
JPXP1kum7KizAr7z+tGFi3kwEDo1jMyuevwVSEEZGf6pJ5J9h3X6vNFvdp5yZzAb
Du7DMCddQeFE8fqgCge7tQzNWkinckZ+45FgrIroy9nmqmMVR3ZcyFat/WDakEj2
rbbz/5v/b4ckB035BJox+uY0e80NFjtRcF3HhmEju9hQeKfq54cqiE1UBNkAFX3/
OoxmBSgVQLm1Pv5z2KCUmOIuM9foBAxwZwl5UlOTuRzwsCw2iNRMh4egOctJ4kCs
J1nGkvMf/XxUfBI8Heo+T7Msg1vWRQCPFwCjM1gR2cWXpSr0znlV2FF7Als3FZAH
4ASm6WXuUBnQRYFeV0M1xJq9zpJ5WfIYX4JeaK73tlLCME2tIBhAajheQzk+5B2O
ZYrCwZktav9A67D4jFgQHIPFxKYM85m+KiEyRHUiz+gXTqkDrgH4THbbpW6DxAT0
YysB6Es2y+aooDsB3tw1EzVoSKjBSq4PKLmU6sAzPfdXVGGECrzKx8DTKHccfuCr
iX09bnim9vPYLOWA3p7h76H7O59D6gnuf61m+YTVwPQhvDRPz8tfoLEffyxuPgJU
yb8fD0bQ3GwUYrc6e3ruVPtc1Ssq7d3TknnZW1v7oaOKllE5h1fHEZ268GGGk/cx
fhcvn/Putpa+Q+T5IpWdnX/IIqmiiKuN9tzHv3W1yBxs7h90SJVyJ07ChNwISAsO
M8CaqJBqHZ24CQvqibA8P37Osju1Q87RwQdnkNxUlaIM0PfUZ50u1RIWyMqEyIRP
hopC8EwJFNL8gNl1fH7vU8GbvQqIa8ra6oeeJ1FYokLpZ6yt2Jx2dR7uo4yu6S1t
wa6XO6fItd5G+Kya5L2JY7SkIurOdJTeqiiet/GsxFqsegFULh7l/R2OjNX1cd9i
HJ/l/hOCzr0qvJFA/Q13RxofnfzMeijThYnyXhXB+9fUtPA0dsQUGNa7bfXEsRKL
RT1qH0Wt31/sWzDI9RnFqZf8U8w+W2/3iKBponE6wlfQvn9pKqGNmdwCFS6AFQvQ
SL8wbekXWV7SQQWR/hPJDph8ryP1ANXYv/VSzkeefd1BKnYfdZ14Oc0o5N8YQC4D
hXNorGdJ2RdZjE+SP1Rz74siRIJhloE0wLsKDK/v2Wv+3LrDcCubqKQuAM6jFIgZ
/GQVgMEE8f51Fn++kIGwuw+Zlg7/CI9trbEpnSQRvKNWgGw1EKhi9Gzlk4MJBhQm
+a44wB0VUIiPLrEyA0g7J+5GEjtqlw/NKmHBFuquhLdKlNjOnlPHyNakqgyXIZoB
/WwFhL5V6/wyeOEQDwXRJWfkN+z4fS4JN6+MzqqIC4AGn7qNLIOBY3oSSRriAZAY
szE798zHm/FerzxljWEaAAa8L9oDzHvQd91Gb5miGDDW2Bxiz7bgy/OO2RQb/mnt
ZtiqZfYbAa6NmiBNoloqjE3HSgv8eYcLU567Z5dY1yEqa/3mTp1AXWPUsKyHO3nR
Yj1aHFiVMErXGzw9OTWEPHCrZRZ/ICEH3aI4AgJVAiIl8BAsNcJLTTOMYjxg77eb
i5RpV7YubaDmJnSif5t7K9r5qpeP9YZ28MRqxSPGca3OSjThriTJzuabedhxnECf
/YxXtqdI0jJQ6pxag6UF82g1REp+bbq8rrqBlmJecvlGcqD1ZD1IwJETQZYWVtdr
uXImaBa79s5YSiRxf8QLu/lup3KrsKwk8e9qJ/UWU1MuKSn2MJ05DUX+Pr7hp5Qq
UENzyi5dGu9/cwDXjd7ho70TQRqQK88kjbK3Dymv37GHelrV+EZGbh9u0SctUc5P
N37YeiHPmyfPXgoa1leUiEPc2SbL605/K+Gm+Wz3j19uQKk5iKnIBuE8zlrZDDNJ
QUpg7HbDVYchTiVi0mmfpEWdFLDgQnunjsiMGQzRRInoCW+xDcByHfzHrjeBHUCo
NR3b8n6QCLVvrpAAv8zAd8+F0BZsDXE8/hvw+KEJhD3+O5pdylhllQTxx5XmVytT
nMD2iqfwe97GisYCfA6UM5cmjPuIab4nYpL5s4hT4woVGkIG7iTz8lv3ZxUo9S4x
wvJNol+MYyh2bVrhFGsdn4eVzMUFennAcFRSMabfNMFJe1xl3H5233IIHZb2rAzD
zTjWhdlJmKheSSAadpTLmT1SxzcgK6T1RrBbkGjwo4NXpIc8jCqeldyxyDQm9IVm
26X8ztqqmP0hHCoQDiq2c9qDsJud4gagCMPwcZCMH46VYktYTS+8MtixIBLGbatp
uqCq94ikBqeWZ+JbTTWt+lfrVzBqh433FKgcMwdIyTirD0fDZM9vFj6MM8zGzKCj
i9HrNZ9soK6BHP77UDurRpRDbI5aEdkPrfPxvkK1muSJSOFBK8H3tu3NhGVaAyon
Z1t5XLqqfS4M0+X50pqb8MdKi7SGRnSKsy9w4ZMoiwvKQsAvIxkkOzu6K0c0Bms+
nwUqjKwa5E/XRD/pxqBR9sIN0JzUffu+e3zUXlaq1QIEa/guhQZ8xLeYFrXTa0rA
aGsi/bPOJLoPrmU3mfoIJWs6NKrXkTtS5I47yvp88ljIY/d6+uAo/u9ofNVtCwRh
0UVtEItsvWYXGkgB5IyQoELbUj0ZTL/WmBk2mnEPckRzYAeoESunPEPmIbnu//r+
ThjV978VFwE5EKBHj9KgEjM6x/prduc1Y4tcgJALQKABM046NSFRwfRisa1lR6NR
sBj5TmASn8Vos/SKR56U91UPuYwnaJmK0Bn7CfzKrUnhGrDvDgo7j3xTob8839B4
axS9jif8Zm4dpnOS4fCdcDkK9EKy9B+GZT8gu3os4J30F/gcVMc2AWTFuskWVz39
TBvUafugRnSYiyyee4+9G7P6HJFUH4c5GBNsApJcRbJHZx4KbA+QZgDP82Bumuay
j08LL4S8Ntjc8OStEE6QvFtfC2DCKTJs9FBy5mSriuZwAcAwHh+Xk3aohRH8ddvq
EoamJzYrJgGGXjyy0ogVyC1niMOrKNmRlZJ2+Z5I0ab3nDNJgS/+eoSDtOEK51hO
TQYDNGFfiupMmEPVu+BdCBUZ7foPf7MxYDGDc++aeS0qipt3V0FAsxa2tSfABFeY
VsAjzwIp6XXboPHZLelUNH8F2nTCYUcS5dzHNmhYnyR9vZ2L312IOCrnVOSba7EO
8gUfaEs1GEg+nwAqUy+2nbJAs2fkbTsBFXzlcCGVGdmOatvum0hddQS6H2gCcGw7
ss0QnEQ+EuWcvhkW2D5iKeFEi67IrJ+RYOfZUzozVtMUOys/08xkQ665WRrw8+GP
wEjErEHGoCdbjpHpczlJgaHfcrjqVUepnhiJSE8JlhHMC5qlWKj9tWDbNU9nuPQZ
GPlmb+aYKxqFcRievGSODD5yeAiNTAKVzuRG2Sz+jahrV9Aqv1iuH/yu5EIKU/lh
pC9ZHiAR8qREUcCh75f9u6fRj8TTgDexG/jR680gcEdenvgA17e1ffy3y0ywwz6j
9aoHhwo2x+3gryR6XkOoApq2s2PLjYAxkFKN8GwVurZ0duGa01hNxVFpFBFl33Z0
anae+ruboHnirnpycVkoa5ytRAQOKiR03txClzJY7ce9ykvorDomeSzKwiQ8Gb65
qSKp1/kmJIQDdlmqzQ60X73+c7G7bmnDrUwmQnsZTOIv/nB5K2i5ViozbhrBSNFV
JViOOSQGGnylJm6Y33rKDR+Gn70XXN1OBgvbNqt6K/0jNBo6tDW/W42B9G9yrLJy
IJbGWYsqLgAFJc430ee5g47T9XUsmsr7si1HP/C57Hi9yk9xtg3jSkH/SzFDPjpg
JIftVPdQM4S1aKbh55fMDb+fZjh16pTs/N/XQ+OMCMJu5nJdJ6HCjMHIdwZc45Lw
U1/Vwj830JiRosoUW4PylKMCYdinPdiw4hNBb1EODgeveyuycNDy/gfZ4gS2BAYE
JgU3IQhJ1BJN6yvhv2E4w6yWWEBC9e4uN3/H8qxLIUWLTgo0YaUjHBvajozz2/H5
bgnSasLfT2umLcbnKnJBLQOBUaTqtVDFt8dRaAYLznOEUb2Jiu/QhLnKY72S4rLt
bUNOyLXFRvrQc+Kg6C19sRZZ/ekqkdO5vkcpIzOdhtOp5ew6YRaogzjrWVsOl4ID
b126NgASVzkUClzvwp5X1IolQg/N8/QAIvqhAU6e+HM+uYJkd5vucl7hJqCGxWRY
0rqXd3XNc0F/D74KXQanXPSxoHDMqMaOrX+SFcgREwhnZ4gmfGE6OG1yno4Fadnp
hfX6y3HEamxu/15uFqVIpKxHE69FzKzI7QSbhrPUIyncudwJIsAag0ghVjWCej0q
Ai9fOHv3v+fxYssLpnoRvVkHIEZe77nuleSriz+rVerZYtJ7XgZm90CESedU18q/
g2VdA4NLRHEoXrWKPl7tlYoUiIC+U0YA8aVuj3Bb7DGXCRtsObzBag3SEPKkG2UU
DUKH494VLGsSdZH2m4SwAhFshrd/bROYUXFbv8xosgS0LJ/OhfhgzXm0hXAtPc+T
kmKoe2IZhA2LVoWbDRX7swfG8gjPRVqydMX85uznZfnIRUSnPdYx8c0aOt7klAiR
UlDVLuiPloNqo9sSHZ2jIDZpfbkKGWQpvirptWNI6Z21dfNF1fsx15cxrHpXl0p7
Zdp+rbssX1GxuHpZc+/B03Qklqujy56bDQSqjTIwks4MLmAZvKFc3WRCqAvuNVWO
Z6mmcHsslZU3nimtH5bbcpestW6v1JPwJo3npZrOf5nizqBZ/awkbUDN7riZZvz+
vkivsMsp/m0Ij4EwTwDFZV1O3s9cul6kgqdQFCfRJ7h/GaiyjqEfWwt4uNekxYuh
c1LuQ2Q1zhO2Zw2cPpqZpn9/JAfQR5Gg4nmpLrq3DGbR82qWqUeH+kby0Ub20wzj
sipP2O3HPpO2QHYnzny1fHnp0wetPhBwF3Z6mCvyE1UQejaNTuY8ZMHW1eV5/Jj2
DbvY3Q6vzCBcehURMLpdgAWa8gubvGpwi5PEGzsI+1k9Uik1PvZ7fNqozpOF8Q4b
7h2wYCXfx0Ggg/ruCLxxTIqeRNzCAWhjXxbGEsbyuMi5J+vceJsaZ8D0G7y04zzl
D2b/wV8pIaTDZxaztesHCWH3kaXhwr1ArOdudtzSMwgji4T5R+vkmQhLG8pVRUhs
vsz1KFytaLrjM5TcV/i9OYqnUZCja/H8Lw99drm2+0fdSQqw3/aAdSKXUCKtgmR7
GrU26l+IcNf7D+LRfiZ0QxoGX5hEdcTlf5mjKxSRmpzYlpNRsEJWtXOey2728AwN
+Zw3GcIofL/KiiFesquVl76pX8QdBY9+UlfYTqWp1zP4QkWQyCpsdXYS2w14YFkg
WjMq65m61AduZkwb0cifjzvWEHrUSFZY95AHuwJunmzLliRwqFC+R4uKFyuIHxlE
vtrLtk6vASyg5ihaGSeRdnfxF49BCJ2gGe/tJQX9lG8POkFB5jeRKlTCEyzW9p9E
+n8dABEuQrmNkynM00BWUCtFGqNQXnUh8U9ltn2yb90VQNhAgn3ZTv9eTas/cHr+
Z3OpKGcozlIA5/GE/bX8NZCNFpUtkKsMEvTXjFwnSJ/AbAOLM5rvePJha84+xvjy
X0cUQmvyLOHqdhn/PdDoyLtdKx6poKxj6Qq+A1oD+mSaSLisOZdxWTFVT6YXOxt1
7UezL5U4L/8u7zTE+8FBWRf9Y6/j1BjpOrEPm8N6yNe0U/3GwR3cd0J+StMaYLLk
tqKRtxpXCsbPx1gm80i2ujXK0Hfnrm1xvhMGmZeCm/lY8RmBdCeYh0znA3M9pkF3
Sxz+0GbhLEWfGBUGOkcw2+sM1I0VuddJbGJNmFyfw4670JiTNNG+WrUwSsULrqE2
BBmlvcGQz9evg1kOxdnAnQYuKtVHllh+jFhz3kTcf97jDnsK3riG97ImJ8HzRHTv
qBvXj4RV6Up/SEUbgCYLPY1/Uz8zBrvglkm/Kopo8Z8KPy9Nb+uF5Kxc1gn6GTyv
4WxgToahUr0NoUmEOPq8i81JV80Mre4Dx3l9xzzD0BjGvrNfn+LcyGerWQZYEfoo
9BO/NeKw/mx5hiMF501wg/1ONm7TUVBePmeDviRqWIzmztnCV+404c4UOIO3OEwi
yzHRCZPXLlrp8eecbz/A1qDcMVsoySiUuvsA0D7ffvcMRF3Z5cPHJiQpPKzrA11K
fXohkoYzJTWiSgXGtXCF4xjO+m6cqdPVt2MtP2eC49cTAlyU/XHWuE5tNSZU89my
5gA+O4wan5oGKahosVT18vJc4XmLuLGs0tPxBibqjQ6FqBOoDkWVSQSdxPlQ7rWP
lmGCDvtSwliwA7jLP5wnEjErf+teGG40UVjaIMRtCXUd/6IticqE9vQUiJZvSNKx
V2gwoYyW64lpZqFJ7PJIwm0XGQsslKCZ7gNKEZw/QhHVjPKx7v0yxdOU+kR+dO8v
w+YDvD26as+QLezrJlrWq2Q9XICBv07kK329riRG3Gq91MFEV/ZAC3NOu2vsjZa2
7foPlDwwo7JzH5dPduVozg8VcL61f6a4EfzKJdBjDsABD39afP8x4BcrB5Zo6yKv
SOl/nLjn0kV3/cBVUxiLa1waJiaUbfD7cj9JtJXHMM9DN9/C3N7oUJR1zHODoLzQ
eWzGgQBToXXBefwITPOGtm72W3ZqtHejm71kKpsaOQ7cNL7kIBJ+QG1XEa+jh3S1
AsLAxSCm4Qx7mghjl1OxHmpIpUMM+dv1vEq2IVEigf5bxZzcgToPAKoktvXWH6ts
rCXpdBDSZfgabTsEDDEN8XncM3IrztNZCxrt9YMIIHUZKUBvv/s8fEsHVouBKnZP
5swcT04SuiHynurlWvLpAYhdUbksO3Wgf58XHAOjbCbKvZnWrqkO5ys83iEVLC4n
EYz5Qns/CMtHxQaqSQzT4pZ9X7TCJ8Ju0qtxa+9cpt+RZt3OXLpzYDL4oe6B6CRU
63QlPGnaLYSp8S89llORzEsjhZlTKFTLvrBBDUAr7XJWN9BgcXkpGgqBt7IOOp0p
cgZKLgnA+0Tr233pVGnj1mEKNexWjYC6TnShVJXSmgMrCHBm2QM6LtZ1EqffM5LS
bIonum0MGRLIE/hT162L9Yg/sG0sThiEQDogTPioIcsyax1RhEOqw/2KmCYT5c3n
btYLoZKWti7Whq4gb/76f8jDUX3dwlKGwlPasLYesouD+pMf1irowtIk290y22X6
jC5UFaZ6fJCQomr9HfPdcDqY5IkvsTjvnjgImjyvVsh3WMBPDTFPfN62lG5vpRCK
ePNeqGNKjRiUhLI7SZ+HULjhNTUZsh/b35rGcevQDaUt3dT25F76kUH4eV3wQDDB
9E6lgoQBFnNrtT2/vT6xrwrMvb+Rt+ivVCVdYxuvOAzsDdRtbLo/3bJuEhpJ8qMC
AIlLAYosP7hQqpKxHxcwWuKQww3l4IRUjXFBLeukSjm5ZlYXbrrLDLGMnofk1bLo
7q0Leea0cRG0YPTO4BUY5fUlmy95vxB+SbSiH3hbpcLOE2tNL7YkZjRHFcfoXsLu
/1eudbDQW1BfwAyoffOhQ0AwvVDLNVei2gFHFpyi3W9SS60arNLi7TmpEGP/XrRS
RKsvZbM6q5JdxyBaWg+QZdLfzmYGb+se+ho2n6MVHpa5kKaOTnxl6gk9rEGquYx5
sBuk18ezRD1j7YPL44izAyYsQdhHPyD4lK+uTq3Qmnr5GY2JZpmvxzUdwr3fNUAz
UK9skr/MEHW6zVQ0r75wZjV5vkbC+tlDx85WZfdGd7yZKzeQZdnJHPazyVtuceXC
Tjbfr4rwkP3FmCSAJ4osMT85cAvIkblSjum6WO6eCaYfltrPNqdjgY8h4Y+AMgS6
9KAAL9OuiVmz8ikLnfT7qoT3Yt77mBbDm95MWXRfClp8Ur1yqThdz71xOAZtMfhV
sbrdGGCnuIX9a7FwZQEqhacFl4AweGY/DfwSpzDxi8C68zerkDPAHmk5rDKiF+2B
TxhF2Dw77bkpcXeDLG/1NTKflKmk6b0N1KYyjv03HTnnJH6pYr+rjl17JNmUGRbj
aqvkGnY9DFHV8iqwhmWEXde+yeLwJMHKLw+vDjYpDE3B2SCXS4QMAXTvda8HrNoK
hnIdB9n8I9TEQjNLK9yTTEb8TVwPoX79BubS2dk8YBzaqeqIQ/jUjt2qDXFqg1dx
0RjTy/Y3KSTGzWa+b5WF0WAOQpMngdIjKnSb/pivV7CAX7lm8VaJ4RZceCE3Ixrm
7+E/ztLyTEj6aTPhuCXnwNBzEAzDPg8NxO+Ahc87rpVT3nNPtCzsMjfpRwnK0ViL
H8xZYEeXBbVB7f5iYVZ6oGCzflfEx5axI4fcdC0xQ2pH0DVeTY+kWuISpdxCtN/3
R0zD1QaLWACeXQZu/UAxE6DN0aMoeqsGdfC9gDBe9QddVnlr6liYplX08gXUr83L
7x+k0wVBpoHanhI68YIF2hsqEKV3w5Jv8fT5UIMqluoB+st9TTFrOK7HPmvRe983
5bLzn2l95u70/7hOqB60y0LT6TJKnDNHJ8j2gwQ2CbAoSTEM2I73Tc3wCTRNnKTu
xh4WaOQKASnI7UqxHkRe2/PkR3ERxQLPM4XpgtDU0HFHgd5JjrEIHlii6T6ri/fZ
76ban60e9ISlu8BeLXVOZSKiNdkvqtj9MXGld9nD60O0cI86eN6NBshYI/Es8Bmy
4kTQZPHOEWjHw9YsIXmD4kIQLbHFr9aHRIwP2jqTSADE/q7ZJHEVssoN7UK6FPBq
2F7o7sVunFxErtAV5sLA86D0p4oxxgvE1mHgKxXihpqzGnt0xagbE6YGx9ptj6Lx
likk6E5BIoh7kJnePKr7TrcBTnXrinU6Yqt2zaymVbI0rtGqojHgJmitli6v3CeU
OK/1KM5iG6BO8QT4QsuPYyFu1dcKjV3PprtmbQpBWGAhhUucTEyeuNWUQxF9iNEI
sXACw+TaTloeSXEkxIFoyifhKhehjI4It4RPnbwv8Fj6p58DuuKqHAPd5p41A0Za
JQIZTpfqBvQDoHc8tVyxGQWhztRGmghVKRpxkGKraLipnr8YjNv272YrX18F1FH8
/0Fgv9RaPY0hFOAjuNAL82MlMdqkkb2FKcOnnmESdC0ItdghHqxowqi7EUMdJj/1
FYfFuQMeYJvuc3AIhBLgE/Ot/cANz0UIokvflHo4ZHgaDV4nhRg1qH3oBwIHR4qz
SKK216BavDoyMV7K34iTaiE6kS7xPVazs7EFzbSIvhw3P1Mq+23N7J9TybTYCE6R
gG/C6PrCUNMBv63bfuWYahLfLRgqjXaxY2yssoXaJdWnwPO8tAx9zgaZlVyd+mJk
XSXhfxBJ22sy/HUZCkrbA0g0rcUJ7qTLu0HIkOMcCzaSb7MgnUdlyer5oX462am6
ctQXjzIVXbtGxE2nwQhSO2XyZLNpG6Xrkd6TRS+17bhwRtznePKkcKncYJ7jaBV5
3fg7M1NBhfBm7uVep52gJVIKkI8PRt/aZdy7JaeT4LHji9wr0tKNAKEU3HtOyrFB
JDL+w/CJPzYIVa2XlqZuuXsllVN9WXW9HhKg6sGe7ezUw1ovVQ+SU+GUvHUNPf7I
I5voYT79nGMfFEuFdy43iqArE+BylyHCPj+WuHwsowF78oZqGd0R3AZA+J0hPXcO
/MENdWq6DtrUs8xmHNyqhs8gxPMWkFIxhbmP29jkul6z3ZS1JvmqY0YPr6gLdoG/
cHMxwlQ5pqJO6Ry99m7tcw7v8MlER6Wu4uDvsORcZR7aGzmA1BEUBAUrOv+Fea/z
VHP8OBcIbJs1gwxdlP8IrJcAUH1B7ZSn8FSxVBmG7WPgYGw+QqFypn/v2BJLB1pL
ihO73cw9jMVwTFNmDV/QyQguI37mj5Su6Wx2nKLVtTUBIvK6eX+8aeO33AMXk9l4
lHeEjhxQ8/psk9whUdib4nJ6/BaVt4opGxMSkW56U48N6NlMiDbhg6Nv9YgQFlkj
3GFjbsSJn7bWzM0xkUuiNr6q5RmcalVJGdBeuKODHpgGOE4Cf6PiDhce2jMOZmM/
/vNBWLwdaZoQ0wOjzcyP5dJVnSR1tvmlVuZEyrxMAa2Sm68e+iOZID3QqZsAnmw7
2yMizrAUhxuOBAtA4jDH1xsLKCHVIRZmM52hv4W5vziPQYrTqfyFo/3Wqz4JhGR9
YtA8kPYL2VrpIUelb3FIsn9g24jTRHcV4FA1iOKP9HhB601q84a09APw/xIJNpxG
aW30Ij9X2H22D1elkZDZTKSdbaogCmHq1eQJ+5vxkhr0kTgPtWeRcQvWvDKV5KFH
xmRsVHZZrEViuMAHinmpUgFRA5fzXQbO20aHYTgHfKzgeM+ClsXBoG2ohcsDnXwm
3nzBLgYMEktlqGFCJ9BFwHwN4K1bn+4yAmSUXBBm1WXCjksz23MxI35EpeuiPwJ2
e+3pJii0Q49V1VIDYbWXm77rBznusg2Qozh5lPb21wOchdpM6GafvDk+vCh1VD+H
ESYL7THGzZTKcVI6rqv59IoUR4/GEJn8bnPKnw3ZzMQV8GoHGan7OMhL5gpgnr/K
0X89Zqub5qmI88X3pKlqKVPiA1G1NgCDhMwgaLn7uvY9k6vgqkVO+kb9ISD0odYi
+gkokuQf2etJup9r34Dpsr9UplSEVxAoGEv+vHBUlq0W8xGfDN9HdnJkUXUx0sEx
c5RA9eTqs6TVER7Zm1awRrAO1bGHEPJer/ZFqLHAvWLMGyx50BRgBRaouwknHqxf
khBP0onnXxFnxpk0RwSCXS/+QZ4xtFHkbifMm0PDT0GtX4iU/sRt6QQT19MiWBC+
APSjvASlIUa/VLp9WVtrV9l5AJMMHc+ipAqClhgBC2ZWFOaSzKkbw71bG0+zK3g/
lT25UXTDISVykNi+mN+2iiamnxOHyVRWdxzuAe2ZDxCeE+weepSOLG6Fqk0iK2ZF
DQWk8WDvehADyzDR5QWARk5YcOb98hBNgG/2o2MLw2ZlJulx7RQ+33PjdNm6ZyfT
9yHRT8s0R75UdEBDmqYYiZATM/Y+dpKV3Wb+yKpopX/NNGg5tcSdqWQoK0QhyEhh
bKQcIdYpbDeN73OetGHhR0QGZL4sW6o4Sh+/0dDCvEY6ceZo+xTc+/i/ijv9iNOv
2DFbJ+dia44iio9Cs0LSI/KYzUOddoOhWlxIttp3jQHP4K3zw0vryz/auxBDQZID
KZKzwuNiPEVvcdhvLGHqT9oLEnVwmxuX7cU4W/pTNI7i4bkmQWtiBIz/pl+zFrUJ
4EF6HpXyfE7Mam+6XXOZmxurb0wZ+mnEvQ0ShgmJ/TlHHOsILYt3sx1vrnCID2KZ
s2LgsKDzwofCI7bJRx2Yu1c2Ep4fwRINtHXyyU7sAKAp3cc4qmnFe1kfFSyyv/7C
8prhNW2GBY7cW/kULrQrMcKCKOtuPcnBpP5guJNp/QYeYc07Nu45fxP0sHQLXxsB
QnSk24scNwSw2HYGioj/izptqRGe7b/OK3H3ZwWesU6117zQoBxdweyVjvoS2ZCL
NGjMhtsiX4bmSN72InkJzOxoKTK+nr1wxocTYXyqIbe+sA8a19vY1aoMmVFHT83I
5kK1wOlGm+XwvG8H9Nyvnx9Xa5poAGX4wNj0W1mIupB54uM+cBHFJm427QQtU2H/
8bYSaqrRHNs5rl4FCxJ9hdr43MyN9O1OXzbyVCpOjI6iVt/1LtBvdMYiIGvTQMdq
PummNHW/FNV01VOnEkPq58+eFdGAZAVpRJeJaKB+lZuVRUaDtcwhNXX8JJb8bvPH
QL48xAvFJn4Iwnd29YaOklCqUsY+xBj0eNRNeAX7PHfGVUoiiVYZa7Y90gAOo16e
ifMrVbCw7abCGIEHJAoV7PtGTnvgqPcs7+mODwKkyxB5p1XUJi+McaHHP8PvQ0Z+
XFoxHoKiAQ0ZrjFrOFgdp5ZYYJRY2+o0rWR04odJdwxwJVsjmQ/16hagCoUSzjuo
iAF94rizhBvFerms7Z5B7xEr4RDebyAatSK7iWu8ij06JDCIRqzX4l97aRIPiOUb
jwRPeMRVUTklNxILkCVGlfvZTMOh5fKU1HvLW6nwdooeocoKh+rjjKz+EFCKwAXh
9QNGhFVdAqsqqzuC2v7Q8MPvGM5sWJ7r9xO5NnJ61SyOt71zz1AU4PnG8XLXhz0Q
BTLglznelTdXoSvGkWtRb021ifUGcfp1c2AZSRtHQHAvRgwwQs61Vcw6U/+sOdrf
AUsJ8E5UD4hjGXeNxnxyvO8kHIGX8RSSj83GKx/nHTsdbL1ayGlCzlZeeq8PnKMh
aNKTN0tOaAfS2iOIbmH/ukuhpiz3C1mdiXCOqUeUEJ4146xUvM00Y4IigqkPFU8A
fs7f/hLQ1OxyVJf07nAhCmDRPswrqN+sEfeFEuVLAUyDfwh8CuX7hC6bBc/3wUF+
rO2L2Apbs59LPZ3VlsTQuMays9/N8mXReHO8UM1zN6EsvRcs+YO3y/tLMg7JseqD
L1/+7xRtxWilF0l5+yRL2kdGMGmTJMfmhvN2MVkRJR/6xbp5m4EJtvVQBh3McNHb
RvASNkMA5BQVyocQ3lqe/BsgBiGkhGYQyTenauf1OEEON0PVvItT5i7ULXVVbq7Q
CeQOn6HcLnO2CdFB0s1VB/U2QWTqnnH7cBbWdcnru6Y4YBE35NKh6J5ba6NpXLKX
EjXMhNFGsUMwRiqDvuUPPj99adsRF8W3isP/cKnjJupC52yAMSkm3G3BP+a5XVmu
1QhgWrhkY1iveSDL21BK3+bnktEIZFPvb01WP+INdzJXRm0M7QfcBNKSy2MZyBNO
eCdVxb/SnPRu7Hn2MICpvu2GjOjgpj/9ZaRm6XNTcpZoOZ6/VbvocMr5diGUC0Ol
+8nqlCu3K3EiDcXNQCAbPSmYGgyq6CzzNxBj1uaEl9ynCsuAD657Gk11b0rtJ4W7
8J6Dkl53OXC5/dIBzbAd93NepSn4vTlmJv2iOXWG6OJuHVMPSworoGl2s6q0P5og
txkoRfsSkykpzVp7bCbxqSST8UseK79zjR+XfU4vlWinkVpHVOCB0vEI85jIqSv7
8c7BIIt4uXTS5GgCED2Qv7Ovd1rVi3C8zwvK+bbSxqu1RqWyU9n4b7+WXhRfudT4
kCWNeRxiyfjswMWt6euESrq0vPMTAZzXE80HVAcjmzAVNUvJlxzWARx31w4orr4E
Ul6Ix4mTexY7VqdwrqDCzjtfw6TUQ4vzf2UYgTCq3QgFvpEkdddX4w1a8YXNwV/Q
OTjj2r/JOFCPVioWO4wHFb4J2Nlr/ysJuZ0j+ACbFODHXMgsxXR/xls9LzDogvA4
L0E9uQa0DkrBU6o8oDiU7qEmJEqgq6n+kHox1Lw3dweQDADcwamo1PhNo9XOBqjQ
LWEvRbjR1jOTfatmAJWomXrKslp/u4XAmqYDX6EIaXqcKhI5Seo+KncTlwTWxEKQ
SHWfGVKluX8lT7eznuySV89gz8xB+7XJrOysJIaU4axOOOrZUMnHe0gYZSjyG+K9
9QtjXfUmpTonboolDKnf8tcXiZCsVCtU4NC5CocXMb+SqwC2yu76ZGlgM8Qni1sF
mn52W4w06E5mQIrY/le0I+/QElVgUU+zscga6JeZIkeOIOky754FvTCFHZ5x4jx5
xxx6MNPjp68/tJeech6E5g9Nc5kFPTUU593PhRsBn1psJcnlelZsdjPWHO14kig+
7BopIIhstLzrSxBEjsaMUcJgTfg//t/3V7IhbbnGilSUPqyb3/qq9UHKAxUXimEg
zD/HAVsqIwebN6TAifRR3z288wB/K1q54D+51i/s7q1WjqIXVUnOm56S3BC7OxbJ
iy5/an+29VSp6zu9awMt2PtqBWBRaHQ06HZDip1ensTc6KogsWGIGN/Ms/nFsj5v
QK9QZ3IjXbhBX2hPKo85HbYnRgWAFvo7QyOS+kTSEF/kvIOaqtuQ/gm9HBNVTwo4
LVml6aUnzXlXl2rqQOYoiMfQRF++QGaR+1Nzb9Taje4YgYxYN6b75FzJx9LOfhs2
06qLukNF8ADs8OtljtoNB48C0MFIAUkuEsHsEYLggMWAbvJDOYXm3WhCr4GPKKMU
0Cp959CXVQ9VKVkhibT+YITDf1LdD4clZgrflaj26l9iSQcGLlgnSTihgUG+iQfI
2C21KsuhVvdWuzRy9lqc0RmHamAfVLhIm+wP7o1wYG4BimPHSA6FFHuwIdx2a7kv
GnLE69fJXY3wbQyqLFjzbnquh3PlILcuhAASoeOvfPKp015VvV609jcV7f53e0Qx
VRdgecOzsJIPhG14/hLLXfgdhkmU/uLITIfBGhGa4R2i1krgMNkRqUxUn9MWQSQH
bc84SA5HwHDkMdApqNB9uJ2PYT10RLaBGGweBQyD9sn8aZXP8o1tw2Q4XWkWGSem
Mh87+CbJkgsbVfFRTWQBC+XXLZubGj7d0mh+CmwJgvjZfpFf8X2T+MOJ/VRcXm01
FiNYMIK70gCv9aT4GBBnVJqQqxZj4ZElDP8d+IiMav5WH6gxr4W/mcgn98bIuTQj
miyi3oQqtHitJl3ouVh97pBb7ENHTG/J5tKa0d4b+PZqyzB1Xfef4jA2zgITJA8Q
Rs+6ofHWhiCk5EHQE+8Qpd93wflorVFZtftYna3n4Ip42VncNcA3MxyO+G2obuZG
PkCcAe8eN8rTznQpkgtB2g0Mhib917U09AWJjRGf92CXICeuKhCQEXjGre8QyU/W
cTsj93pJySFfubS/NpD0dR85/duIRKrjkR+qe0I3nZ/efvecYNypguhiVxwJVhLE
7kWRtZDDKqRj0i3GiTqtnbTD4xfsD4DZzCNxRf1Xc1oI6o14KGAsgiPzudLJ4Ryc
zUuGtr9fBBZyDBzHPLwhxGxspeE5msHXJv5li5r5WmrQpYkGhoyoXPfKsBVSIVE4
P0FQ+aaw2EFQWYT6qXZ4TmRmSdipIrFIV3FJUwDhJbyZ9yG4w7qoZdGIL9Pum1XO
/XEx9bLIxG/lw3fj1SRstqKFNNuktoAFf1HBe/jkB9HsW9pfTKVzfqugaT5rBUlH
hOQoRqVMxh9Pvh4ZHIaN9BfTGedzwVP1H4ITa1Ukh5ph6WXhIN1bSgvi4Vmlj5BU
YI4k4Zcj470BLqOT+AU7ct5JpUMFiY/I0MvwYXjvmO/zO900DOlhYdn6DdeQ/0mQ
pipwUhWcCYk34d0w6ip/S87OmNQzoYYwkf1XIqSv4Cud1iFSsQZZ6nr7LfxQvOKR
hF020xrmDA9hOfupSgBnWbKMM+VWZXb8uDEb3iXAcJ6GgKANrBE+Avy+ptvRfQP5
TXC/ZCWYxYkGCasmj/U7iKrtRDw4piq5X6/5HA0keEAJHNWC4sNRor4cqj5hfkJm
TriUvB02/F7JjD1jfMrWEAchMPukVk/GDq9jDrUTIqadGaGx76Hy+U6dCdnuZuJh
kgP++TySdXk4zqxpBjdOBLNniZmtKyO9V0T3B4N3fk6mHANROrv0SmyiuwvzPTML
RuQTNZhWSmKqPNicOHF59MpJB/WSgK85Vgc+64oH2CZXjDGphSBkyttkoGKxnw7d
i9Jn1mZCKVHcdDgJgS8Zd4/xutY0GxwQgnkfKB7bdumE24KRPGsJJ7n+25ZKfuze
QeqGcDz0Xko+iC5EzsiD1JaIczAksidOjb8pb6atdOUbtJykG45tMczwnsbYDLBU
5xnyelWqfJptL2GgO+jiSzFEh6DXbB5xu7FL7Kh01blfeebboRh+6uVPTSGRZllp
r5jv19WdLlvCZD18K/I7MTLZCvLJkb9y6U4a/oY44/384Iv6l0DXSWPY72oqEVOK
fBT4WukCR30cXiBsmp4dZ9e4hz0vCA6tqRhLJfgulVBcmitszeZPRjXH2KtgAxZQ
z/jDFEIQEMSIv/BQSJ7t7ueq3Xs1nJpvA6AC+xKfPhLrjILtXWLLgCaQAe7OY0Lq
jWS67TVyj9tlpiPNxZkWN8pu1Df1Qzu3g4UixLT0ohBCeMCezvMthrZd615Wc91t
6N1p4WtYzkYsmP9STR6Y8SY8zhmy0LO+ughOouB7TBqxSbTNxll0pjDsl1T89ZvJ
p0emCm9rYZO4CcnaGq0k0ACY0pUn60kFpRCBhmPuKBvHXPq7Rndy/MM/C4n3zXjj
FCIvw1zod2sRcMPTnXwdXk9a36B+hnKLDsDxYchbP/3OA0uWYLd2v9BuIZoTwzXM
2S4Ms5RoqJGydcp0FHAgXeMCTWYQS+88kLuuz9qvt8cjP4lRcFERR0AYsM7oi9Rx
W+ucE+Flkk2O7G3ZO5MNO1KrXkfOs5AFCsciHDu8aLUkjGIwa6tiMg5719h9AVvu
ROc15jrOZTwCDB11/2t7UlUqim2YA68u5P1uAYFTq5CKJ6N1TWJoxZYTRvU1OA4E
JFESItgpunPC5g5+gpCR6lzwDO9J0StbPIY+NgI2dA/Y6+zYvt1Y9MVoHUArgTaC
98m+7zO1lNtcAkER9Vw4RMkLF7Uc6NOGUJh7yCV9x7ax+OlhFSHTplMjepXeTRER
EqupcpC17QOt1tQXOXeokWuHHqxaQ+2goAd6R4UDP/3yrtRo95YewIsKKzYV5Rue
+bKpKBTVjSnPPmTjD5RDijdNdzjlv6VB7tnFH2DMmCoNpO6WeYFT1ZYW+i3uHlcD
12gd4+6OZWJDNRmte0W5hGrU97xCPHmDVwkxNPKsNOuieo3JcYk7IKIK1Pa2/aFp
DIpqqsQ1n2s9B85ZFtpid7Ux470b96a6aPEDYJwMAm+lShPX+EBatLF0RyXEl4Jg
3j98Py57glSlo0qJxzOP/FXBgIyxHpZqSUknriyD3hKC4JigkmOGjtFFaIIQgmEx
K9TIGQ1tMktEOfmXwHknOT+kYkFbwifa9nuCCkikRTHf0aiKPH5JJ2dcV/V1VtAR
iP8EEFQRMFMqG5bIBBrC5ueGEghed8NkVZniYoMU/KH7h0bHqk1Uf0dKbeh5qeH0
TytiFCkIZ4X5uAy16/vIbSWXt7DL8zug1/obGoZPEIkbwOz+gchZwF+heLJSddZk
iBc3I6eJB6tws1wsNWrOS3NkiXqa6CWjQV7/daiymQu2eWJWjuGZre7wbleVnyie
dO7nP6/AZaMX8i577iFcpVfX+7aEVRf51mpTy6xAQ6PfsKNmOP0JXLK4hKP84wZc
7GJhv3xg9/R3CmJBBe65vGGN3PpxEIe6gn9pnQdRVQenFg+L8JqcrbmXZcx793OV
5x1fGI0lRtxgqrXqv8JbeG8b5EOmpAKbbAodVT+BHDygF2NTJ02XavKMNpW8ky6J
7EniyjG3nAh3z494p8e+1oSraGPFCGwQ/Ln23CuIxp2k5IbD40EfvXDj1y9QxQ+H
991/7f82zSfLPTABHzSkD/Z5eTpoIrmDAbj8LSSPLcrboP9F6gSM0hXiRcEGyNbY
mWe+OTzd3AsxJYo6BwVJqtRycVoDOpKXuTENQ+oSYfQv7+Xj/MWQgT2MDTA4fQBI
w9pcF6+jt5SVMvYhV4Nv+TETN746Uw3jUeo1LCjxgK3zKy2XW4mEF/4gflKwwin6
ke5OsD5vwO3JHpoA+W2UyI2TQ0JZrjb8bkmrNEtvXNAmxjHrF1yprnA8UxFjIFBq
mTtxy6QxfCbV6iksbr5QbC3tz3DoS8ggRhrQ0iu2FU5J1USiIHe+zd4bG1DdCfmN
iEI7wouHPFhJZKHLRo9Mml39ffDSKLkNgLIOGy5C7fyxHhRQzMT7VI6ycO55g+iI
yrdQIBV1t5ZSLT+EBxIRTzYjc/auXGSwVIcY/ZQzSWzniN7SWWU2e+42NbhhMVYV
tGNUVXrEZfolKHdeiacBma9w96zHsT7ipxf/NB2iE0DQT+3qusjrjxM45mtI+2cU
J8rUBO1t+BxR16xQ83Sc+HvZ56bypzOieLFtPCsbcKJQV+/hqbzuN03vpNJDbdbc
TPlBCs3AQKwkLH3A7Y3NLXqpMU7OiZ+1HfY2AAdtmeb7bn2+G4b8cq6ikvjp4p+X
HtewKPAq22+4DmFwAU/8e6qluR6SBaSYnsfJqZ3yfzHy/jjlFmHzZCnz/FwvospI
I9OYm0sFdeg3jSV2DGZhcfmKsAD+FszX3rLj8mzoIzeLegmlb2zI0JdVlH9zMC9J
4gcYGHxMBY/g++ZwVfG4dY7hWqNcw22doho+TCEixRlBD7jZJf3JzWnIZ2p0oDNm
2ZNio5dW7oM/vDyF20ZyGq+GJAFSizSpOTrJU4hahYSVQCVKKkfxgKFKZVZY7pIz
u1x37Z6iTrXNW34pqfg+qxAy8EeJUhWd6Yx6G6Wxl5iCIrixqptOMquCwhIreuie
kcShpIjv7+3qtXL5OQaG+Cz8yQl/VG+jGskJ44GG/MBGa46IGqY1hk9SogZSnSj3
8BPCre8lAkQyEOh3d76J4MBVnnhbFaeIfRmIYwYtTYrKqUeNZS+M+PhpLCTSuc7h
Ee4fs+knN3oKDFuWQuaSoPpA9zHToXxrG9YUJ42vPOwbzND3j/a4DUaE45mypPX+
pfvfrQZJjE+Ic9ixZ+3EV6fFGTS8sfDVB3q8w4ls+HS7WgrIHX3m/8AdhO01aAgm
2jf9/30gS0dxpnvC4TJ3T/JG0TBtTPUlfarqMFucqIyYNkHcPu9cAjOXUiz6eFq9
VTk5AJDf2HH2MzjosH/0YBd2zZxNJRT+yIOTC+SO1r1EZTtSHaF3cKyzojyFRXSl
V0t+IHPgOXEPJ8lvgvG70DC/xQmztdmek+Oa6Ro/yGUtWUcTfwM2O19LCK+0i1Z+
F9IUJebHZkc24jcGErTmOCAW1MF1ma27Y5Wal4DrUZ/xKpecIOQuwhQvhnQ5t8Jm
KgVqGNmT8fdhCdaWwtVRqAYGA2BdLkRm/kcrBI1BZ/OozEkOp+0SmqX5noLkLOd/
QMrMyL5nwCrgGa78gD6W+ipxITo+fVo8E08z3hC7oHVCecy+DA7NMbRo49oD7rr2
0qVb8V7AxySvEMUa6oxsF11fbcLwweX97xTIH4BpT88JSrAHrchK+noGJ12hLtGT
JzZURiLg0wtwe4IX8ktMcNGU2B7PuswXY6hsBNy5O2pqFDLUwlE5H52B7B2OFjN3
YY3sJww5Z1+jilDpTM0IaDdyPPgwjB+VzNKgVKfrBPK3/zK7Te9NTUMx7WZafq09
5fgKOfKoejnmrX/xIbpBuBfLK5DYZp2CckVbcws3dVFTHpKjr5F1SKeV2lWP/5SU
3o09lmrCqpEjoHptcDAwtxXsq8GtRPmO3rt8NnrO1lP7xekO4rwjcMWWbdipeHQH
H74gfhGf62ENMUzGjI4PXheELwXYIj5Jjqtyrsw14sQeX86sECDD+/6UXKiv3vMv
55KApYJ2+vJhugQ5EFvFhRBsqxEpYLh5TR+WZyuH+OBMNsGbhsCfUnFzyZZz/5db
NaEpoBTJCSIcsDFUWciChPWfDBY1RHTTibVpLB7Di+dtwxXgEmQsCwZCInnIvp3I
braeeed+cx5Foy21c39KvXo0CpD0KI1uZaswH9TY9LSAjJgTpLl5NwYID5hGRQkv
NK+6ZFhib68Q8tULG6ZuutAgoIplsnWD0hb9CN/TvsRT3TeRulw0hKJ+4k0VtrDW
K4U46NqvMEHpUHR8g8gEwU5J7U2kivGfBZot+6TEtGnestUZ7ZyP/5M1oaQ0SYyf
BPldC80LhhmSH/gFGofY5QpEIgW6FkGeytXdR74Ch8Lz+JenojMpUA3YJ1qAlnWQ
/8WyDH2bagtV1gVGZMsp3tHGta7dTnPb+/47qjsBhTYm+IBkQcZ5AnVsfqK2c0zW
YYZyqv8R9lHpQItNfGZi8f0r8AKh4hSH+opA432taMHLvVcCrB+zfI1O7uOUU2YM
J6YIsObXbc7h4vjlvT2/LvVKwXIbwL1fY2JJYkL11sH2yX+VQfdWFNYfDVUTgnqu
ft7Z5YYG8V1d9Ig4D5GWwTjPdB01QV+LP3ghAXDBl3dRRyVGcv3SlEC+DOMjKTP+
sIIwMAZvih9Eh5cA//KH7x2UHQzB6d+X8ZGqM7JBlYrCBWzYFptDacGC5GKU6w6n
2GL6M701w6D9c4POKYlCuqd74isFNlIHQT1ILzIvwGhT+LCZlPni/NeFCI+9kQNZ
kUbalYD0MVuMObfvgr+O02InwrDdMRrPwv7np3lUhnilhFBHegRIZ80oVUtmIlRt
/4/pzDV7uOF/R5o7y7xOL53rDk/4/nco17zOT885CbdUu+VVo+jsDfEoosVcz9um
6t4abKRug56FaQ3BydMVSfWUiRA0JXEOTAMRE4flQUoT3wzDLrhKz1H85wVV8qnQ
Cqi2maeb4zw/HGkcLTK/kWCi5keK2xnSefg68iELM/c/jYf1vuwVXd+bPO0ROkWU
aF2HcyZvDYYQw6U9gHsqZoJs1XBRKFKIPwPoMe9X6LbsRmlBJ5xIfF1QrI0KzkLg
P9J/uFHwLwnwWEkKETPIFBryMkiJOgiex1t8u79YutRywmbF4Y2toiL8N14vl5KG
Uqz9dr0mNbpy+agtiwFL4ryubBiueRnsIXoaJXcPqr5p7JbubvMNstZprGU+493U
D+FoGw3oDwAQxj1vkgpWVWigXQM7dY1eUukPY1hVo8+tajhANk44Xk5TIUD3iZ4F
hdGdOBDDoMpTqLPSL26gprZ/v1XOLTGeey8ChMDA55d8N7mIVZN3fJi2sad2eEmp
LrZaK3E+YIeILmjdJDXbEwzzUvxRVLDVtIT91koe50unwLiulZIDXtqY7kbAWicf
tKGxtQHdF79GxHf4bJcjUwkAzxjCaFKY2HLmWcX5F4iP3phPvxQT+XPRdDJzymFM
cBiu/sC9DNNxevWWJkjz4HVMdyRyho7JpidL2Gj7ocFEBreYoa8PGZRNtHwjzo9n
YYx7j9sl5uzzp6sGuCAsy0ewV0OjQgNl0KG2wqFSIN0hAN6LLAGIYiVY7fYKi81F
SqVYZTpUW7Jm1KNcrmB1KyVABQQ+dknZhr4qmGa/rPBV+SPbmrW/gAn6T9sFqgEn
vWOb/3CNGGt7fqWcCazFsiSEEsrn40IOmvNpxm+z3Q2U5xqH4j+mVSI5QGIwCNHc
bNbpkHZLFLhTIKJOkWccPRYHM3NA0Y6ZZkPWJ2v0odbzCKfaIahZJzwyAYgKNpCw
YEfh+v0w5zSbHqcanR5xLHuSzRtC1DJM1pO8S4lw4RkG8+7XRDOmYAAWCd5X6Zld
LBME0eDFHbP6SIJle44hkq0N77LjdK8DKoMZCFo05LCmynFyFim2a1myq2Juf4KB
DHXzwyxgqkE+LbZN4QJkDWFUOYWMPfbMZWqxAKzxDte+sAYyHG/4bWxHB4jgWZZN
Fn2FEhS2dXBA6EcXPQbwfL4Zy1cncc2IQjyJBSrVIvkKUDZaAlbSecgS0P7XRV/O
aSK1KDzpiLnNQ6gXLgHoPDW44+9GfZ0/d6n3oSfruDvuKluebWqFmvkPYfehDysT
qNOaXWA0iscHqW4v+K7fpzCv0hMHDqtu3CSlqm4pWnKTsCf0DWvbTfWO/U07y0se
m0Kb85AqK0rVSTFnhPs95QcCkIC+XiktC4r5jKdzGF4tN79BACmQ+sjN75XaEcMO
qzieRCCYPs9nBubjw0pz1Yb9jba4ak9iXHnc5z0MBVePmAN2e1dzd2DLiJshHqLN
71afPl8srFOkMSlo/R8nkQ7TA3hPNhqIgucoMuu8v1MNr0M2XIY6dunjrX++NeUo
kXAy8iw8K6jBTkYPv63qLQJrdRAXzUPmahyljn0gWZFubXSXPxNtI1lYQ9gbB06z
8Z09wkyUVJPAgPEEXlhO/cpjZP9k11+CA89BFnT4uan608Kh3jV9Lc9jpjW1Vawl
6AK3z3kHtRN9CwHVJ/Xmxwy4FiDTKOPZheOMpQ/NcuTzv4PY3CloXcEkRQcGAa4F
iJPHQRCMmd+W7AwVzhc8R+3OCLrqmoYvkjrr03XNsdHWTZn1IlcGjMbCMbpwgkxf
PO+ktd6bNvLX6WPnctgYW3G6kUMwarhDf7OEvL6rmO0K3Wo0o6cph9gYi91kDpM0
bQ+8MuJeUAAJnkkHyQDsJ7fOPrXSLABFtCXZ4PP3eIwoVCi80F/fc6jSoCBAcHCk
eHdOkd+jJQOu5sFZvbiju6kWulIsVbmSJGk0bl7cBuIqzkZ18LFIBBhbSFU+URsF
CymQGDoxdgEhpY2P66Xrq6uALhh/CE6BYEi52KocH8DV1qNx729HcT2yXZq48/lO
r0Bq1tm6liqN8oU7xXczgf6Wed1ru/QKsuDsuzf554TrIRV7/ZlAOvE9Q7LW8ntU
w2FYkjEFtHNzeCDXDhRqupEVtRH653vC1JhQ6qofakrr2OnN526IPCe0M+/Uo5n7
c0WDr80YQTZFK3yswoew+SBvR1sLXMjxIlFsT2yi0NqJkaSZlSycqjsPe65lwfYh
dDuQb6VwLm9Isw8qCKgG8ralBdvGL7mspTpaSjoed6HsjPbdASfOyj+Hx5cVTasn
Ol0AefmpYZRPLv6yIpV6L3frOKHoewYJ+ZYWpNFe5tZQPWqbjFaM71yV6drmw+yL
6jz6jIwWVe+6H9R2kiYS50Ek3Fjzs+UsEWXZrnNzxOAvHWF6dxF/APVXbIIegvBX
iFYFqiZl2VuaCXSz+9A8V6SDOkIIDkTlwNkRZlYxfPE5w5lAZMuiS+1Of+Ofv97O
5ekrjoucMETTe8NWdMIf/zZB8eQCQT49JTZ8/dOlHlse7q5LMXjWGDOe+GqpoqBQ
FRvtNPLrPIALvolbxwSlbb637+TFl681eKYEOrNCIwzVCyeUB4hY5ykzBWZBCW/m
6ZpLelg2+q+MQ1+KBvHuo0g3mAxth4eCwgXraeSWijKugw85eKFh8CGEn6a5CLZD
H7LyWhEl3+sbXZQ91S3q2vGNBZvI+HgfQo8h82RREP4O6yZneRkXXGy1Ndnu8v6P
L1hoLBRuulu21fUyk9NazZpi/whcLKyGva08utbKoDd/SyT512czaFIBkgLq9P62
sE1+jGwoMe6nORmVwc/An/7h23iH3L7nuJbV9N/QkwDbG79sZ0BxS9xT1Z1ejr5i
7vvmUkPBM/OEogabjSHvrwezLwFZnBaPAKPeAy6Q7yZrX8/gnHGvRSMIjaKALmY9
sR5RERCej8KS22gYxzseTFvbLSLe7Z+1iTLAIxK6QG8iBxKQ25lbJqmWOV4d9yqp
7oWndLNBfwm3PgRFWNZ3qzdbQdSVxiUy8vaXYdLfK+ABc4QAxOF9qaVlVcsCY2NQ
ar7Ijddn3Yl/RLI1ZrpmusONMGGWSVvQUWIuLMJR3fRwIoz58CrD0n1t6PJjiqmp
S4SW4f8EbG3EasCh66NWD/XlmNWcgKo6Am3pDuIBfMhOIU6GQee7Pu48bW270P6O
N6ET2wQqkwxnWqZ8pp8PFwviqT40VPVlClnbVkFKA9qENrBxne1dyiAKv7juckfZ
57JFfBJRNoNyl/FKRX9IGnIRhHiohz2/N25R9G6ZYHYQyawd220ziRhN2mbwo3Z0
tT//r1P4JEb8ScxPkJjK46HFURRHn+Ba8K6ivQKhpDRbY6G+SO18h2qWsYTTv7rR
asTIt9SOQKCCi3sxnEibQpRRpATLE66WhGUk4PNPSSo8Gi27shkzDKtG9GQEOTg6
Ld37MucaKi/hBZCpzHV2zhCk6o63RJW2JRYgsFM8IUCnGJ8IrfDKmVwbEu1Kf9dq
djDQo8io6Q9tjuUV/kRuBCsOMTEZbWezYHJgXcxV2F6fSbFWlScOHahvQd839iwV
nOw+cdeu6eGjLQYrYStOPTuQm8ShkeTkotHJmf1WUuG7i/CoOZeaUUnwbdniSiSc
kztjZ0BLwjqDdeFXRIT3UETXM5YjnGhJPSYXeuX10+KC2jQ8J9unEBiJeC8nelMw
CWpsQax5mjhyTL7SXHeWKKKsJQmTTh/9tA/gfoCht2NkVc5ayssq/oCAnAp0fgvo
XRghG2VFqI1wyjj6n4VXPZQVIxfCnMSTrbV8alTD93/hoyhxRVHvhdRSEnFa+mQ+
btszAm2OTp1FjLAtx/lptS9Sf15J/kZ9B3qQYmCtrL3woiLl8zx3sw/XVZli1SPG
zdFtzdVYER+Y6NcoTyVkKEPjKgruoH8IUlRknv6Iim7/pxkfm9SS5D9XWISbguQq
bH8X1GGAnvP1ArDjpV0iVaSz7o9jATy/fBQUVduuB8s/RUZq97VtP5DjOsX1X5hE
F2KqAqwlMDf4ovcMQ+nFTE7IyyKZi3EpSVxBmSadHg/HtFmTNTJ5CnQ0FjRaBvmH
vJHC2KDorC4qOzfNqBIigXSIo9hz/Ph1lxJaCgREncq2Iw3jLbtkUWfUPZnDhN98
sHYKAMW8iQyyjD+RIGkltITNeHZ85PKwizRyTiGhT+8yTgbq/r2pq9nh38J8MbRK
xK0WC25gf4Grkouo0GpoIGbhLy3cVstTIfkuhPBpqt9d417VWagoKGG9zCOT/lZ5
aRMKGXR2gJccJZZxgk8bsXhJv0nfjBdW5zcNYbL5WD8GTBQyBI4IeKiQFPnQhYsr
ZmB2SCH5JntCNFP0jsovjA2YpVIjIFvO6Nswzw6HIQ3/deYmmpP16H6Inh46wQ9i
UgB5jpAbaUol//NG8Ca7pxNlrAxV/GlTdvsZUtVHjNlk9b+Sdaon74YPE+ax4VoC
EJifCDUH2eytIvdaaqXjO636/PvjnRGFQBeHsH0rgOAyNLKsgNaH4XMI3P0t3Iie
ODmN1spp9afF+t2o7oLXEuZ8MCxWVV51kZhFTombLE09SaeR72HZ1cBv27oo0NIQ
rv4r2+Km0UQI9rNT5KYAa/nRH7E+9l6p8HdvxLk3A9H7t3izqznMnERMVVMkekmS
VxhtFRuK/bIy6IILzuwtVeOgiAbYtSMT4SOilx8bqpGdZfUoejhT6t33UUcGHuAU
pz+Cab0NN7GRCxcyB6qpCCAzr5SebUBBnzMPUbOLiMLmmGSjRxyQj5frq5qihIF2
LLa5pKzMlILfpKwq5M47u1N8xu5W34Nz4Qaj+BD8ihtOUECw2zJeYVlBYqQLrK/3
QbcjmRikRCH6FdzsoY1BY1v8uiQVBcorPtifT6hakrbz3cIQnCF88BlLPnBf0ZmI
xk1TPIN7oYGmokouHgzZ5ohMT/l619QNbcsz78VXE63my86KAh12rn1AjgeoVcmj
P++KcQ4p+UliOBAEmYFKm9tIQ1g9S5uMItYaK72hotjK4fnCHZ1qUrb9a4+lLB4w
7EC7oMU52yzTIR9Jeo9Q+4xAJKZmUVpA2bcLfPUE0TPLbBZWxcaDQs2jYQ4OdlvK
eGLkCG/W4zQ6r6jmumDvTp1uk7CTivy6FLXTrgAXCrytR+KJr5DEQTa9O6ZaJT4+
9AsSB6QuonhVsFeggwnplKebnUg4sRJQ/E8+txjLczwhR7480CEWcu2bkQStg08u
TxOTl5ed3YKQauAqQRvzckvdogKWlbXX5fnIh8NaM/zdiQFDDrrXPhjKTOlpB41l
28ZQGjZhuX7HrfzaiCRw0Ywrsag3JAZIk+ns6M0HH8TsIVFuqlzxA7jJQGWDUWFw
anDBTtXuxe/Cg3jvATWoG8cqDzxOJf12K3+IWe8CHvN1zFxn8vMCsz71PC13XKlB
tlor4h8HYLa9FGjYfIKkx6a7Bl3rDd/MEJii2ZlZazY35k+E36T49q0BE3sSRbsl
x2NU4NuftXarofIw5Is/nEwIdrz2ZLuOu/XIWJrNwWW97lTGgIZqVlRSw07HAJ7g
leEl1MJMH3SxCrqzfc8QiE90OL7KX/iUsS4Q+KaIP5X8gRbcGkklCepPQbVdg6vZ
K7GyvpjZvZYhSdC0tFx4bMGpw5x6nmy/Au9lM8NKogHOPjlHdvD1+rpBY/q7WkF7
AyWJ2uuhYb3/4DfpYlrBzDmdM+9aaqYMXE7JSwISbvL70NnD9Ksa6nZnaCqU43Rs
Nhe4kF73JB6axH+LGjKwCcZj3r3ivSaMS99snHM45iP89e/huAYd0lYPbXC4XwQ/
uv2cf7QblRphqs9hyz7qfnsImRqq51Ro+sg0eY7Y7GyKEiSw4takaMvPuaJGyQRF
aHx1wc3PlES1qCZiU+aP/SH4BeH5o8CSZXe+7Se+UjLsxe37jpdlTdvRwMMRHoS+
KDh2itmex+I5sa+ibX31pTSVEaG+8SJHntdyTZu+BXq/sH1el3lYx5Eh6SfEG3zh
cx2P94tnMjF/cwz0jmDqcr8EjakIjXrYPaU5iPZxVc7NZLXM+x3KR5h3rHnZnj/Y
zreJQoJTJW/uc+Dct+TfAItukUdi6WuA6du09EjJhR8yKep3L69Bi/Yag0/X0L5F
zsv9fk9Vg3O9mWK00bzeJ5Gw4g+GrnvEqlLvJRaNpekdskvNfVzNOpS753UaDtk7
6QIdHf81Yi44llj4+cZOpDhr2+MSdvN04PRlDuER3hZoBPpt/9AQdjSOUaUDOthT
alxL3kCSIvPkZCudy3WcLzGu5CI9MARVoKIGMBiT++lwn+URCHsvOhiVbd/pZnyx
9UGAEf7yrG0sHfNbc7sldD3BMnSC1nt03zKA+TTrL28hnqgCkk3KhRaT9MffT6En
cTzuwNmpMMVULt0cANj5Rd1W1aBvqM4Q3eHxTCl/i+uC3RmlZTb2T+tOla2YqbDL
vEzqdusAQ9rJtjbv21/FHhZaHHCzIL8l9/5AjefuLRWFRbqVP2kV8/vuFoZ1GSwh
hCmcB3gnXQ57PsS69VE4JEhLV42kSqeGtD2jpnEoIb7o4V3K9VhgxfChvjaGSDBB
yw7PouBlS8GLWgv1KXraGwiWYkwa6g9/dECe2nCqg/6hKotvi7VV/jFORdVVZZTV
XDHuOpRa9PsQxYLrYt6+fmPuKq6nA5yAKo2RoCGXYylf7yWUS7xWosg0/KCdXD/Q
eetdHXCrdTnHWyR10LWU6wK2kM6LIj/2TFOpG5a8shCaAI5MAwnekDhePhFM8Jic
qgg89FE9O/sMhCSEBWvUFSVY20zKRyluoVJlQQJIV/p4FPjKgsFOSl0RUivy+HNT
8Iuf5eTlUatZtmu3y3y4sE+sTKFQ866BKHHKKys2lqhYVN61mpX4hX06TC2Ln/pJ
hu/D67z1wydoaPoinvNw6u0AEkOjowA/wVNPR27YAkjnsgtrEftUQz/RbhaE+fhU
IDVmBjqMPejLGqMfrVQOkp1i8vw+CVP46doBMxqxgoDFwX6OyFr1GGOIqL4yyIX3
WhZzs4q2j58SGr6Ef23OE6m4B8Y0e11isISw7g4IcyhwyKkviqmcFvqHIj6QU5J9
FYzQ1nv0xPO4ghy+wzHVGSm8nHZK29dKKmD20+rskBAY8a2tEWuN/F3pC0Yfl6x4
7YQyyC0PbxC0/yfJadgXGG5VDVFzg9kE/QUJhG+lU+Ss1LlTxeo4bioYgBR/A0RT
m0GH6xygRFnglD9B0cGB0PyztY/xPpNUH9No83LDkJTMgHENBQXsJQrmLOW0xj/k
gpC1Gcq90R7qBEzaLvAW3AwmoMG2aqvrr2aK/htKX9sMjdaomL5ylYY+uQOWq3EX
7ApiUZmFA+p0VFp1gYMU1LKavAs7/SP9Gbf5WSXa9Fh5M5mUQYUGq7JrAqNal7Pj
eJdPy4if/GJIgWRiYYPtGqBEAuKHuqd5eEDMoi9GsNkSl/KMV5RXQ3XWgdNQWlHQ
uPcsrS9dWHih9SeVRnXdsFMeMtD3IFnahynhjlKGOtIXozqZmAqO+n3qW6Gh4bUq
H/IqxApRIEADqZqzFr2bpZnWgoQzeb/yzM5J3SdYtJs1X2FzItgnuJ9vsSq5FXHx
yjVi/mmJYnHbHReHDzAI9foH4DUYoPNlmRclXOFq6wZZHESz0N0fo+Z1GL2nx7cf
JT00KNAwnCRh7E0QhvGnlAlNVEyBB8tXAtJpo7H+gMtbf2ZR6MdvNoh/i6dSWTtp
aC25Kt3YgM8Kt5kEaRqdgYzNn+C5WPmpaaON5YgF3raePVKa7y0GFWB0Kz110ILR
ykvqgHem9qE+oEnDq5weyl6E0an6Y3tubF0su5mVSOOPmZxKiJNt+LgFvg6Xw0+K
iqa8BjWrh2Cot49aCcyKbYF7ni0OqmTFyP55SfAe0lxOiA1QsRVS7LAI+O3PGKEv
dL5vjtWEJT7sNeazIRLbNLZI5bQV9xuf4bhJbIY24eCooWO0XgoM5fG2ttu3gK3T
bT3K+YFqKOUQ8vnTfdGfj1UYRdqPlqo1l30NNHDIfQBSO8DC4WNb+Kkb+074d4ov
fkbXGn/Wc5ZEIS+c1XGaB4W4OnyYUi1l3yMIbeXMEezak9A6gZkDCmCGeWPded11
CkCst1oV+h0czv/CS9vZjGW4tpPMDlDVTklL55iZyThyXGu1IRwOdmUeEGgKFE3B
mjBbLSJtfrDVbLZzIMJya+Iy9vBVOarCsNOmfoRV9A1ixu1DsAIf6xKlTZqFhGaH
h4eIqfhytWP2qf+JzDC4CdXdI0xxUMRPeki+cvZ9woI8RWJWlWdcQyEyaGpv4N/d
ZxeT+FiL1ncmZhxiFKOLXmaNej8NywyScPNYY98rTHL1GZ6QHh2iXpy7UJN1zZw+
Ydgam4d6/yedWCqP0U6pGI8cjVIirLjYZ6SwWJStYynRrgIKZXSGqrT0EX5BDYPM
+F9XhjUn8ALD6LWPLyL1BVKaEBvUlj917DNxEvDIi9Q6sjjQNLUEQG0tk/J41j7A
eTqQD0eMn4kod7RwRaF3Bz3VKtH/6yA99RFDdR7cYb9GzaHsQ7A1bi4AE3s2Os2R
qbXOHxcY86ouyEnB9JiTEiYdOJncNZ/FpnknRPdVEMtm/rMSfR7baqoK2bBuxksa
SEA+YkMwy/sWpCo+u9MbGgxeYPySmrpQV3SaI8JuB/etl7IyTjQTQgFDD763PrmS
aP6ubKpcguhbd1RB68UEXCA0F8l1tEJjSKw6ql7vBTgtl+kqfNLHJbQQc89L0C4o
31gle5CvR7kNaJ/ZUWHj7XQEvW1TtP3Qzrh6+mW8lMkTdPzQSloTEbwRpc716IeF
t5+oHyWBYq/mpHBpcxhJuqep8IAw7SlaJpvyMjo17O0gtDAj8RVmSXKGc3O9o0k/
PALBItMUSWAL3DUUlK9XHPplQrnqKbJPv5TEkxarDsn6C7nCe7f3PzkmlIOtChUZ
U0hcuf8wIe2CYV8NvYQKwCT9+GC28gqGgxfu60KBNzOsG+EyS15rb5SfDBRgcpkF
fx7WF035htAG1zQpSMROBnqgJ8ZNs+Fv2kp+um8MgU121Ke7qgT2MxNgJtN+72A0
oAmpwGleRPL1vjj+YNmHbe8NVYMUXyx/u/RgxTkMvqsepdJDaRuaFJRJth7CLLGW
Y1FWG78t1R1L/BRxh63KjUuRZwNuHaJVvkeR2QQ66CzoRjv7X1NzHLn1ihLeY5C8
UvAKeCphXBuPCiY1vYW/8DOp/FfneC849yPP+a2ATHp8uYvVUBk2Kfcl9s2jpjpx
IgBaCxRjQOXxBatBJasAGVBgz5tn1GVtj5ZzsCP3viift3m3geb0ZnAOlyaOezPS
E4T5vMfpaJ/HV5Ey01MMCEyasZfVJal15jA/2qnt7CPlE205uNl2u+9IQHykySbl
37CWsTWop7VgOhnpWRsN4cWf+jmEH0jGCkIvQA+j3CcW9Ehup5NiDzE+fM86eCio
iRr/lhPivOT/hWeQvYyEy8UTfX++vnPIYQWNDvVQRw9lUaBRY1roRwp70lenSmX6
NpA8GLzBFguSWwmC3SQuQMzOJcHOjbwpEb8EqfSSLTANNvyJd53xJgiKw1WdIYGQ
GGCuVST6MnOKHaSs7zqgGNt33yyf1a8pjqBqZdMc+9XXKXUMWMImPrPEjxb13qT4
fznIJteBoKPSbn2Td5z/PPrRdi/e4u8qUFPBVUjwHnFAEUU2nM6R8hNQusyoCgNx
WQ2AFF+nlsOxT9I1RB9WjDkJEzVutQTjXpftwy23SrIYCSksqnSJkXe3iCFnWiCQ
Gb/Nr2ftj/otRhpn60P6Vfs/9TI+4F9Sh9Tt7nhqGrWKEigrrIlYK5y8t5Y1IpjW
Sr4+SBnESXpGr2Ht/8JO+TfanV6oNIx0w8Vp/NPJLdGbwQwVk3hP2jEl8BNVmBZ+
tglCAkS3QHobLico5FFgLaLdGRMiPQnMRCIHt53kbMTGubaNEMMztMV4NZW9+oHV
/2Nb4bodtpYnCA7mdG+un0H/t3BB/JiFy4zcYq55jgmq5FhAp8U1AbBLKglfNAG7
GXtDpeZ7hB/sHXUBgzKsqVu/xJd1N0We2wb8BAJh+rb9ZJGzDKlHG7iIwLjg1fc4
+nBAkRAl5tLPxDn85ruFl+tJYEZD2wNsg+u8KpCRVI5avCqQbgXpXkXhkmfXGP8c
AH51mYpmurug+nKnMU3f8x/gSAacn7N6Vbi0W+txAEbEag1jBmPgpSr7Y3MutEQ/
UjJkTzjX0JwXDBwoXE1sQoaoNHKW8lvACzuDEjpNN4qCavGAVirsHjg2e3rCvn29
R1dzLWAVRAP2RopcY3bQ7OFGsoXbdGYYXy8OR5YwgpRG5MKgheL8keVJwlRORvBI
ce7akzIfp2POKQudtLC3/nipUgw1qouN04aucyVie3SQ9cLM0SfHlbyHG3ge+8Jk
LziXk8xVkavm1KFXvFUI+K7ocr4ZaJ0dPZYQtIFew5FGWq9yN2nE+mmwKXM4U6Vw
/kFNL+edQmXG8EAvEndz4kA90LCiiZdA6IRTcMa0NzbPylyOJ8FL764xFj3ZhWtk
DbY8yp8lqutMMkHmuHIMfbU3n6TudBzYYG0aHSpkdgJszpNrGtQa1yTQvOuSB5iZ
d42Uy8sGm3jdgUAuYbZDQEnNDKFUIKeCDD+tvJUZTOHv8g/Fr6J4RFYJ5tchkQLV
v/vhmIZrzgIeCPg95dkg/784ZsgfJDqx9i/BKKbPdq3Y2eNL5BMMvzZFfYx/Y0rh
IGNDG7lbEAuMqpV8QD0Jhf3IVHVL7KN/Oh15ZIQb7Dw6jRZJDxlycTPcAUKEuRuL
Qo1N6Eym0VXcaPgOUCJnhC3P1ZCJdGDqrKgapmaWVgDFZN91q2qvfR49TYNVTWL9
76Xmjgud+3wr6qRO8pXxpOWNPoyJ7JUPgon1no9oxo62aD8XyxhBoc/Z7nXkN8fW
niovW5OwetQofbhDCgi0Vp69uEUVACjdSdPzq/ATlKOsKcURedaM6tx9uBYXHKgB
ep+WNTlfbZH/09iE3yPnvgSMZWG1OWhWD7L74NSMkQKisB501/xUhJhrX+Q5Jftv
hzRv1Jv/zdkGlps/62YbQEZ82LydCWBnKq4m/1FmivuazS49t76HFAz29CqoLB1/
I56NpISJJYxYhaqMk4qlHA4QmyK/pA1+OFAjwLU8cUGlricVsgsimzmtAB6wHB72
EPdqA0E1lOlRntu7IG/2bk7Q9RiRRMZlBQlt9Bmt07w8leRcnWyMWOSNi90VRtbi
ic9b1UrBeH0RWXHFtDcyTvIQIsEfNAtFvcwp6f13ssk00D0ZiEGgUB90bZ5GwPAw
1nB3hS3fYe8H6Z7KS9R0yYaG0FmGYreeNFaZfTbs/c0J6pgtTuevxCHN/wTNL1Bv
kUxm+3DBxS7pSARWOQrdSyXCc0BQxiEFp4iWnSgcQtOONipLDWX0n9vHgV2GlpDj
uYMrS4sppEQLWE74ea5JJGtWHJWv+OliuD5f/kCZsKH3a8T4UU5QnOgk4kwBfmef
l+E98CGDF/+00OLj2WCxFJCjrvMj5gogyPu7zkg+fUgQsOa/3qJQ6MKPdQTJyczq
36nEgNIyTqRby0B/3TzEzNB99QC+7ZlfZ+azbsuIipj8cggWudbRbgQk5epjJ0QQ
ZqiigOsHqaFerXE7rjhwCPFDFrUsqcNySywAL4SMuwGiWKqhCaLtGaczCVuN0Dhl
5n3SRJrGLzLANUCPouAMxKQdqHbY9FfQ2wvrwY7UTtDFFOINI2qKEZwWpknDrUQ/
KhTc7egJOph0iiYom+mfAuUD2fTJI8nwG2n+k7ln7QEsPKRlOgWcLKgaaO6T5qdi
oBKI8UikQUj96d5cjb/ftOhNTikPEc9xEvxNNOtsaoEvg88GiCWPVEhjVRgO+T6c
CGzzDZedwKWMStrCUxsV3oFHF3EPH/tuVMXYhxK108DO9JnpPFkAPTwDlYerUKqS
SnqaL0bVArRSJ4kvS81i1S3ceHUO6HryMspofSwLK8F/zKFPP68Ta92pomhuMMtJ
YgtCfmlIE819VRL1paIf4GX8N95oxHX3Xk6HITvyivUCDXprdr7CNqdDHdrDRUp/
lfffuthy2BzHfqzX8c+XAFxcCR9zykFbDVOxhx5A8tUJLNzoisosxNyTDdp+2eb4
7+t/N1EV173qOo30YHjtbS0CS4jLhC48JQQy7BHCEwAKOIYsJYJgmwobY1Jp3i38
Dy2InRyXdXpGmCosCu3siVLS9M4aw463nPU/11yecxIslBCGrMLHe2IqOy7L0aak
lP7a7aARkLcM9ELcTTTREtNSn/3vygvyGdxW9rxKb6TSo4xtf8Fc1wyAUXTA0NR1
snYW9FYhESNEE+yq0ud2UPS/rL46aqm41foU5BlPgXqViIADJ5S2+KBqa+BaOIzN
kTrStogPX/M9OVxh5gWWvgd6IZnR15nVGSXgRj87PID/QMcxlKDetz7SuvZLD7SR
MtHnqQ/2M+kCFJGDG878xVDLM0wST1NCIJiJPWfty8t/5b8XuMpWn78nTsUQ6C79
nGVmFn3hpclsrxClmoRV+pPAEy1t5a1SqB961iLR7REtSEL4NOe/iCp2twK9U02V
bC6aSjpEut+MuDwOu5FOQkHhfr12TgTsU5balNYo70D7kbU4jzuiTA8RPXzYlFv0
f4U8nrrLcsHTuCJQrklwAlBjX0AnB5ohOH0kuuRmBISo3CaHBOe0lT+rpXAa01LG
3aWyfy4LBdNeLDRT7r74BGgHQxy0r0Dnaqwlzz1/B+knBlmjfb3EDUbxftpxqLz5
hGnAaLRYBF7GytA/dISIO1Ph2xXBfH8CBItKWZvOJTA7CK9RczBA6jk+lmqoNmJ/
CwXfSFp2icODejgA4KRzSv+VGxDUAB7WvE1kE2whu0hI43Hm0bqnUgfTtUvgeQ4W
ZmH1cTeEWl4lEx08P0fsl98q6e2zGo0STYzvWB7b6y3Nm9/ojmwWhCCTDO/j/EgL
oDYFE6GAFkQAVPc2I/ePekOo6tM6ijwbVTWtu7bl7dVJRByIdk0dPDZtxPeay34Q
v+DwjBZMQZb60pcOf38qKYim8JBTsfqKJuNp4jBZU3EUGtxHCo/USFQPPacVcix2
k+DGEWIiEHA255qKvLrKaiW6zsWUqjmxK5JTZ/u0jhFYo26exFJRba15hfxc0B4v
QxqTrtDKXpLM4lq6v34ruvlPtY4SjCJPQY4Qg8dAnleuYdp+F6F+ID4VDnnuCfTV
sNG9YtWuWUTR3hn1groKf/gf+VZS4382y8bR0lGuE8D+9RYZacxaF4rApL/bYtNE
LZOkYhe3DEJumDgLjeZV6okI65mxhB29qlkJy8eKsL8wAOX6ASmXZk3wVDAK8erv
tRkvPjnvq0hAmQqq7XkreH7kTlnCwnRKHwZ6XNqTKveCmSe+oAzjTnjTApdjzmfJ
x/eEIpBoA2T0i1hyb1ocWM7JQS4frD+LZTX3ssLpE35Sv4TKfijl0rg1WrFF/Qhi
jSgrK3DBc29idFntzAhVJzzEiIgepv7wilM/Bs2b3MzckHlcmRQNtxuQRa5SEP/x
LRHD/QJOuC9hXzZeq7X5Tn2hX9HzIi+xPAQ4H39mn3Fx3fg/BtfODJEc/10dBRM/
WxcZFnCioQStyilu0TJJfFLWZb1QCFLQ2Fk+Fxuie/GVZXVqzwFnmSFMLkfOcHEe
Fk3zF0bEWcgn+jj6F2Fkg9lP8rq43RRI2Bx7QOw99ajEAdwPRVWMDZtBZdK37cwo
cRzVQWYvm6LDL+jCrsBDDKzyDHyGtezXMdS1T1n10h9qVEjJ9bNBNNZxiLjMAe85
6H+IbSgLEqar904aPg7d/JNuZeYiY+60JH6rvVOivEFn77K7P4ufTFrBShFTAtsn
OE2XgVdaUXU6uBv5fmyc26yXmM3Dn+aLpowy8LYq5przCnn9MEfirwp2qiWwP9f1
uI/JsrWbZrUruw/qpk3O9dfQXMJ0T5J3fPeDPYw2LYlDR1coO8TR2HBhtWOjiER7
kQLCyOOVrylb8Y65QftdPhzJLU/hQyyvZE1Sw4QbBSmKRytWtuQPMWunTWWUrTYZ
tPOrWGALn/8wCrzivPUsS2jvlv9hM2oL8f8chUubQrr9sSEHlaXA2DmJvR5CJMPw
zhYlRUkLwZErwngxCMve7yqvIqlI0evGy8EsGq4UMxHIiQc3dJ4BfE7CravJKhCX
firDuynGYcOHKtwmO35OtiPZZcnhJZ7BhoIwQJQzZhWOYrBgLiUqA5wTyNEDeMH/
AI/Cnl8cxHyrt7ol6gxinDw/86+ViW5hkBQSo+1QusECcN/f29p69I2ZmmX4TEb4
+GFzieBunW7wYp55MBRVfIG/VOJCiaogzGRck+vA0qVt6UlklpLkJOxt+q14zIvP
2Y2GPlnq6JyrmdPEwcfvdwIJi5MF/qqqobpiFhRyW3LZKjixsUevJxryBVfDKPLd
TlLrj4lssMnvOKP+chMGPrkcZSsNcUx04ikgL/SCZsfWCpvHsUDewYK0x0Qq5fcb
hbVDA/Vb07Rx+oQEs2/xAhvhrXb0BRgxStdygVB1KEvY7Zw9jSmrnLtoX51pj3tz
7C7vuuEySZeEBOG/EtgrvmNsRldFjZhDT0myxjpH4neJBdxJioroPSRnvAzXmuHv
q2IOIBsTNs+kDJwXhIH9E84Ehp3gDrVqPy7j36ls5+Y+44Lur2OWwz1RLB96T0bl
wr8FnUiGjfLbMK3OGDD/CZICSFBT2LHg4fhCDf8YAq8/BgNaO9ZuZ8JsGdIanxP9
US17/nm5ghPULNpQrJcftniCTj4Wu8SmYrq9Psk2hXbV9+000liZf2+h8LXxuH7j
LMpLC/0ukZ5lqpr1uJ8HzrXRmRjuo/XevRwBrQXD4z1LLkPlf3iPISe6K4xz/9Xw
mgzLliKq8o2Qb+vIfeyMK4bFVPp5DOKCuQsKd9zxVl3KKKd2oM+mavCkcrZqxkAI
6kDP88jAOl8NLXjxyQho2N3WchJayWumzuYR8LomKKGLp6PNJzXETa78s8PuQWRV
R/W4UNbPBtm+mKQaDYTtLhU7pGOrKctWsYoqv+zin0Rw0rU5YmX+ufRjsQWeTWqK
8TerxtyYzpxH52Gmy5nqaH4SLsoYDN46NeOEq4BG/eyY/8IZQPKERkx27cW2aDt5
Wq06TnVI/riGYCcc53hIGf5aXCoXb6WKG/ZdMHkFTAg+8Tffopj5cVN9V9DLISaM
P69JJHzp/0nqJoyKCHfTTYu4mGnjB5a/UvQsYL1zckXKNl3gLi8pTnuAjkuVsBOc
z64TqBhezV1p5v2dcyJ427Bot1/Wvc9X7RQ7v00GoVa1qgc4iLVnje+mQtuL/PXr
eEiYAAsvzrhZyiu36lPpTlFSTzcEZ2ncgwQpTabttpNySjLbpGfKRcYwEOkCfBQP
CuxfTOpF8Qf32d/FFEZAhuMTqwsb3tZ5AslL0hZz68TDon29KcMB22n5dVqJefBt
eF/AnmnGfwpqdMo01pyHGJUB8T2HxeqroA01jUshG3K3xIrz5vnIw1Dl4JpBKqOq
2RMN+YdfPU8YlrdeS9xmrqZz5yRsOJUm2bpRtzlhp/lWeVggfuzemXpwmoKwyl0/
morUhX8dT60yX3y5t8GyxzGgX9s5wRu4JAUw0HIWhWgILQUt27WMihRhPOHGcDYk
Fmrh1v4gTviMICBDSkQ6UrYoEcEkCUy/abe5SNRx4ic+ZhBG29GCYbenWvSUc00n
E0NG6UWPHaFyahUcT0Rrh1JDBP4huR08h5O+J1UCfdYZJEhLqb4kscg3YxcOt7fb
FGasuoy3HYNPld4dy37fQmBSiGu5VwV/2F/ehAZD7bjytcpv02B5qqf4uOy+EpiW
HdwXlVUfbaVO6EkTuJDBCEypM2iUo5B8JxM95BNsVIExgIOKcMAAHARBxgGNuvEr
NspCMOnzSa4VFZUiiG1YId/EqwNeY+nq6HZjpAL6PkmaaFp8U6fRlx7NG+detE+S
KTxV0brl4O7Cn+lNq819hN2TT6cJYjr2ATsRZ3Fb8QJkhaMWoQlbeXJQtSagmKLs
wSOxtHRzs/5/dlLDuSIZxKKlbZxkS4KWA6xX2O9VMDh4eeq/Z41p3dRS8jilZrCw
SFqPBtg9pLBy12OCjWmlua3J9PE5qJ8FQMlpmHKJvD9Pa1K91s2YctpUpaZytfLd
p1VravvXoMMxWRoqkWANao/msk4M8/RSlmRZvvFucZhJYUn0SzOmRqYF/Zer9ukW
`pragma protect end_protected
