// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:01 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JYiQK7WkCIXR6UiIx0ngQodFDPju3RW+G1osE/rhun2Qsr5ghzvKXPJz1j77bT0g
pypVct/D5lmEkycc3qpJ/HRZDOTJfCNv5sjiYhl745mj/B1h4zWflw4FFW0D6YSU
HFFbRTCky3jEH+vm+fdGKBpKblmtcIfrp+C5KTFqqfY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3152)
kXfEK3xDGv6n1oygpO1RhtmVgynFpLV7pmf2/8MOt7gMGs5Zppvfe1yNyO6kJw/y
vfmoHvusSAhRsbMkypaFYWNj2UjRF8+DWEsbZhOpeIYOR/VElReFuDK48sRXXM8P
1CdUyNW+eE2SQI6uA54L2vZSHipOGDMwIFXviVKvRQbMlx5zv9a9QU4dwFWdeiGj
olfGynB4ph9ihtkY9e6if4mSarNCDy1GE+JtzPVi/mvUKQQJsuKhjrgNQKm8nPpb
18rsq+XyHAYiPjb434vMfSoUlIwGH/mBE9hoqS28faCB/C7Y93xFGkAGIjapUmlN
5Xrc3JV1d3KuDJv+5BvQsX3FbDGBl3FDT4UTg3FHBC4yOLRY4KoRQ8yYOfEr7X4w
k10AsSBAOAPTO0F+Ei5ppoEvxFH2wQhTs/RZuEBMjeH1wZHe/Bw9mfoOMrcbg1mi
18Rn2NVUtPQilNWXyupHCJYvFZDZbE6eCtmPA+y7nn8lu/IC7Jkg6pSt+zPaqJCl
dTFA/3+1E3/YasUIh+fEGpfgOuJczjdgOhFckGIQijr5PLrZ4QOk2mWcBbxZJTG7
m81RQoaJqnohTt33Tc7jU4mCpNFMZBzUZOOnjcoEYh+3lP/rTosmxxmBc/a9LMqG
2bjEhaRvCu321eJHzGpOHKeI4cMhXNL5LCDfxUPT/v6o5RJI2AbSPGjSaLB+E1yB
cDWRuDiyy4EK8DMwox1u1TRm0F/V4ZAWrR/hPBUEnNx3zSkP5bq9/vbSZ0ZbeOFA
kQPicoNgOuxicQ5sRSar4AFBLLI7crjt8w1zhSpsNkH/WJM7MFHvHRLjTVTfgIIN
yMxomjah8/O1/zFi9DDGPCeTNxz6QRLBllAWQLYlPKv8Y7z4AEHuGCG9cK9nIisj
CNigR2p3yWJWCpAqeOkqXJhim6oINFUH1yN0gxOZFgb2n6/5Rns4CdJK4Oj3D+qV
e+RVQdJSxsk21MI9K9HjHlmleSEst2/+P3L1JZxRl3qPfmxY4nAqtfxMzPeP/51W
eDplf3zDrAwjf1E3xRYbsUgWhfjgbuuSftCrn7xXsxgDxVlBbctUFu8UfYPOnnOE
yyZIneTQIFe0j9wa9xJqSiNsx940AWEfe5pGhiA8DpJ7HmZYqnkM3bAOlSVZb6eC
d+j5ijqE3fmEX7/VlNeLs+DZtKWDXA3TYJiLHdIcrQlafBQaoPkodoHix5WEeogw
8iosUQAiPjDGBkiI856dJLus+AVHjU9pV0TKCa+8ie7oBeRQOGgcRh2Ecu2A96wU
VMgXHoGG/cZkBYoygSjs0qTlvkF5xzk9/bTnh4yTW+fUBfOxZCKHS3wsthMk+n5X
PoC1fnOmsw9WYUP51byPH1m3VNMg4CUnOr7plm2uZO0hZWmLRTmW/gVUMHY3J3tF
hFJiTidfWovaEPdlGwiGbPL7esr9DVCaz/1awIoyeYMgYhPeuV1UcLylaHSBwHHM
GKCeHcnaGJHYHiKUtl5v7e6qM2y5+Yges81rQ6kCbtcEvWpPbDEJlWTdcWsvQoWs
G7GpjiWpAsD0w7zoHhXNdW96yxkbo80Vu+U1uEvwGnKj03OxyiEoN7jucyMw7Awj
gr9JahHqDGMVkaxxp/H8VS6oYwOSgg8xqsqZIn0mScc473ynIuEMvsJg31Cre26g
SaYRiT6i8BhMhB8rwf1UWWl9k8l+7As64Aj8JYRiYXyEvGJH27i5HD3YesggNzNA
H/VhrJV8fezSnfldM5jIrkt92oegWHb9lMsKonAS/+oKycbeClUsR4MmaQbvzhZP
9lSflAdEwN5lrOFX1RPsydhrYjJ4uZN8bWaNvWoH8ULQx/0PxMwKkQFXOFdo0BO3
0NHzNOyN/0pIY2dl72Kd4NEkrJeRK7k0pXqH7iDf11uBeL95mMb/1xW2XmnAziRD
tl/kPNThTxCg86bWCl7EN1LLStbkC77nzB3fkFy/gn/K8sDWQL0XRFMwfDKeb1uy
+1jvlMeeuiewu0medhHEZNE/E/6Fu6Fkpeo08Yyx1ngqcCEWuD4FmWgJeUWAEvSy
kRmd48e3xYfKTn5Tv1bfgS56/W/EEbbDssE1RpWTZZWNnyrBd/xX2AdkEM44+nWD
XcWN0vPuymBcggOrDlb8lYtY7sbOr5GftkEYVEk4JU1Yy7ef1ZbJXO2JauODI7B9
MgIwykEoInnxQAJz+179YchoYafl5++J7gzkbjJ4SCjvb6WPTnhBZji1Mf7FqYUS
yMrGMAk0ESajnZbg9hkArTdUr7UVy2OsboDwTceilE4pgRHt6SWZvBXlhlc2GVik
5KHhIgI2S3aJT/eSAR8jYOU3BAyQW1c5NpqEZC0HYIk3RIMmexjAxwn/ibIZchMH
o3Lv7BWFRdmwnKIxD4FQ9LYjaxHOCr6DTcj+tLnlNKvMx4cR6xE2ydq6JdcPED/E
39SGwbUGSKtx3dhxnibYrncY4W6R799fYe3K3Zi9m9OvokArvAO2CYEX7FoSI4RW
LM2MVAFDMXo2dAC9P3cU54bQdd5tIZX5MtgAJBGLLyhCvw7fi86vpIRbBbfmpXx2
VPytiBjZBehqBLYiW3ydQZlR7kWfd0Uf33r6uZ/x1WI5lRFe37Pbcp1LU5i1GB8s
5xUQvrh6vzflbvO2VxZt+/EQ7dxJcUqTvlKZSWWSZEitwOogu69pZcxoT+FFIgAz
XHYYfSpnCPiOz8h511s69gY8hzeV/0jLc5BkvVC8fhSa0eZaT/cI4NbY7I519lYa
OmvoidFHNC5ja4ICNzN7wMf1iWWXz3n5ZVZTs/Paax/IvgicyA91gA22FIyJ20Qh
DH72Ta5kGKF6QS6sDS1mzKgRfeK4U/yVXeLxkQjbvP8uRDanHMUD93+SCm6Cw0kN
N8GCwHqJ7X+vMH4C7lA08fvgPiOb3NBLdCjcqoAY9qOmlBeXtVvU8LO3TIeZ3/bR
z6Wx2omC07DjgxUMKWEO+Iz9dJ8OZA7Hj4HEztUDGrxLiaVN5AZIGeqb5thbi9Gj
+fBTS12ZuuJF+pmpVyxIjdXtu9gbjk5G8FXnLzbVIFZkeYIqLp+GN2gQqnfME/fb
ZeQo1JzdUD9hicKOApfIWIvfWl9JU9q/3lLoZDCziG5b0Imd1uJ8GW07MTkSWKdN
OPYgRkFh47cT9QHZG84rcKtqclZehcRnDVzku2v+Js7vqs/UJ20mo5Wsmx6kRQ0f
ReNabq1+0sioaPKUw9ZbZlH63FkeAFGuM2H/r+F5UlC2aMB67OB263Dh9fHljRfq
ig+5ARsjU1PqulwI5vnhVHMjS1HXoMwolMjg9FPPwvYKF19+sRtbyPNiZqkV7lPV
b0Zs1yU/vdfBy5E2lNJ1xkHs93a+vaY9qT9y4rOHbCuMj2e/eO5tSpHkTVWvplt9
GTQjC6a516l8fnv2rweRz0texJKqjzFA6vQ4Am5YeZgEVqwygf+RxqRBHC3vdI3O
gIZG1yRYq3OY7Qhfk/+rDN5cwANfLtm17iwQX6u3k/bwRa7V/rhAvCKzhkGn23gP
AS1mazOjDxnMw1NadXZOPEx292Oe84y2NxJKNADFB/Gkb1dn/47dzWkAJUjeaZ6p
xYUin0A/6ciBC/FYiSZGzoIbtXAxPyi9zoiiuLCRHzSvPpIWmV3/ugpVSKwG/7Y5
Nqmsr6JwusBEMo3qdZAtNzQ4Rrw38782ble0gnXRB+S2R38vR2Hrz9OFaCpT1VVn
SHNd9Fo/2i2EemrEbpHQw893e1q4mrx0Xv+Hod7pnrYBwrbmWZDGCPxXTZZFc66g
mc9qKQ4cxLj50P+uTLWa7L3YRug669Xnyhmk1vlVqnMvb4C95ra2GFIE1VX13N8q
xfORSTHn74j9Fmxql/cX3niqhSTn10ps8Pd0508upT7SUowuTsCd8Sdw5NS50siy
oPkNW141C3YLFTfQkM9UEkoDyhwXYgwiILsge9By0CIveBmfUqy50Esrj7Dk3tYQ
mplKi8AxxxMqhmZO8+3yNFDApxrnElxb681EjVFRdSi5E/AHzl4jhMWxlYGHaHIs
1fh34bcAYfXpoaJHnd2/N3uaijHiFgGcotU1b8t6igumltEisdS/5tVo9KTr+iI8
trUA1V5J5PaHAWqUSH39Y5J4/Yk0I7tX/UoV/cfwpfO5kCxhnZbyU/S4KSR71ivo
3T+l4Frm/iLDj5KAWItcIG0HySuCOty+07SusRmDbkw=
`pragma protect end_protected
