// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:28 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ciMFaTF1NRvpWAeW9WtnyMblacGPB8d5nYoXaA7KcvSQaOlNDbV33CG6a7USeVwp
kWDR7GirY7K7b7OXWB0w0kq7yXLYvKx7m2lSFbtnJDbhFxtF7ez6s2ILnYQrxYB2
CslKLIq3ehl1SWX3BeAMOuOu+yLYLWP7KKSGPkAP7V8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35312)
LSe7QyDenC/TqNSlvqi7Y4WNjPK19CKuS5ZCizfVxqcMK/PP//jFeBYEpgyK9z6q
IhlaHASWV38uYejgKX7Du709FlwwQ6U70v71A1eXj/XtyNfNB7hl5fYZ/m0WW49i
M13nHdxNO9dA++CxskHumUBRbhgRftMGDpmULA96nlk0G90z4A+Tq4iXhwOAv7Qp
pbecOrpj3Ay2kSDL5hx+qOakptP/R+c344X73fSVyarUAULzff5lyIzX8+6QG6cf
14pt8kofjP5lLMzVmCrsaFPeYWtfVzx0eKfWVyNFoXTuU3AsGHiBSuBWV0JClXg+
nhttZqKD/zY8FHF6ropUOESAERebhGCUAOV83oB6RDWM+fXvlFEQ74jY+eSo3CR6
fZXQtxLT8sEU8cwn7ltD3x18ea7Cowp/4st8kFemvv/2Axu11hc4o6UcEcpJsa0V
uERL4iBMtgoycZ86Bit/z83ZSa3Q25DFunSbOInDQyJgcpXZr2FcojST7AVmLeaH
R35Mnfmen5L9rQgKhlbYQPNl52ieKc9j78gF0UbmxFze6eTPak0/aHEwGQQmNrt1
7GesSXlx1M7s/apBlDgmlFt8nqHCAdjxZwY3nXCnoOh+RkIv9HKl8jWQJI0vI1Om
bFGae5TwTtvkRRTwxVLNsErpCz0uM3e19gmJvTj9cqY2kLRpb+nTlhN4ck7k/Jc2
S6LtML77vLkEs1FgTJWLnOzCdK2JuXjzNwe0LoOaLVnDtrPWpgWT8GBPwFFlr1yV
Zjswt/qV/0etG17efpUgxBVivWWJ2r3TRLFlik6maiveqmsXYrwFywAkjxyYiJFp
u14M1XdbdtfxzkqJsUhIXLvinGu/ky9s858IMaigtaujPmbsS3iI4XjLT69VNZTX
pmvpCAd18MzyG3nMB7Wc+0qC7nwDoXKq8qHO0gQr137H7NMJyQJYP1Puyfw/T3Q5
OHcI6At3ip+GwUqwNcZVnplUEKPj+ZYdw9MrQSgdf+sn9p7MOPU9KNjieVhFAl+/
UmVFguLVr6+bvceS4Vl4hlNB3BiBKbY7E+SjWPavI0kd1OILfrnkkWT5RG3g1MMv
itlpxzD7/R3IN6q5Gxb+BjEZw3T4aGavCD4Z95OOz8zoccUf/CHgDyBS9h1Ryh/K
pSjjc2LWuA/I10ogyWQPq944Qf07r173jkDAVk5p9+iJY5Ihhdeb/1iiqHOsoUMx
qCGRw/1YiUuupgl5UBFdwktwj9KTXQrAU2AArpn2Ae138h8M/2Km8F+MC+yeYqfw
JYAo5xuuppZvEr8N2vECQn6Jb0Inwg3axFUe+PDqb7o/JCP5P+eXa9TH/tYyGWKg
AioaKEFRt1Cs6M3ax6gmj6IS0J/Wx0bJD54maLNp8oEL/FDe1TIiHPLJ/NQxtSWl
rverjPVM1blDLW8B5/Kx5A2XZGE7D5Y/QAwB/5CCVMvt0JxON6AHcEeuv0XCJ+gM
nAASMeY+mE6RQrMjDMtY0AA5d/zF0ZNqN+OK8qSqsGb3ju47qOhvVWpDQGRfTELc
L6OWCEUZ2BKnDhQyZVc3m//q7QHQFehtyqcPhYeZScJ3yzWlU8YrkbqXzPHF/UZk
IEFfQWRpm12VCtzxT2NxtGL6SiOWxwNm3GBHCJtWarLnp5h3MUxEEhb1N7kcoyUm
OArMpyP0nK3Z83m5Ulb+cJFup66CNWgz1VZ1kulnXuUm3lV5nlC6SvxMc2wv6cXZ
bYo8TR5nf8xry7OF3L3XK0umUhpqq7p2dFGlfcEmOHRvdgSB/PwwFOV7QXKS4Gp5
D+8jSkhOFwjVXG4zObX9eyWV1LG88DdE0YbmGcTM+CiSdaGZr9GcfVFn4xo4Cnb9
UEHT+Mv2meGzSY5SS/135htb8zTi6dwoBBSXziC+kZitiEBkZxSrNo6qq8iUKsfO
zXf+68sqOe3VL6vRRV63RKSzt6RBuhhqwkIaJv/mlgiVwnM+q+4/yvznREw1pClF
TDGKewev58nQfcLwdkLanTbUSyZ3ez5yrPFmkiyIWD0ZwhDZF1hxGqLuMCztoSTU
1KN5NjhPXwVXOZQeMdg/+qgBWFwOHjT9oFwQ38yYBtrRcIJOJlTh2uFStIyos8iq
23DOgfA53eAObIph3FcAxrIbZyyUUZrSmwtEj1azSy5XwCULT2sW3x/LNu2ZSseF
bWe723xFvHfyLDTEJ5ltzasolZm+hHFdY+rAJVwMvDntukvU1f9Xh4eEuLZG0aup
TrH4ysezOhHnUUTq+yHOM7zfnpGg73dW/8+xOgwCATb21toWiZDKx1H5pJzIm9uc
SNc3JR/OCONtt9P4hI2+8lejsQG6jVkT/oQ4PdgXCeHHSm8Uun4NSkOyl67Feg3z
tdrvodXR+o89fDsuDxC7Ig6usHZO52qtaVv9QAr5L2tvlpQ5L0UMbD5l01tveapN
bLAr25TVLH41xHl3clXpxNAsGFhjELIY3c8HyUZejjoJY9S0ZsANbqxrbJy2YdP6
ZVtbzHkovXu8aMDFviE6Pj12sF2MANB7c0+eKehJgegHw/1EkOG1zNBTlLFcbdnq
vGRy2AAkGjfbjl4PTnY546/pqTJxCla8m8tocueCRcG1/7WGn8QhHdttnNMGCm/J
G/waPT5cPqjewnvlSG0KB7rhS5p9zuUIV2VLF8wTrcV8P0Eqrfd4YCzGbJ0GtV81
zT6tKyrHBqtKfJh6ZUjWm7lm37HowvBbJ+8reETwssqDv2VNnQnjxckwGEqT7X+U
7/tVTUF3EKPck/BouRTMHQeL3HjpXzEAahC9pO8FUuEM7ByBTXeDZLTmq/UB45Fx
eHhpn4Aw9ibIFyKw1ww+0yVz96IxbfiXoPYxBDFi6Q+8GCWXeWl1PqOCPABECKR7
Sl0ivfdT8gihTgGRLMNardK68rwvM6biIFXzENl6FOzRS/L8/6+rDgjC4nnS1jaE
/U8SC7YHSlZaV6XiBKm0upkE6+N99YaDrfxJJsTMbVS4Eri0n83UZtNH/gftqI6n
ql8EfRVFwFs009FRuGjII6YMOI9PX0sH5qwPaxqMsRaW5fuo0tX2Gom7HNMSp4d+
XVqrSC2sMixW9TslyyK1cJloUDQ8pcMB53RkEaYjnwo64jsXv/LttQEi54JCInQx
6gBB8V89oBEP2zvfiauvP9plkOE1Js8d7hKUryv7nhZColzDcdQSysHfdEomRLwS
b87VZTqZ11IBSCkyJwDvOVHFXfI2hxe36uKl9MTFCAefmGw3BVdSqYee9d3DGZJB
u8cF/GyDXCGiU65+p+dRh4/KW78xp2uX3e8w9I706ZJ2TbT2a1oMZ6WPYDSMszIp
PpRLR4NQbkm3nC9Bfj4z+Wco6/fe9QaciJXN3HF+a+obd0lIsia1yDFz12Qu/CAh
j5uX4rcsUlpBQi+RjEP26h2a4yW9b1rY8Ai//6RriyCKllGXGTUTAxzRw58hBBni
LkuBfhB5jMhaIZIisi55X0qpDcwlxjRt87pIEosSodHj59jMkvWqPOZcaRCFqE7r
qGqWhpu9wbUQxbjjOdu0tn9GA1Tv8p8VGUVPtw8tNE0MNKgnzH3RRpEsQ9scv4un
F+sIl07b4yTKFry9872CvYH6UmunxuGs7wejvOv/ffHVJmwtVBDwvYN0t+LZJdPq
dHPe/Grdy9S2NoUtBhpj9r1Bh/VV6fqdSG18hnV6gBavf88K5RWdkjwhIecD6YKk
EgWljDJYYLE10aSaXcMsKwVp/+ZLWEyOHzn8wqH4jjMroCpNrWXEMp72v0nutxZG
AepMQehHQnakD1BVnb8zsSkF4AlKj0gHdxI6A5Wv6MNH1EQX1HFYo4YUWBuWi4qi
BG/vgkRtYa9ZC7/4GwSZc/4UnPdyQQO3VVxLQFYFToqX6siLjHZODGKTZ6kzL75+
Nvly4RA1xEtOHbOXUC0AXdUVjFe34cBOcyKptRxcPKde45jKv9tmhgiX0E1R4Zkq
8Z3SmzBGQTDHjHHwWag2DTP1wULX+fDZCO+A+YxvfwmnpzdmH3TqhbQHjJ5Di2wU
sRmvDhPQuNiihme2bUEIL4JZt6nBsOfoZod3OqFJsDwfldTWWjDFDAkSyP4yuikW
lvoAJ1s0FXbY3saicPF5Kk9F0/GRRadaxUWe8xsVkLlxKyyvCfgMKDu2r8r9Gm9r
dQkLvejY4smOdJ2G3LmqUY2cZf9XP5btbx+Db1AsbL4TdYZRMMrIlWog//lKbtfI
OqPiBpI0OPK1q/vUBioXfytavPC8U2qlWuphwViiEji1R9ttK1//LDYLxlxn5xmw
a9BnbvLrdKegKi3oxd/q34b+GIAxgufSmfkADs+rsyGyl9weTSyiabecBigIS8/T
LJVFQWeZjGZxK0yXR0gFL5fpWbjJhM7JFH3sqZQL0aYyRvln3zFi7b6aoaaWHnVs
XWriq3A6DmDy5X6ml4TKpu4sWYz/YksxIDVrMEv3evKyBmmjIdPBoAlSujXurM8c
mrXww9zXiMpSQ3WUq5gNz8nDMKF738jKWx2tfnirzBwqnX1eNmtzRzX8WK79yhy8
+1sgc7keWxv342yl2k3GZDN1Ci5oOUcCjU1rpZ2M1jfeRQZc1Y6skU9RDPN4OODN
UFH7+hrrVkZqK3fi8dEbU74Cjr1QxAZBXH6rVLT1stSzCS1e20EMTkSi0HTF22cb
zI147N5/nR8ioozDwScs4RAaDZTgD7CzC3iCg0h4W5C/6J8fvWoOiRcAlHMQOBww
It4ODF++qqQGuf1MIQ2HYR6PcNhXJ3ME6ywTUsm9C7S5H1tObFB03FzW1jJ5Tg3G
E8v9dsLH85gTWyvtYT0VL7SGPQv8hDN6A3C0eYzfs9XYmGWZAaeYnhSplwxiElhn
AvwFb4eoWwh5mOcHwXNevf47NsRyDAGwHyDQQyHauhMM/LhyAfLz3b13sToQDD/x
MR9ctgzbWE7c4T/bDDNK3eHoerNxNLY4StbA6fudw9R+kHkVhUaISHeA6lUji4ni
5E5KA1tBpiitDyn6wMO/HJ1fcrao1pT56vyLAO9/bpDj2C3VneSw6bN6XEjinZpi
nwFayK5zyW6uATxY785IhgZOSpU2/aM6ACUiGPSnJx/nnfm9zlYh8zt0xaR4U4/D
fgcJQRDTcRSmegaKjpnpwXMuR5nYtxpysifdo/OtPr4trDwkWLBwklfIcp4iEHn0
GJJ7yb/CoIoFldrm9viu3pIsClvfL0LuI5GW3SLcck9OpqbVzISMRhDPvVxSFjLA
XvGPIQpJi+Adu71fQHfnDODM3l4ZqirC0fi2RhjalpsAuhChqVfNLtfU0aDn77dv
qUhV8dRNeI1uQqb0SKlXSvNxYvnSr82kkn/lW3JCSHiERU3NM91f4+dXSpWcgjQR
DoRVfGMxOafcWDZp9k1jE0Fizkua1K2z9H99xrpJPriRdvbj9TWGv4f+TRK3kOk3
5aH1eInRR8NcX5uCusxBNuH0KI1WxfzrLmElHesu3yiy25C6IOmSdERnheFqMUnn
vO9XQNNRwjZqsKCALfolV33U2PFGv5H7ESxcdrT9DLRwi9ekN/PUENVZOna2YbHN
jwxC+ylmTaNT4e5aBlB4OrQV9BSJ2bFHRdQbgmEKmuC51WbWVAA7GMCAAUQsXHFY
0FV2FO5ciwivVG5iwDtSf/wH68XE1mwo/yR3AMrFFU86GME9H5uWMnomydb/8Tb0
d+N0u/V+uHXBHY+Thg9ihsRrObALsEDAIXd4/usGUDlRO0Y47fbtJybEE9r7ISPm
mk5XInFWaDgq51mbLYAs7MT8N4sCIvmFnIQl5JEZmPZbPAyU6hvoaJHeX4trMDNP
L1nRSq/gcdlbZ9IUhjx2hG1vAxefq67w5cMuMw5ImgrbYhG/ieddRMOuGXC7947L
q4KIAgQuAS9HRbNaZshLEI2xvRJKtOpU2py3QvTKWmwPTxzPp1jM6gsIrRkZFQ5z
j3qNYImsRV+lvpck/mK0ZfYocjTvKC4O9Ze+kXXdGKTra/7EuRt8OAQov0oM3mh5
/+Esd40lcGrURkqonwnA1Vfb8bRs12U11GGrXyg5cSLgx9xwbFG98Rre+Qb/hppg
beCUjsAr4cqiRdO2h3nvBJkgRtHTyy/oQUuY4L4g9KEf60Y8SkZeSSeHtIFZs0R+
KCQMfC+BpL0B8xsi/GNrjwc8nT+CZj2BvludpMmDiGV2dsO3DbSXmRyLQok2iOaO
bWphdOF82/FJvSGqVZrFpeNHOdz8oPvRWRZ0CdmNrH1QnUR13XY61KvyBpnlAI6S
klX5aL/4AYF70njS2I77/QzehNoWiJXROwUD+8yRbuuim7vUrpdTD7IitvRcB40Y
0EFd4CfsH1LCxJVnt3+j241DPW5sFpUCQUMZE7x/vsDOIN3ljmQrcKj18Y3eOnq3
mjp3raTlVy8YrEbP18BVe+TiuRU7mbtFkJEbCz+Ha/HrI4Gwz+JRytDAMDzf1hnh
7Ik3xx1lyRy7pW4Vrra/f6uQZS3aZle/aMvS2sPxfyGA7B8WqF6WG3uORRb410X7
3igTDXZc2PJSKStL07tyDxy5DsbsxAZGl94hfEeISNoYSmVDB64Z+sREyxRbZJv0
UcmmeX5pm9dVYN3Ht8A/WVe4UnwUyZHk84sfZKVKxOLDSkYbvmcvTfPkoBrVn2Se
D8MhMRdYZCjUcg7jFvChJc1YLnCZRmGt4agMr8WcWjunPy1IaiVI2zenVWvI4KbE
TXWGv7zrTwiwCNqYTcQZctCKlqdJwg3XEWGCjEfB2935TP46CV2omhoErQG3UMAF
2881RCMi3HROVIhdp9NDbTyJMvbyLKUUFPr+9ugWT3+pixz6bBDar8ge3YLczDr7
Glel+h5bETDzHwFhqmVSY/qtywGtI0Ws0gwCZJk4NZP+O05/pG82iP9SlARJNuNv
aQODVg2gR7w6pg9q0K1/H31w431WnuyF0wG0TeWUGcsDnpSGuiNqOpiCmfMa9Bdm
R5lKctDG/UVdRpyKqlebunabNyiwr2EBd0Kq+oug3WMB36pnM5eePHCn+9SW51ln
wYY1AHAx0cT+kRx9ax/6W3+mkEVCwOwCvYnCwErM5i8bHCa4JY/3jg0PE9qIRVAO
nl2BgTZCWCxIH6CsTRbOsih9oM1PmP+UwE+PFSmGkxlQ2JUHM5E4gsskhgm/WJ79
qv9l2MGf563c+5CVgKt5mY3q+7+oBQrGxTFi8PXF9HJpY6Edosw9P03nfZGXrwsC
9gYQHwMXnHE/hce0hummGfIqj3Zh/BVEQzrZjREtLOeD5w/Bdk7ap89/dYNo+QOR
TLFl3r+imUHlcfj19m55hYmh2YCbCYimJH/E+joUeoCzMse9lItjCaQ6S+jWL5MN
RDVSLrinCl5x8gUv4uprYuA5MKJxaJDT3NzKqqLiyAwDqkkhIKZYCagT7gwBuyev
6iD6akD7opbDrKI1u189Qo4z8q3PNGIFMnZK+TPKjey1v51dgsTkYVn5LEgtOkRY
GZSnB3XdJXH+wsDkaKWwtYNNgkGdHqvRznzpR8KMFzEqSd2GSssCmtgyGR5lK0va
QjkSWDGt2GRSzXrEOGOxf44F9Hs3nd1TloIVTWj/eL1llCxtwjxguGbk9A3tDqJT
TimHQHry+J9dcOG9B+I+dviWKB26roQXgYBB/PALRvSu27ZypMzzmzjboS5vgjrn
OKVA/xedS20DyfMwFdUzmwrbT6WFuoC0/oXL/SbnEcNY3A/+mOJa0TtO1vwKcHZ0
WG4Fc9SdOW5FblyBAjMKDcLFsnf84WphuKCFddPl8mRwkux9V8zE4BA1Jgr3A8nb
tBUYdok2ZjP8kOaBvKXCNEsXexpXaGyC8qYjdvZfFsjVw1ojxEdBI9s5o+4CIwUW
AGiBLsaEoAUCgX06RjOiNQm0G9kRsknvCooJxJAfhPc11RlG5ZG5AOfGb4FIAhyz
JQIpqw7v4oyzNseiOwsYSrmhECfz792NBVV0n7jlI6ewwPBW5wdhrETqPjsYaQeL
GBkfK32nbOMdZE6/iVBpTJ0WnSxSvQ9bs0DtWEFpbEmlYiUiF9OWrOLpYJs56H97
e/xF71OIfAaqmQrIdbjpEUG/ik+TNsVc/O/QotsU+wY90U810xtJCrus3Ki+c9vn
Qf+IbVpK5C6BPHaJwVNenmi19KMYBGzZT8G6vBf/Wo7emwDrfoLvNnsyfEHZ/fia
rqoUR+7mm7sHvwQySjt8CVt79of5qAXRCgtbQ/hivU6pk5f79mlqmzL7r95/Rmkw
4OX3Z3CidR/I4qjHmyMhgY0h/tTGbaAbG5vo72Me5+hjQYR3cxNqVYitg8O7fzQO
4vHduUZWDYmhSMsU9QE5R7jB+L+Yl6AyGVGVOBO1oGAuUnb09uhR2OPGf2braRWy
26UD0ERTp8wlNX0MN1VuJ7/90TbzrKYfJ7DzsSOKsz3yi3LNcuVCzeRJljmGIlvd
SpSJ6nRR4T15iOUMJa83r+FNNQKy2ZaJHfHH/KVYjbK/irGaURyCcMUalhFfw3nj
0Ig6vfV12fVLP5IxOov0k6s4Ue7DiCkQeBxFhSNh/UliuqMH0zd9HxxzZUT5SiQT
FyNbJMZMQJoAzwlf//y/IZrQ2KEtWSgGMDES9W/ZzBlfQEA7uTmfSHweAhwO03V4
Z4DvyWhLE9bKjqeil7NvJjfnI4Axodx3SbGFhNibKv5Akvw/cjOdGSAmfTQPpv+p
0f6B+wtedK67hXckJvt/j31nrHmC6eSQINFdGuEYzHC6cXvzNvaQNBDalk7HeE4L
4TLUK7ST29ILlYndKbcEXjNC0K53bYq+Hmwr0aUHnNRvue8Wp8JdJOpYEYfuMcC2
0B8pia3eCyO3eZJh5a/KEcBtJHmGjy5mGBpB3N2C7YxDXCkqiZUNW7s7CcQRC+mA
aZR1IRvzOhCUyimRn/m39gJL+Dq1cKvEYp3ucDxAtM77AirExEjyBCuJEIVoyjQO
s1aE/PtrEn9WvVV7/vcWDiTszkOrNG0z9MH6h7uwiXNH7FntsHW6dAoO8xSaAiqU
4bNocXerqvpZ8zCUP90bDbrBSQY0ZCmOCHpmQ9L/uE8TRVNdQLHQfy6cIvibu6C3
UCkn0ngmmYT/eXYPo9ySGFw5OeFG71WhidrAWKhtcgVnuRo+Ew/BPaQX4XwZIy0s
wmb88IYl1zdPsInQiZ8b65NzP3qo+D1/2aIlGmjFxPfldaQL53xTxxK0hcgsX0LU
a5Mb2SNTs+viSxIA7PqKrxvRbmmk5irRzmL4w7AHK8S5gruqzBB9CtxUavnUDp6a
fS7HuXI+x30ZbooAFFn2bT7d22y+3l8JORx24doKhWzJfQe5fBMZakOuA81P7DRb
VQRO5MCtSjixjd8VdvquRMKdoS9si7J+YOHXhH6yRJ7Yfnbfn5JXHqth/ifGOTYu
WXb1DCTETuC0Uxhrw7kBaHj+5Qq30UeyjtUGXuarErLA/IcKniAJYzhBYewSW2JX
1OyRgIey/7J6M8dSPCiU62qN6JMWRegixHa+Yy1iPP7bHfcQB7pmCbTYEjVmSMH0
x0MG/jMir1l/++WpQfnmt2mW7G3Xb2pn5IjqgsEomGqqFAC8SIAom8MZk9OLP3l4
b4xtqadpkkel9/1Pwcit40gIt9KNt4+sM+beSt7cJJDG7kV473g1fQDcmOfynWY0
qVT8gS3dDRUPpQhBORWcVuzvPy4Mc0wLtjqcAvnJyNC1R+ULQSaQibjuPclfgO1F
/QgcIu8OOKECcwOujs16k0SZHKmb0aXjASLnHg+uh7cVN+TqsV1lJ/H7Orr/yLMt
1b+wImAgGfAfj4hTdkONKPQpkpqL18qNwnZjm2HYScsTHUWTyWuOI3nYZ6RXfEcm
XmzWcIzKW3NcLm5B/9tbRNGnz2OiaFHrK7B24ZmstpsyMnUonEJvnKDkcWefYFak
avgpYGgPkDvU3B8cQc0t3Dd8wXBDgv9WjOGP46L1LQnkLc3+/Zgr25V42fZ40M4h
IDv/QX92vIj+R1KB3hTO+30+p+D5+zP58MAdGth6Be2AiZJ0JpuyVaxDMPOQB3mr
SG0Yym+jWG5KD4xkHXdWtrbMISJBrnZeObhzuT0pnFfNC62WSDUSHH25U7TkEM5o
RN5CH8kVPrs2LzibDDBjXvVubhj2EWrPTfQ71cl1tKxaMenjLwP2GMBlTNcep5V7
GkXIj3GF8EKrbdfbHPTDLL7pnmrYBBPnSPcGmsUGg9zos/oKj384Ve72zpFpFvze
74QTNAfBa6cO2MZ0h4ymO6I3u4KmNRxRzTkFtXlvj6p0RwQBRUeOGnxhNo1svvnM
t7gqQH2B1lMnyuSGUtglm3U2qc9Ooqnxt5BnkKUWUpYKS7VW5wYCx3YxD7+DAthB
RUqb+IfKi9drELz8nQ5QMmhHTXSZx+9rQoy3RlSvM2ON0EELFvj23e6XDviSL/0Q
mBDvgznx7Qkqam9vYZhaSq+m+gxS6h3sjkBeJBM6J/I40HSpY6WuYr9jZF6NZzvC
aoZGbShTCjaqvod/Ti3S4cvtmd7h3g5R5Dx6TjVoy987ygMWon+WAY3szVNaa0F0
i7eKMqBQyMkgHIhtBf9uFAEPM8ByLvyqV3hTNvxI21HJsIYTu5bT9GBcOpgIjULp
CX8VOnuhmmxCJvvAwuIrkWj1A/QoNtvqdDTvByBsUvNIaPD/2FRZZhl7unvAhi77
1kNufRjS35t9BCJHkokou87vkWd93MHpHKcTH/DRuDMMT65ohgypijwFMQ60atHU
LPnnaOlNGwi7Ui9K0W2m3rBs4rh/eDwo451WJUq3Hni4WVYPaYFEA8fstVf/2zQ4
TT2yZnWjngewR7tsOxsx2E56ZeCBBXFA9lTvhXwORE2yq7Uu543fq1PKuCuaBaqF
RTyVDTRP64axXtxCvCz83me6hVQU94uQGPP6BU6L2dPR0sGgaE2yg9fcHjkLjKwG
hxFhbXzEIkJh+NreIZmzuGkQHCU6YUZIkqJlzASBiyhw2QQ4QByOGhbHS+jvuWAN
PtTYvCwwsNjSs6bbhjJg9g7fVRhHb7J+XZRy7XG8/UnNwcy2G0D5b+4AT0Ex+LiK
eBOTbSxnuJ9eDvC6lad6tDiUd/LvroS9oZC5SUazllvWeMz1mxPcUfTTTzZHWoCl
xS/NqbKv3QBTQPkDKWR2QgiDP1+NS84x1h5cbewvZDXbeTAyWx2inVBn5Z1QC+l8
x20qTcUltRrOpNfqW5Af+rsWriGLtxvVcoODmKO6xCrWwtDedOLB5CIC6d4Gbc+o
+i0Q74/X63cx8aV1w4GY5rnRHwANUDdck6KLR/NZNfI8GVqwRyh4+rcZi53l0dO4
gosbMSMUeG6Hs6qfpF+lRrMuH+2AXInNteg7nPLNRuvbEOASKPzP3JMy0fzg8d1X
mXryAB9yo/cSh9SpmyE2FoyGI0VaeRjw0tTfwQi9zLUBtpjRTzdU3aWfLI6dckEt
3F0htAWAuTJJtQ5QAr8aBfgmH5ezYf7EuZ2KcZDfgsZsleY/XH/8fE7vL88uYNn6
O7hTe/1imUDQIIyOsuURFiRVug8/yIMBSY1wkO1b6jyUcuPbkKCTgW0wvNC5bbAO
bChofPSZkfCDhGdQKbvlPNN2CBLxa0DLW1ngjfGa7f7EfwuD0/onNvz7x1aF/f80
/0AKLyJnsd7kNikCHmHcS5zwH9q79tmKTLWk5jpugscrjs7mvxRMNjivSVJIhuU3
8wa+iYCPYMPlqQssEgKVxf92+w5Gei/xalNLbeRzAX5stb4tFz0bvvAMok9Q3AuQ
3zb48mubqqCwnJGpFxPNBIbzSPmdJxnNvBDEP6ljks9xkJ9rkgx59uxrL6HGDnx+
OmJENeDb6plikVhpQCAbgZ5nve6VFxz6v7ESocpv6R1GlyB/LI6ZeNrBddrsi4Mn
fSladONodNHK5GTFUH3KG9XU/dONH+su15q31LIBTkTToQWvgnaYbuWMhX4cfT76
elT4pRs9pRzAy9rtOkC9p2YFgq0NfYnT5Wu6dfemerwMNpyz+vav5+HUI57g4jmi
+ukhXOEdDoWkjo+Hoy/WhlsgXq1ZYFkboeeqYJK/ov7OxFXkKNPUwi+MRCzlOxxL
ropmuEeqvyoxtD9IG/9dLHaHgRYXRdGbyq5R54kxdBtwQJFXMDFDvzP2vLXvRZm+
iVRmAcwa/d3aJTJETEwNjOuTU4DJ7YW1mRBrJAAY6WizqNxs0kCiFiTezBJehFQJ
e2nRBT/B0QRPBjzS0FDVqEEEMf9ZJFKgIlrutzvxols9dHtI1ExuYN/yj2qIZNsj
2FL5pOVLxe9A1V9XCaeIwYfCquCgAA9EliYpII1Unfbt3FAzL2iKOO2mWaJmJJ70
DOnr8cvx9hgMd7mi+33K0GxydcCfTlGG/d6u6aiYePKDvu8PRlFJJTRMRP62Y/ut
gKPTXUkMGwhljlUCoux8bTgvkNQz2XgvL6wE6VYbUrXYpP/SUsIMWMn56O9UIUIG
fFxNNLAiMGmnDFiDFPAfJxThtWRkDpxAzysL15N0KxGzeq7jZW7KAs/2ank9P5rF
+fgGjsRaZM23T/NdoXLzDIp601d5pY/aSogH8aLRSgmYi/FsKN9X+E7z9+vHT3Ll
1WxqqcUXRS6/xTwJBv5U9gM4bS8jNY4cf7+5gItDtbWoArBxLu/RvrdbOyli9ViY
iPUXFMQQGQLKODaBohoc3q1eKqD6hudHAKCkenjhao/JXSUnYClSES5AcZA0Eizh
CI+E1KfIUvj7uzbZjV+4YqRtyqN7EkvCgPsy6QQelCHdeJLzqd43iBgmMskYkw/M
QQHUZdEA6nvYNA0WktICFOoOquGd2DwXnAkF+3I/pIyOgbEFnwHfiojblKM1M9Jn
krzY6XhLmOcRbf8co8tNLSa6aklmCP3c9nK05n4pPPYqj/KbL/DYg5LhBAkxpiRM
BkbDmyJIsQWQ9Op20bhLMUWYNGSsC2xkMS1AQtJXJfULltn5q7WP7CKBP3usc/A1
jEdyLAFIBvcT1qp4AIO+K6MNVVgCOfZ/kHQ97Z6zWf4Io4p2//29u9My6LXcfjwm
d2KtAZmQAjoaj9IqMgLbe1KCeiZrWryyNatPPF+/a5BZIwqhSRc7zDXBKeUeaTNB
N3xU8BZCkwyk+AGQfujwz3lwtq6qPe7q1A8RGtmo27HBJLY+d+QWUmTjxUbIzg5V
AgD3131raYTm4vsRI+apGmbkM+Y7xsVravjUzDdHvj9QuauuVS83QtcAurfWwiOW
gXKQ+H9k3u3LMpDCCYgAAqhIBNJVY67H3EQv/LD/nKxeAG7DIlEkaYkkmsBKGxHI
NKlX910DIGDRwkTSxgSFSSCbbnPqft1FLNKlD2G23udMAPT4ysNVbEL8ph77ymim
d0aIC/N7n/WSOUJK94N+pOqGspat44PVwRsEpUtkjZkWp5H3gWDa3Yt1WLDP/99P
K0SgkRKzB4gu0En7JHoteNu2fBnjChUI01YGmrl2Ga2O95YG0AzWoxd05uVNLGNU
qOJc296iWtxwUxIVg6FZX3P1+gxMTTkyYxJ9q0FjpjUTFlB3R8nwSj4nuF/oCU96
hnuCHpGWrXwXhJSJvLgP1OCC8+OUETFfdc/lIbrF3im7M+uLW63dzVJbcTSPGwHr
SSsGSjmg7bce6IFtRwt8YGkn4gn9OGQEXT+BaPN6sWQ2+SmiZeAFYzBkn+asTUf8
Wo6d6DybnpsrIG2/hbN835saIm9uEuk6g/llyv3g/uGrhqsk+lib9UNCBp9tqUKR
fShv6ZLTRLPaj1iRRxVBZT5rYEmOsiOv5kNoMbof2Lvv+B5cNfncMJLsS7lNs+vE
oPrrGyCH1fmszzmQz3FW7pZyNcX2EiRjpssfN98pmZLAFUmnUDnKXfG8POfpwy+/
Dblv5NLdjsI5nWUnZ7aeODBfcVe7cCN/B2qe9GacSJQLD4zryIkVZbWxB3MWcSqw
j4xEykOBNxnH3m0q7yz6v8icQ55tFdSHVM/8h3La0Yc5633jevemvt29MR54eNCw
ZXeYeptsKftmO40Huz8AexdNqj98WlyK28dCwMp/S2hFfMs+Ixv2vE7JH596iglz
SkvBMVtLODTiHR2MNgMxqNmMdURT4F1Vb2DizTqx1yYyodH/C2LuaLfIzThjx+fq
xi6/Dtpm+Z0fbyfKbv3PlxUkktwRSLfLa7bUJiXIs/ZuFwLLs6Cs/+udwnbzBmrZ
PyCe/F2Bh8Jqqh3RWUHT0rhu45q2dk2lTijzoYEJg/U97l3hRn9UMCM+Pe+hTLOb
eSMfuSbdQgZN065LIXmyH7Z/1kVxvQWKT/A9wLsxDiuscaR/iqKRVWr1/x1e7N+E
qPHNdvwzD1L4VDyHVQe8PHvjUzLbpwRKMubFC3ZDG6AdrCM3aUPP7l69Lz9wj3xJ
lDgxokptcsBA4R/8vBtEeIyIawpMNynZs5PMpR9hWVHF36bqfLxWEPTebvKS4Tpx
a6q3WqoLlsPgwicexxwkptQmY422WwrdbQ3qrczMt28OHBgW18irR63oEXr/68/y
f9NXMskW22M2d6PGpdeW/5VErWdVo2TxDo++Ej+IwHhpm4C+xKXP4wOVCWJzhwDz
Q5CKyBY0Sd6qWWWWpfmCv05yLFazksXLQy/mYFHKUuayEbsvtB4eyEADYZhdM0Sy
Se7yONLuMxYWOLg6IrR6Ld+hVlwiHMHcOHF/MpBEsL1wgZymMTtMPEzYzg7880Qf
sB6M67rgEEwRDwUkHPTCW8MSD7to8O9webAAJEM+fVanB3HI7PsRJSThqMX+DPfT
5q18f9R9RbjO/VSmRGgbr6TvadAt1krAi6y/aRK6T/D8A8sY0J/Saus7wW1rCI7F
cOgU8l+POBxCi+9i/3UF/mCHBeEdNDHxriPev8JetvzY8Ot5SIDsvpDh57xTkNAX
p/IIfQqwd1dApwk0f+7we6C6P5neDyfeklOubApuAm2It6Nkfjhjzb5ZA8QEgE25
gRv4CqwOxXneH/Xopa8YxzdQicfIDxaj1WamvOlqtXh7LF8gEDs6G7uqH/bDS1zb
P4RYkTxqSgw4NcyDByFnVLFM60+0mZB75XbAzQIRqBzyDzjQex0Vo1i0XYUN2QEd
pbr3983NcxiI+R77hnitVVNshOuTaRR5OPzTQC1y4PZSyZkvCumB2YaBvJAiSvYX
wF2ewJQn7UJFVee4GFKn0W6B5QrtjiaCHlukPMUAbr5DrH+ukgQF15GnmAjwn1bD
szKKsIlQ+bytrGeptQ09YFYSFJdOPEuRx/nCF7JdTQXYw3DbnS6Xonuc73uXsCcR
KqMudzfZrT23qQxHdoJb7WsyvGnjxYC1kIAWeCr1dAefF+nQ/dGOhh+1XlPEOU5p
lgExRNZsJLeuVmmB9x2e3tKM3XZOZ9x/Ge9U+4Bcv0fqj4pUDdmQS1iXXouctKYE
tz0swW3F+3uqEZzLRi/oZEkaly3cOXzivcN4KKehGsyiLGbVAR1XxBrzDpI7XcXh
wHHo7Ybo2gv48OaVOO+YOaop1c4Kah1xv5EqKKIex9X2ZRgL+HUjHiXcxZPfVjHq
51y1QNnQuZORlp5YH3zDTdyHcPIAVuyMmR+m/C/LS22UIIYK5X8har4TeLT4aKGs
Ap/8vVbLkz2k0kRbqbkx5hYuc14MFbj9yKHvC1hSYWIAcBRfsXLKPEx3Wv5rlYzx
FHcy4r+nL8U1pR295euNN7jo8P8qvGrveZNgmlf4G+2sYoSQMAONi6S2haFndUmm
L/HZi9V7UN23/YXVnFvx9Q7s2z5/bNIye7DtvW98+RkMlMSfYxVKcGwx83QIOy33
bi4jrPeBF+w6Pdhm/oIdpq5Fcv23d94AxV21/3WwRdBagbMkStCSFYG37/Tiiqg9
V36QcS7zGAS5Sow1Px40tLkkXDjsABYwWfaiBzGLqTVWS3zVuP6e3hycLm8q1M4B
wPpDTuBQI1Cp6p1tvDaB/ZdvvGRq4qLY+F9J3N3FxYvat0AWz5WKbwkNWAKzknVP
qKvxdL7kiTB7fHh8Gtli4dS5anZn6JQBiXvslZk5az9nfwW62Tqnzg1UToGSUo/E
10Jut8nfUruS7NefESAMtp3C7I1f6jCg0VzG12cPbiV+xlPflWD02zshEjE9Gl+t
lU9Ws93kmtax4ZYPOo6P/V7ZKOHfPux7bjjH9KMTrHaKoonj5zN34bioVAFrNtLM
nDcemhn5yw4cS2lf7QjoUeExFUNpJ+9Bf6nfLMwO0D++TS7yCpjGFqd4q0srS4im
TgAcaP9TjJvEl32YW9DRjBScn9/5bxLQKrtYHBKfmqYa8ZE2mxrtByDJ3H5ZHY3Y
Y9HYOPTFP4g6RE5zHIkU+OfiX17NYzN1oiAP7P/zeCHd5mOGMwHu6uaEIxrj7EFF
eTF/bMR2HT/v8AOaKykGFdI07TZ/wPR0xVu0ba70XQoudYcN/K0cdNPwbW2In6Wd
hw9im2cMc0sNvRLAgiTwOboPHlS5NyrR/xJ0jAfnGWlRdobUR3Eju0PEUGplGJPP
u1dW+lmvOqofEgm+4Ua6pkwQA/IX1nK2ULhc8xWtMxtPU2L4Eo40HE7ktvGiJwf8
l4w4JbAEDmALE/zsoCUZGujhMBgPIwYQc47KVUH/C6TQ4VEDOzBBYUU2+MbViMXx
5je8YvhpWs4H7jsdKIklv0ASAi7/5PPOjhyPTtOjxnJ0jxTidonhVmodV7w1o2PW
Pxr51vNp5cBqna1bwtGIuncW7VtRcdIO6mfypyomwL1FVszZ48N3wDpoJioQy+rl
xJjHVSpk3arnsdU0af6Jghv3m6LRA3VdyFYYvWHrQRAqSwwNIY1fo1kCyVXD/ydX
7FUL1vRoLXxkX4OMFCNSTGNO46uwKA9m7LJRxawGfZRkanTASb6J9iEuswFGtIG0
N8t0Y7teYaVXE9BFAA9uPuum+vn4sGl5QE5HOHrWD7RjjkQcxcuhIcTce5uKLS0R
8VW+QnJM0QsoamtMWvaEPAURxo5nyVwqCga18XV/X87l5Ab6TtYd4HlQT+fQQ5b7
d3meOwsGVrxATQtjTGLL42ZjmAQxuW33n8ij4x3YPpMd35sm73YbW+2G8ZqOoRqZ
K7/9B26XjlL2Dw1PxLenh6NuAYOu69zCrEOzLXF80AtFVV49L0JgBTCaTncFFAQ4
dQ0DHgSsbNbz3Iwlm8jHK4p0f1qogbUkJEP/9+OEhLUF7R4b13znpw2kqjLRlmeN
A0PwiN65NVjwjDann369nsbKkhRAhwE07lHnF2IcpGJk3jS/PFNsD7encambInow
TWVgtbrhi1KghuQKoFJBBep+ORuF+nM37Gb1ftFH4u5AV0hWkdDZjpTD57peT+Nr
WCLyrW8dnhm4Gyd6ftUNWSYQ4Xsi21XdsYTDefPZxFJHcK8rQw5zHwzkj5erwvpQ
V236T74tsv7rry7tZjUrhSByGAAmeXAAm0UTlEjKXsreGOTnYTukZ3nimZX00+PP
3/7++Zq+uuCRd0IC1JTeN1J1yFan/nP1FpugT/e3VL56vuVj+DV52u4DNmg0+SL3
Om0u0Jngrhxshu67g+mAgOCmyjHPjJo1Rkk5YZ+Q7C+lv4JzBI3f7aHSMqlV6t/P
PHHzS/5/YRrIh/IrWESmOK01vbGzkq/kmj1o0Y5fSGk0x2ezM11hhWAwsv/A97og
l1GOoCzLipDjp4l7p3rY2QluyCUTKlx3KUtagbbosFB1KcQAllD7AHLoSTQkI5TO
L5CTGNrw/oX1W2f8mEhmqnnviY+DoXX8YeFBYhTie/cHuXT5NN40loDhfcXA/ocw
cMiGfZ/QrlXhkT0cWrrWotVszxygx6to6O2oovaDqb8XBGNxoxtpWXXa6E/IDIet
Zd6xmaEfPB+t0nO1J8fKuvtCGaOldJ1TdcgcpOGzNfWgNiY1jPI0IwXdjc38nNwf
iZxFjbiRiCiMeIrMNpcr5ZSNYFnunIBS4IoKSgkk/MdZ9hs9i3RvN8m5s15hb6VJ
ZI8MOl2No3KiUQ1gB9K1L3RmLEx/A8U7kEk/cZhM3FxL9pIHbDsQEhn81y3VNoaw
CKVmGbjLfsihvcwxQTcYT+3knpiwmJuz0h/TPzkil9EQyb7x8rr22wuevzJC7ZT+
15NGzGCLjG1mjxbtG+gzLovI48DW81Jfn7RpF3aCNLhDVK1n4n38CQpEz28sVYm4
f030YA84U0QionMa7rLNT/t6Iei8kxswF5dSd9CTAxISG7RS2eliE+q2QSu2VACL
FgSrsDYoExrgtHAR26ie9b4IhaBMvpLcgooFE3+tHMifs3lEeiiTLUuDv7y4BdX9
w0qiOcFqvQUmx2r/tHLEFkhbnY+jcJzXntPCf8tY+qzsj1cf8benGpgEZwlTLqXC
RCEqUA9EidNI3ZbMOBO10Sk1+si3OboQH9ynlk+G6B2lSPAzFAS0pZhV0UFlzfpj
Xf+cXuiIWBlfui8OIFvB1llRytSv3xTzrS4Rv79mI+JIXDC5i+3wp1LZF1IrwgnB
lKaMqlcIXsvS/zcXSad53/GCJnHjeeQZ8IMmYoGGsbWFmFUsxL6v2Bhw9/H4IsQR
jxDhVxhxJmDIlpv1ZKWt68J29sroNaNXijP5W/GycWTkQtS0OvKZevCOtfLKVLFY
wjqMhaCJIucGIXenAYpLjhEzCnXER2TgZ1Qt9Q6lK7NyNW4UCOcxBIDHFRzmCWbC
4b4BvXV94xu3j6wxV+T9s+Mc4Wiu+2yv/G44Ghe9TAbW0WSjJUFoF3vGtcGjTVp4
cU9utNXolTpf3864vVH3z7LaomCzOvMZGv8QC8inbP6vL/Zf40Zoeo4TCddQ9L5J
1k+f6vsGKY0qevIh+5wS+G4SZgaglNZmctr+DufjVIxtAJjGAW8FXoQpGr1hS2VC
pc9uH3/ANFAlr9Dttq0915ej/7FXVTgyXZB78UmypCZvD0zJmwxhPTPquAXoLjch
4Coj4OfTvb7LBRa9WhDLVOox3Jj84Imt4lxbLi0+gfWlG+t2nDJUpRrv10PvRbJN
SVhyYx0Ij8Jj62nuJwBUteZd6LvbOZQF2Er93AMyPLXTM/yKGMtRKnBMhjxjfa4Z
NBxq+t+mAmI58kWnsZ/hji+McTUrJpSPeL/yp3CEuRrMwC7nrdtlEN37IYDHXfi2
kwUQXtD2d051qafXPQ4M+J79OsxJda88VX9n5+Cm8hb2TSD7eX8Su3p2oQFsQUV5
6jekuS1KVgktsTEifsom0gvk7NXUkbgM5IH+3lyOQKO9mEm1zhG5SZplubRt4jES
JGncDggIj5lrHdj/M9biPART7UBdBg4c2IKJBI5dteSlawkklzupg/BLtpwH3B+k
kUFJXVPQnmBq3aWC/mbVzWbLmGGP9wZHomofMF1xrU0LODlRas7nRfmWmnvTiXkn
ngYtoJFGo3duVn8GCcRDoAKMmwheHNgNyndepfeDDwZWZp7BKOGJH2wefrXi6dKL
lgAVwacup5BStlx+ANaJ2ERAmjjiS2/42/hIRiBTzzkK/QF1YGYIEv0SA6FSeBDe
ZsVec3jOwPa4hSaKlGc8y90cmu0zCceqNE7pKI594ApEC3prH8KgDAg8NO3X0Ji5
vp8CJaq+cCf5UZNujfJkA30+U2RAr2Nall14bcyzvwLv8eToYM+lmHQWF3FtbC+4
0DZ6mh/+uUKBaWETMH67ANxTzJqmpTiOCtnd5xlujcmWpyV/OY/AqcpQq2qVKw6t
cbbLAHBt2yLLL/4HicJoTAqbV97lg0FRN5vYyaax1+eEYg7XzRIZ3uPyxQnNcArN
bDnI6BFHjebN2UEooWRl+vBirbty3McP3A5ecLB+sD7IBnuWA79scOlxMBKAe8YC
CIiuSLb66gZe7FbG9tH/m4jnI/sGZMZt138AWXUkpuMSmLAlp97jtTl0ZqY/VDGE
A0Gol0f5a0HWGu4pBcJ/oITOYK1F4ZzAArdRAERaknQKz+aRhW/UuImR3rBMgZHN
mciRka30l2vIFKbPhs+gY7GFu7g50KRw23xgP1Y1T6f3veVdkKPRkoYhkjWhrb14
vbRyFgAwLjvrOXihWd51cuCJeqSVGs+YpL7f0WvbmYZsgW7edaZcJ3H9rqHyKDhd
7LvrWER8tEc57t8C82OYXxd9TMl58yByHQRcq2URhRyyIcdWJKU1RHXaZ+WOuXkj
GzAONAij4gl13/Uogw7a/F6PWSCl/REo5wKtvSQsqtuy5SMgJf33o16HpMYuMktO
XxltabIoQwSzQsmgG7D29kXFNq9bTwVlPppr0AsbfHM4m5s91JCPqyFIQRkEBk8o
5THRuK0LVxM/9zjWzUM49Qrrc6LUBTmYtJ2W+krqHCVTJDTCU9mpQ5E4GXrpjLRK
nO13/ozVdCVUqXdTo50gP/5WWz6IxFnhrOaA+4HW19qmVc/WVz/PDmmUBqom+bdH
ucUW7Vl+V8SbGNNnggo5rXjQQZPYiDjKLssl6XtoRAv6bwEMHvrKPmk/mkH0pZpf
qCBcCgXbny+Zz0vKmHUt9NbLJKuSobDvGYGfGUx5BGfKH4+9HoO9X+Wc4pzIpYeo
53oMdLWBcO9KyeiU3RB8/Ap8mb1cP/35iCBUF2/RhiFM9QV23zIIN9wEO21wOhU/
87d6GIizXcfHmlhnSI60366FJ4xgTLX0GQOZtXrIH7DGM6yWTwNe2JUJp0Q5PsaG
DgfObwP3GnbG86AF/IMRDuEKWFbRyLYU7JOwTqDDhyyCyDRjl9+9RnMrm1nEMlos
OpaG/bsK0mRqVUSq9pIlkHBZoZmWDkxI0/iiXjDlok7/6zEjq2tsnnGY2OpU2tRe
QDzD8ibhQUOGT8Ig6PI1d2ujjHzE0kohiNZ3BdYp2TCQwpzoda5WQvSbiZp8pCSt
VbPoHdUSYCKWMlCt/h9nnpJ26jMUSBL4VtNe0Ez0DOE629tNj5+fGMtq1qPZki2y
4EKczMgzkCd+X4vyt7m+BvIpi7Uo8lVCHxsNGLyiJFY4Ti4kvWjx75UpKdNd4erJ
QaoppDccZtoeyINJwC5MT78rogmH/e3wpImmkl2SitawniUChq7Ybl2Xe1QIPInI
KaFyi21oEWPuxEuRY7MO2tbKpYMt6HjdhrCfleNSjtExFD6haLZfDas4nHrjDZa+
Rvik5woSbNW+h3lH+Xcue8VW46/9ZQHnTqq5aczkyD6dEC4d9TgYbQLlbgTmhK26
+2PJ/IR0f4t+stgJQ0E0O6aToLIxXl1tLMO5Kk6LJ1g+gawGLfkxagqo6OyZQuem
JrPiRP1yqAbblS/yCq9VqsI99muhHDeJJqBnCG2PwJt3UW5IXOSbOCaZVIgP85jh
dH4lCIN4M3+s0NTFHbSOzBPLAQlUw+CtRd5p/JjTp3x5ctIAS0OfsZwyRzdN1ZjH
JHNdrKY2Lm/ygrzLzSHG5Nh7P214v+CPPK+ii/wzhSvOL3/z1IK3rnXLwljdmtvn
rwPCN6l9pTN1ZzqwGZm1OIwe/yDF9sTIX3g/uTA8IUjzJPTeTN67on9DeArVYWXl
XT8WgreTPxl++RLZPnrNplZV8SrgERrT6oB4S0CAd280quf7b5EdyE20K5gIdHvF
9HE50Fl5UC6vMLozrS8587Fd5DPZtiUjiPF7iJclIgH2xikUUMeOiEni1RMlm421
ryq4GO8+BvkrE/2EGvFhox2j4LbiJKGiVYJx6RWrmHb65oIIFYvtGJ5m0BlFvcpX
4e7oe/WGv/DUoK8wrrLkIIzYH8abr16Irzdp5nPtuodDVzLNJOY6/6KHyaIAQhob
fFr3KcWFJBeHYNCnbURBOhdkuj1hsL++UZaXsG1Hh2FZpek4bjaQF/LFVCAIeSpz
fQmrOmdP3cXV7LmzL753L/T8B28c+lGcr3ACHdoyi1Yl7IL2B6rn7yXHhSIbjTuO
W+Nge1VJAqWax8dMx4zPRUBhYMfvH6AZ6CjQU7aQ5DroDSl1MgBKzuKE+V5P5bAk
S9qMS+O4/UZqXcdKDP9wQdA0BcQmU61RGHJKHBKJvyYlVpRC7Wmq+uwOm3m4FOwQ
roy14jCO8jk5vowNoarF6VRw5S5tOK3RMsJ+axmlMyLcomKc+3O9jd02NcW6FR3R
yJTM4ho8RM84UzCrVYX8/xmcf46f5/z5fGX5EOgQmDcbsH0QqU55FKdVAY9s3bGk
u52T/6fjRDe5aov7KcCcBOmDs0J0jWq75277xaFkk+O43el9gFiywTSZWlRBYX5F
VrJ1UyP+XUtbPPv1izGRiE8ww6kwA5LaBG4gpkVWU9UFhExo3G0bVOIQdt7OE5vv
ZsKDlHX0+9ijbzTqE003usFn3bmEUXf6YgVCH1irq4JxephZLm/cPCDtL/7smMJL
s4Kz3XYNMHpAaM2iZRjWcFl0ckBdrQ9x5ENdGSzgCj4Z/VjNNxA+3XlpbUPw6j2U
Kb3/I1UB+U/A0doqZTspuUrQwO/P3P9kpmmaqZYXPxB4Uj0t+cCwIlNKMLnvugjr
SXwUBYwXGzo2zZT1N6YEkzA2Rh7eER0Zkri7fo4KSzdrNi3ogpfsNE1tIptN5LT1
k1x8nm4W1LEM0z7/vMYP3eGtwl0/XGTfEq7AlHtnbR0tChv+/wygs6gBoL9Ixx5i
NraXwCmTWZbegy35tobaJCGzw04EisbtSa0IsMej1/PMHuiSAsfsDwvFF8ZVwZ3j
jOajA/lIK+NYrf4co0MVjLthLqKuv9mFOo/IeG3SqAy6KC7mDGxdfyRz9s497P7Q
Bd7cRhdEJDdVSzGVF2zP9TYHuuj3pjE7anrKbzYVkm5III0KKCvPgmz0HqsYj8tE
z+U4vfHIcJ59k91IiqMj10wZ+Be8XEyBcyRA4i8bzAUhbYQs0J3unGsuUwsdu5Wb
AXe0Lv1B2d1HlONWsr88lqZ5xnk0OgL3YgQe+ROUughX+7r0osRUluf7XRtwj10k
F5ObRF4fOu3lEO4ZjXX1CBK1KjqX5pFbpMzHwDPNa4zhJ4eevq0Psj+lESxLyJfx
PQJ7ukMRUpGtwk6L/9B8B3H2woUaLCwfjWg+YHmXegTr5zUG3H4DQ4+PZFZaIvZg
/gzE0iGRy2Di62X8wpO7m4xoxZ2/rs+ZzSTfopjyoDKeaRlyFccfvLKRDwJJCyR7
5GTvrmzO4Php5zdI206m/DwCPe8hkQ0MffrBGgB4RDJl88wkiPooo7Jw4XTDE1bt
LLJVgx190qMeRitqQPFafOBQz3eQdRkAy/E3bVLiemZHs016/qoLvyEku0/qHPtX
ufuc5taCs4nfKMMnX3crGWQExxsaGYn3bw70oyM8rCbWjzLrJza4k5woS1oJsgy6
7ZFw9X8GKbWq7Dq2TNQ8kbDWjnDxyEsTZLMeu5fegRPRuZGamgcSR/8K4zyy4XlJ
HGiy+WFR3JqPbA0YMfzMYjF5lEHCvMwf7SowNu5H/Ogx2qSH7AX70rb+Juy0q6qs
AzTBo+Rgcq8U0j5GW7SefhQHXV0x8pCpytzBw4NhvP/Luquk5kbYO7M8Myg6X7WA
v3v0VtXA2rSTZNrb9UirzO35zxDu0L7JAEw4lt6FlOFaYhgE54kDootug5kFTY0D
S4zt+/9q2w89vWHq5Es0ltHq8dkuByCSySfJhDn6kJs03pk5azsgRgLoAf4trZaJ
fBLRQqPSm3+kYfk6mvSrdDqsJA7ofZbLG2GEXuJyk3gCu3PBheKrJrun6Y4vJLzr
Pm/sDhZHR5ndaNEqpLVjKliplGuoCnV5eVczxRsafilSPaU7zVlr5KaTOPP096X4
ELWRlY8fOgcJNmVvMLF+ZWPlDiG/Akf6jPJwRviCP4sYlLCxqFd6xGnm8bHrhxqa
Rxcw05YbRZ0lW3vNkLnHdTH8ivoQioqrhZNruNVGsP1YCq/9sLuoQswvHYrNksif
/Xh8ubfUBh1/TeJX3QoT+Z7yBNpZcuefZEIxpeWavD6S9gizY6YXnvepBCbO3doq
EkqcnXPPwrv8SUNV/lx61K5fxTRZYZdgYJ/CDVeunY0dCk0e+BEtRL0LhgFyOHGX
n3hrMMSC0cFiQdjuq7P1jwv8GmW/cHxZy9AQzZME6Ak3d+6kbVwrG73pZLyjPQin
mZdDIBl0dtqoXg6Tqfgbgf0KEKBVF4wZOEp/9K3anZiSijoV8OvZDbJ5Qrf7QJ8y
+Z8JgcoRFPJZgBY7YUqlQ5K7r1TfJV6PGgqeF8y+8mCjtmA+oKrRceeE0DseT0sR
qaCC37HRLvkgeEOy43BsGgXOvg1m+gbBEeKUiZeg2Jc+SrUbXfKMDtsQMVh0hmmr
HPOeUpBFuUITsTWOGfELcJjHHKqz3GXJob1J2OB7h/Kzsw0CLytIGvmYPIY6ThL7
3yQgt7OZXG9EbqjuC9v5Bd8OmwJ02nGCM73N94GyTW3i64UXGHs1uVI0qH/LVuZM
SOUz5IrgwHdvGjeJFCB+IVKdmK6sFQTPIoI58QMuuqrIxZa+7AEiLoPEUav1TxVp
T92kZAACieSuvz/j2B2YGmobP9BS5Ib3B6dRSK0GhUg76KzznF955nIqDs/VJHqG
qiq2HPSrXyp80pX7C7lQkFKMxqLRHqkwOrzl9kufjeevNm7DJxt0nMSEGFjG7lvY
rtJ1wrs49+YLygF/FYDLnesMp0vkv6f2T4DiGJsHvl+WOcCNR+Q1ON3FA39/UyMi
NRMgulw2zJZal8L+Ll+HhHNglybVIK0+PYm2bQCRpcMdB4kGVmolqPUPv9Lg+5cz
tifzoikzOj1LuRSrSTcqaaOvl2aEZjYwBriXu+d9BI3F3DR1rSCzxbZqCOODjUFC
NZAXXUxjcuvXZllE7p3uU+X6kuktqxfYgOlzbraLQE2ewaqm01hl29qklOt6pgze
xktoudmTFlQdjJlzo9ednZq+K2GRZLlqAVosoS48TbbOB0F5zBY0jXzSoNPKrlVZ
Dyt7WgQIb6EkKQW01SbJZKZBLsC/dtkclcTg3HxXab0/63YnkPEETDQytUoSpfzP
ExIMBzyPQ6HxeeuDBPZmWzWepkIvOTYa5mG8nIDtH81WpKnR/MLKQFtlCMw4U2nX
qBROxbnJfr986XepqofUNvu6itNV5AVriFJpyV1nENLD/gwnFuL1OIkk8gsrt2hM
TCc1uggX8M8+YEYSH8yo28GfL12CPkE1Oa18yUr0Z9H8Sdc3KFao4hn7kBV0ucmg
yvm+B9W5AWoeaixbdHWdZhtF6doBL8pomF4QpcrvCmSk+9JMYK07dhXt/uV5+Y26
t6R9fOPM83zzYfmFktmpgdi0SahE4FFV4MM0GU30BvctPDVFjjUGrocceypNSIWt
UpGHbfpj6cPrcB9kBIpXkXhdE6Nb2K58cciNUe9CXmsegXnPPdQq2RgG2HjlOSy7
WjFTPEYro9Jn2lj0AtfTO3WzimAmiIYRyf2as7+RhIf3/GtdMGJLH5y4G7ThMHkc
/y7Nma/GPwqz7XhVvYpcpMlqEBohhYPbNgSV5qv849UbHK1ktNIv0+UOSmhxWae9
ri3761z4PMEdM0+bNI+5ww2VAZ6EoysfWWOyUzVeZ/fPYBGK6O/QmyTe8HnAHPmx
QzLv6F4kha5mNvouU6palnoELGwHk4/GNObyO4mVuFGNo8C6DXa0FC1SRtgjj66a
mzbTGsC7CCOh/6rAY8D+vfF4kCCYjgLGjqTbToPiLP4krXttIJCPv+yEToM+8YKF
BBftqjxlEtbQ81Ea+wspw5Vgk6l4CcmedzSGLJ1sjcTxsKAlD9BggoiQSV7uXxjD
oBA0bStCBDvkv8HC26SvdeVyHnc8BEz+107+AqcN7IvutcRnumzul/xODIbrE4ng
IMSfbdU+XeY939ALopYuJ2hz/qynwgvBERDFDdzsQZju4TsyURMAyVWq+TtWS8Cn
KbX0+PXS5LB95QJEyynDZQ1mDxLk9fUyYLFnVc1gWOnJKjVHqngohKUSu+qthkhL
Vi0IqEMGPPUaKNDUNi6SnJl5I564Gyf6Sksqt5p9KOZO7fGczYu8Cp11T9wpBqnJ
1b+vtY/oSA8vVJc/eN6v5AiPq9uwYcgA3+o44zIAQiplgnfYVZ7S95lzA3YJBApA
I5PF23+Kgnc/YvCFFKk3W21HdPNG2wrQCqNLuNMw0NhlcepQy6ddXc4ysPlh7EhY
QMLaWv/tggTO/x2VlYV4XH13xN06PMxZ63DlkY+edHDMBoTw4DYofKVTwrIFzTpM
4NpfHoMUwH0BeSHX5ZCCV5BaxqJZjGQgfLlCP6+j1FFjWCXo0suZ7a0Ji1CXkafL
Mg6syy8uUe6fsHhJfPyaaQce7gqSHabLnxNwUc4ZhmGjnxEK3t0/p63WTykYUBTS
+Qqc8WphoFv3GQ1Co6z8yLGGRm4zRBEiNNzgaYirNnP46MO81WXqBDnENucQ1aK/
2LBHljyvJptZpXHKoc5HzmCkXBKSTJj/DoeWxan/NLu9NITOnWY8B3q9gwsV6aDk
nPUWb1E5JBSEmDm/SyGXUucse81Wi6mpyRiQJpI7QsdSDKw/L4nNPIBQkJPYK8nx
vlAGXn22cKpVDQwK0ydiAv7MCSgQ4r5sCohzw4MY23Tn81uJRuygesGkoofNjHxX
X6HjpXyVNhS7ioaeJDD8LeVTg3TpP49iCRkXg6dVSKcXRoZ4yq///qrlQxG9R01i
ChqCujzOWh+mLC42g38aWV2RiEI9am6TmIYUbW6BMPFtvufy5NRwPglHvCrHkp1+
ubJ9fuzkHqUBznFvjR/idRJ0Pnx+UreBT8BKUH9RLSgvmyAMRrvtbNec6brkdRnN
SHtJEcKf2XKP/lAoH4sdHpmR/IrORdsSckmRYsFVWWs82Fe54jtyMkwuC+rniNYf
2FxoUXttJe+EG2pxlu4bufPRW9u5sFLDq1p0koOYN/cC5hw/xu2jiiixYiVoWck8
gz5HjTIk7LNng3DS+aHYbC5PvBIjeg7rjN/WOGTm8hcRz2G+3BuHsLndQcZyeTFl
rP/d4RGKeWZ4tYK/MVD7Luw980uiivTB2BeLQJCwz2xbIn0Itln4axWcn4jALLg1
VmJYwcn8tPmp7V8jtlXtFSoCkjFruiH7/3j2LkkLVNAb1jqJVMpdS4zg7tnLrASk
NBgjGPi9cL82I70XlKNBhO6Cz5WFsqP45PlPikFDCGQpJ6R4MSMl7VFwgnnit49Y
higplt9ubG8eXRSbLylpqmlTl1Fj0EUfK4VsOuXP2fcZELICdbz/d2/1TReAyN48
2pMK7nn+uN55gY9objtpjIEtEqCJn4RREQJ6xH9F2hgxW5oCDmxHR6ajFO3udit8
8EPwceB9bITVXahrSHX1H8gwDRgziW3RvhjMyvvfSys8A3Mup5mYe9n4eFRSmiO+
F25G95X/P9A5Qo72ObeNzP3JiZj8mYreS75iWqaIk0+nS1qpmdZEz9cbmpkgmccD
2wCteLJvyE32gjVLnWdSf3gooAwqkmLHbmdwKYoYqA8scvQbcEl86+HBek00hCDL
MkSmfYTUJ0Nv4XMHF8Qt7i5X9ucg8nhW8GPSlffudwCVvf97vq/VaBfvAglhuyPf
35k+TgFWXJMWRhQA64p1BI4HWuo47pwAfxavmvMZBCRXOXSk0mbY8WDhGM7rGplO
+obmSsSe0t+ox5db54YC/U0c0RqOqqhs/pecgwT9lnpAOmliUVbCv3WogjwZyBC6
WMs/uMsliPS5MupxTpz5T/CidqEQKHZq/TGcYk1RlpnYjC1Q+2yQdMvZJknT8/mK
LpWnY6RHSatAzyZfnu7q88eCYvOWnUhYPPkQA1a52t/ajM3rjRWCYaWDtwegQj5x
WNCzzOwhs6qI5ujRPjUzSX+M5991IppsgIyUyfX+OEiTIFsn/wSbU+vvu9Vo9anJ
stPtZcx93g3szeV5hs1KIdriaNBECUVo/UXluVjpQuNvxwm15YKZg99R0vSqfQqq
FFF6cr520CzUx6F6n9+M/KEjRLJHuCnkMbQFICXK2orZ9t/Sw/J7dv78hiFEGz/a
fLcC7x+XFQCor5nnGyANj/8OkP03AGpPvcvuqqOP5wpZ35y5Fs2wFS3HzZjPaOY/
Kh45jmFKOcasDjPJ4ZD53jCzLYurPxVcdzc5wyNzTtiPE7crifn7BqUyKR7LTaid
JA8imtqhIo5LxOJLTCZbC+3J5qzXZvDmiPqdWdytAjWa5Q4RMjwiwLeuG/EztJJt
0R7itN8qwBPsP+woAw0uZfgmmXkcewHq71XKYmRxB4xoVDwJbHlz1o7Urt2CD5OF
IXYv9b+O62pWv2v/lj8rneqiLQlhL8gmkm8WoaT6VLxHSB9updQfZaVl0zWIelDt
fPZPBJA2Kd7Lcm9ax9RnDUG+dT5GWisI88Bm3IRw5XI8mM8cNhozjGSefRLAwj6u
q/61oG/5Pw3hbU/XGWtyG6NqeSED5O633DNuEfF2oCmbgIKsIahbCv3tF2/miXvc
TgLO1EH8Fpst5uCM2aQzdpk/dRxWfxrHY8fED1I5q2sFEiAGP+u/QKydaFIpDex/
xfAbO2xubZ9gUeDvslo7oSHaJpwzuVpCbLH3Brc9Vmom601J2Wt4VtkBKvQCPdIH
5weNUu2odNS2umKvVBYSllKRZjzR0i6V+z0+wT7ViB3ZVmT51Oka72Otap/ALBrb
bEozHp9VttTvUXxIOA9COHHIfDyNVEBZCLX76ifewpP4M+A75To0kFW9/dzxnRQc
AW3xv2+Fbze3OQJfa6m86JZRu5v8SYuOFTS6jMRl1BgfD6Qlg9WizUH79Evf9s4k
yvl4+M2ClpoRDJNAmvZm6ZNKiacpoage/J8jzQOGHgYzPmQbHUnbfkSAuw5HHvVX
MXpXvAn29MqjCX29YzcvjK8kgIaeiFXZxP20pR0Fyqqq6FUoCzdMqhwF9N2mn1HM
+Cxmusm90uBar9sGV4aSfP6PKKmO83s5sYUD4JPoMIghhTEoTlBA17Lm/ADs5GSQ
oK+O59mfEoW7MWce0pLFQLpPUDp3MNJakrdvzIk/Oag+JCrWJBgJZVflbvfHCDXk
e9oRVCe6/pPgoX2+4GXNiJRU+5OTgpXUC6YyIuHExQjSvxY000ueO5TYpRosKqD9
WhCZdzGywCY4zN4rFzEec10xL7rO6t5tezrNh7mCH60ZhWnBht4D3ZTwmliC8ZXi
GYavXZVNxR2ypBpyCePPzyGEsJRm0xaMItU8S9Na7yc45Qwp/kJN/kLHzUt2tR+k
D44UvFSwDTzM1Fq4Y3aD5xrtG1jnk+XRS/VowvhOC1NzkBLpxZdhAdTK1lRdkByi
HGGnfXkc+tyXribDxOUMy4XbdjrOLiZmcq0bBKBmCm2IUJykj254YYbWo3GM78kg
YzKAUdmp3kePxv2+0+ccPGaRSrD24cZyzhBTCsk7BhOe+9Te9tusO2oSuLILmI7C
UcFhH4VKZ+/qhDTvjQn1zto32ngmZppEB9j96Fq2/kE7Ggluy8OISRcpD3FQe9Bs
nk83RCYk3Rz73ZukyLQKyCkjFzFd0yX5nCr/t8uCaLCTPVM8gVeC3FH42IhPNX1r
dDcSVuKqI71M9U8uN+nU/eAsKFj/aX88dXBcP63GJCXdk+vt7JC8Hd0TAxhV61i1
VcwzyjtGn9yhQTxgIZ6oz+mjUNWVmaZsGk4q9xf2L7Qd4MtpfRljFWl4T+aXhER4
TtcP7zJ1WfvMb5YGI0//VE3upci9b1LSvirwTPieJym1pb/3AH3Uvj/JKQe9k7Mk
duY7x9OxtN0Xb21oHiMe5B8dc1hbqT84XJem/jOuMQP6CSv9Dc7xaubtfBTIdn4T
vu/9qWRdz6/C3yp/0iqMywzDW0amyQouLZJ0kb5A4xEHhujvErwqo0mVDW5YWCEF
jNW9grDdyTfpMEX+U0+qhGGK6Belsz99LtD5/w2nMPPyM9V9vqa2GqBFIOMc7NG5
OkVlQR63MoEfc1X44WU6ej1jfrjv6nVzCwDrD/mptoFujN9mDT1nVETOE6sztiIm
HID+Cf0SXqU9e30U005V5UE1DmsdeKFnYzzKq8bOFc7lfpiXtrJ1RowaZnpjoqAz
rWa53N991P6E8SqzpG1IKn0mUHFcVJstPJsWh9b86mTrjbwux/6wi1TltR+59aB4
+HSkhhOkbE75gL1M+JqlRsoqvAJa9VV9G+d8D4QRs2j2BVdWqfMEjOCdH4aRIHnZ
ORMZ4eErsiQ7wtRvD4Qlaz5FM9RBM6aAEBfmspvk7Sw0tKzGHHqpaocLpxWRoXDf
eqCniGvOOwroSgc7nas0ianscXl7w9N4INelUvPY1X6gFdFoexDQVQChgfehRf3d
hWPGfhEVB1ulCjFiG/WvBoGY+Cga3KHUBXLM6dznZOdP7LSmSif9td1lVPMsblEP
tptVn+a/mSXjcP7CMg9KyG8jUkWtlQfgXtSe717FZXfh0LMOJLh3j9/VobySPeZ5
PzUr9LtSuhDIBBHVv5kie7JZrdWO88xAMNcHvDUMVjb78BOTuhOS6Xph1TW8fbh2
9cTYd+3OP7pPJsdsEnNR/pYd6TX0jp2ngU+8tQeJhyo+kVvbUlFulYUl9Ka/l6Y9
LprtlTSmi8mcgxJU/NZrsa0mqbRBpKIkFIr/kzHNtftkHWCurGW92lf/VPjhTl2Q
GOx0B6gX4Ws0l27xO3L4mzQCGOPCGOCm/cwo3GG4hF/XTD1OL2jWexreFCbNG94q
/ILFOMKFAfP1Wcq+nWUhcQEerUv1iqGSruMiCko0eI1+7DFhITnZvUq9RH+n4Y3V
AYrViBV+NPmL+FnUCw76kck/wFLFG1CuWLMurSNMEaYoqWkSVxskfGYOemI6TOCR
RHTf1mUoD8TiEaiLhTaZBn4uGKHP0QGQJzKby7XJhOeUkv3UDd3m+KNV/sH+ig0i
8x8/2b9pZLRKdraFL9Hv0PzuadC+YLoFHjXO+ZVKlwYsEZAsVBCZXD0AfG7LEgPO
MoVO6snV3NEA0v5+WOJ6GwaFmD1Mm64v0Qazfe5ueOaeRb3kMJ32r1ojY0fBrkUK
Uku41+bFL4y84cuplWo2uu7nDCkB0AWmSH2NakWVrockJ4r88KiL8ZaJHRgBUCRp
OMqak1frj9zl7cfUyCY17g3PwW7sdXjV3p2dygBWvCBqJz4IpJ7JEHJIgjPMAx70
0uYstxX+F1cYTw27Dk66t2iq/uJeGBaTS4lT3AAPFYrTmK4S3ntg/06GZnGbf/FB
6jUJEn2jy1pkBcVWTB9khvRMdmp10uA73SZ+N028C90KYMLzI18meiPZmHZxKhGO
BtUtHiXN9aAQ567eJxy6Zps6xnehp41A8FE5Im9HSxPJ/qpIlwa87lAbpb+BKx1b
aMuWAtyLY2N1v2fhHgo7j4P86UyVlm85uWO8S84mxxbFX1zux1S1zgk2AY1kyykq
/KbQx3qJECFzFfP8BKVuARwkY/2I1JolXMzH97P/J8e89PJog+xg7qyUEHzcEzAX
kAvxBC5p+/HCWu09yidco1emZLaGIyKp3PSssKEdP2+Fl7Vr/0/yO7q/UPtil6uK
Z5Y6icFYUGxfUma5IxYNUyCR1Jnvomqwfg4AfXXMzVXT/YQ1IF+YLwu/BLnELz2v
bvSpdujkk1jB2vtbcodDBVleiuP1Q0KHxmESrLeXWpRCpUstwnrDQQXDnnzL8pbX
LdQQfEjCjas5eLbkbAF6TKVgJZeBiWMV4Ek0BcFFJnypdLEsImY3dVFPZ/ztHTbS
8UsC/vdoN25ct52IreThA2eMbNihO5aHt+BtiXidpZ8tn2ZtKy9RF5AxgEaXJI9E
HcQmxUbgsCDAUqPm/G8Coq3y4DdUezo6fblZeR1tvTLaep4Bit9tGXA+x/RkSRdg
VOLM2PwL+3zh1X52Ty/hfUBZ4htxHH+RzZE7Ye/3b5DrFdB+jSGJ532MenKFf0hc
ai0o5z9LF0hBebXNepDhKcb4jJq6tXNasO4mdDZx1eAySbBvlBBOgTxyd1OLSIyN
dP77y2H46yv4HpWAoKLtla5PVyahm45aufswBqq4ZNcDrILGuha5nHU+jvSaTTEE
LCbnDhxe8aUuo0lbUd5w585AeeWVHbfwOC5bqGssDdp95Nm8mab6HnjMMVrIMd/7
quMuNHkDYS0DDtdwNW2z5f4nqKDM/imu/bZmdfmRUQ93dwbi5mlpqTcRLGgFhL4L
AihflHu2TNil5uZOJlroLI0GZX5eeNOCrJ1rxYWi/0sFThwf080OSHD/90HYxpOS
4uK8c1LqHm9Rrgillm9HXrtomYrJupNYNAb/jJ+yijkCgV7abkNFw/2COSHibmIf
wfI6oJUvcwwMDpdMPTFARoFO1UYoj9EMnZbZ5YJbkwv/iZgSuQUpwSxtL+YNXXtl
kFAS/UqXMFjX/GTYabzs7o6E8kHE+AatGkjurSjQS6h27eK4OZutUeGpeZFQenKE
q0bDdswIX7ZigbWBrOCJ8llCvRAh1PaV4MUoGKF5kZrQmvERYudKF0+LDxIGqxtl
ou8G0jqY/xMLrj+IBFbPx9qKr031LUQ7T7ZATW3N2A93OLG9u0IdOKT7fZuK7Dly
RFFcuAnD6srwrrSxZZviYt0epf3h42jTT/9ApwsxOYgL2nmDLi+K9tUFsTRnFRds
Arx+goL+rMcg738c5TxuIogvscl2bFYXpix1N3AKS7QJM+rkMAxUvlOUo2I9GXqM
JOQoS2kfMe/FyMV/gcySgkn3oWyP7ZIkuX8HJCbTqDIhnIBq7HwkBXXLeoXXrtZ7
WnItzLy68ixFOshYL8dLnJ+nM9DVowfu2E1d6w2pv5jDJmSStf2uPmxvIee8VgZ3
vd+j/8muZkr2xy+TiNtEpqBTVDitrUHbteweN7LnhWQkGlvBFIfqLE1vwwcVPyhs
b39mPCBNnRSRyA5a2RsKypBN3yGXsey9aTkRwZsAlOsiSno6AmZ5Ivs330DYtsg/
XimUJDz/U6/fRv3bYZC0hGUnUX6vchugLibosG8xXvrOAzrG1F6hOhgICdYkaiRW
aL8UHO9DKz+4K99WGCYadEyyo6aiz+eAfidUPd+pC6TSh2XSAVuH8bJ0ACwSlj+e
6ZcWXyjWTyyA43mASI5zkEN70HLxtgPsYc2tynCwogPh3hqAfnuuCZtYxWvA2nKx
AMFFEEXTM7OIhhSFqBr1NqmBN+kJTmrcAXStu3iCYFVeEboM7OLI8MrZBqV1aHGt
aq2BXCRPh3yq8SGn6fTgMwd77SdXWFLl/YGwzGMtoyYvcNqyAq7wNrxMAMEAbRyJ
a3rcD+lYRcv7SqhpJJ2GHjr8ce6qoDz7pSjw+nipphlWym3ZRJQxakQcwDCtfzHj
kxhpaldtOIBQBPlj9MSuK3zK83liW5Gmp9+9ekNq7CzlOx9Ebi/Ceh6r5O3/Slgr
WnzeTKYUE73zOqd7u+fPY1Z9jYYLPDs0tKMz2prvfDtYSzJ5SBCYa/AfW/nKKKzW
3dXxT4KPEBaR/eSLCJV0aOBmOB6Lr6VOAFIcaqKeBpLQ03aaGBXpfXVowRBovj4t
HG/RtkVnWUEibEpcJKXcCDgE+x8Ez/BwoPDtlEmWMopZz8kkHR5x+Pq9I8uovFiE
kPjtcnlwIK5/tvdXqCnqrd2gqZGgVxOBlwR39xiMtJf/Pp7LpRNrwgSqsYXN/5XL
N+DCXixtHEcr2WgHZZWgueT2myz1yS7Olr6LYQbww/a6OLPFewA3tG0IJL3nsFXF
ktbgby3xbuYMeKwu6kF+wWBQ40/FgYboRsifafkMsGzONsulatFEc4Wm0LXZuSR4
oAs4CSlxrwmPozx4dh1FMyDHJwjb6dsdQfdVDV5/CO0KcTpihpl3UxAWmUb3vkFV
hmVJzudryZ7Zw91PvI0NdqUviz5BU9n1Ukok7YK8u68EEv/63lV2KSLh7JtM5Cva
p+e3XfKkwZqIuB+5B9TJML830dIIOAAVIThF2HOn6eub6zhJk3CANebGWwlXGxkF
iA8t+eGmLytmomT47DcQRWccjJLJSfPg1E6NztnfDzonjpq+7jZHb7URHI+6DJen
WowZGwniqN+GcC7V5177B5Oy866Dgr6FXSvLZhkzs28utVyDwa4NKx5zjqwjkM7o
rhA4VvV+GOkSsfKP3XN3UTtBKwYd6eokEyFpyVjWCN0l6WO31GCY9/BP5rILeejX
FdpDxyfj7O2Ph3qDfObqJmS8uZ3/cn0zLgZpIzj1Pg7UEsUtZXGxPNXxyIn0uwlg
aRlS7RrrGkKs7uG9oP5n+62NyyLYtExVntJkb+FXas86aYV6sg958xrfs54Mz0nY
vYowExvkNpEeifEpHgUtsd1xxKZ3ZcKeu1Thx4b676gLFBu4pbGLQo/63Td1msP6
VqXPc2w6KgUfvuC3fo9PbUCe9ohm+BRclTcowl6KBQC6eYYSt97E8PyBDnrUKJzG
8cuM+oj1m1ng/aFBih9C8xqdxFcMhrObvpt6qRWpV3e325wa2Ipo8igdaXydlAau
2heZ3RjQ6TskfB55bmMYhY1N73AT0hHkiDZeXf4/S8lLnwSumOrouOc1P+oBKD0q
4uwTLB/4ANWmSG9JfANa3EBuIFMTy8qSy2rC4ZJjBhLwlu9Bia+mezImEkHbI0dV
k1mskvnzNtqotikf+5lOk8wj7YI/bRyzT50H57NSz8p1WiwK1ZI7aKsnuMQMjSDC
0Nc/qdTLV4PVON/+JziNH2Zau47KjgueOJN7WMMiTcIyqfux6Jm9NTFLt2RljqB8
PXBSfhbFL/Fe5kqjR9lN0/nwMWbUoIpiH0zdHx0/6y7sxtiQ10se4fslFD/IdwCA
BeBwxuEBoJeMTGaYaJ/Bpwf6dpVUeJlLfj369bxcZf2mOmea5Jpa1DPBKrLbqhzY
MvfBE6hAlMjpKOJCu2Ro+KDgr/CabRkpfuWtFXWN45VIYZ2mOiiROhSIZRY2v9gw
n/Yf2c/bU4lgzhBnZ4x3xE4hmXD7dV7odJ9DwPRF3mICMXA/HSMTuYG14+HM+ZJ9
15BDmfYATTHiYy/IFlBPuSkRGvEaB2VzaPPlOSsr4li6wvN7G7j2eu0vScV2F8ck
CvaNHmUnawf9jgmmSqGiWyDrOYbUudZO3g2OT74pqJwGjWsx+/f2dlF6WYeMKMPt
dAOMQkM8DoltWqdBl5N0BIRBP8F8Ns7de9W5MPG5mZu7PKlyka05U77LiLGWYmgZ
FB9YFQNCRUfDIU4/3vH6vbdvKYv2srmyEv5H4qp2f0/ieMok0imoqJBaKKMqC1WO
iTb9O9Ro4XgOd0s269aLGMBYvTZ2C5m3NQoN8Q1ofR3FhX1p/aobn+iviMPgZo6U
LtJp+aoWEqutnwWz0zi3YuhE6A4n6fH7Cik1fRJeVfmOpyHMSQ4kP++l8uzxJ2J8
h5/rxzHLYKuQSab1Ecx2AxmeVdzD0/c7A3C/Pt0qYMnygDtdb7SL9B1kR4Qpp1Yx
OSiFu8U/b3uK3BHoNO8UM7ooOZzLG9fF6gCYOuOhZAiq+1UwuTSlnEqvjHZBs070
iqG5wKe172EQ3RWae/p5zAwahu6UyuYOPlSisSiTGpO5TjgyGsQmhdlHBjN2TQwu
Cnw9Gbg3Uq3KdqJsaFhUdwNuEY0DfsfX9x1p0mjR6UI6/gFIPgcr5ZK2NYdH2wcx
WKqruj1zqiojsk05dOi4Dp3q7LCSD/08Ns9ZglZ0pMWE50LkRjp/PApCSTUKHl/s
R67cTtcN+EKl0ZZ3OkeHbs8suoBXWjZnUmsMQNQgnv1cpSaymOxVlMsua7PT0i9V
s9f9QU8sSTrlInjs2X4JBd4rmRyE8qp8OKiJjuB5f5ktfnmDnklfy6x4ovWUfFqt
IluGkwKv9iUFvUD+3/oNXWiJyimsu88JLe/m/HhoyScmxgMgzb2brc9DaEA8vUsy
XIg74XiQIBKV3eZf0lysn0oTszkCDuex2pYVs9Co9XZsuqYIesqEF2KlzlKUHh+H
AO2bnq6mY6Y6miL9R3r9eHZfFrGs6Ke+YlDjL3YgRXt6SPO2lLWSRsmFA5WeqsXy
Ewmr3U4GToYOBYsrP8wrPpiGqPwNRqNfrT0W/j20DsdW4icLWpjGl1B1svVMHDfN
wERSX6F3vyrqpBB2+6GEzQ5VHWIzgVMupFqtU0odLCCywslP+KtqrPEdue0HhWuK
71aO1QbdGElWrxDn5A7o6/rLq55w6f4RcQIxqFoDas1rX1Bg3d7CKZu+9WCEu2+J
rkF0XWqc/9Dr591kEFTIinJjAZ2LBPGMjAqfRHcPwKxCFvkpbBxGLF7ujas4DKJC
y+cAik/4Lyyuk9J1SIV+Dny61AldCWzTKNOkpy/XzXKhkzCqUYowXPS+pDoPtjHi
DVpAlPvLiTq62SmlY0/U6t+fvS2hhCXD6S2vCxB0YBOMN5KjuVW9q9LD/4G5Bnc/
UkSClMCl7epxOAaIdVjJNe2HtBhFcnX3pDfIlTLlmUlMS4IuE2+1bPjf8O1qd8Bh
2XNiGFqJ9iWb+CRxAxDW65q0fpFPF7LpMDGoDC+GqsUFcDUFFXZd5wWXmOoH0Mn3
IwSr+TlDlGHST2lqs6n0RY4+/BcqdrQuYvnrr9dFzaCHFtN/WXwPC7nUU08DkgFw
3yAxSuuBruPPuRyOTshDow1fvA+RKDk7ZZvKa7xW3RwkBQcT8zKs5NVStRx5ZDpU
wQu2xIll/8i4P/OuV1kKwnaNwOjfmqDaiPW2Wj6N58QZ0B+s0rhyi84P2zlDCyMV
seTogLlcmZdajf5VXSLhdepGz75ORexnsek38RLfU4tmMzoZ2raODAUXcAJOQXhE
YHKAKJkL9sL39RGF6hMh3BsOJoM+UKItvRSb1NfecDhoWQGBxOLb+IJEjmyFS7n2
GQMY+rybmLSz4kmE/HBun305fesBzKjh1eTYj1ajkJmW1brQ+X/9IdURbRdUDnup
cHwxlgvveMu/XWbvIli60bLCWOEnCWnSOHHQzspTk1SWoWG5PN4FtOjXyqo3wiIC
lY7je0/++uD9oAoxslVI5X0SNzNNyYj9bHAa8SKm9e+/C7HugRClV5KaJUZK7oDY
7y5slbRSsYZnoZh7C4Ysmx1Wwot0iMZLbbiDt8i8yNoCkfe3xNt0N/DpvSNRPLNJ
vPs9NSE3sN0/nlX4KJdcJn85238QJxC6XfbJnABFiFt5m2HC0az8jrmZ54OF+OVK
sF4fBx2sv5Pedx3dITATKw0SEcnMc0/j9yugTQXb3WDg+9l4+7QFyPxcvHOnuJh5
B8XUtG0ekmEyfqCvPexcoJgJdbQUJDK8IMreWsa4q3TAC1d4ofzrdI2TsUB8QagB
04D1pUxUYN13llOlvFgA4p5jL3HED1hxRlKdU175oSMDUJ7tJ/5cai4VvWcZrac4
E4mmDNmPvAWUnnTGkUt18zF1T1KZ7JKJ77dPqKB8UlOpv9zIlti5HjUrrL0Owftz
mJ/LYGoBnOMxECgDrjkPo+is8eYjR4vH8B7MkLpTJVo8uN6N5Qkf2k9Ytn94Vqum
fLUYFp9aFNJoP+sQu3tG3eLjQtjkWr263sIkFVGW8l7SjoVt6ljom0DcGXHQJlHa
AM5IAa/OHqJGazcRwzJtWjXyaXAD1YQmEaKbZ4+72Yc1RowFAttBidEelKD6/jNx
eU6/cecfpD+JiMxTCY1LUD2ZsAFb2JrMWm8HJebX2sBOJachU/lBpHXz3l+tJ672
WpBB6dieht1adTy38KPgz3YncJd5B+qshSUStLmF8ywcXkaBm+PitUDPOLTjoQRH
Wj/t/wmtbugQg/xAr1xWUtwAS2+ch8lJexzUVLWnQ7/WhcjwlbeJMI9CWlNEhTBR
TmBA7x8QA9NGtZycrTgCtemuz2ZotG2tvsMPekIB8NSHZVXQUjvYgXdATDD6JzL7
jZM3H/1XrTWJTmftgdn6sdbUcOlJEVsiLwG4uwJvzhVaLay7TmqDcQDPlKubcs38
wKp8r1TLLcSw1wkNsqRL17cyxh28qC+BeuQV210sb+kKpfDPJvOcm19F5sl+isTH
L6nlnUN8FqBg0uZt3ufHhDg7ranPbkBLjoU3h2ov3P8xCh0DTJxxbzYelbPyRZhL
EpHfABsw2s1RVMeGJs/dKgUsmSsIxUzDrQ0qYrVKw9aj23SPAu5ohTpRJSlaoY/m
j8welM9Shnku/2vl81jiR6jpBXD4+XC4EZIDDZDkfDyzpm5DAaREnUMg1DRFTt9w
MaizB8T/uqHXWwgj0HFkgs+GUpKhw5UtsCgqCFPDJaiVkyFUFBw4/m5zsu0yYAVs
A7plmLVYhlch8NiOCnRpOxwS1NIlzQG/r13Li9CGqzIuLy6y+aSm4J+780hEkCqE
9HLo8vVHs2FZ0qQODJWU+8/YhEqEihiOBz0HCC7aJ6YyIkI+F3wxlJWqkRzdIttI
Ey637G0yjJzM0v97cjqAFIS05s+UV3nBIfa97pGnC0Pc0JNJG9d5gt4vzZJwrwAT
W2WKkqkvZpJxw86WXlQXM+22PU5eNsOWybP3ydb3whRpi7KinWyxaa0/L92zvuzq
DPBIJzp26iHJr/bSfB2kWpgFZiu+jVgRvQ4+YUhiRKUw/428yNEMFDWR/043H4lK
VTh9F78XzanUiuXOXJJu7dVtC8YLyv0DqZF3komyzluI8O11QYtPZCy+6r0J3G3c
cYawyu30i9yWAZD8TZ67a8reYmPXIFMbmlV0KRe7zaHKk3U2FzanQUu5QCjP0VcN
+XdW5zYD3mXqqdqVvtI0jnJtkzAuLRVrlxiYPdu5ks1VCp9Yej1U0V1K2lBXmxRw
hSVsvFg7byt/mGOMj6O1tr7FPXxWysjQ5KJtaD/ONllbiUU8sY/KEiH8K/LYPuEi
QqAg7WHhoQ503DDAw/QlyrFai/WbCcMJTNmIC2n+5+OJb72hQ1PPc7Sc+pQiUzVg
HQrOFGdjJdovPOjt6mVp4OCT7zQgkKjVkURRDwD0Yh9C4BFmu7p8BYS8n+I5x1A3
aHwSwei4kKodJdYZT8ubYmq1h//+JdqxI01I0iJEWLcl+Lb1qxRhb/FZ8pzlTghy
gYomvWDT+nblmSZq+L+lkJT/IUbeE9y/y/yzOuG642hMGUfHvG5WJerdp38vev8Z
5vdwHnXSWV5fpV3t9AjgEthR49uqoUzrMHlU7/oh84jT9wIm9JlotqqiGL2q6Ipd
4KDLj8lpwZl7mTJnkeO8a5mxkNlDRNJjjvXgSJaRCOgSYs6/04/8x0JF1GCSLyO9
IEwa8SdYUfAQ2OGOJbFd6kij1GP6JpD9J5K8D9yUgSzewjGTQAuivaW64yBePBjD
dfcHjoj+q/Hi4tfshPlnlJGikovlqdptebAezRren1z6HMtFGa0tpKA2m0/3atnd
bANdUjLg5v7OOvSv2YKzwWyI8bF6IKyheP36v8LwhGeK0Z17w+DMt8uzEmRdwAgi
Mjf1N/W7oKOa88vqjMajm3Ph/f5aapU/bPSPCbc6Fm4FQWoKACFd2gTcplVrNFjN
cIbfIrdnOjcUDYU8u1w8QXCiTkFytisEgbEiIijkYhf60JX4EqHh+/QXVAEkEpbt
EIILOWhxA8LHt7/jW9kFMA9ggjRoOzwVtnix/PTUJ/c5YeUdW7tpkQaILOzpRprw
5016CetT55V4ejpCXaXire+QBg/rFZn14EI3Bynsq4g1GKGQ47q9vQO/w4lXwoaC
ZvcKl0aFgAE6FVDpyLmrGuFNrouj+E6cde+zL6MHosAfnSPC6dkVJjIZ0sfytm6s
O9cyX2eBfY6GuLjIU/laGUAwegSxR3cAUpUYWGYHRocspIn8I+7MLbAdgdYTRk/z
odLua7wIEhcEunyV1TTR6WO0aqI/sUUyzwVIiZd0WD5+IYGnxIc98i3imboTXi6j
MM/XAMT6Dh6i4mNeMWJTzzy3f+I9lKxj/0oiBWTEYGJTBiyQIgW34nbL5og0SI4y
CxHCK5VqtnJS+5vvg2mUpliMrikRfEXNlSGuaLlNm10eI6wZMx/ZhTkUx3H7xLLF
3YDo7G8kM28pus/SH6E9sENWDgp18UB9Q5INi+WxOooz3Uj4cLbkC4/UHEFKIxEu
yUKnqMwLlV4SJLeOunlklqzN54l0B/pazRzPWtNjijcB8E9rSY2SS4rFoRKbhiNf
sCLttO8082GtJWwkgnZZzcOl6obTz85GHNcaHecKThxBSOg6dMehUzmejLKCsqRr
6r8Ah0mqVYwszsazNZt7v97h+o0X2t/hzLosBRTqlRsai922GopvSJo1J3kATw+8
GmmT5k6IrDoV2fZIvjiOyZm6AbB4fLRVcZqaeNaX0QBUfZozNagM/4VRflld5udm
DvdZaTbEcsODaLyhj4yN0iS5aZ/Iodh/jTnQnYPFVDt6o33s8uOqRZCr6L4QFEi1
0mP0CJ/Wniwh0CpNR1YJZZbm4TUd02uzQelxBCvYsTb6Hla9qxbffTJvFyxznEkz
Jrn2/SNfvR0SmpRsixTJYsnpBkImk+GbfT5mRVMDQePQnpny9+EXhEghgX+N+izV
biY0zpTBSFcNHwegiGj91QwZG4j/Y4iZ6zcxQNQorhW4hCp28DIkf36Vj3Bm9ZJ2
iykNcLK9mRwTsuuVNRybg9h/N+r0ksTZC6oSk4SPIA0otphp13cmTCk4DzxRmsU6
KGUaqtU0j3zdFJK1MjoSZYDnLezAgUrgA43ecwDoA4VQ7GKcYX9n6pGtNeUXBtaU
guhXK0PcD5wjYKe7tw/3LZbomVTad1XtNy1vIpjhPZsWuJZ/mOAVOVp+4ZBHNgdr
JxrPbfUsrpTbEa6wev3zX3WHQQdF9G+J6z0AelvOeTI3G94phYy+Ch5nzvyYYUVJ
7aeD/9l3BxJ8dDhlbgi6Bd9afWnKdC5blnfEUpv8wdjIyKQpih7gBMJaO1VORM4B
XsXvKZUVqXr8Ar9LfUB6fIS+Nj7ThYSOC1eaBaccUi9EhXecWNg07yjkKm0XwJzi
tFlbdER+NTrqJNb0btxuuixThhyiGVbUQgoLr1RribgavDZdu5wA+W5Hxqmfn0c4
YTqtP7yLkHCCMseof0nCklOFw3XjT+h12VUwUnuHNjUw2osogPiwp3HDeWUsO2t7
6gF7yNHAIStjgiLzKTSRj4e0clfDDiEsil/yamGS1Gj/QWnDRiiLMwNpWxNdKvoY
VY7eiS8w2SCCFPJnnlHqrR/saDApBypx/Z0RtXC59l1TaFAI3leXPDNweyxEFnmR
g6YyGO0FnXr9iVxlq3iaXz6hHlawgI/CO7qlKWwMi3+qUqkcMKeTlKIbVh9WqNy8
G6jVv9943M5fpMoPWefMqwFwuPx6tvmaJgR0akOA8Um+ANQTA+FVgVn4nzC6Sj/c
ADi2k43rNxYxiqnLjag1KiCEqOagtGTp3/1ZwEUgB0R8Qc1Ugn0ttmOJoTkw9JJ8
RJc+3rb1NPiTDbJqJCBqUBLXfywUqcuf3pd/4vwbovgKgVnYnHfQvRkEO/GbKZqR
aE04H8BGfz271fVLpAndDgg92Omze87qF86fHtu6B3M5Jl0RhJJtTgQrlnGJIPen
0K4OJtsLvjmwCWxPTLH/W9Bd0w8Wg4m8oziUM7q8W4osulQ+W9AUJ3dEq2jrjqsz
iO6Bx8Cc1sS9VX0UK1yPPQVlUloDCEuYs+fHOWxKKnnncgRltkp5mvaSVgUOkT/G
sIGKNp97vfuTJ7AG1i9PDnVuf3e1VOxTiOd/gztQ4mNYvF/0C2x9JHzlGiKUnATe
5PlU7qfF7ofS52ZEPj43z4pEB3p+3DBTovqj0PknKHyHpNQ+WGJyklWyJhvb21aU
r53geYolwFtpDZNJdVi4cSmCeRzCQ1RqNgfSWM4Swp6Ec4PkYdObBVjRiwowg31L
NsxQsyMlEreQ4otK62z8EyPI6gAve+ucnbZRaV9+tfRr7BLs0O6N0vwvnMP39vgg
KCM2Vp7LGmyFRebP6r7wfhZn13+mcP5bG0pd6rJdOY5hNI8jW2wkW8fadM4BJvVC
bYHjwRpj7tDSNQ3rkZHvSCESVZh7FEH7c0GCnvIBxuyPeEaa5KPxHMeRxTsBfdx1
W8DSn4uuLrQA+v8N1f0WPFmpIoHuazQNIBKcvfu6GmMCKB3wsI0d/uU69uvL5z3i
nRsclArhycf0Z4dlzusZCQUsZ+eiNhM2JfdKWfxImi9bIOPwC2IWbNAnxQhxUYoR
dC+lvcrOPhwyutw0GWI1Ik3Sa+1gV8Z3z/HUI2eQTsKiU8Saprq9zdKVcV1e72VM
N6TX5cIjQTt8gqF96M89PUgipC887y20clDYp9JdfUjX6uZV9RgiO9BYlHq9kbGZ
oqH7b72Ufwju0IoxpIXtK/v3rc5AAIydbWt4dS1MZYtJWpguWFP1mKMnv9AybJQ1
7ex0YgRQwXJI0tq9Iw0F+cPKy0g2ctGEQh4AFg+AztaXXB32MvNXLJP00kgvD9UJ
3zlUiYHFlrFvAIukAvMdrnyOTtJgb99yZLoHr+x95LPa6ZUonBvEL4fMATQ9DV3X
9XJqiz/Ww+mSW+jakKKen6aoLEa/lxUM5NEQn8E8loXtkvZ3nrPfY+oEVdzv/Fmb
6YFpPVFYDxzSgHZnB/xp5cGhJJfZQ+CdWvbqFP+R6kr/oRAJp71ynPQa9pVQCCP/
RUriXeP+jeED8AIyOHiSG9vPBCfA5LyMHkUG9GzsKlS7Ie96FjmoBKL/t9J/pzN5
F0Bl2nTRtI4RBANdiz36US6oBzMu5hLZHYqgfUJ6Tv0FOBN8Nf3EYDvKP9F3OKDq
4M45kgcdDGmdyGi92OSAgIntLCAJenPY9vTc7Ew/b3ad8UEJ+3U+bKA2n0aRP8Qy
bTp3MgBSBQJlEKIo1MjPXj0EYh2aVeypUddispfMxqkfDVKi02QKeu6KxugwVEEB
0C3R0nDx+KxWxoQ1CrThcYMhGcfGtZphJz9TynJgGuFA3z6ySx6nLj1oHUY92squ
TQ7eEuL3d+/iH5FLy1W0N3Y0JvidEkC00yxurWVd0rXuCdJFh9KnRf6fZfhw8ngt
xT0EVG7at/rbZLgLyuWlwjb48Ydfc0S3nCOHeOuhWVCR7TsTfqpKxMEONNe5yQAf
upuW+1GP+vhE/wPl4hikFod++2KbJojpObVugmXjM/rEnYn20TdQSXM5TbxHWARS
FbeY+d/LDbqXtkhMZ0pZM2Gw7164SCxhklK1h0IzydPX8xMW6ExdUjXiRZCcmpKz
0lSb1da8a4CxXCBXeAc3DdQ6TnMipusodphNq/1OztXjHNB/tJUx672J9mgfmbsJ
S468EDDCNZk7f4EAicLCaaGjKN+HL6oleqSsROKvi6OJzZ6pVChf8cG5mk7eglqL
YzMfApSdThDV4GUTJwL+EqaC2qS5fp/fQLKTe7oBChmggk3HmFTVGEsUq9lV2TEN
yDBOCg/rRJVFav8/SBEUwXg0hTXj5sa+sGzJpcnWk5ZNCTs98PZ3hjCkKRLX2q80
EFSrLTtA1afAf83acGKkqBC3ZKV8hekwvu5GoMhD6U/8tgn3FPb0CvCNettV4swG
flDkwPvAJ1hfhLy9EZTEEPdpVq8BbMN8yyUbWS+5lmywDT94y72dIRrY3y/k9wie
4nuhFvq8xgM83nopwHo7qICteqsEomlO5BnFpRTyVvudjr4y2CgfHwmoeHsj/t8l
MKvGAKeTpfrot+UYjOID4iEzcS0oTDp+CJIo9+ipMtdrwLR0LNfpSojJNWWqWmaN
nzSXN0DIrY6DmAiIb6gtSv52mZTDa6bGbToE8nepck5SkHcNHfJ8IwW7mcQD9JIO
fapAr5KvHfg3I0Ww+pqHVtPHk4tyiVF0ruxHA2NxE3WV6BnTTFgFq3doToIRnuBr
0Q+ryo6o+Q3JqevFj++qPLxSmOCehhYegUgD6BCoqydvxMv/OmIiENq5imAi/rKs
VJ9Sbe4kkeNp/V+HBdqK+DGddPfR/u1bn163cMv+3kSX6/NDP/5lv+mx+9QYLWUe
EzrjryKCYJFmiIz5wmOd/DbO+Xnpk1dTvQjwMaK/tQawalYRMvU2szSFSk5qsu/5
xM2q4LpXJi5dZGZN60s8jxb9UvSlhvD4lNd/ZAMM03xTkcA5+qdfQUzQUXNCPSu+
f+KgAdvJkGKcBf4CUM2CVn2CPInkuhzR8jHuaITRv7wHXGnmBXY+KtI79UOCelGy
CpDyFkS5dKgZGghMI2elmpqnZ+rBDeguRxwT6w5HQxRm2q+A1QGq5skNEAlmPewf
0vSV2I5NB5DNrRHSH/5G20Rl/1hTJjSWY2pimNjyCixAevh5qYIAYerqBB0CLWe+
ChoIw8E6dzCiT3LjNDN8tMXTit0mWjDK9fRmf2TP4dzWcnttzKzcbJ0ldFs0EKIv
62q0+nUELNYqkd0mr4aGplqxbrq+Q74eJBsP4R+LquqemygLpvCu9DqqCnKKjac1
NysRrOu5lZg80GsRTnhEEF+VZfsRd4huChK1UVuOYIeHinU7jmC8UYnNTAP5zvAG
rHYix7XdVMuQsCkjXVtFM+N8bDglvC2+tBx6IHhaccGRNevdM9ovyccfY1JLsSjV
W7evujqT6rIPuF/BG18+Tx57NlpI1OlLSxVad1RDgNbSmQ4/ytEbSO/TB+HrOQ3y
U9AEcIeRJ61k7YhegPt83sETTnjVK3mGJWA0DPjWQM2KsBblu8I2Odae5ScjXNJ6
YFqUJQOPDoxwo3Q6UovGL8fkmx/3lZZkicWN9ay4tPmx2ZxlMCinCOt+6SRN+lHt
kClswN1CeKpeEYkLK+PmQAP6kLjDGK6MpzDz8ovc1Y+2gE0PrWF6KIfc0wGMmkDj
lQWHQVLmEdI+TsU9ovSq7XYAlnSjJ2MPeUhc7YkM25A2T8WAqC6F+P2BYL9Cd3fA
MpH/Hymb5glwRN10O7Gakmf8BEo48CXxm3imofVjI20iFAZWSXo0HUuBJuBICgb/
fPyIv174wa9GGbnFhi4HI+whgZ3eH+S48sI6MBN2t6o6QN6SHEYBPv4loFfuowSc
IzuIAg5ajP3WAreTjuuwpDWQ+/vVJ4SOtITmu5IejDqcHszOqxRTfb6+HUjEDEcf
/KvvfrkIdTtKq7rJVAjNM3fYol/Q3n/zbuF+mqkhvFsk4zVqiM81Gh930tyAUebr
CFaO3B7tl8VIsS4T8LXY5R2RT6qhm2zJ60oZEnBPZJltzevc1ncGJvfxtXIuFfSs
Ei7Syvn4CHtBKE4nvlpuUnAlXTqAsErzO+5oviU0ciFWEEBaX+YavjHest6TaL0e
H98kEa+T1ti2ySVOPQ8nVPOlPGNxJLXp8JB7fSJwcYQzE60cTDol9mlAQQcGiWx/
QPAfqPpKzpqwLgZxGUejTt7ZIIpi6jxX+jtDzWl4vMoqqjP/LMVs/w0K0fmqixSC
4jTT1IaKnQW/Jd5gyf/ZDkE7BE3DNYwXpS5008h607SYgwZnnT63zuNeFkqQChaH
vfmUMc6T7YY/gz9hJ8GANWPRIWpM227OfrESy5zA4ffwy/tUxITihMibzZ8jjUtQ
WoPdO0kJ9kQ8aYmg4zaRg8LxgxNJIqjX0afTo879uGMTOCSw77+wTrLhnPh5mtaz
LwaawpoukeMtZTJ9LivA8VkSzwcJByT1aK7+X64tnXJ//u1ZBg4aOzfBbGYuTuMJ
rZKq5yjeOMK5qVFPlGjWA0fuXNiVCXQ7J1zFbm2MryBch6RAmIJMrp0/lWtmO2MD
buo9otybrkJEFfYouEjlEKI2PbjDCtfzxDtZMINPc+qdBAkkGD+w3ZPSs4VL0w7b
flDbIU5l6wfYh3W0BMzDxYOBt0PJs+fH7sPs/jG7iBlFqDRXHgoS/03n8brAZ5KT
Z+i/jJXguwF1XfQahf7UmVbC5zJ/woiyrfmuPwuNSZtEcktibVLWkxQbsfBESl0m
j4g5QQjSzDtfpfH2MIYA1GJjEAZ+/wrI63qKIAqEZpYivEpNut/IPAg+wV/fGM7Z
SULSk6fC2ScIRwobIWeRQInJ+wiOP9uxv2+akE2D45qSYr1ySec87aSZOCoVuumy
4I5W6PBZdwgwJMq3pWWT3zCuD2VSLR/BYsaAfFBCpr5Pq49g/zvufd2e77lDtXdM
m3lTFwDxblDUa6pEvZYzmL4AuzowWsVC7HgzdxTieuxvO5Qv/cShNYE0AUpMGlA5
Ji+BzbMSfYIF51ubt+AJxnBMXZRsiW/xWncfSJS4ZxJyoX07kWlrNp/uB55WtDjR
H3DO/+ok47XdGdFd4ilyWwJCsEuuligryOGRbATVi4uvH//Z+WRfIwKauUkF7M0D
qN3VpN8fBkdCVjNpue/uwuUiGuLoNqHwCRpVqX+ZuaeeBfV84xYgbV6dJcUcCft8
qgt56V8XHj+pIIeSv6to1H46imlIP6VYkG6wuhXaOMlSfWqu09wD2JvLVyNdBvf4
tKrrFdEiAj4eV4GEGw/2KGTMHR1l3JeQz1rmzUOKNtDo9F6OWc5EZJz11Od5GBJ4
pA90LJI8ih1Ib/Fdz520ai9S4pdYwx0WfcMAwCrbFPqfd/YBFbpKVw3Va3p9uFfR
frqdNkME8F5MGpFeOAgeaLf1QkRkBm4R/wM8dR17C912qRZE9UN13EsjSVolylOc
pZpstfkoyiMJmFmYUbljrbrAFDFcvQ0qAhM1eP6gsZhTo7RR0FPSdohRWw/ATzBd
ejCscuqQJPlp6fVABOONAlHj/cXXw/nR65p0IvOMCk9BEnyhUMSq6dBCUmTzHPyv
osgZ1rlVkDM8jE0ZAuu8vSDsrBQWUJUMWiAPO/tjPQ8XMAVn66rH1YYGXTruJHJd
5usQRjZ5FqME/dJ+lz7nyEayRW87Kzd5s7SgVAMGXeqp0jZNVsdP3v8hGe3qr8UW
hS0gdk9ZFi+jD7E8Oen0qkWVIcJRqMu2lMow2nhsurB0ddbKxZaIPI0jFW0TBJyc
8txqgyLwdIcVY6XG2484SOuzpmgy5XLG5j6Qold+18yXx4wUAfc3m2Thjue9ysCc
wuQu1y9VJm6dDhSNW1pjJigpiwTGk/lOo/0somTXIeWfDqjzYQhP3aOgD1Fo8BL5
abTzrAuDP6QUmHdJi0FfLDN/yFdLzWPk01aEZFndnHS/4khY9xpzsYK/F/81wDvp
V44HaKWcE3n2p9YsC0J/+z5y/kOU4Od1zSBo5XrlcRY=
`pragma protect end_protected
