// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:59 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qt9r3g+0FV+fP08b9XluW9awRNsZRv3aKbaqFnMSMkoHrRjR3qdL34JalvqoCtqG
8AbeprPTLtDai9766Ruyj73BPwxUPymy9QOQaWb+TaIV2MgV5EjyeBrcbVTpPuVd
ijrNq03JuA1Uk+DDX9Oj5eO7wJBaV6s2dI/EhDr7imA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14992)
NUU68ytSjiFHX7tbsRnN9rubAs77E4cz83sZVfPEfbzbCxyu17SMyeBFg4i+43q9
ALZTKje69eUjhXNO+m6Xpo1fEcp2/eV6kfjQo5WaFx0tLxEYpbdqKbc0wnZ0Tbf4
9ZTu3v02z/ZLsM/S38pHdqOk6RZx1vSsRmyFcuwp+xOhOcxge4BfHvYgU/UIY+3Y
PFULcjDL9LzohvX7IKdErdnIQA1J2uzzrATGyljhA5Il/R3eHFRoWNyUZ525+6Hb
PZHePnLm1KsmLmiOg1U4ME1VLtTjLupwczr8QPSBLUOk+hMN1xfKXaRowseGZ3LY
8+ZMgWy4sWLDcPIeOrPjGuhFYnWaM7l7NNyApYJj4lsRuKkIevrZhv762DTnRcJL
9cMk6l2IFNv/BPSuau68NH+SM2MWTg/N9Fhv3Y8KaMOnNoQdzYRtRGaciamtZu0G
sFXNmg0dn+4awe5rCtLpG8vKlQ8p6641k9nO6qPqY1A4iABbCrYcKzDH8OAskDKx
Hu3OJ1G3wHvb0J8LFYN1TulVyv/OtIlHSFsbVsTOhRYg5nZdlNfyI7dEo+q253aw
SWVtIWLurHITRiVBD4iDZ5y7O5q2an12ub/JWgxdeg5QPCj7e2Fyvb3Sr16GgiC9
Uq54UgXs1xi2zils8rRh694KxOMzLZkzt0J3VOe/GcAhnOY5gmXvj4Pnvy5DJQu2
njXAFwEmaPH1DroLfTJAdENREiLBlJ2kafUlMy8353n30bA8s/lEffckGnST1rsZ
67qtNX4LBx2KWpBNmav1i0Ig6pHnfHrcjaxZpNmAnfqqI1iKZUxPcPK9J0bJo18x
C4IRlC9+0j9pz07zmGE8ZC/U6YaX4Bu/1OXhNMLRSUn5m8R2H53iDUcH68+aGsKj
wn/2GmUVOrFbblZ/0UisWzSjaNpsKWk8dwxV+r8lXN0FhGwfAHMTfwKKPZIkwTsK
rdsT6KW9y/LecdTMiGug6A4U0OfRaPEB3A59nbOoM/SOR7QLZNtt1wQGw+h4SdSn
FvSPQm7eEgT2CS0HWVG6uKU7dbBQyqYcKctvCjSJUpwKk5jDPFvwVrjd0xunPSh+
gMz3ltFBA4XxALkfxZrDLijncJ1x/a8tlhOPfQbX7Vs1Wug/pbGiAWiHQxi5eNlZ
1vT/u+8dFupIvWEm5fyUmBcfGETsQAly0LgZVw9qDXznZXCwGNJbJHrUPNyu+2Vd
tOpIVynJ2neNbZQV8nf2gyMkH1nMivPmr/ecHspe2xdxbB03O+TTzpAOGMC7H369
/QXafQsrB6rgGS8kAX5dSyyPaf8Ron6NCIi81aKexJ2tVLeW+tpwKraYjVtzUZRP
wOxHHF60eV1gm2qvAcIwpuArv6qrNlAJ9Y/FmaQQz6w90k1p263AgXIX8AyaQVoo
tX4s7Jr500VXbCsIqtDpsF3anKiTqQLMSvvomTWAMttLgApzX8AQMSXdItLpkL9q
citoiUEcli4K7TtUzW6uv2YwwPmidP55KwhSQW1xrmTh5/AlMU1GbuAe1vA4Xzyj
BtFtY3BxP3FuOgJ6q8eqfA5U221uo/FyCvVczKaC6eiefZoeYqEKEPlOqMKdlgMs
QOwSoVjbIIWawARflph2hoURt3/Iieumvp5cNRQgBqfUh68Mm6gQZVxNaVUTOemy
qKqt4F36VNHyPkV34tRf9eAk0Iqj17qS6VDw8JveBfdJaW83dWgO+3JSWfOXu4LD
Y/eu7spqz/U6J3Dn78002PGkUWW4sbvCfPcL3YvQiH8qFwHntRMHIanKGeKB3GAz
PLsNfFerrels1R3tKYDiv0BeSxwRr29y3JrhFvd56WlNQEfqBUF0cusngTM2m0+l
gK7wyP5HAZFxN4hY2Ez+1kk3vEG2X/66idlVcm+Dl1APZB8Jn66xP7hjOfegV+Jv
Tql7bjhmdkt7CTKmCc5KlJ1G5UsO37n8+pwjOhw5QUzLaeOkMs5QOvjxQcTAuG5w
SKcBaGOBpHINT+CwkusMKf7W/Mdsz5BWwcM//sk4UaSFH3DCh7xwH/mRkzHWTwE2
A4c9/FBZo8cYPaZYdVcjtjPLT4fLzy/0lAI+b2iev1qxAndaboqUGfUPg825605G
0CzthDEzrSdCSXHF8XNKX/1f6oH1xGLypGQyzsZfQtrRIZe2c1y4RcVHbddhqF4i
CCtlpAXQRUOmr9tgcoZiIMGwoxIKwk8vrY08NykfJpo9rgYZUDqOkGPNkRDZRxmF
+viq6+wdQ9DZ9UcVDARGskX357wyI869BrfZEvghSepMQYf8w5A44pa/BQJkYC+j
n+cxnGsDPoTH5M8SVslgGyIWGPsMQkqM4VhKXxrv8kEFNSEcH7gJ27y6CFK8XONq
4T3MUFoQcFrBm3Heey4Eq1RI9O7w4d/8+rWWjaaSKIgADe429D5O55TcwxEbhtCk
mSZ5L9EkF3yJBtQLxVRQ/nSIuT0qH8oHZK5XfyHllq7df3Kzo14+5oD/b7vZcIML
6R/Nm18werve9QUjo7CpcEjdnc9RGTSR1ElqGzO/+6eDYNX6QxjkPJdUEGOmPsis
9zOCzuvqtop6azDhawSOEI4k3QHftN8bNsJaQ9VsyR0BD0grNPgAhznsPQLF25ZA
f9/d03xTlEDZycIxwT6RLeushI/BzW/iR9Uq/IVSUWBg2kA4hHjgLZ5Yuaknvd2V
cidRyBMbVZ7DetuIy2Yl5SctugyLeJ1O0GWkYowSLQjsKRkAsgNOgMfwfphZxMMu
zQN4grwCuOm6Bj3ExU9KXPlZtO1uaveDIuNwdjwIS6t12J5mMYFJX9rv5m1QFCVA
GGdlIvc9vESosf5YrZ78FoGZzXk8pjz568t0QlkEOxErYbEkSnqepNERD2BNlD42
zLp0+YlkanfBD1gJx/sOaAbwRu57KsQ53tD+/yD+o5ZY/4vR3LjAu/nLnJCROtsQ
2X+arHb8i2Ohi3AEvMweLYKqTr9YcHi61WPHmEOvUYTuF4O3830dLqdwA4stCm1b
Exvld/vGrZn/plXB5f8ILOC5vICNlS9tezxdQ+hZ0kSo2nctYV17d524AkMBpfRE
pP9rRTsA/HITUXm8uwOjeuUXXjccipYmO+xtaDW8gCq/7QK0m40qoZZP2Rr+JTkN
7xl/Pa7qaye0s2mHFhR1Ak+xCkrMCulK4QqIaSVzKSUJ/nZf4N5NSKrgzHwr3n3W
l9LHrT9xLLbpcSZ4HAcvgISZWI3UTmbaPOEYksSrFYWXAJp6wo7Jh2BaDGinJhx0
zJMTeRMaqbeQ+/Gi+jvNrPwSo3NxKgW8yu0I6V+2F/a1ZHB/fsrtCZ7fUbUHdPjN
5cP8ei97ofjCEhOrhf5jRl8TTvJ0ygQVsV0l7JfF6nqIkZcxnDJbyMPS1AACXEwQ
1AQ9KVfV3sqvI2B3XzdREExiIrpxBaN1Wtdw5Ht1ynL0FhkPhusMsiXPNgwgTMrZ
hqUCjSIs+B79U5XK6p/Bl4qKfehsOqU8j4YvaxW580U6EZHgpaPPYXVjWTBRD3PB
N6d6CNmVv0aVENamlsc3/h7wbQidnmqz/Eh7eC3RwxsiMO5dsNh/l+y6JKUH1pMO
6qhGSSSqH+SOSOzu97QPPtriP90Yp6kQjsTtHISaJfag9KafAUXK14+y0gYiH/zx
qlAPuuP0JKMbFrS+oFyWwAm/MlskWdmhGgyL9awnnDaATygg8DKr0V8eladP4GZl
PXNYxGS8onGbUVglobVTgmlJOTrrA5tRtUb4hgG3KK4azVlE+yGZnj21wUZ6FqZB
eLJDB4wD8qUw+oISbj21gcl1jn63zFa06Jogs2dxtAyBaPbE2+6jsA4+mnStnVRH
8bpoFmOTOXIA+Ccv0NLt57fHEMahB9xj26uohZerjHlmeaSzZOnmPh7htWrBy9AJ
k/CL06B/EYx+F6IypYkDZIReWrs0x+1/QjUfi84cOnhOgoebWXAItoCOYHlb1faS
efU3Ladt0OCIITQ8O5Ujdnt2o4fVaiGghpGeTztkmjQjrwmjAsc0QOLWUHdFF3wX
i03DC2wDaRmVSGH9PhcWtJYk4KYP4C4p+KHfNSv4/KuZQ5vBQNDniHFeyycv7++t
j6M0+tfJa9xKLU86qFn2y1C06MjjMkMyfipCKNa+/kqnmzdB6vTsIwdirhdUDtzP
pQ/zW7Q9thg95JoCnGbeCReZJOvvRwrCgNpbZu11UQ7E9X3szkaZ4l0BN0vLBZxS
o9PnF/3wPhoLBtnz80my4H5eZv3lM/ZtNqnzHqhLpP/dizQEYL1vRpYI/tByoaav
JDU7V7Ru60CYSj0c2g7nJTsU628B3rfra6pgHoypZiKla+Sh/+Uza1zd/OddGHSr
shzZOu3AfGp6zBafEJd5FCvqChvNd88LRSjeSZjAdCEK2VY3GAXJU2bAAzkuYczA
mEPTyPz0ycDCvcI3QXtdIo9ZeQcB6nDuHXNeXk+YsTNNJBvs9uoIuHHIuDGINn8Y
ffIYVtfCR3qCirCcxvHLY2rW+Palovq3Jt6QTsZWkq9jHnrCdxKJiURM8BoPUSNh
H/gjl85E+IeLMrJQftmPe1aElcQTiwlKGPgX/okao3uU2ScHh3V5pFQhp9ygeZHa
wspq2Icek4NTSN0M49WftJiXIN5aQTxRka99Gx9bxtGoJb9umqJ1ZRAmUCXLx9Hj
Jxfw9w8B5K6yhZQk08RlkTDA+arIxnrn/nYXi14y5qxIxXZTyzxy0m/v8JPUEevA
nhIa2Nya3c9jdtBL4cCath5suBmX5JmIQMqV5KAnr+JXtx3V16ZWF0PpoGkE2S3U
D8OWEwdGkMxBovzYmzdmFW4bqTvrR6uKxZ3temKsWsUsLbMfCpXvGwCfNEDJyEmH
ZsVvMDHpYilGQuoKzzxg/Yj9s0E+e0NvPGyzEGG4N+XrU+ppuLfHWrnVnSLyZOId
lyhPq1qn0Ueb+ehAxe+wMtwlNMIjEeIPEt4mg7EQ4q0aTXKMmtsGN+cO5HLADtg0
cBnh1lBvY2bEH4D6KV/WpZMWTln2dV47Yr0gXDmHP5BFEu4Se/ilqorPsqzfuxaN
vP6+GeMaGg+G09Ceg+5GB4epWU4N/o6ojq5gzhC/+mHvRfJ0I/CgKX3PWYO03URj
iIrUZhkUVTdc9wxL1TMP+B9xH905Rhf0oHVxFrnfXvFy1IboAwwLlb9JwTeoU080
xEJLzCopFOmSV2O5naG3mcmThYaNK9gO+xlGFSfJzugX+bOiwUMpDoDjG/sTvDxD
qOqYfQKHtPh7X4z7K+IT67AwWnc+Yg9m5RcCS4onp6AmK6IbqPpTeFAoVJ1YOLue
89wRTcyyQz+udzU+isgcGGk1lZuSATqG294ORmO1BZRgNKfjuDT3fe/DUCvO3NuR
oWtAFsOSINieNY1M5H72IOh43zpXaSi0nimZ3Hup1AeAg4Is1jRcvlA/eGqeFv/q
rPdaRdiiKa2TzVp4SW51eK9ZopO0DoIO4XQe8QQxSnG2c9Cu4/E/ZqxdrAM6JEx6
caXyon1CaKJIrYcJeYn2qBbrvC7QUPL+QIBpmGok6h2yxmmFpinBhmeVyvaS4fCC
JmMiTDlmE7aVMdzp1O/5vU2zPIm9Zw033ZIbUVvpPgHe6qi5vfG8ncCfLTQG91pA
bLXuPOL9+Q3RPDT+e3ccz2u+w6hJ/eNKc7k+z058ji1Ch54tNmoeBL6roQ3ar7wG
+B6w1MOEvy8xdjNwiu6MDL9K99CIiJWm1/8ouaKelmqFWA6q5Azm+7nQqqRoc49g
slFnh2+RCYlzZFzvLuicN3eNkzNR1l8eeikQthMhrvDVJhjHDwMRoyz8UzJQqXyw
JpW+9v+QmG4JeKcU5c1a0bB04rk3g2LvQPLJ8h59CJR8WuOgkfUdavpmH/n8600e
cRZJS62fuTisZM8tUyDaPymXPR6J3OhiU2/Ll9GXD07Yztic9NOpVbef3ggntxma
JljcdLqixLaL/tcXVPnzNCvdu7WzjUUArSLMFpxOytF3x/Sc3Jr8ZA89UVKMb6N5
sh7hVTxflePzPAmr0FCVNesE4xFzCYZjc2xTFaIucdjIulgolib8KLL2PBMlqPv/
NB9pqfZ36BV6v0WcQlZEo0iQ2vg2K1zaXsChpKDz8NkwJ1gezJ046yacVwRqJfUh
PVpy4HJMWg3VuL7vDFM4qs4RZbm5g+3xgVtifikOtIIViyS/7Ve3/6Fbj+fzgCqk
VEpirpB5Qf0wmCcFOLVWlrQeFQC8GOqK0kENV6T3Vv3otFzDfLkFvBolba5asVNZ
CQYWFIQfaDBEYB5iNoj1BoJ5qElkomAYokaHua4yG+bcixAvhmvkGPSgL39bj3L5
3FA76JxlAWlLYKFbh1rl4Zscslc8BBiQomyM3sEPaexFFIOz+6J/jyfJAW4MawDe
YI9Zt/Dfg9QmykgqP5Gm3NmC44HmcSneuSSlLyN43dMsaIfAVCOoLUaMN14gOWue
JPq1he4tj7X4yArI5MBgq6sGybA66ymtkVqiDEj+kwQuUso1o0u22D/bZc1Y1Xkl
wlnuOrPeD3icw3F4fo5YPJbxm2vCVzY/kOm4QtIgj6TbYeeQZW8I7/3axVbG3oAj
XEKVKe8lK8SaCbjcjYKhcOWFeN+XkipI4dCWpg94fxA4DWipJY/jT0hiblbv/MgH
gfworRmOyDWPTvHCjdrQvBeT/tKR7REdEyjfL0UNlH0W3rSi3JrBgsnOf0wpkzGa
fPtDLn4ihYfpZBZkz1/l5G8pJLqRkutrjSFIH/2+RxTeE3NP4VZNIXxGwo4qLUbI
584KaX7mHnBrwKchB5iCsJUKc/SNzWg7TzC5nSxgt3BfJA3V0WSvSTgTv0XHOgZX
orKqxfZ9Uqcg8NNrfq4AzyTsZxS9hifcT0Pwb8RitIaATxz1W+DvCanU3DWSku4y
8AqZpf3NrkVDU4oWXphs+MnjFRw3eFLYQJHkhyd9rWTe7e8y6N3UU2YKFw/bZ2/V
aIPbgfC5MX+Ho7kgA0VfeYmrvYYVidXOxZRhNoPxMlu/sJIE7BziaI2KTGBw6Zuc
cXpQyZSxUQ9KjYDzqiSsO8wGYrfuBHR3e88xTsvmTh9niZatFv8T7hCPLNy6K+bt
V21lCBxwiGmD1BCtV2YOJK04QrdAz2lccqvWUo6g46AmpyFdCPWefTMRY5HxKYfe
TXqUY2Zw6et8Rs4/PUuITvFAnD1Cl+FQ878MdnDQBNenCdp0+uT1u/AjPq8qCezW
J/ZdnooNDzbmgnsr1p/wfLHCDkpSxdYYm/uREWGQjPMrd6FzoX4FVvpOAS47NDlc
Vnmv+5wbifTRKq0VY6xMuRqeEjT6piAeYuD3T4chCJ10XxBLgpqZLHAUm+xmpWi5
XdofGf+7Ry3BA8NhNkH9DOGJAy1AnzpJYe/Lm0o8Jq43NIXOpEWrapBiZNQGjqlJ
MbolLeRLnUdUjQmG+h2gT6QiyTBOH/7eBoshLLn4EqAikIWpdj4jMcVh8IpNP16R
eFJr76ECsc26gNr0lUjkdB3UjLSTCGyop1nyhL3uvGjQ0jm9QOV367cv1/Ulq4k3
RjavBl/qJeFECzK45AVfmC7B2r/I2pGy1ZmaVTNJtDrie3NyJwREDvg7Zl4ujpZM
tHnR/qT3b34qvz7pJjlDmdnpDhQaRwrlVM7z39Sl6MasW4JWMkBSMTuuvSSJhFnY
Tf4uwcsOmXg/iMEmjCCeIIC15MV3zPEpU1CnUbHvh04suhkJ3I88Dlba+0qrDExK
MjM0auHx3v3TDA9QpQrXW3yUiIGXdyw0GQB1nWpERfEfoXUhXttJMrNV66X/VZOV
UyJ6RbJl9wURB7EZiov0qyUtaNtao8rO3D2Ubheghn4XZidXq29N7UBiRwMt46G8
PN8JDAlm8Hdb3UE8ya4wN04Zb3vKBYqvSbXtghFuAcyukr9cpIlblXyuqAzkWrbL
0x5jsSByAFhuZeFJvRC9lYiGLyEXFCXg2jhSSjjhuZ0F1TjOAmdZ3VKqFTI7FBFa
SDs3kHYfL8cbrU61uidXWy/RM8YqHe54iMnlhPY/5xXTlQkxlYU18XKNRUTNgUsG
NkzgO71ho53TQGM1hw609i5Zu7PLZWOsmJzexdSJ7EZgm0kFxABZa5iKeOeTeTZK
DbMb2rCTM3P8uqI58d/4XZdmPTvMEFFt64u70xOmPxAbUbZ65kHZu+sH8HHj999Y
tuIvbL+FDCBF2kPaclLVywBffjf0CohryEimRKgY7dZetaE0P/q1fowiOTG0iAQ3
Gp+qPAkqVdi5kbK0IAgOoeEi0AIvuXaAoM2ghMDxTpQukftLyKcMHRtPm+7LyxvS
5x7z0Mmyz99Ju7Q7U86wNaeoud6RrljR5Nk74ECDHNm6gKWMhnnjTl7zFr5vDBzB
KfdjjEoTPvmmAYJ5a8b4ky4dudAsFvnUeeQpRm/r1tzXLCDG3ek4mYmyOjbdZDr2
fguZcNROdN7h81UpjytBq1U1dyNycH1XhO/FAjyrHsMjCFBKjbwFSMmSUiv69qjq
LMrr23hnbMkhHBF4GzarCPOUOHxioXTZRdpghLGsGc5QbtGme3wGAFrxFSoVn0cf
HSWKwNJRVlo/5YjCCiKLwCxaf3DWRBHdw1e66JtnuipE371EAvtzpNqQHYBn0OIr
hU883zat4wmgm/Rlf4AyPcwSw+HUVEjLVWJ8D2qR2xmz2zvI6MSe0RYkX6re3869
mBXMPGCLZJskP/DbvHOPYtkN2pyheY2DUAI9wgFAA16/nPh31UJZvHdD7hGBrHB+
7BztTgADNoODX6sJXwdjtT06orxtG4NuR3YUX9EtwQpA/n4E0dhfWAmKkhXJV7rg
6cP+uPGi5+TbR1CIvrc/OYaPcGm4JD4OIcP+uwUc82KoekkHk1P8nqzNBzTLBEgN
GqP7jLziW0W0KJ+IrrcaZmAPmvR4NyMDDHqchE729F6S/G/jPAQIbBH0VUbPXsvE
qhOMx5eFSNbaM06Zsoe8rGyCccDh53ns/zjBCS7wEu2TBgXDoW/A8+u2Usx4meHs
H6o3UkoiIvkWxeRxD6STeZ6xQvy0tS+VkmeTr8QsQQKyNIAy57wayAm9nlIKKOHu
Cq50U+d27JZXFaDLuv8g4tB/w0f8lQg6Jzc2auOk4SOFnpCYLPYfIYwcW2YfkKI1
k3mJ5pxqOEd3/Gb+hZrY0NPINJ5cdB+x+tyh9wVeoSsbR6Nf3TGW2haYKnWghFA+
EMPxy8Zcji/FnrG3oT5HDzj5Vknb96h0eeSMqWs4SzOMl8DX0ws1CDZ2WPdSfZ6k
YGYW/kWWATj1rYT/bmn0Wgb9CjmEdyH12PE4YCJaJiXQds+mj0cn052cQE9mSFEj
ws9NJG5o3iZ0nDEP5ak4cG9CCYN9UT6I6VMFcMo7w6p3VMSwF6ItCjB6UHxFwvVW
P5oMNeh7ez8U4Bc6Btmv+w0VqTY0OsVjpEqh/KvU1mUaqabKymmLqf4DERv/Q1aa
cZJASSFvMDwQo8qws29K8/ZP56eHr5tGcU7Tg8ariHskYlMQFRwsJg9dnBRpFnJ5
Ev0BwmM/7Z+2AA5e4B7X1CPOde7viPh7VcsKRX/K8BikIgbsGdyCN9mSDNcin6OF
WdhWVLVWGXyaPqcMUlXuGMn6tOcDAZPbGlRX8KPQqZBJKlIgiJCF0h1sEEGmekQn
UPDR0HdRC3E6G6Hx7XoSmu5QmbGOdcTQJYy0MNiNr4w0F1tfQwG/Ntf3CEFfAxQw
LX1EXPTPvMehHIHOmSarCL/+jb5vg3Vd3DUITi3m6pcFxCR5pJ716TRdDSy1IUfr
BOACAvyc4LXO8iU+X0X76ENptfzxXItPjp/FZPBifCelMX+rtxFeQoN/+2kycmMx
nEbsT8T3DRcTsbfFm9LwOKl6LkeP71B6r42mTgERIniOZUhfTfEj64zgUmuFClSY
L3OlrkRLIMofFxAUpHMrT6flR0u5ds9G/YUabgk0Rp/byfllD2Mmnb3xCHQ9pq8f
NVI9JfRsqxG8lWfnKPTTyBfSTJZebG3T30iV0NWiXBPHY3hDoxSmXb22nC/tLQCx
Bjt/ei2PZYveH13TmnKD3rVwxKf170CnTx9v2gNyGlqXSpSknyOG63QIfjZMUREH
B0YQs9lvFwHUzrdoYG6phFRJBmHb1xQNtCvudh+hXZBm4iLi2Vl6S9KZ7l7LwSQA
HckZ/bT0WNqyW7r5/JdyD1xLaxJqZL/Aq+Ti6iNts8TDCdzXu0HpMJsSdxSMcHXD
2hrZenPeAFOA7zpA5Pwkns8lNGwNgHD+ymSm2GNa/S4QAo58byTttMGIN0HhDIms
arR3kky1kDWvgO4sNBhao318k/gg3eVftksfW3wKsK3vW4jnvtvCbMfHDsZivu/L
miQb8/niPdMtfofJBaEZ/5GJgMswH2K1IC+r8bv74rgLZ0ZEdd7+ZAqH1LsRsEXY
23zczDPWXEAX9i8QF+NCOJgFVABhZsF74ETEWyPYdT0Bi6/yikhGbehlKpL6C/Vv
qWq2fy/++LV71vKSZLEIVwthl8NEfGQ9GOL6JAZ2tTVr9UdAESHJB5eEwpIstXau
n153y8S5SHnraFqCCLOTB77kxO9jMSU0ZyiUZx3gTlx+9LYFMSS3wSEcM33WfyOO
8NwlcOobzqkV6sHuKQsLFyj69UNsotMRypY1Z4xUEgpoMljLOfzKpntK0hJ0lkwT
fftqM0vsFnyoiM2w51rV6hHyUSqU7ccAPUIZ9B14HYbJImIWvOxxlyYcKgKa4VWX
jEl9HuUAH+kYSSRpaLCTLhAjUTz5NyfZhS+bzV2gbfeXog3ApzTsmUqwPr+0ewLG
XP9Pe/wudlMlqnbFYlWUXEQRKMfrCi1/rZ3S8l/c+3ZRWVitcPsj61nHloQPRCZX
vYPoyTExKH4AS4Pl6PI9C6SputQ4o20TMCCdDuElXNYsGvhg4v6ZeaGuxnsmEPM3
IrVwS+L+6ODHMUYAjNyI7MoPldqJaDnC5pFis016KmVQHZTsCNwmkq8PpNKSVHgP
mLad1Zb9L52iTqdp0je7IDBwwVXQTWwCueErVh6LZYBlbUQ5Eh5/JIY/e7T9RgHk
DlPy5GhfOCRdFniucBPheBt4GBj0W5JuHWEBSZ1VHLQP+0NGmOwKmv5qKleiB/S5
ZIK04wqJ8Tda7il61PqpVrMzrFpiim7JRaB/i75/EVcSVWEV4+s6/hgSfzk1n705
5Ksc/Kz37K4vzW8KXitYl1Q807N+pgSQ3ytUS7hkHuF2G1QUWlJUuvDOmsIutTzj
ISampCu0eQNcfwkiV7EgAz5qHEmBpTGYdAavteYEmjagBY3c2mYnOU39nnt9UTva
JIsInA8LLF1dLhsIEgnogNwsv1OcYhLjMWd0XXYgXGiISUeWmh7TtV8pl9O0gkEC
h+zd/MwnsT3UmS9xCwE360pKmyZpdrfQ9WR8QOcPsTnSeI8u1Dihf4ibJYMTXI3W
HkniLD4aadhIv862bg8FjdAdE+pMkUAphp2WiGb00nSzJFN3E+1NJziMQMLs/YdF
sf4awhqv41jhzEEdJWCL/CpGAQoEZZvMuRore1O/uJjB4dKxtOZVUuezbmTNsHSf
L0aDWMSI9W0XLtpl2oGo0IF0TEo1Z8FcNd6J/G4t1tDXJJZv1pxqGlVZ+MjQdsYX
LJZU0mSztXXWZVQ9AYKgpZCuonAQBdgK8OV+Z4026p3b78bw86jgSo3iPdaAYP4S
n1RKSXYIdR8VhzqMopTjEETG19hdPSWS2BAvMmjWIXyfFKsJSbuAZigjrGzwOQQ8
VaIi/iG3Ylo5PxHYfTFu841jtppRZmxUkc4BzblOo/OY2mhWhzi8s35pyuuaUZ3M
g95n9N2Ue7M/BRWLIy+XOgPiC2PBuhwWV0zuboJFnt+btbHBpZ0lmB8A9uV+hbvj
U68LZuRIWAnPFu2wRd6OrSdkrnNsi9BFeO5gHp6HUImltD10ZgHO3fXIsZAn4G6H
2DEbi/U3+Z1/tySU2aWIn2xwM387M7ggs2JV1Qg4g5xIoRTu1s/CmpzrvrxJhUx7
DtBNcBLvU1La5N4n3leiJZ+6/eH6TvwwHagkKBz6Xfce6NqShI7FBzqt9SuiCpkn
ms6ZbKv+Qgwb/n1yT+/g8hljVbUzqK8xFaFBXzDf1iyW3d7S6FYgcjiK3naWiVQq
YWbXdtd88sxmLWX+SKVYWn/qVjd7XuIcjKgVSfjTsEmUK4bOYrywJWfNNAg1i0/L
YXF20lnjBlXO+N/eAgrlnLNOhtvmiU+pWGtSplePMnqAIzj4+ihpV+wGrE5t00XN
erQ4WzCFyYBDw7ABi7L9mTh1WF2DWt5LORi95aEEJNqySpToY6ht066xN7/QMKos
CRFNal/GJqwy3ejQ8y/CpnnjvamM5GDk6+Xj3sqxAQMGZfd47/vCY2V9tTDDBrDM
va0UnwA2d9OcZkIlQmopAIK9a3pUxEnx9vUy4Mx0LLkhrWVUoggISn2jTL7j6F12
Qd+5bWeuBvFUCjCTU9Dd01OSs8cQw6yZ+Cb/4JDPNQyyaee44cLQFGqIXTwJ/uwN
p5/6/7JMpbauWe4bnpmd/zQkXWyhYyFf0XS59DZlvUIVTjCPKk82L15n37jp0Xwo
W+eyBmb8NNfPyhIEIARa2ihTgd3tAU85T+qEDC76ZZH6jgCAodfI31ox7a8MuJop
2OPRVwSu588lYrCHA8IswsfF2e+YRThJ/CLEygdcw9QYFhHkMdo3S57JcXXjJQfQ
/wD2G9zW1/68lP6xzxQw6eXoj3T3pRYKl7rtCnA9+AsCOyCdfUIca5LrDfH3oYt1
fXk9GUXRTBRrKB3+I0zQqWz4f9JRnlzM35mGEVhLhCo7mQYWF2SIX0/fakEqVt1v
OBwZNAvRWDpHHvBR8XEDE6MfDkyJiZuOtYCqOFnkPFSlBeshLY2arOpl7UgTdJGE
bp/mxrscaoC6uogsdlO/JK+c/snEG8n03Hy98skyuPxcloq61kFaDADWA1+9VY9m
3gXlktpr/0GjOqp4ViFk+KZt05VpeCPSq2Cxdfn50l+UxP1z6FFMejB34UFLqwYV
NtGwdsSJLnm/Yy4GWYzHtc8B/Ox+iPxLmvCQvtYFSb25RLn9ENCo/AM2EVkHWe1f
DHyQujkikPsSRrsgG9yYbJCslG2Q73rgz9UJ6z/5jKafnfy/v0P+gnTDvD+CG3a8
uzfMhuwtQnSEzh+AkYS5L+fHSwXpedNnb47F+4L4mEpZoR58NS/X2BBavv+O9lfb
6MC0IsuNOJnS4U7nR6qPnVudkErqNfPufiJMdjz7eWXomD0kVHmMquVf3KvmbWQg
kPvt5VkdhkULckzf2V01tY0J9OWK7VeIwL7ArTLTUZO+hKcIzfP1ehTa4MCT+ueR
L9nhZ/CukKoTpzx/G6V5VC7RTLtvIATlgIBUSf7tmvIA/urKK/OAZDiNMhv9w9Rk
tiQqWmDWi2QTXJfc/peG2+6K9D1cRrdmQVvBTEELHowktD9JlbAM6NxSftU1XK9Y
nZCS42x6PiIK3BYc9ZWAZT2ZLL/GZTECoHanwGU59Vxnupdr2wOO0Ov5L5vUvo69
zOVBMVwzZ/lmoiiIMUxhQuQ0OGybfgYyokmMzAft01HOVA14h4sIuR++6EBcaJZw
9hHzcZzl7TZTxK7ZNYk2hymLs7yeDd4WHDqe68at2lCH7+HtwCKcc4GvH3Yk66/I
cQ3ND/gKRMSxoHsL7Vg97X9H0cC2KelI71nmMn0ePZFUbpCKpDcfP6fQOUpp5+LM
aPtOODujMI78eBaMWtbRou+Tl5Z+i0qeZExQAQRvX36bPOOBS8fAleImV4uAIgng
qkpFG/gX0uMMl1vD3LVmQYonLUk5A24M62FtVurH/gdy+PF4BTOT70MbwLtVEiO2
wRmdwQJcYPFl14POU3ROG1pdvsztRz8XGX7GOjgPxBggSU5IjGKNx5GUBodBrqMN
6nwIlu7EfZT3MqSCgpUQEMBeWP/O0WzS0JtuiXdzdTgGkpshkAxNn8USIRHwopM5
ZRij4NUeN6bo3GIv7xkoHf1LX9GZrvGf1fuNz45cqoIVI+Kg80z8Rhb2mHDOPT4d
iTM8sIsj0UP0cBh6NF/+BEaMS9nqc3QOBZcqt6ms9flZdvR1/KY/EmaA/QykKwos
pP94WhhWxAmbhmdkygOiKFoMvkMUmYQwAJTYLuNqimxVTmJYSCUifjXNc/U3AoiN
K5G5Z63ne2Wu4X6aFqL2wnWHI3ru7UAz3A8w/5Kh/wqa8f5bEZgS6/XJeOn7EkPN
aHpS+OS/p8d53noHqBAbTImE+eGUtv7XMAyemw1k2rIHabFv4wp4ZBcoGnS5hHLW
TUgi012CZE4gmD30r4QtlCeZ1Svg2gvgL51O0XSDU69PFhlaxoui/V/XQQwbjQuD
6AsPcO4KEcZNi7cgK9+w2C7COUIZ3KCWntcAg3E9ltv7d/W8XFUcd54JmGLqstAi
RxEyr8wfzD9dyy9oYc3M5OaIphhAi7St3OCsIJGyCKW9ZpBCdKEPQHLg1ITWVdUA
+OnlOemeDU3zsO35QAON2zK0/1DunoOa9KGS8/YVYniIjRkwB9rBJDrIm7wRiSr8
X2T8ix/v4OQKp7ulJJ5/OX8/BWEh8q+Uiupbfi2o0ieDDRTeLTs64jJxcW+p0gV+
WckfgsuHR2kc3QGgDBSC2ZXZkQFWQY4HuxdbCbIHmpcLqHju30w/Rh12ayoKXmzI
UM3ILzeZUDHb/v9AH/SG+GTcxCewN5wXa6YeR6gzff1rOjilamQmg6VUp0pGirx1
sQ6EppvmrCIsS8PJll8Q/1S+0jtKk7UtSGAOeXWtur1ekr4vRfCYqfrgNhLC3pX6
Ekb7NsUh+o3WvoiFn7dVayZtAzgeU64MTi/jsl/4YfRRMvUSJzSTuzmGoZ6x6IUk
hOYRElSA7+wiyO/eNz2fpHRlBYaRrju2GPE+hgAnR8xrQfnzuyh1cNFh7Xl0rI+q
6CkxVvuksShrlGDaWyCiyOB5X80YEW6T8SjNbph2RaVl9+gYH/xhqjpNV8qlZlsQ
laZMzz4rUfH49ebAasFblUd89bpP14CeqA1Npnk3MqY4WDT2M9/jnBxz6MB4H8rE
RMtGmdyQOolaqNv/82cmL660q59i2SLeoovtOJ4JvRb0AmjukSKf2schl8QtsxgW
WkuZ8ogCdLIckJ8dAIKw2cxnaH8BeFdXMEsJtiTCsTMruTp221XZSo6HveTtvKFV
9TvM2MGGxStKqC9+ijzm7nR7LIh+9VqxPHT2YdlOM3bGzIyS5im6uKH2fN9aY8zd
Z4oCQriu5rBHEmHWeOAbmwAPbnCBRSkS1H4ynC5gSM4Qm2pt2SgR06bJBPEFE6Pn
wwzrOW/9zTzL/DbqC08fWu/zMMzGQYIi795NSp/plMZmBygOodBHIV+bUroexS4L
KgpG/SSylBe32uJpIYKnh+nDp2c5p9fZcKOTz9sEqYcKJ+TW43HHrHZtYJ52NvkZ
IaXpCRTsWjQyq/BCknn8HiiJkDC7YwjkjVQpNJ8lVEIcUDq7p6Cn7yFwRv8/bJ9k
gcGRGpC4BZ9nXBH3LLt5+pVcEgLwNHMUmXivF6hNgo8nv2qATMXe6qLbd5lTCsN4
MyLO47ipLYZaAW9dXPBaFmBYLezRVG4G1H6f5aUrt8sgr3QtzAQ3uXohi4RSjfSb
MsuEAa2AaOsiHzYcqre7ixhlMUJnmnpjyGwT1dzXNv9myuCsZZJbyR2kvszDvZdR
2rZrzmjdsP/l2cDkMFpPOyc0tdPXqy9Mh9astBw8zMNlfqTdczz4MDutL0lUQJlX
Ga+d4W1VX3IilXt/L3s+YdTHFB6x2fGPlaAZayAhU55wkIQgwnTOVeuNnYve7zbx
j97QUmbzaEjtEVTz1NiQdJRWZzXwsQD7TAHlmTPY5ATGa1qRc1uFtl1zfmKWGcZL
n+Zm84PqXfutTPbOAVJ4eXWXRUgb0AWessBEWYIwtcJXJOygcmTZGGvAbxurKjpe
7tu5kHcvgmQWyxfqz+0/YmzmoKJYFvPI3G+dBDVufTj2wHahEQtSt1GsOrKS8uMD
rzfnYTPB/7v7p4+iGZLF0mIQe8U5at5iBA7fu4x+MWMyrAD78UeqRZ6azva8ZeK3
c/c9YX/u/u5p4NpMc361USxssKCL7TjCtZ3/yCijyc2I0dzWaYux6j5pl5QGOZIW
6Ac7FPsk78lGTqAG33HbmgRhw29i4cKDRNyW+ImvkePNJQAThuWMe1J92UefrALA
fFHhI3x3jig0TNkYxHVqyo7v0nQ3W5McYkESIlIY8PJA4YOF9iLx9m+BTcZO/Hyg
ihkXGum48MIRbu/KrbyYZz0hXXFcqRyR5gn9URp0z13bi00K4PYCoXBSTEi3b0MN
HAQ0bN9mxM1A59SVRbv+24tWIJsTO7NdQkqygiEze5uwriIr418SafXT0QG5hmMd
Nw86yrKix9ukEFoQqQ5pqGAEB/PD5QhPm3BclRrhKXESTx6TDEM+SWR2d0q+epbQ
yWUuX1N/ewQSB0u/y5XlkNyH4+SxE6pUGs1+8/rgACBhqgZjhd/jmWdB5y+IvrLJ
7Pv3yGDB0+1e4MAq4qdxgMzgTtcnqLNjAw9lbqHS/Tdp7BaWB+9GexgQinGeUH6J
CkRVVtfAxHMk06hXOWDvYflqjvDUqSvNWHNqJD/7DlTM2OXuoLovIEHh7Mi7XYdU
TfsnMWx1FNstEltNzR6rzkAPWpvBIrw/yLFC5v0PTMjJ0K1+XutnxCXf2W3F9EsZ
lnyDSuwavMYlZih1gsyJHa+tsf+E+DC+yMYPl26ilFC662dr+WYytGJ3jodrpcZx
gL/rWxtXwadgfjZsobO0ERlfhDpV+qlYwTOoZ0tXnUlcekOwEaSId9A/dplHvY0p
odL83lXoJ/iUlLvSk/JHJruToybIF56OyTNLcyLGJJx1tQtpyVErvaqj3sIsLZoI
Kr2WwB9c+G/YqnuZQFu/eP2V3SjmmVduTLhifrEbcfPPGg9SxZVe8KFk8BhcDchZ
zI4coooMuQ6/QZ6oOnn/RN1ZwmXPmLXjawfQx6xQEt/fn9Wl1W1eWnx6f2C1xu50
o0vmkFc/97reInQzdZnF3UBkB0lvojpmjlnf4uqJ7uhG5C39DUpraRftklLuYNgL
QQwwZQKmlUREynRVJvnebEc2t78uIsSfZHKLls92DolM3CxKdp2Xjt0+GzoVvyfX
qbmuUr6c82UVp6rWuKn68P9iQG3Tu4utoUsYPAFNgbZ296Cwv1P0W7kUumUsqEpu
Qa9sC7NN0GiBFfVTa/jQewL307/u8FIXn9QadKzM+xwzgcIMyKwD6mY0m3cdllBt
pT2fzB7XBlQEF9E/fWQEE5CFtdjEJ0TYpXqGmiTgTLGbsbD/w10Hlix1V72o2HKQ
9VSfvTe2DXU2OafdRUTzXIjVoSnItKMV6Ak7BuNmeYiXBmCMR5gRrjy+QYrhRQnA
vOUAMF08AREMB7jRAjj3fKHt3fc2D3WK9keUkMhMHYSBiEhvMvUdIuBIj/THrUG7
peXPuUOTZxpua2FiWjl1x7vrE81xOLfBojcs/p60DzyxkgfWuLyQuhTlbUn3Cb2K
e073EypNBo9E2JxOJIyTNAlofAA/rHac6I+22YpRC/V9c9aPRe6L6ILqUkZqtWfN
0NQecZ820BAJOosI6vWQ47lywf4PrtTbJbxWz1vJgTCrijZQCT+nAXmxByoQP7pu
utP7jLHOn+v5/Vj/z7zXOsEMhlre3TlqmRHnXt23JFAJM8EH9G9t5hD3GLBHvHjj
ASqQS8PxcEq7iZ+iHgiN8PiW+5o/7KfBCsWsfV9kMmw9slzKbuZuAbzH1AWmZrxz
tb4s6qh8IbBXNaEIznvP+27egAnEhIgxzljUX3KL+lMmTyX1SRFPYMEdKuib5jHl
wn3+uMRj16jKaoPogiP5EG08lfRrdWdd7V/CFVPqZ7cW8vXc045/n4r8IjvkFxfp
QL4/YBoIroTN5Xehp7shLTuXCj9TfwnnHEnOfAXjO0MdxrcAVZB/SoKMswfQNhH6
inPtLzN2dLPheAcDgN0rBpgJdVIWK53WXTUSoIw56MG5RIT5MBv0meFTypTUVwpt
Xi36hBW7KSWjCOCILBEmCxPlyaAd9/KfyvXpF1ZXrsQYhxionxYkwOdqaDLNZyhF
rkYPg7dPYVPAAJvN3Tp9AWCwvxGyyShCFYIQWhFIEX/X2DylXZ9FlzHgJ/Se5Vse
ZURkLiztT+tKbVYqkOuMlXCnfPY1O7oe4t8SvpJ3ylr04/vOHyJkZ2xy/iKXFKED
WLg64ImO0CfSjz7BmxRpWt9MElAf18nF0IwMBuK/w1BrNgnMcHsbbyoycnAj5avR
e8vs8ZxIe9qD2IZoMyx9Wy7uxX3tKs98cQdjp4GFIUTI3y5d5L9aphM2XPwVv2Fx
YDGGBC7aMItugomh+6dEPYSSx9UXcGLntdfPSynXCVwfmJdXlhJl1mjjX2MBkN2i
aGaBHnqJoy71c2UA1l2TkYTF7VGfBF9EkbI89T4DHhGeCoH9gckCZ8S80jL99PU4
MekJrnzd5lAQdJsl16bZsEzT78yb+T3yyerXXuTZRkoMJUBYEBygvKrpzrpXxM6h
UyFokRcKzaPdrBpp9/w9DVAQuuaqjp5DOl87uYOig/dkwgUvZ6zFWtLeC52PrwuV
z1A5hRYqHsDk/YrTeZBT1EO9Uyia57bU9BS4ykNWXM6MLptNOcGhtoyq7ZB1ovXK
qqDd8Z+6nEXT0z1mgO37hXsOI8rvk0wjtH9MLE3Mpr6dgIrMADaWM6bSkXbse4dQ
5wyOAds6NZXIWzQLpI/aSBvAnc4hvwZCoXsgQjm6u6ULuipAHGpzshg8SJnN6aor
DPZ8UqgK3ZkZSGuuYfjTSCGrbf2xKABpFG04x1xM2FPVP9V5QqHYFW37OvimFRov
FlEKyaa9DlXq03OVTzBCGSSFC1vVTX35IW3tQ9b7fRnwC6qm6QBnqFOGPVTEkj3o
jXXUruHuIkVqGTIsT6RJzCCl+mUVETGjVNY73KTn3hoL8jO48aPCZq/Upj+CMAyc
ofitNSVhLG9lwM4p1I74DDwTRbkvIdQTh65J1c636MNBF0bjvio7yzNQ9Wm046Nc
bo+F466tA3IhGjyvRMorUU4+GxwbI3vl+UVxx66SFieFWvH8cpEZyTSkMAEI6+CQ
bqSpInqpP6Ji5yttxkYNuj8i+JHuxabxtoBLL9BoHcyM7ozbwiiDhKVDlccRNI3H
0KwkUuoRzX4j9mCrq4h8xgH/WkD+3OFOO5JSJfJQLpsapoYua7pGO0OEt8Iy3gXY
pZUfxgd5figq2WerkRq45z7cOQOhWU/8hnSoVqmgSIpXunDkc3QkYkEXXCV/HQ3/
kYiYIW2XfHOayVdMQSe2dwG7Qnod/osrp2wdcPPjHrP3xR+nQK02vsfxqIhXa28R
YytobeQl9/Acy5m8SXHaYCrhQ4qLD6dBqFpmwJc+mlssptojUMD9T4hH7KnhMhbw
nPuuPMfcKh6d+mVBCq/HyaXRB0lVq7qak9fdp6/fJDrOhYhwjGawn9wC3Hc9whGX
crWQnQ+/NdPPocyYdgSuNYy26Cb8mDUWxW75LYzOpcX4No3LuoiEyl0f0Czbm1GH
nDDcSTEbHryukHYhjJCkUpSk8ZCJOKW57Cw0Qpik5+mRkgUYu8FbXo7ZOluvNwfM
HkmjzRGjmQ53WSgX9FrMTjJg53c+q0uYBTk7Mq6Ulg8CQH6AYYAyTucHK1fEXut+
Eyl2DKricznB9fjOASaXFUrDnsi/bbRYrn7Fta3m2oAE1ko/bX5LkiEJVx44k/us
7X/G3eU8zTKrjThCVdt09PlBQybsfEsRxXc/2ali45zmlL00Yu/C3Q9+n3z2Ictg
48rKqPkoqhp0yoCCso/JBSb0iXt6I0HSkOLXmXJs1c6/3A0EEnxJbknlqWX83zYR
EQtTyMDEpp1Ne1sfv2N6jQ==
`pragma protect end_protected
