��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����Ղm�SF��Gn v���.����.��Iq0W<|!�έ��m�ŀpɚ�մ�����$Yc]9�Y���?���7T�SJ(�V�|jt�/�e����-1�~:d(Bɦ/�3D�$�?+p|_{��	V�;���:��7�Eh�-j*B��Fc��6g*�MC"��e��Tl���-&I�֎/3�O��sz��D��H�#�X���y�~����0�b��a]�t�T�3���Q���eH	�?�	t�~s*���O�mY�("�?i̦��S�G�9^�}?F�����[�k�P8>?h�E5�쵧מ@�E�s{F�w�Aݽ�h�W�P��auϕ@xn��_�kD�7o1u�2�~z�[}��y���.���{eO2g�jc���}��TpV���C>��e�v!;�&Az��F��[o� OȄQ.���"k�����FsF��Z>Zv4������*���g
H
��}�������]�E<��?9���ε��Ӱ
��q�!@Q���a�V����h���o���v�dz}GE44�����Q6�Ewy:98|UX�_:R�3�70��9=�?���"2�5|�Ъ�wH�$ow�؎O�0�o4�*D�����yg�a������V�D,k�*�[����tiS�h�*h�]$�5� ��v�\^������	.}�h�? 4���c�+����)�C�ّ��#���3�A}�ѕT��D�M��H]�������Q>�Β� ����<D���C0I@��/�������P�A����Fm��IlD�GfZ_����M� ��|#2:���x�Y���۠���3A-6�3����`41���!��5���=�%Q$�,s]�Rd��u%�̘�ԓK���=�1s��v��vv{-+y���"������XJ)m_V�J�;�-�B���JmD`4��3�|eJ����:&�U�>G���F��龂��˔X޺:s
�� ��mVŪ8��W�_ ��Q��8?��~4~淿�����ټ3�����95�ei~�*ؗ����m��;��.] r����`�G��Q���W'�(
�ݢ�V0��<sp�R�5��^����N�'�\!��̪A_�j�s�=O����Abs�V�U[��J��Ј���UЮ�F�?�by�[��>��؃���A<ǹ��י�b}QƸK�||q'��n��g]!�4���}#ZU[���%כ����.��9EϹ����I�O%�c|���#������ow�V�������'$⨜UgKa�z�Q���j�b���ϵ��%�2U����Hi��of���=�G��	�L��@0��%�d6xG(�(��
V�_s^�j�pߪ�Y���/��5B}hB��L��~�MH)�m��.[Os_�����Ȁ\�w���_ ����y�����C+=.�޺����"Kv���v��δE�o5Ƽ���9�����H它覾�=Dg��ƹ����[�}��4zu��4>��cV�~l3��`4 ���\�= :�@��s����<�7���Ӌ��J�0@M�����ӎ[^ @�+��B�-h��[�����%>��=�0�V	�������[�2禁�K��8_�T�e�I�߻���r�
�Գl<��cfQ�ʥ��<f~�P� 1$P��t_�&�Kf8�`�O%4ʭ�ha�6���E���E�Ss�o�b���e���F[OL@ج[EA8��u�C���v�~̆��K�7���b=TL�4O_��b~�+$y� d} ��mU�EnU(���
[�iu�I/�m�"�	cۮŇMnXY{	��wR���.��u�PW���!~f�)$A����gы�����$B��X�V^l�
3vf>�����@��o�!T7��Ǿ�>�-?З	8gJ+���*� ��D�.��2��<��L����Q���Sx���Xm�;	�Lm&���ա��Z6Sً�H*����XK�t�n�#Rߝ���BV�u�9Ş�6Z��|A�p�r(\r�o��c�W�KB�k �4�7AՐ�̵dT7����s�_��K�Z�a��̇�W�'^-����*`s�5�f0h�_I��y������B(�mG��@�EZ�"�qh���h"�'|��J,6c����E�S:���)0M�u?Y�w����W�5��$Pp��Ӫ>�=.{�)��-���D�K���+H8�?�Pf臠-�$��~�iN��h����@���XP�U�]�,��$kH-��u�v;|��x[�]?;���|[�����B?�11wN+�����5��W�D�[T(Ӛ*ī:�7�A��W~?��:%���+q���:�q��Uu�{�Ԅ.�]l>K˟n']�|�h����k;G����s4%+���!18�ۀ�q���Ń��<�v8t�{��Ƥﱑ!8 �̘c���H�˃w�trŞj�h$$Z���@7J`�;e� ���	.�F��9^�E��8*��)�J��\������0,_\�� �g$!����<��)z��zG�tÈ�L���k&�w�o-�u8�0��9h3��a�hH\��"5���^E��Q��R3�5���c��&�vjuJ/�����͖��iE9�a�菫�팽2*_PQ���O�������?���}}�ݭ)	� Ws�Eq}�H���|V�h�����)a����w�Q���.E����L�DJ9��M�a~��;�ڳpȁf��M�F�UE�*��T[TpddQ]�/��&�Q�(X��?��a�/�� .[���Q�� ����s38�D�2�
�2����7�ڪ��`�95Q�[Ys6���AOw�j�5�'l����炙�
�gi	9�^�A�Q�q�A�Ѣ�����>ӈ���\/��	���:�2��LM�b�b����2o��[=#�����.��^���eS�c�O,���[��B �J��MX�I�����D���S��F��o�w�����F��|> ���UR-r>��AX���v��6'Ҽ��|�p�O���P@��(�t�b�����������mG]A`��m4����3JA��{��i��ϛva5�['���B��8*�px�  ��95�䬴4t�`KJ�1���*�뀕���ޠ�B�a�
�7љ��|�)3n��������?�	Hl2�x�x�E�)����"Vq��4}�$�S��(&�H�~�q3q?��u/�$�l����x_[���ZSPM�RU���ֵ	�}�@�^ٿۢ����K�͵B�lEp�=��f�˟vL�\�ed!\Z�<g�'q�	�fa�g9E����g_F��-!( $�Q6U�ź�z�R �5��S�I��"m�h�%�(l��c��J���M�~f�����Ir1o���wɍ�:�����U��Y����P��D̈́x��0����E��mB����3��PzO��۰��-�Hn.�;`��>P�|Ǌ��Ȋi���a\����Н5QB#�"�H���# �,:����p��y�v:�!z
�	c�рVQ=�@RNqA���'g�
�2�ev�nt�7���	��5Ү��Q����l
TJ�O�c�]P�&h�j�͈�2��ˌ9�u�T��%>�1gz�v����?F���I�u�H@���\�ȕ��܇e����I��:�Z�0��Qk���b��Z�|��EuKm��3�5�b%�C?���0�23'��w���mI=�gUn�ZV1W���ׂ���x�k˺[kM�(+�%۸L�h���Ֆ�CI��X�s*��;��-���t��^E��F�V������_�N�N��J�A�x$����*zw�M��l��a�7mF�)�y^��+�$���W0�܄ҫ�렄ñpǑ�_���^�0��jo,�ܼ0�AIZ��	E�6��D;J����^~��Qmv��e���[�L�I2��ye�{�1���O�b�1����L��$�=s��io��*�96�Q����Ҙ���P
*r���	<Hr�p'�ʊ'H�3'o������@�3�1*���|/���#��祲c�Bg�XC�1������=������u��!U����3�&K�6��0\����!RW�����10�k?Q�	%�#�aK���zR}�	~z�Yl_�!��<۱۽�<T�)��U�YkC��^Fi�S3"np�ذ�j��q���Fdy��rhL��l1&�k���x8��C��7���<��ky�q�KQ���&��|ݭ�fþ�D���K>�ȃ���S=������͎��Ta���d�|�c�&v�b�D��+3g�<9�"�ၐ}_9`few�\���a/(�����GP[/`l?�E��+�����xD���hF7�/�u������4þ��?ːB^|�T��8G[�g�k�o
��`3����qf[p*���F���z�6�(��^�8I����ӡpĂ3�{�b�B/TrB�x��{��PD}��rݺ��~l��	�e�%��H�8Gy�	(ϱ�;�_�����:��<f�*�f�3��9d�$�W��Zp��8K3:>���_�J:���r-NZ6��䣮|n���k�W8���� ���^�	���2p���ͽ&N�4q�Q�Z���xS�ɜ�4���`1��3/��q�i���s̕]i_�ӡ	������Ǹ���Wi��B�ϘL�W�݈"���n��❟zL��L�Q�4� rϖۊ�� �	�3< �p���h��p
���J���8] ���N��i��g�H����w��7��P�Rxy*%���05jt�桪.F��ÑҌ�c$��By�7ӲΎl��������ed�����H��rd;����ɻ�Z��a�W���ڐB� �������*}�<5K,�-{���o���mn&c����x �c9�ؔ*Iut�N�9ww:�FJ��-���~��������{5p~��Z�Y��sh'Nd2�?�7��k B��S�7;o�1��kЪFVR���� ]7��f$˫�K��){B��ҥ���0�Q	凃�<�Ym�EN����J�^�Ϣ�1VJf�q('��jAl��@),�Ѣ+��͉�\����[TI��# �_/��N�r;��J�ZK�1�!+[^,_�~�յq�u\Apa/.رK�\�ZԮ�%h����0|簏�h�7]7���!���d�8�R�Ё~�7�=8�]�?9f(�d�W,e��x�4��T��߼:R	�Hݑ�wL�eI�?R�{	J?
�Ĳ��cTZ~�3�ځk�?p~���,;!{p�B����V���$�{̓f��?]�V.���3������pWߞ���#Ċou��H7vK��4�i����^��wuQ"�o�tb��K���E�r\b�aY����\.(5wk��,�d��y�R�s7�d��B�/W������{25��0����ov�s� 'q,��#쬗�6(�?�2S������t�c��	ċuT�(�m��bzhx�p�����%,6x�T������<X���}�5�ȓt�YKi�9�d�ew���]�h��&M1S������Y&Ԋ]!�>�1������v
ڞ�	�*�%��u��+���!@�,/B�!���~��� NA�
bV�-��� ���Ɏ�g1xd�DOI���n��8�C`p�EOdy��m�$����1��������V�X�e�4ep����ɡZ�yV�\�4�Ze='vd�3t�a�����~�H���J�Wi����6�/<.�^Z�+@�nm��^�L��L���Q'��`�Q��z�ꬉpՃ�,���$�A��\j���Aì�vxb-m���8�o9`
/BLE{"���$i཯5m��\��ۺwŢ.��7������.��5#-(�
Ձ�O�%�GkC�8���$������H���^F�����D���o�y��]@J��W�6���@�V���ݳ�)CV��.�|���`.MSY�g�`[d�ao�l�%م�9�xޅl�;@����\�ZU�٥PT��?���®����ݚ�~��z#�f��d� �Dz�C���\ӠR�O��lgf_А�^���o��G>��!'��	|���ګ��:���N��0i��n�@_�+̠[�Ӊ:���7����6E(N.����~�F^�c�a&d^?��x��Q�(�!����Um��B�F"0p��lb͘B,�٤������T���!�VT��A�"�r81�^<N����i��<��W�޾Mm�qB�9���,˰�s}Z��qf��o�Ht[�k	b,�m�e|P�z�UtY�5�@��y��B����U�#� �\�
PQ(�V��-��I2(��r`�^1��+��`x��
6�{Gr�j��H0�i5Z��L��D��y7���c�H"��N���$����P��u�^�a����K���a��{��_�/�yz�a ���=����mH�}��%oGM��26qv���<���
h����#>mB��z<�s�O�-}�V@ɮ	^�M�y�#��5ce@��n��܅?�` �l�:B����Wl���Ǘb��<�7����a���A��wAC<i�n�k,i,@~�*ʽL�:B�G�+;s��!~��j�"x��}.i�h�;���E�C.3�K��KQ�2꜠$�*�"Xo\G�I�Z�
�V�2S l�\/�k��`jaE���wBu���1�KL�#�s�K�";��*�C�pb���N��^��r�����_{�:c�z$˰t[dߺ ��F���f���"Sӭ���i҃�h;�}�p���d_'t������Y���Wއ�a�Gþ�|�:n�P|�E��ݰ&����4�p��^.��a�Hu5�������g`D	�[Wn�e2�}�1i�A�X�F.�X�9�dcW6��(�ҿCeس���T|�qPL!�H� �]b��1B����Ѩ��ʤ>�肄�W9�����5�~>o�kΎ��v��R���ys�#�$�	sA�I��Ԃ2�+[�#��ƈ�$K31v6��s��,��m޿�1�Ɠ��u��l�QTI_��73Wz�]�����u�&]�B9���p����>'-�;��� ͉�c�P�����-E�D\�Z#�=�\�Qd��K�&�ݖ'%<��]�f+b���s��S�\[ʞ ���Af�br��M�Q��
�.���7Q��2�SK�H�uѮ\e�����O�hԔ�N�k�����6!$~m�)����w�Sf ľ���z�M���o���B(3k}���?�f%��!i�Pg�1�U���h��8�g����6F/�>/:�6�;�;�I+KX<^��s�,�_�M�]y��Q���v漥���Q��Ay�9i�Y}��W��E`'{p��E�Ӑ�H򐞱$�&���\*r_�X6��I�	Ǩ��onm9��'Z�"���A�ut��N�Bt�W�PS��'`,��� ���I-7v?c�ӆL(��B�bH���u��n�HZ%8�E�Z�m
*G�
���aۑ��_���r�A�%t&���,��F�y�WY��|��R�5;{9�J;	�t0'�3¤Lk�z�V�%gԽcD�����:H�rc����3'�9�\���ˑf��<-7����^Tem�#����]�a��CV_����;��y�G�Go�E�o�� "v�[��D����ҳ��)�$o���(:'z[\��8��'?1@-b�M�,��SW�x���7���:����3�M/.�U�1�'�7��`%[��0�Y��������R��?�n1�*~�/����!;�쁹'��<����|{
�6}o�g��<H�~��_\-�Wu��N �lf�5�����OB�ٍ��r]靚IbtP5d@�W`�����&,�v=��t���B�⣄E��.�w�uߑ�*�N�/�v��bXra�soyIi�|Mw�9e��l���W�"L�u&VbNW�h����晆b)^�N%��w��}|�� *�i6Ȯ�����.����n���¦�x�4J1���� �?vN�,Z���������!��yV�dF�8�>����ڣ�G���2����s�"�ON\��y��ZJ�Q��S�\6�<����:ٱ+���:��nVC!��I��<=���#��3��#ÐS=��u$
7�#ޖF0vgy)k��ǂ��$A&�·t+��}Oӣ�e��VVx2�>�+5���*t��2���s� �AU0�4���N+x���J�|��k�R�qM�_�\K��ķ��DBy�UhIA��/s���b�X�>V�#1\⁏����2�QD7�Xk�f\�9
p����7���[�?�����'&��S�	B#ZA����m�F3<h�������C��Jq��v#�@��|���[e�}W�n>I��I<dF�[u��~e�P�I��L����}#�ɴW$-w>�k�˘����)��63�&�
S�BT��ER{5ɘq��%KwՇ��/$��}X�]����.��t����F۷+��U>�1���Ź=~�f|R�E秧��-��!�u\��[:� 8�B&��d�����lԮ�rcnG�WUG���[��ћ���ڛ���co��UWV�:1���j��6�?w��~C��Ŭ�E�G����E���M�ǖ��*U��|pJXB�b�*��\��
�O$E�̘�M*������H�[7�W4zT	�q��������u����b�{�2Q����L1/5�&�u�E�E��]��6cՌ?�X�ÁK?�}Y�ܵT�E�J"���"�%.}{i��]����&WB�Hh��4$M�Z&3�����~��GՋ�t��\e���l�;�s��PB���$CR#��U>�T�E��YA�d&z/�C2	��Д�����\d�*�d��)�݄�X���.�6
�m���� ��4V�*�J���S`�)��@�P�֘YJ�<Y��q�s�]Q�#�;�:r�	U��᠓���\Q:�˰�:��R0 ��v�\U�B�-���2�s\��;b�O�՟���@�څE2�E16�ݳG\c����	��(暊�]��翕��[^]7/��W8� ��Ⱥ��=�9�
/A��qITh?�M�x���ӓ�A���j�f�C8I�)�9,=K��q�S�&D��g[�Ļ��4�p�L}����-G�w��:­���쌷�MaP�)"r&I{zg>�yǅe	���LœY]67J�~8�b��9�;�|l�RJC������^��B���w ���n�X�+)���x6N  D�G��_%�*�c2��lZ�\��sXr���|��R�ҏL9@T3AQ�Z���T��@��zM�V���U��u�Zuu �@GŢ�;tx���i��p�)�j*�T�n(���I�46��w����[��Ѐ��a�h�uP�y �{�O��Ƚܥ�Im4j,��G���6r�_��ʟo0�b|"	b��dm`�U2͑�rɅ��Y�*N����8T��4���ϥ��pTxH���+�&1�.%֦�Ѣ3���^j�f�Û��f2e��Y�<��vI`ɽ��Z�N��G,�p�Sȷ�OV�(Q�U�'�7<Zy��h���c�O�X�C8�-��ŝ,�����t�����e;%5��mY�>h�I��ba/Z�]S�j��i)�~{��pӽ$���gO`f����~�'	L�F�A�{��� (4ކ�����n������LTC�2W# o{2��~�횓����Ԁw�/����67[�Zũ�f�>N��r2�d�霠���^73=LEߒd�!��Nu�����PA���&�ps+�)��.�4��M������#�k����T��~�0� Y>$�q^d����mR1\�|��H
r�s�Z����D��+�,��j�[[�;	�{8ɒ�(��3�Mߜ4VBD����H����ARA�Rmm3t���M~J� vZ���(܂Y�Z|4�?�׌�J9N�����Sd<�_�\�k��}��/�)�POy��0��/)���酪T���K�=T��r6QW{��A�X�OdX1��=�v!{��Fޣ����#^&��Z7��v �u��,>2f��9bn����N�Y�{�\�sO�p���՗>Q5j۩��G1�g �� Co^�������Vp�M;��eY�\�1M_���V��m�]I�(�Fzx(%��a}�l�.���Ews�9�^w���@�x����O�6�t۱�w���<��b)q!+�so 2c�M�Ϥ��Jr%F��k{|ϙ��0d�qѤ� � fm�J� %�;#r�I�Ǣ�~E��.����|	��ř�=z-�Y��VH��M��F�R��+�J�&�������hi��:�T����P�c�+��rn�%�q�U�a�S)蹻K:>M���g��]��PH�#�rM{�%���{(;B$u�e����R=�[���#��9�v��'�ٗ|�#���v�Ixt]Y�I'�c˺��C�lY�E���I���T<(R�j�1��ٯ��G���.�ʌm�9A�`d*�ȘR�G<�E�SL�hV��6O��6�&�c�i�=n���'L����|_8|L�9�>]�o�vm4vm�o!)ü0sm�7a��/�qB��O���UTO�g�� �'�T;1rT8��Y ����M��CV�xo}/�q�b��>���KC.�u��ƨ=tӵ��ٵ�M<�D1�ߟ��b�`��a�AK�4�ϻ�8!�#w1�XE{xF�>�ړ�� �N�|S.}`�~�7���5��G�Ӿ�K���'PD'p0X婂�#�F�Χyv�<�������F	����-l�M\61��$�Ap�P=��v·���s��D���E� �(�0>���Qp�+�s�5�ZONȩ��lXC��7D�b��mG�H@j���|�Ѵ�n�}��^�?�+�Ip��7���A^n�~o�Kl@ig�$В�������pH�� ��P�����jW�Z�`�����"�����XG	�}O.J6�N�,�=l��Z����(�L#;���L�yz�|kL!� s�Ŕ�w,-G��3P�`v>& ڑ6���2�ӻLK���a�� m#�.]�@�g�^�4,C�5�:�c���T��p�����ž����C].�j��M�~ec��$$P�钐Cב��=��C�ݲ���Z��w�q��֡����
�`�������*/��� W̴Ex_
�fb���}6�DH��~�EkgV�:-�^s����k�"UU[��ʖ����E+PzK�q����v�|Ϧf�$	�y�v�!����)��@�G���f��ɭ���q_�l5{O�%�p�V��$t� 2�p�Rh��0~FKm�a�Vve���sW�NH�Q�n��<9/=��71�S��%j����#8 �����s}ޯ���y�Ţ���87&�$1����h.��]�AE�/MŨ"!K�2hdU�ZR��w�!F�44�z�)��,�̓�S�K�@�!$���ß@|�Ǡ�4�$�(e�hlp�|��BX�o�HE��W�EESo}v�Lڜ�vO��O$�!�������쯛5k>���5c�$)�h�6��7��8�a	fvSxuΕS���CO�
ڇ�g�J��y
b߸�`A��	��O_�q�< "A��\�*E�\����{�����lX8�.t+34P̒�>��ɱ������X�swQ)�άPY(9���t������q�j��fh������u-/���N����~+E_Nձ	z[-"\��%~�8Xs�T[J��^��7Rl�:��^rzTa�Ƶ�ej˳<W����i^��_��5ՓJ�@�I�d������]�� :�z���ȁ�aM�̠k9�[p��}����X��c�j�<��U+�\Ud���N�����P
su�F�!�W�9��߫wH�p��E����ΰ�/�Ϥ�&��\��Y��8܌vw�U�ƏB���#j�@�AO��O���\�d��^�u���n�1ac��U����<���������Q���xm�.J	�atI�P+@7������O8�b�U>��2����CH'7��2�B�h��Q��+JVo����w�\�:�SN=wPmH Ȋ0>���QB@p�C%N}=ؒ5�"h�C�>l[��M����9{�Ԧ���X���4�Y���<̏�:j~b��d�Sx%>���q���@�!|�W8�|��Mn���D�N�;ꈡ�4��_\��!�;��g��^����hH�$�_��	L���@����˹��ZX������"��\������$��I���yՖa�����g$�ɖ��&��$�YFj� ͬ�z��1��=-��K7����V�I枟��)��k��6	�:�զI�h�M�X��B�:���0��6�0"�q�����I�[��1yn�n�#����-I��͠9+�a_��V6�K&RC=EIS¬�^�%c�M�e(��2(\����$0:Ƹh��D̙׍��]!o'�L�Jt^�RY}U�Q[�6���֫��!lЖ~}B�Z���)�����Ũ�3�n�m�_	%P]��mf�&�M@w��\*�s�%���2P��\h���h�p�z[���A�b��{��P�lA<�l�`Tw5\��B�A��AZ�pS,�`L�lȝ �v3	Cfx���^L(eT!mE#{�%�N����[4��C�"_�8�	�S��p���F��DQ!iZIsy^k����Cp�#=��6~�d��Dc��c6�0���bwf<��$O�=�at	��kw�_��ez���h���Jw����J��v�a/���#���\�e�����y�1�!g��h�8��kf к��uWÝ ��"	RS0�Z�j�m��j�/�F4I�7<VsS|�d�Z� ʯ "����݋���&!_b�o��d�%21�O^l(�=p
���aog��][P:kF����-��L,G���_o��'���<��5x��[/��7�3Ifȋ�>����P��T����91&J� L ]FP8O�)y�؅,���B���i����s� "iզ��|�Qġ����l��Ò�<}ݜ��/��dn��H��k��0����k]"�E��o�7 S�S�A��[�rq`�u��x��בY$��0�>�Ky��M�����3�!(T�4"����i���ꇵ�2�1#E,w�b�]�>�8h�E������U��
�b��"��ǆ�-{�{�y㧅���jR��W*�=L��Hz�^`0�������i���p[ulw�X�r:+=��`T)�׹,LhT��&��t�	�P���
����������@��!)�9�e�|�	}�&
���÷�~��Z�'�GZ��ҍ������F�|+����nJt@�8�ҴTsE�k-�$d�X��x�C91j��ۙ�b�XY�Ju�p!a��Q?B|�'�g�;V��_���֒hKhs�Oe���+�{~dV@���8�p¼��IX� q>Ák�XԺ7��q1�II=�2(2���JObR��ML��d��`��O9��?R,�Ӱ~`!M���>��3�������D�6;ѫ��2 ��u؏���8Z�th9x���K�P��k(0
��sPR��Zu�~0�/}���>�/Z��\�V)���g���cI�8]d#�N��"Vn`N݋�5΄,�U~~������O��d0���A����ԜBӲ7�nA4C'��T	�W{�-���:������w��l�~��A�1ȴ��`Kt��~���b�i����G_P��F�9\bڤ��1���͸b�,�>�̈^�v�/o�x�i~\�@o�lu��hF�$����C������m��������$��E?}0 �"���r�>�~xv�$Y%�*�;�H5m{�X�N�`5{ ��G9g�M"m���/ϲ�y��p���c��)�D��u	R�M	��{�-�=�j<a��31W4�(d��%LBo�'p`Ņ>�Q�y���&&��	�X�H4�Dot��;S�K[$p��d�,�3	~���B�y�V�߹�<�H�?�("��Q����B�vύ=�ª��Y�h�WN��J��i����e��MO���"Rs�L����_}�y]͊Q{Ro?��ď�>��?aY�Q9%�R��\l�>�5���x8?}^����h��6��R��Bׂ��4̝Ho�[1�X�F�����Q)�.$"����؎�ʘ�	�U�K�E`�)Z��u>���a���Е΂r�.Aj���b>�_� ؗ����w�l�9!�6콟�^)Xa��4�Ij�I,�6(��%�1Z�:�G�����v�&�.��hK
E������SԠe�/5��+]v|�!��V|�e$м^m#y�)qf�<���]�o�Ⱦ��$A��*��r������ʾ��w�(���wz�_�˰�Ďt���kC��h�v]����'�N��H#t��S�9�ݷ 9��׫E����k���)�`^F��q;�cY��,�.ϳ�;�?�_��o�6��ׄK靂^iGj8`T[U�D�DN�*�q��ӄ�5����(��`������XHb
Ԙ�U{�D�͙G^Eɒ� G�u��b��4(�,��Q2����\:�z0�^<4�>t�]�3�]�7�m=^���A��\��@��)
��Ϯs*M�wJ4w�Q:Bro KuôȆ<k�������=|����i��\MM,h��%j�0��X��஛�n/���~׵;����E���K3W�`�؛����w�}a0��y$O���*�3l]�6W�Q����n�*�I��?����ޯy�!����$ ��uN�~8/��>�ɡ�hd�Mr��>��B+���p,M�����b��d�)��:L��f�r��F!��u����7V
|��?�K��(|�xB^e+h}&�~��W5T���������~΁d�ϥ{���Put:xi�����/D��[��lk0��	$�]u��%+�6���{}�p���
*J�?�V��#e�Ҳ��s�61@�^Κ��{W)�&����w:+��ֳ�� ��������يٗH�=���U�ј��j�wV���k���S�̐e�5�h��Hh5��?��J�:ޚh��-���7�_�j��s�6�R�~WZy�<�C�G��j�']!m7����D����:�ө�&=!�<hzI,�{��jsyG�ѧ�i��������{}C��^<���w6����/�ln��{��:Q�,��s5;I\w�Ai$�*ϖ��x���w}h�H�)ܬ8�!�x3.�R�$�șW�?A�F���zHn�D���o�KR=4����p��lK�������[�j���s�����dn�n�z��M�בR�w�XDERS���ZXt���Tp���=⥞�D��o��+7ml)�ҕ���Qڵ�Ƕ2/Їn��7V�@�����`M�pW��w�6��Z��6����R=&ڦ4��|�I>����ى� ɇ
�K��5�����2�8sPfb�Ntʁ�����6�e��՛���ST
K�_a�ď�+_K����H5䎤���,1kd�I&�����
2&�a���&v���(QE��6c�2��S ����L?�\��K�v�l�|E,��1��=p���h{�u��L�～q]a�B�ZL�tIxt;υR�`)���F�*NU��X�9���/ZFN���]�[wݰ�:G6�Pt5��.���eԻy)Ԥ�tb�����q?F�	n3�P�8�f�)t��N9A'ۋ��1�JN<Q�����ľ�^��۸E�;�
����4˟W�9죮[s^�ޘ�VT$}���:�qD�҇�5'?��O����*YA�+����o����Շ�t���t���5��敨�pn@ �s��sl��1ŵ�}��r��0>Vfʟ�*K�-��T~���%�qZS������N���H���x�����]��wG��¨g���_$��|(%���6�"�"M}g��^��!4A!�]�{�YU*tPM�)nY���-��������R�O�SK�P��@d��hV�~���'?|m�`�Q�%����C6�EG�,^Al�樇��n$�r~��4�h��������1�5�\���'�~�=��4�%����LVoWjXp�Z!䅚Fc8��z��}���՛�	�%�2<��m��)�=�L$[nE��z��N!9�瘝����� �
;8�E�{k��ol%����0"# �GϪ��H�����sK�?��ɋ��p�9�7�?j	�7����w���E��4"�abUg����7��_�~(���Z���V�^�)���lA y������Lw;��HM�FK1p�-a^�HukJ��0����C.��J�T	w>�����2?	,��>�E1���_;���9B\ϑ.��F� �8��~:n��^�ď�(�/��J�˒(���\>��\	K�+5��+D�N�\E#�8����\���Z�1�����k�<��y���c[1��3�w��lM�,;L�s4��5���e���|s�\5T���=7�_��t�%b����6�*c9�a��/%���S�aMB��Zl��!�
�]�4H	��~�Q�� �u`��"D�y.�;b�l]�;��зx��s����Ȳ��a�Q=������g�����3FA����Y�1Tٚ�{��O������Gq澟�hqA��<�\���� ,�)ϗ>�J��Ԙ�e➻f�]���X�,9���rK�R�^(N
�T�����Xp�?�{���SG�n�Ux}ಙBƟzޯuY�1�g0R�F0؛��k��3�.3Y�8 �1�87� �>B��2�Ջ]a�G�kJ8���e�/�� ]~�?�q��/�h��^�� �VvQ��n��ט�>�Z�\,=47�:�VA�y_��Q֜#CYя~����8ޫ4ȏ�o��7��a�\5�9�s����g��^Fch���P���UZzA�3,H2�.vyO�#�}~N > @��|�
Pioے���1-i��W+�YMW��"	s�����3����3-C��qP3�o�6|D;�9�uI���K͍�4U{?g5�`�U�ˆ��b;TƐn�+E�\�f��8����(j��������_�����͸ֱ5���;�f�����[��{���i�܅p���L��p���D�Q,�+j��[��ni����؅HӨS�%P��>"�0m��K�v��ąTv�V_4x�I�+p�{vc���1Z�i�Q-m��ԉ�d�(l�C<ZLuDy9�:FǷ�� j��d��/��(��nH��+���1�v��v9�Y�w��J�\�~^�PI�#m�ɔ
2Ύ��jk�K�{��UJqx �,��Bx��ujHs9�ecK�s��&���.vj���'��Q�q�⺒^����/eUR��UX��s:'�Y���T���ب�f0��S���m&�>�%��N����te;��7����J�9"+3T�	���9�g��<T���l!�y=��2yo`��*O��b��(�	ZLy��$�,�u�ˑ&�7�:H���,�6���D��8M�6^G�7��ͣ��%�"����ù��N����Ġ�L�  NBN��5�R$��i��X�ꫝ.�ly����nE�w"{�o&w�;����W ����62?G����yί����D��LdX�A�7��J��$�q0_T�mm����,�1AF�}�ȿ�:2��ޣ���£� h�y��3ұq]�w�r��/�0��ٿ�V%f�G5d)T[��)�)�!F��	��Q�a�F����6�_�q��L�B�w�NkF��b��S/Zg�P�]���0��%�*}� L��rqOvM�)?`�W�;�%s�ڇ�J2��}�Vo�8���\�MM�,��z�c��T؄G����Ƅ�+�X�G/��ۀ�[%�����Q0�g$W��=4hE�zbGwwƿ����#��?�0ϥ��T�#W��)�;�w�=G�?J��j4���7XkYbH��o��ӶE�S&�%c@@4�́�;Hp�8�=mНrl0�@���oܬٓ�g��4\�x���hn*5y�OYq��g6�����Q��ĦI���!����u+"إ�X�k�sp� 7�'"����\����ub��H�lF/ʟC��]^B$�o��V� �_P�@����_DY`���kJ)��*��xbפ�:��S��K�L��ۘٺ;Z!���xc�G����6ԋ�J�݂<��l���'���btq������s� ��l�J��3���bǵmU��C	�e!Dɿ񰦶�w��cE+ a ђ��Ƿ��M�+�
�L�ӧ�M���'��U7��mowh�@C^i�S�t��iC��~0���ڥ�n�Z��!��f#]?�������1ge�q�U�,_��J���B�\�J9����Xm��*�Ju�ꃟ2u�/��?���:9S忯�T����n��Eo��6%�q��w�"�,��g+�om�_ k&�QJ���?b'*�M���@bV�w�@�������߇rU���f8��~}�?��<
ɝ*�� ����C���ٮ��tI�w�@wl�"�����hl�>K��CЫy�\o�����O z��T�M�洨�K�z�����%��&���My̟)3�f$Esyg�F��S�@������BP�Ǖ�<Ou،\�^�4��nɵJǛ��7b��Ov�0�Q/�#�n�dm�qr0d�")��XTB��ד��KIJ��_*)wN.;�K�$�4Qf6p��놟�E���[x}�Uk�xG"�[��D"z��5靫ʁH�o�� ��0=�̦B�A�;��II�{���ד���n�K�u���)GC�
�lrb��b�6��G�3�����~u�&SC}���ե@���ӄ��پg��0u ���]��9�B���՝�HT����.����Pۦ	����]�ᗃ�Z���'�b�A��Lm�t�5V���ѧ��lh�����d�2�=�v	����'e������oz��Cұ`�Zau�#(0���7���a�k,V�J6Ҁ{��__/�o��� P�8���J���3���D��Qb���a�i�Ԡ�p�7N�R�l댧�]Ҿ]��� -��V�����d�c�Dzx��7�_F��NWC%�A6vT󝑫J�p"?��f,ږd�&�%T'l ��� ���'r(�����,\��X��[ .�j�f����E�B [|�B�4g������`�D��:X�-կ�w��ОQ�ş�c.`]��+�I�3��uyvQ�~8�ه���G^bP�{�Xm�ü�hG�G�>u"n���Q��E�]=��(�+2�ܑ0�,���C3��4s��:�e^Eȧ�+V�NQ�Y�4�\j�g[�_s�c]���qٌs�Y���&��Y.����v/o/Ḁ����d�W�VT�}��ZX,��N��U�@D��������PR�U;"E��_�%��7�j$�m�=��h}��V_npA3_���p^�,���Ab��+�~e]����,B��j�X��\o�Q�$Kd���<A3C�^	u��A�b��i���@r���wb�;�x���8�o����^��6`�խ�#�]��#�p��-\�$Ol6�8ETK�KB�_���OԻ����^��e�=]�(�_���E����ŉC���mh\���`���.������v+�W]ӓ�]
Z,��H�Ƕ�@�l��� X�6��tP����X��9��M�M�j�0��ܸ�ғo�Z�}B@�~� ���i��	�7��H���vlN���Q��۸H�!ŮS�WY���壽^�i����t�JL��}˾�S��93����S���ՠSq�릈��@z>��i�:>d4��I�\PAx�������tl��2k�^J������@m��g�D`ndjԼF��'�W���k�e��x��$W_�ձ�e͇Dk9H�	��5���q�nwU�oTr�
��زU=�e$GD"}#lOW�V%�����E�bЌc�!mՊ�?͡I ��P�kKkR
�%��b�ɏ��z�,�Y�����x28f~�)[�eX6D�R�7�M�h@ȫ(�H Y$�\@q��"��z:"K���?���l	��|NA��B���xT3��噯��}'�
?;<�������ˮ;�K��d�8Zbvw��H~�M�ɓ�p���+��R��7�*c}a|��ݹ�X�8�e��޸���!U1n����20;��p�u)g�  ;�������r$����U�e���n��������n_�6�0�W��}T�!�L؟��Hn����GF�g���3]��y�P��.����X��jݏ�7���W)���j�1����*�Rb��=�E���`b��7�W-o����E�<����&6{�C�����/���sY���c<C\yzS���������]ظDX�n��n�k�g��tT9P=�<_[��}��������<,��<�Klɻ祇���8vmH���x���C�NYN&�ō�� �n�v��@��OIߡ+:���*�`��ɞn�6�w)����>3*6xwD�K*�ֿo( �g.���w&�l���z�f"�F�J+,5��Ӌ�t&Q����H�����+�|E���-Ca2�1m�~|4�iR7�-��&�Ϭ\P��Y(��1̽'P3�@��ru�}V����-m�|�w;��ʗ��R����&".$X὿�FC4����h�X�C�Ď/�~S�����n2.�d��O�r���OXq��F5��oni�)���#��Nȭ�Ǉ����o�gI���J�3^�E����aܾ1*Nj���G�PJ^��M)䴑`*���{����y&�K�xt%���+�׋fe3��{q�Z��G��y����*�^`�OB��(��!�+����+E���ˁ'�.$�^�j%�;�C8Wޑ�ЦT��(�1���@7�]�j-#?]�,~��u�a��Nh�imϞ����JE>L�E�b�TJ���W����W�LT�?.	4�kkc[	���&�UG�v��}!É�bT��?�-?������9U�f2�}U�&�>��	�U��mg�s�U���1I�����R���i��%��c!�m%&�U�ܻ�����8fG`Ѝ��x6r���Ey�����G�K��߈���i���z�V�Xb&���͑�*;���O$ަ��P�v-�a��6� �����yZ�[��4�y@��f����x^3�P���o�sR���:A����V�W��t"�R����Y��3c&����G��h��H��E�u�{����O���|�<zL6xK��\n�&h1�_�f��q"�;C��.��Cr�i"�t1�xf��#"��!�\'[[ݖZ�Tˍ�C��R��v��Z�?P�DPjIl��a���L����= ���?yq�����@2`^K{���w��	-�)Z;|H  e?��>(�^-��hŷK ���]4��嫮u�LF���U�ߖ5��ǁ�B+�gWQ*��A�T��Ұ
�j-�{��O�����7�:[�Nv��,��H,���`�٣����̰�S-/c�T�M��v�"?�� �m�����ٴF7O����~�f�a��T �Ѓ�`	�ŋ6}j�����aXn:�y!d���H��d�~���Զz��ὴ�q�l��=���g��!�74��>Lt��q�5�"�osq���sw��A���i�g�r���g�*��$պ��~�.�r�p�_3�����C��5�i"��X��;���f��w���F#�k���>�(О6N
���G�5��?5E�Pk:�/�o����!v�
�ԢyΧ���U����jo���`�����o�80F�܌��_��W�;��N[{t����tv�Ϛ�c���mM��i�4 �:e���(nq��X�.L�R��T6�Q�d^���/R��
8~rr��e$N�\�<n�R �a�k����սmE`��$K���UGa��>Vr��T֥�9cQq�@5��΃��3���I<��K7����]	x�����?���Uh���NaPӀ ����a��j�=��a=�[�$%[Q����^�M9���Lki�`+��\#���@�Z��Qz?#��b�(��[�Ş����\��3s+V:K-绹�"SGH���(@
~{Tz@2����E�Ԇ��8�Z�����p�RGG�j�������x��IL5�;-0s���Eځ���@���X�5�E+䈍�0L���L��%49�E�H���=-��G�~��+�_�h�
_� {���e��%|#�F��)�:;���,�;��ȓ�Z������m�z��%7�+�E�����r��[+oI�q���4�b����8Kج��^}�����oH�5��E�0�ֳ$���x���)\`=�涎�c��ӳ3�j�EvF%[�v
	0�q(3�n�p{��~��e�L����8�8|����F�K�4��I����kМ���k��=���x�;�_D��ܬ.t�*vN-�P��M����4�M�"~�X�b�� j�E_�V�ߒFy�[d��V ���`�[��h�����o�1�,ʀ4�7���|pU`>�*xiP�͡�c�1��`�X��E3�j�Z�����>��?���:�7ǿ���j�����/��4���o>�.\!�gE��[�<�h��6˞*{{Ai�`x��|h��\��LmC����-�g*_Q_� �Vy��64��Ew �r��R4��,���FG'��b�fwv!R@ג���kF��#�*� 0?�$� F|A�;o��HT�mਊiy�A���!Z�xZ"����;*<j?����	�(��>᭰m���~I/��?��O��TŲ��-��8!ń��mcF�B��#ܦ��b��p��#�Xܤ�'���nb�/v�Kϸ���|���ĺ{���/��3�?��I�Q#��\��Y3���p�#����D9Ӕ������X�}Ar&+i֭	nBL
�;��Y-����3Arٸ=u �t޺&�EĀ�佒���WA�ʏ���\M$�����0�ÜK������w���xG}��QT��c�UNm���d�~�Mj�,4�'��D}H�hf���\;�6ЈҀ�^J��'*�b J�H>�IHu*DB'|[i�����"
\P}�O���o�f�ƞ�*�n��wSIM�!u_��۩�(/'Z��l��O�J<N �ϯT��]D���r[�F��c�VU�WdO�: K	�DH9����G"��ɂa�&���}8�d��L��{a��X��O���1�E��=k�5� wDG��%��	aVH�����un��	���m�#��� �Eo�7�~�����0>�=�u
�_��!��J���@q "Al�p+z��s1a���L=�!�PG�[���2�@w�&.�&ij5g`{~�4)�t;{.�l1W>�
��J�\ёH��(���0���ن�p���?��kO��C�dzE��_��]��z�ʈQ��?�= _�#L!�A.e�_�G���j�oZ��hZ��n�G�u"13O,U?L���\��u�U�����ոCb=PP�d:63����6�^�*q�9Erv-SvB���y)�)�w�`���H�8i��rUp'��>?!wG	���Ȟ�&If�q�_��/L:��ƽ|��Z(`��p�������q_�wr�l��� �!])����oO��ֽg-D��4���V�ߴ���՘�g�Ţf�l�G���	Y�I%FE<�e�/��s@�� �ƬI��#�N��<�⥚�@S���H(�E��g@��j�����X(?�	�^�;����@�a���`<86� ƣ?���\��L�iE
J�k~Q�^"p�[�S7ȤD�S��u+�Pg|H�@���Ә�#g�Nq���	�_s���ˢ�q�����z�ӕ���vk��K�>N?�x�o�/�t!k�J�o�B�H��oE��_�����}�b�-UA^�U�"����˵D���&�9iEZU�m`J�r]�Ty�7�X��~��2/;�U�)�����jԔ��bDs<i�S���;UK����ds��Y�ޓ�3�_C�6.��"��)O�]k��RZ��d�a>��U��L��>i��\���^��S(܍���7 Ih��6ŋ}�h�=A�-��3+�g$�����[&�T��\��}%�:��z��p;���
�-0��e:��sQ��U��ս~N����q�:8ì�R�ӈ��Q���!�L|��g�0�z��7�v$�__b�	{�+��xE���^%9�ܩ�����=.��V���%�C���u�	⊈��ÃN_� �� MV�07bU�Љ��e����!�hbp
�K����>�����Z4�\���q���/��p�����\2�l�t����G��c��rU[P�:�8<]�?����R�����uI9�&x�#KO�Mh�㢦W�_�/�(�'s9��.*r��J��P"�y},��v����|D_C@��S%o&��H���`�	��a��&u��Jk6E�1`]	��=�-��D9�)8�B\�d�ǬF�N�F�'a:=��t-�o�I��:����Lh��.>Z]kͼ��%����[W7��yK��7vk��3���Lʰ�� ���xYs�z�xc�D�
m�+j�,Μ�RhOb�
�)/ з��W�90����[s&�t�t������&"W�,j
\M:+��I?u��T���Zq�:�J��DY���2�S�B=�z�GJ1k6�� +iˋ�a 	��V[����B�����������f��;�j��<�2K.�a\�4�Vj�"��<O~ͩ{4`����a��WW��f~�Ρ�U��f��(�)s�vt�\��F{�v~c��˨A�P1�dL�i��j,�Jy���Y޸�Zo�/�	*xi&�.�| ���� @G)�^�{\�tܥY
G�+^����ص��r�<L���v澓���%�k��1Y۵dm���M�}OҲ֧���p���q�W2b^'�1����义�f��j,Q&�򜶷!���q&^Kx�Po���m!����.�&R�KMy8�Q��8�P��>�d�B&�- V&�Ue��G_���X��[BgG�J!�e�\��߀�Z�a�K,Aޥy�41v�k��A��wʧ��f�MP��Q��b�I�q�>W���B]�Y�hXn�158Ȩ�T!��Y�q�g�@�M�R�6V�Y��'��3������:P0µ��|E��$�J`	.xx@!��t�B��K�KKP��Lj&V��
�J�ԅ�<t��8JJ}�K9���MS�����%t=��&�K�,���_�f3U	��ǚ0�/'(cU�;0Ԩ�o��v<d�D�&#tF�U��;U���E^�y�|��\���� m�[�R��[a��+^E�~i�`���aK���~Hp�B��]�?�������.a><!�'$C�y�.�d�n���A��NDǸˆ�y�IN�#�2,F��$$4�qoi&o0�A������Z@0�)�KW�����
/g ����1)��6'<��mXmJ�y��Ng*��\��Lq�լ�:+NH��r�Ƥ���&����2�]�J��p��lX�	ʙ��m�e��A����� =����̈́�
f�>���"yy����!��fIy�?�y�ې!d��-�Q��U��(F������u��K���2/��9|K#?X�vdI��0��ƣ �Ȩ�P��,�����Je/NxF��2����H~0���2W��[;~T��r6��c�B��i��
x�W}�s���!C؏�Y����僕�M�J�z��6 u�8244x�:���А�/�J��޽��d̾� �Lb]�$pNk�A�J4O����D%���"������
ͫ6��P��1*���A� _pT;2��@1B�����x����'{\�
5�
� �"�߉���+���+T����샑��]���0$h9!*�0��K4m��,_W�J���%��䡆/��_X�WJg5���;����X�g�h�`��_�y���*$7��8U?���/�E�|�+��@9(�&6t�:�{� gN�{-r���/�A���w X>�p�ͧʤ�	�T,����?���,7��x۟�C�ӳR8ON�<B�x3�K�U�[!\�������R!��A�3��B��Q��l��m�Q�O�$�e T#,^Y��/�s5�`�����p���F "����֜+y܆8�%��MF�%���E�s�/�S�U�7*�)����50IV�=I)��>���LeJ�
�%��0�^�7'�6F�2gfޭ��KY�<��O0߆
��"M��$�n�(�_�YGTc�ӴI�qs)�y��\�w�px��B��!y�B����N8"�M�l3��EC�J��l�'���.)��c|+-p��*�g��E*ZU��C���Fh�˔��߷j|�bN���FQ�K�u.��8V�n?�����p4�YC/���l_�ʇw+���v�!����Y� :?�%=�G����L9ю99�i[E�u���!�&d�$��)l����_��x*<�����4�*��R-ͧ섖�^��1L�� ������D�g��#Ǘk����|L�NY��x ƽ'F
Ƿ{C}aL�z&��ɾ���v�e$�1�O:�ҩU'�Hs�;
�F�y5��˶,Z���fi���n,Q	k��%X���=�a����x��RffP6΀�׏���s9:	�]W�e�V޲n�6R%����*O��GQ>�9�tq�e}��;=��\V�X��fs�3a�ٻ谫��	��v�9@����@�{]���Nz%:mt��{��0���De:Z�@g1�b��3�=�o�<�Wݥ_�pCQ.�z�͇��{_���K)��QyW�⩱���,��f��|��j�;z��uz�|���� A?�80q�\��\�_��rZ�﹁tQ`T��/<�hέν��Z�&�$�����?y�^��ӹT{<��3�J�i�o܇_Q�6C�b�n�qe������@�����C�L;�X���>�Xд!ȸ
����/��*��wz�?�籱|U[�eYX�_}��CpZ�y`V���]ĉ����f4�$.uWr��j�W4�I�,cK�?|��1{qbz��L�����M��n �&�݉e�W��K�᠌i[x!k=�J���{��5M|hl�"��R��}�������/d�����"��zQ����:���`SR���OwM�� �Ħ�N1Ĥ^��9����mF���:�Жg��XAӫ�)�b%NEݩ#qb���<ޞĠ+DM�[[���,���8���Z)s4���ê�	��u���]	�s��=0�(��jr��ވ�k��%�P�8$�̓��b��.�cJ���A�{������?t�)~BEtQ^�w��k���㟽���Ao8JTM�Z����-՜f�E���7z�9}E��x�~����,�R�-.}ȍ�=�9��n{g�7�2���Ѷ�ֺ��+�����_�8t:(:� |�����cs)Qy����S� �?b��|WbN�l��5j��:*'9\m�ݖ��������٦��e{�:�im��H
]|�3y��u�&�IƑ���_��1{Z|b e�������õ�4,���Q�Z*W��܌G�|\�e;��8�ho�p�fe����9��RA;�y2�k1�����슮�E��#�t��k�]$I4�{1��u��+뺖��R���+yh�z]�S��a��*� ��/�?���t�n�rp�R�xr}���`�F�|�¨)��E���T,�f�J��V�&_G���9��Pݛ����
�#���k�v��,z����E%s�p(2,$��b�\��n���"�Pq2:�`�yEִx��k��r% �X!dk���j~͗hۙ��:��$P�����=��eY��N��&���G{�to��L��
 ����yGR]b;�:j��l��eY�z�����ᛈ-�lR��wy7du�45)AM<mh��;��C�];��a2�}Շ��xL��~ �ϢY��?������5�c�I��� ���RڇlA4E��hW�0i�$p=�A�l;��)�U��f�2�e+�r�*���S��I��|���6h���N�R�l�=�QB����Tгg���o��Τ��ȕ-����U(/���YK��o����:{��P$>�̝N¡5�8
tw�W�x�E�"��<��s���O�o�b��c��N1J���G�w�f2���f�9���e �QSia#��Pw%.��y����E�W߼�+����@>�b�cuDҿ/�@gd�!*j����Pq��I�?2"Z�TcW�d�~�pY�(Vo��2�]��%/�TO|��}F����X��~�b�%Æֆԓ�ʭ�i�jz\-�}������t�z�N�.��_�_�u�t+�Uuj�u�֣�- �O����;��v6G�p����@���O�N��e8 <�v~C�m�
8�D����'�:�czh W�__�_F{�9����r��i/�`h���r��lFJvZq�!��}���T��������r)�J��u�`�����˷�h�q_a���҄2i�0�v�(�/�����.�~vaԑ���#U4L�c�|� ����K�
k��.=�*���?�����sr;h[�~�F3]zEMp�k*�3�澰���g焉��
q�����Jx���l��w(Bx�ډ�|~&{B������%�������Ҙv����,�" �g_L�l�gBP+��^���H��q����d��Ay�ʿlp��ue�|E�����Q�}�L�Wd�<�Y��FN�.XO ���\�4W�%d��2H&�hD�hCju�}���(������O ��{�5��&��@�/��[�{Q��aH�cQ�J&ϟ��p�=Sf�����eq���>�yQ���J�~�=/�?ҝ��%��lg����֗WJ�cg�ߥ��v	9�;r`}��w�f7z��#�t�!2k�(��"Z�� h�(�S��S�tbC��g>J�>�=�`D�I�H0>wD�pVm �}C��=����9��� ���#N:y�)� "�`�JB�@�<�ƑE�M�' ]w�	c`��]�:L��-� ��}�t����=��돧�觻(q�s��7��#������Y����3PEI?���M�t��h�x�-�k�{ƽ�E.�����KC�Wp?�����,kY��rPc��*.(���tϐ<���$����>�c"ƽi}E󓅬X_���_h��q��D�{�i�ĕ,Ԛ'\	Ě�ٳ<���P����ծ����rc5��+�Ǥ,�r����Ԁ�K�:�nߴɁ��D���k�Pa��ѝ΋Ĵz��h;Ҩ�;�bgw����h���#���V�[LSs:��n8�|b���kx��ZY�I����gJ�@���J:#sa`3q����̨���p�Y71{����1*���M�E�O�I\e�Օ̞H� !4���,��A�H�n��=��|��T������n���U�J���pB3�cI�\'=�P��������i�>�eFm=��
8/o7�Kl��5������ޖե�&�cK��(
@^3{�i����WS��_�$��Ƿ����)ĭ�\�t�G4L%��[/�h����:��9	Pb�5�P��?��esrC4D^��� �X�?3F�W�����G^��h�w�$�]/P���J�_2�h�qT�Su�q�=�z��}=�����5C��&+˕��.~$�A��:|$�`���dg�( !ˑ-��@@�����M ��ʟW�g�&��3�� uܹ'�`sĈCɨ�;��:h
�:Kɿ&��3�4��:��~��S.�ͧ��,N�Ы6E�6?�,&�C��?�ՠ��O���_�'���y�=&��F=s�Y�����`a��^;��"���� ���Oڪ,������P���q�P��ּ��X���Cf|��k���|k�^4y�ϵ�;��`��͚ ߐ�ǟ��I�v$���	k�AgAy��*��K}�L��g�_�ɇH$� ��r����4��M��@��Fp��i�6�$=s��S�i�v"r1iKT�����$R�@���:R��1�E`�x�馮�V�bgfU�-xu!`�O���^�R�A[>}�pRf��̭�6˘zd>�<
n<*��Q�±Xz�
�B*K.W�	2)wv�����,GjvܝtM;�)��N�2
��u�,*���櫯R���K8�_ͬ]���7�x)ˈÓȔ̞����pцh��Ou9�����#��:ÄkO�8p������
ɸ��e�dE�%�Ӵ|�0R�(�;���A�.)s���#�~��w�0A�q�o�-x�q��@�t����U,�>����$�?�$6�+7X�Vx̀�µ�^�{�, �57;�SW^�����)YR �6�Q�)��a�hJ�)��w�b
g���:��>�!t� ;�Suؽh�moy���u%�$�p�O8��m�Ը4j�zwIUW�(��W�[��=zD�}9KE*H:>qP#���&�~< m��Dm!�_�c�pN���[�(�K���9�ue9������c�c2���nxKb	L�2qk��l?�m/�$����O�-��J�T����̋�����l��b?h�%)�z4�p�B��DAOWT�;#�g0��c�~��/.7O��Q��r�����s�;5Ծ�x�B$/�ʘ�?����/�o��}Y�tE��"� "\ @H~����Pה߭�&:3��;����;6EL��,���x�I�$:�t��&�;�-�0���k�����֋�:�
	�,N�o��7�M]'��f(����J��%��Gӯ42*�W���h͍���Vq=iVF�O����)bv>7�By���)����n9��n���H�TcC�w��a�4�������	"^�Y&����v1/�N���>���{��r-��R�5��Av������YG�he��,��a,�:k'ē|�T)AĲ�/��#�O�迮���_NN�}��hC�GH+��XTMK���aB�&Tp�s�W�reA�-���y���@�qnf��f��]y������fO�� ���)[3Nn�<=�o�iwR�z<8�����R<��>�#�v��3�c�� �ҸDC�g��^6��9̊:|�3s ��c�H[��m�^]�U-����; �V���;�µ�Y�J�+����\�W��
���䠈;&܌�-�o}U��B:	�O!g���^�u9CH�r�`��{�2���5#���Ο�����O�HjSoܩM�p�O�{ĵb�W�jz39Tv��MU~�GW��,悗	�5w��`�@E���ii7����MZ�wx���"�0Wz���SX:M���"�/�0�e��B�|���q ��^��e�l�_nd��ki�_� ��D
?� �
�M:�\O��Z�\46&���"�q��}S�l�G)ί!D��˄� A��h��q���\�� 0 �ܣ���,�e�yq�
��V�!6,�m^��u��TK����oHk:���E���	��%	���C�Y���߅{ډ��hl���bYxl��I�Gn���i�~�&���Y��\RE��.�}��|��@t��vB��`d��d�i�R���
�,���P+1F���q��mp(�w�1 ����@x� >o�dn������uq%z��W��Pm�_i),N���[���^��f�v������"Q(~���]54�9q
�d��L1P0���yX��~H=�mS�Ma��|��R�v��q���H�_�}���L����:g$(_Ґ�����q���6=��y�Z?�L/<X~g�e?�^G%��ӟɲJ-�� l�:?]����{������ҙ�R�k�p���L��BC?��#�m���p��Ky3���Mp����>