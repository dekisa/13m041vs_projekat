// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
zuy4NUPyg5f2ej9S8/ihqcHXWTnxaBbE5ZjN4wVQFeKnKrErfala7CgYLwS+8FaGcnpeKdTYT4XI
EIGNM3d9uHW4uYLkoBCA/jsvzlCDllvcXAKT6m1LzgZcWb3B7yVEmC5lYQgNSJ0PBaDfjLC9s9k7
OEY8+JvRvTpG4bu8whHvRh/wpu3WCBwqUXls6+pH4+9bD9isVK1Y2ZoQ9y0zhKp0HBSoDO+RWP/K
84lNbh+oHjIqmNsKD9GGnNa+b7FRdRX14Xa41dbmintzDizLe7R3DWih95dfzQBD64ryo/GxAF4v
CCwe5S5/J/G6a7/KnFbgajRYJEAFuax9JAqedQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 110480)
IWL4KQownOc/b42SErQfv2RfKrY5SAuMVNdvw2Lg5LQUaeCINn9HhGQ16NbKgJKdflN1LgmUtSVV
MVZ4l91JEPAK8kUmDyCWZKNg5fdR2PsDq216f51GlCHdzUYoFKtMGHDfZ2gfH0LccHhHGhWzzi+C
kjaFsca2zGzC1ppVNpVUpoomCGOYmPod7P4xNeXdzXAaCaDzY0Km+46B6vqCB90HB6csePgRhrzd
dpHbOLqi2OOwFHeVRA93hcO03LbKD2skGd/SpvtEUtIiE951d7SR1VOXHXKdr4PKo8CFDLiNzLNH
X0jsCGvRI09CSZj0MKtLbVBM9If2iniZEYp67fT0Q8lYJeONv9thc7IN8PYFXmlbXmPujRRwGrVk
140aEYAyNDh3UqZes/dtG7/wmkoUl3dHCpMRkEWmeMssx0cVrLzA5rJxNQNl0l+0O8DRgwLrFbDB
bHy3UXAtvJeMdL5NtRsJUMq2GVzalcubzspyXX9rm5+OgzkbR/yaKHhSbvXTmQqeAr7G8aiEPRQ3
V5hpSLOqOaW+A5w23eyFJ0uAj3h2a9fOEN/g8Z6RXFIVL36M1dg6zsvHveBBqGHdMbrp5FX53a7M
tj2uJPZymGPh5mTnI5YantOGzU9ggFTzCQgVaTGSALzf+rhIROGAyBfwXnl2S1wCyDTx4qGOrrJK
/93p7K89wxVvMTh64U9QLa9xFs9w4g7oIdh7pa3kll11+8wrEMokGxSfET02QHFNKX58P11sQYvp
B7A6/Vz7gSD4tS2UwO+AI0SUWrIaEJmUxRY8f08CKWLXen0LeVh3s0fd36ztMqpkH2y3K8dZ0P7d
yv7cLOPwXKMvQCszlRf7XSoyR2anPT1Uql6vNv7LlwiV1enfAsiATDDchR3TRNj1SiFTaHuoScDs
YvMlkMKmYY7BMywL3u7uRulv+i2A+DYgFZjgxKf+PP/2lhfK3KwCqqxYrE6oXzVD2mKkf3hBvRs/
Z4Vc4yEA7N30VwG0BsPNO0AXIztcnw6MeRonkUEBGetzBZ3Wh7d6immvRQxp3VxSLrsvZ1xsjE5B
fiSP6xJj3vIvp4JLQ2AlaUC+p/u9sMF0lYrLVN8QEzoC/QToPLO2Cs7xfs77X61Deak071/X4wL4
REOYxdTsEZwxSWjSiuahgXs/kfBAm6H0TSf4ccnQdahqmML9dNnI7hEGX264CdKussoZT41/nfo+
04/8ZqpIzR5UkBnz7xqqcW+IyWBaVf/BOTCwZ2wNkamzHqM6ad1SvzRctdQ1WaRHGdDPU5P9/seq
Oa9X0Fhe5uGFAZEsdK8uaWHZozVrkcHP0P/Gu4lPLjcrzhP/p+LE1fnUFnBVwi+XkYXyTyNq4+m6
FkT7GKKsLYmz9QPRCLB7NHixu8D5Zu5tbCRluoJ73o7JuuntNI8KKbRY5MKqsF+qBsqqcSQy12jW
0U9mEgN5v6AgEjEzp0yOw8wfjy1VAhO7bGko8zzov36WPPQeugyNPhIcBZAXDzO+m939LiiWfpj9
BUbAnvleKWRnj9MKsLsBbnmzmfUdabjvR1iDTKNu8wfF4T4Lz4oWvVOyLV1cNv5WxfOyNTgQkZi6
zqNXgPYGXAhaFMk54Z92X46zugj3beBHR/JmWH/JiZme8FThn4so3kvKkw+iiPNQ7qFqDQu1FNV7
jKr5wN3uNuHF9uKmyl9y3Bvx/YaUWWy1pVlhFRUisdMCy3NvKHJpTA70CpdFn1dOmwfmgOSa/+gO
G3Kwl6csz4FiJDaDUGcllKls69OIL8HHJP4JmS2lwkVATCpRDqyQ0rMKgIcItWTOKY0b9tpiLvS8
PSNYtcgY3LlIiTdfBjO+oetLSlbU2f19IhYbjq4THUZnBFuPMFW99waN7LUxCp8HQVmygaP3k1/X
gHLC1LPoxmjiDmZ8dmdKnTdWTIfrj6GdODqNg9shviWP3SZjpHdCleZPMRkra5yvEav/ZJ76ZZwb
Wf4U54BAXu193sVnOGII6LKhhLe8RYS12GyGiUdvN93lmSjJVKia7x6BH+T5X/TFH06Rjv+WdOis
8OjhcbxkO6Hfj89H+U144tSODfUaq2Ih0zFC64tM3YD6zU4c03OAvR+OSIccmzLEUTXRGvnEloS/
GUdtAlkW+VHDJSiyt9DDb6iqLxqxx5iUWgIY35/6mRHqI7bYx7/M0lfdgvo/VYd1Rqlf8v8yZPR0
DKYw/FxxrtigV+3VGoWJquseFNbD82tnie3VuaDEXqk7ZwPFLlgDiXWnC9a65BWLC/MG6dYU1zoR
eFNn+2lcRxupqXRlUmeHfaVlzvQO5BDYNNZQ9HRqsvDJNkVETnxe3QY/lnujwFgiM1zXCwRIXh7N
jn3jv3CACVdgJdlkM3DMLYuSgor11jh8/Ci/iJ3Y3Kt8dU5jddZPMuJ9m906Jbnn7eGTO5i1GmF9
krVBzFxm7sr/42/AuvhgOZvRgE0dYBl2SkOkc1qTN7EpqL2OXa+gY2sN6ygf6g2/LStJIR9d3T9G
7AlXb7nhws7x36+9c7u9FhaWVGcoWZJqtn/meURq2Mcxu6aT/kr805lUJCFhJRsZesNqF1mm4Lv1
tghYxG0p7NE+0QE5T+ZhfXniRpU6HPumwiRAB0QVZ3OR1jVbXil8yVdve8+23hPAnNgCRKzkvU9J
jqVs5acfCAjzhnHAQezwAA6e0mXmJMi6hOvbghyjZDMEMW4UJ6gqnr6oAWoulJtUPLdUIYB71Jez
PkHXu0PwN56YeW4ZZ3W4x/eq/cJoL6QGdEolDEu5MZKBgBV0itZuojwRmy/dQSriicjS/7HZQ3dE
XaQWD6VfQIx1JS4e/HVgmaMZnP/nQqrO4KjJjHyj/NAKKwhZiRj9es9oJDexb2KshSdya5TsduzW
40J9Y0cuJO1iL7tShi3BCUlhpIV6ol8Y78sU2vwjvkrWzUjoPjH+OrZm4ZVEAo7XA4JfjewXnhVt
dyehxrCFpxgN16j6C2z4BRHMZgZuPJe99D3FKLdRXIhUaAuNUZjpI9VV7Q5j1iq6HXzImk3T7WpM
kWyQhEUulYCjlA9zJq/Dig57cIWdhGfdbbxU8BLb/rDPeAggsoJrIqn4XGZwRkQMx4XeCFnzQKM0
XC3cepCQ5iBpF3YXsQAYZV3q+olFrdZ1p7L7VPrbfC3+LY8IveY+XUHX/PQNQ5sI2lrd3QAokpjK
KgrCZsX9dmm33rgWhfSTKO1A1d/BT62lo3/akCTIEyMldD1LIJ/A+GOqxgm8gJ5x37HmWJWOgdR3
MzERfCBKJ45QgBZnXQ1S6bAo8VlOdmWw5xUHyrb9ayketzb049pxsfPHxw4z9EUjO6jq9Xmfy6HH
lyHVaAk/WGYTAKwrkBc81STqzBGnfII6uzFT92cxZGG3Dx7xivUXIMKQgDbb+QdK3cbhFvYUuF77
gqSMeqR1ff9czjYDu99WbbC29RfbS0Uro+xoJFKkds9xCa+rHiwnv9XZNr1QYPaEmNEYUIVeJs9W
br08e+mcCG0E6r4Gw9GW+HxZCeK0f/4uvSOo0eJSGlK4E3m1y+SEyL56LOjoRVTuUgb4Sd+akqaz
a5N/YDsVW+zvu7PCl3F5TJLrL6XWwTpeZD5yxZGBy7lk3FEuPh0Aozf7FuNFMicwK5bCwN1idpkV
Q8XDfpGYdfK/f0WwbvcVw/xEPh3ZoZH78hv3Lb4FDNXj4dYzOIT1ucEI7xDSxEhGQHSFS3e7gYp6
KSwfsOW2hMfP9g7R0FWE5Y/0gFa+3Ovy4oDWxnQWIq+lFs1KBx8MO2jmwNHJfaGUYeGckWha344h
9zqKx7uR+ypzvJsvMoHTAdhxqR+XopiLR1eDKHZlxHsyZs7hvR2pi5003YmdRFOsVtNgWQacbylz
j3ameqRzKP2aVQBB/HUlns7Vc6gfsETRi3Q5NFLBLrdllT6YlBSAD6+aYlov+JfUUoWUFWlx+ecn
Cvt2riZNhNjlZ1tAdRMDMlKxb7BShLC3r3aM4ejTMAWqtaXPNoR1Ynj4NYO2YcXjkgJBU5NUXmkU
mWoYBSNVL9TLQCFN8PhSak0wsjt5qzOWcZFANfeHl905Ti5pANzztr2pLSVKiBfUfqzAHMqeFSEL
iyfl6VK0OsGv7I4MjxopL4wtXDMalKv414uMhao1TmgsXdSoOlkL3EAG6/6HRBrTmOFvL4Jo6NOF
twMv/1TG9q4IholIo8uVC0Z8lPt/3vXzjj7UXOi6onPQRsxLLGbDqQ2sV6m5tdbgyiqwPqz0zOA4
P3CTYvyB39NAHeVFsHUcAJjF71h8KmxTCf+nBFuVwJgmJZaBTxg86AGnONWhHQ9ZpxBT5wl37Tf7
qKwoxnSlIamsO4D5otILdSsKVU6lf61AAfr6hNM+VmWRIcdRK8opVkwbWVASrOLOgzhGp9ydmPxV
zRaWF+2yfFhvzH1khOxL0RKFN2y8zmtOsQjQSzW3lVxhGNbQ/USe65hpzMsrKTtLYxHRFlFZTtH5
dNsiCrgRmldTUMpy7oV5kLY6tv2f7lEsAYcsJpNEppdPEXrGa7u8B3/zXZawixeQ8kFeRHCH3LjK
DE32hDMaoC4OP8/Y0ry0HY4r/t0oKcOqdYjMRk07XAmakZkyqw84WYGJrDEVDSrwxC+dq21yEx8b
cxHQG2uuoHDQ/iw9x3FbieumuaiLlVu2yVgYIRVmY4UmiheKsgo8PVX7HZflTKmu+6NJZ9ByCv9K
Dht9K7g4aO7g9Yb9wZm4DmwpzY2ui7uQx/bexUccKm0MadI09C35GQAhBBsfAUx0/7suXHIXWREe
fb4x/Ql4a8vsRZGRxGujKs7UrNBGQT7Cy67/YIqX9KHuZf8Wd9fp0PDyBy7PocB7I5uvwiCeEnbz
oriOEI7Ej8OisvuYXzpmhytlTawrrVEk2cuc2OBquzaHvKkz4Qo7gS8TfHFQdJF5arcBXTGzT44h
l40P/ct6d1ExmhVdNKyHHw69zEKKsU+rrSiGNbDL1gbQH+o8WXC/RHpOFGjeUn1Q4rJewIBHJO2O
vR6FJXgPahTSOXZJcbinsswoujCeoG04mVGDzU6lwPI5QvZnOirplKtpUyt0q/JsZjqJ6GWB6NtA
zMmmgQ+bm5kgEPGzd2lcoUqRg7r2y99zAYX4Obk7BRaAFnJ2yFyqRpjkDhYGLIqUfLPToCeFmpkE
x4O8AJ85V8TaZXpMjoPI+BdQWPPC6kPZ4ksNMtraWCZbEIEETHEeorSz76L+XLRdtOyF+HWMuRi8
8B8cmo9dWn02iizctKyM6qJ2V+Gg2kfok8AXgKj/qEidgz1D+GE1gUfVJr+prIcgTYd//FRlpR5U
fwMpDNIocs6V9jheHYkEbpPKdVDaXXT0zLvnEP7SbstlYpEtwqEFhZIWAVx0vHVPQIltMUtdt8MM
TsWyM+isY0tosw+Q0QfYwkJr2K5O/yF7STp/9cEEKr5v0V9deK32Q/bVzHqmlEGySXBr09qHxHlm
8KY2JDMEWoxBbnOMrH0eFR8qWOYJakDSucaYLYdZ6puhF9o/OQKg+8yV1dknLP2waZgfgAtELwWa
jLJkv4aqvKh0Ijv0uZFv/SGL6PvgoV9FZuLwxH4U1/n7mQMGhTbkRhLNXPe+DKxKkVf1VbuHqhri
qxT3yo66MwyjkzG90V3DjTPml/3xP1Z03CrV9Q5vcLSPUk8sqEU3ujDCkkFA7/sj1nlOYOkHutvG
YpnQoy4+ef3hQTyEipO+G4s4ANYbx23kFbeTHJ8KX8w+n8QYfOA26IyXdjXlBiwS+tUkOXc/l0Px
53/h5U155LUwInsYXbTXNOBmqQ/UGg3YNd1b9kq/jwlW/rQY3J9JqaGdchRxQ20It8EwGi6VhkD2
Th5KMZEiVUvQTEhVJGGwIlSbAF1F7jQclIo7NaFE4H0zoDg7XsG3xRcY2ekAeIt1g3dSJ9OvBQdZ
+2gi0X/u+Ppivj29g2gJrGso4apD8tGC7CeFVBKecgKzv/g0T+xPXH9r7qxNXKRYGYaOACs3S0ib
kzTb0PBwy6IPRV47EueL/MHJ9BOf1kgXXUSGnzws3TOoZ5Eji9BZA/NQoacujAKr+J7wOQguR2vM
JxHdGM8V6DgbfRJCRqo5ic8Tnu0W80ZfHLpOI6eOnjHPCNdrtglhEncjVdC/ym5XnJwHLwdALI5Q
v68qJEi3v6EEViaXWgTiMjXenKh6L3ILnYfDHaxmP8oDJ5Wlfd5P1Q18aij/bqWOfYlwINUf4TGk
AFIJwMR5Vq0mAbYIEKViJzNCBgMz8C+rI1spDN4K96doa6dAmFAOBZn/KZQ7WvFXhS7d7q5w3IVg
fJgevXLRK1FY/+6JXR4KWdXTX2rK+NGudLxxWCqb5TtxS0GsTXcEXqlv0yyno1eAIugxYy9+owhL
/3daZOtCRR6NNgLDH22hcD832kqVAY6a72BdeC85v/K4UY8XgnRv7GpXJMmlDgSbbNbtt6f0hI+3
TTfioNQiGDXsxj3JiET7jrAiJefyegAegTFG0KjLuQ++iRNmerKWSuWrInjS9HTO+p0V6ITAWg0i
kIihqWKcQq0lSouabG4SZaiTDWwyUmnMv7OMg84CsiDoBqR1KRf/S/6Ez9blDUcjpC/zN3+hWmEO
KmUSIQ8L6hhM2ysKHdx9m8w48yZvC2OEfbGuRbV8HZQkW9tQgtp4D9+xBXK1evOhfXvpDJnnwpK9
l8efZi/lxfLCsfcnKqZIbogWvnrZJpBe7ywaLOhbOdZI9+dzYzs4vDlnfPHSWHYwN66p3a+8lwxy
9aMJwHRjdqVTWxUzk13fkeJFa1toyfgQJ4aDkpnffFZ0AOd/ZV399JlH5zZcToHK2GLffEDSIdfw
SGCAku322/S442gsc2a3S+DWPQ21KtdPIotRVLlpFk7ZmQcznqtjAJoQw7ENL0TjRvpgBL/ITH+4
033MvdIWCm2GHg2yodf+akofwmqqARvXBunpzVVzUcuUQMprGZIsgj/kKPR19ORwI7MWEIXEVQeQ
TDLND2tUnRytWz6XP5p2qg39kE9xRBLT1VckN5bCkQbTp/T3FsQvoSs6S/cXh2HnwDvC5F2oTxoL
ghLzfpS4BHec3AB18zYtgDHPLZyWawA+HUSrZ9RiAe1MX9qt+FBB3TJDoPpRGRGwO5ee7OOnD36/
ROSQfPUZM2AAiBJfqINXJqns0crp9wZXieZSaIwaTkM4sbKeZD+7K0/DJHpeHpfgwJn5cVLjiNMx
6Yits44+uBLnsvkBarmz6k8gylzdoUI40c1lTlO4166eAl0GdloN2EQfuX8zKTUD5uWrmHf36BDK
fo0j0MxIhV2YkQvkpgHFbcNzcbBKdHUPKdtJPqKg4wsPU4OrBC2NMhQMwoYHc+B0m1OVg6ASnsHe
Aw7B0tWN3xnBnKQVU+QYo++nhMAzly9rGzTK4ECz8kZ0bvkUdrLvgik5pTdzMjVVuTLVf+YJR92c
Q1ZAflx5K6k27NFFS0ITjz7EaFMoaVyR+j9ySH5RUTO/mkHjPVWr04yYp/HY/DROgPZxmKKBQ+oy
FAUXPYkgo4+SGL/00Zo8Uix9iY0Oy2hotQPpxgf1FEWG85rhmTIAOfZfZLkIqz7YkwpkZ6FjmGpT
bA7ItKdPowlNkJldOIQqDhGdlSNpjexScTJqopx+WvhauV1TIHnI0+2gbe721PN+FR52wbccF5ut
oXLj6kDKbSbL5hQj2vskIJZo1LqfbKhwx7q9PWi1REF7BT7rd8PGzjkzU1qpkhv9kkdIaJyrOwuk
j4dTCHxs41DZHSMi1a2XvBkFlfGnZoNlQ7V4ytcCt5dL7GRZxLQLBQ/VAHtj0j87F6kfDS0BnsBT
Qg7Um/CavAfL8avjPmr5fuYZVH8780VOyl1q+Aqoaj3jtDTDAX1JNwfAuenZJI2HAhShFxYf0MLq
BlZ/PgnxFtz/BX1f95Wt/P4ArAWo7B1OT4ZF4tjgibzy3ZcY8jDCWxY9m/3UjXB12QO59uNb8iNI
t5cmIrq8Ibntglm2zihodBG3O25Ir0xdccYPSbRUIVBD47+h1r5UM3Sjjj3IMVfzpsxlxIoQ9w5J
E3h9L7+gyzRPfgdBjKdH0C/XifHUG258D6Sf86ESELPvCece+sM/WV1iQ7SVDgxFbIfa2Fx3klZY
NEAAXxCDKFQ0TIDzKF8QdrYpa9xIcnNbQukOSmNiw1rBtVt6LE/6Z0EjUo2wMrcWZDuMt62+jHOm
cefgKKiK6NdO53LMBAprTr/Drn5XrJyE4BrmkkuQd6sV5P8nk4jwKzj0tf56ts2M6K5ajhIHMsk5
680/1UoUOiiaDyI2gEi04h3qZ8mlzEXvhuwJ1qmDDD9PFPDvK9RjmmpOYxOrZiWqZVRx+y6kbiDu
v7XhSm8xw/AhCGE+ceeTVkFFXdOHn8g60idbVjTU0AtugZMdqtELO5tHZVqOBTPqS6mNxaEP+LK6
3yVtzjtcStVwrk3niOJbuFrQ38qb87gnqJc5tUSwPDUVPD7M7wgBKHkg8PQTbmVmkkHN7bSbrwRX
U0FEHE8yS/H1OM7wAaKoDEgZpkphyV90w2u35MA2lYKS5J+yfRk3QE3sDvoc5lOGvNKt6gKkKwuM
9M90hSEngW7UkaieT0XwiC06KQfdlq6AgMZs3TwKHWN8bwV++LArCiR9bmbbMFODJT+cwMnrd3nm
Y9qOGbUaQPms5P96thj67zZcRkEscxMoeRnMlEBEbdhFE72QLQWouLWziLaE0xUV2ARDJJgLJdSZ
+kopumattHNsPhk1hu5oJMyeBWzQPm+JxK/5CBjogDO2sUIIlPZFbdR76UYorquv9Nq0riqFex5x
HV1E4zTwjvYOsn94ZFuggyMb8RFRYm60N3VX7vjoHbSfult+gVmKdfhvpGguwI8FJhTH9GBxV707
a8dd5p+OjFQDpMDSipkXD2OqvMUtD2RYNpSfxjB/D3BR119urOpkjV+mF10KmkIrsQ6gWrdJAjex
Q0zbhlfg+Cae5jB7OWGeDeE+AY9yqrhrLglpnxW9ry9MZLxWFu/eStwQJ4mgrZ8r65xkJ34keYoA
q74++PP1sW0i/1i6hQA5KCFV13lUmiS8YRTuZLnGkOsDztFezJcH1z4+gk3qwT8W8imH5JqmA9oL
EjDnbPE8T+hmk0z1MoFN7gdNe4JPgS5UoRL7uNtZVTASZpzpoZZT8O4rew0939eT3CoZHlvJVpCx
THjRjO+QbuemHWExQzOM5RFkeLcKQ3xq3zvEdGUHT+4q3PYaDd9q/YxdzwDlLNCMxuK4RoTeEX00
FK8+7/e15vyzbHz1WvrlOf2+LRz7+h8GGV099bNB0+o2U4NgwUWk9fbKolnbL9oU6CwiXCPzbtMe
SidpSM1kiMQjIcpIOnYQCXW/Jkqw8cY21LLDZliehqB+Q4jMralWoQ+M4MT+DItF8p5ZHSdGJzMq
rNRqqGxRb+o3v5I9XhPUEavKuXnHV4sQVn2uP78TU5e3jMaH0UN5ZRwYshT2lQNuNlC6hqMvmuDx
m6267mNPOdS+UPsk+XsOVANfqYRmS9aID7VOF+9guHdw74WclrdwqBPpVV3VJr800R3EBpcPvui0
gxEhGtYTlsAFaShNzSb60OmkeS46ISXMEqhedKzH67leUX7uXyodQo++C2HIrZbsNW0jRnHjHGsg
wW/7Wbi8p3BIDqJS1O3KamxlnJcoB0s+fRcREwnVZYT3fhPcn2Cup5OAP9sExOv8PZCls3pDFdKy
MS7Jl7yUt9TZqlDozUmu38IzUm6DAoVEnKfHuByA1+Hjm0luTugnnPiG4Dofk0w05bmvDAJCYQMq
nYizT5zykKdC87GwovetXmXDN91phn1SiCdJXe2bbUTV7kFza+ASr3y4aCAj3V/s/dXZWN5RyVI+
pvfLDMXzh02vRSl5Tmpxmpw0zLKnLcWc74cG9oE+vu7zDzEbU1aDSXaYOAyO6f+rUVUx4CvHzR/C
QuhjxP3eJSVR/K1gouzg+NqSbt5vliQxNm/xm88lXzGkKtD8BUVobd0GMvURgIhLt99+JPo+nIz1
tdm/s3+9xODtXthXnLWVGE8IKqbjz0wNRaUHDOfL3uNAbBes2EsjxShkpvKZDNdd7tl8+kWZMoBr
27chstbQz7w1CrR6H2SLJvDFNOugJBMoZyW1Df7mTE93p601u8uRMB5ABDt7zPWMH59agR+m/MnT
1G1JwgyjbJAPHtJzvZFVibWjG8xE2tzwZrvFlNS7LSxlMr5aHXHjFIUfLTteRuSaBL4qUCctXYnq
Dr88b12W6oCZDM8ZwBY57Bzygt8pvWCKKxpCesw5bRs9PB6xEo1XsDCPhs5MRY0Eh+ky66tPQ24s
mgNu/EXFd9X1q5HUmPbk6U4zV3IR4STk2XPbNycKyj8zr9U672yZzrUrcxGtllFHjJHgW3CS1aqL
WF++Tw0gDFCOjyPiNdfpsvQtOHle1eiwuxBGdLBemhZd9bhu+UeY1TMVwrXbK1j1SNzU4QUek9FA
QjY/nn+Z6QCipTNP5gB1ziuo0eD5KBo+XVHCXjwA9J0rVPx9cT12NZMZ+3SwlyxlviAgfd1bJbL/
qOQNOA3fm5nWQDeHhyDXkMftG+qoFrk56o8BAbPEbZvKtsSKxCYsgRRBgjrPHMOXBSW4IJJOJYPM
fjJZrRPIyYxJHBCrhvyy55wrJ0KbQTgpL8OCpEreC8emnt08E8zc6Sdenbl85FYxKMqo5I3zZVkl
2TY+ubI8Whenm/3ibpm2mAk8nQVznPNgFw46CZXhksCb1Aq92K0NHDFykKc1/uyj+0kHlikPddCQ
L+hDKHkxdJeQ+iynUX8GjzeliHy+uHN5Bevfxgnq/v1LOjBP1TSyILjU2M1QPs+FVzfHwexKyfSh
JeWhsj8KBj66x7hCm9HlKOYwPoUA/t42ouZHdj7SHOqXr+33TJxGXRe1ZQNfDd028imxTdZQrKJ1
a11Jp72cZzaQQSauF+5ZbQAB5XWdVQqHqpaWVxy91tMbky4kvun/voZ56sijq9m8uxG8BGarjfxV
O8Rye/U3FJVUmmIuGJlhnw/HIeavYrn/ADcxSRBrOIuEjIzE8NmZh+U6X9pN0z4tZBc7S1uo98qr
GNYEylXNmAPOJWP6qJ1VW72LUKK5wI8ey4y3VzfuCYBEn1Por/ryT5bjzgT7bsb3IMgWDra2zSmd
zuHP/q9bfb5EVlxaB/FL3sD0C3jCW+h62JRlu6//ZOPcETd4eogUVJFP3ry2BMVukimY5SgMpKUQ
F2COOtmVnE6Ycq6SImUhpA3/aJRpvKsmytHzEsU8c2h37eddeBWow4HSX/bLRcoh1NKUwOSdQxcJ
BnE5o+p5zULO695u+voHRH6ISBR2Dw5iGm/gvAqoEsiteqCnFtW3UjVeWCLIvDES/biFb4W2jd0Y
Fth9ZLm/qcIRBnuM7roGxVHXFmd84xopXbGafVaVHca6THv/TWrwiWI8pbrTxZbk3is8FU72AO4T
m3DrSPv7teY17eHmbwYcx1toHK8JvKf/bsdfi4iZkLw0xTUDn3XLsg7qoG5FNE/rAiNqeZZJlBgt
f4xqGxHKEozHFLssiM2RNIZA7uyYC+EPXBYNZnhOTsUdzJkI+IjjVO6GE0qRWMY1j9fGKy7Vp08U
iD6lsVHR4sRXpYPiGePTmiQbpYMRBaLPakYltouUdMCBo8BRSh2VFv9U0ryyeUHXg1nmasYpls0r
F2paImA8odcVY5wTO4SFyb3LQoTIkfopzmjVSz6JHiSdMX5aLgeyQ8TEqwvHGsrW13kFm+bmKInU
CPbtqXxTHIwABHVe6VkOP3I+uL/URFdO8JkPnjtgo7A2UuYPjzhyBSjUtEUVGWmdQjO90uPuQBWj
PSl7Rsz2RlaoP1ztN0PcQdM9Hsnr3Y0iL+DWiRS8tUG/huh/0pIpO9m4OYVouCWiwGFfhj2z6Z8I
1w+XRfVvvyeB46AnAKsWBSwiC5FMNY2/FgLVVZ9Z8MV8rejPZcomN9YxNIF2Yk9kZIJjk7cBCzs4
GVZ3oPi/1LbzhE9Dde1fnBp8yli/xilcIu/IiAD6rJmlETD+JH4zOuZpcpXv/GSW4ITZSR8h0w8u
O4DrRCtOKF9zw82bHgayEpgAlGPxD4Vt8uKIEkwpADgGREeLJr0H0O/dlTymIfJuPnorEmVN5w42
2vWbLxpfmAHHgyv2NVNyI6MaAB7wqrzD3rlg9wR5eKFTIvn9JXsOu5QV6gj3SD5L7qnzwJQEd4mJ
QZUl934fUaZon5DjZoSw78U8xLUX6Iv9N1HsKJoXMT429UvZyuS+1V2dNaE5enQWh3cqeRXq/ATl
K/VufVw/ZBm+GP1vDeP8AhPXA7EvhKWYjwAFQtKT3IypdEDtblwG5iCaMAkAO1aQ3VblnTQhU3Y4
fQT2kzaWxsL8+0ZbDRiDvLCDYwVzwl2+iQYQoW9viz5OsiPY+EkmeHrKJExxUYH0GW3apyx5JSmn
BNDCL7GiQQkglrhYvRIiVqKz1sF2XamuuruNTJlcIoTjryRB74/HTIt9rT6MlzgOY64wAy1W2JcN
4GicTdaV48J0KGVctszYOWhXrGp+DsmqGykkmO6XOKOF27KmzPmjL6BtxH8FRbDmSSyxXmH6W3Zx
yP9Ds1J34gHXVrnrlNi9S8zqKqzTdho3C+FEHlfjgZ1p5uG8TB6vzBsOaSBsnjklCD+rTpL6xhwN
o3vpsVlLRsInvjoQZBudHa0bvGUOlBxEKHF58GVIl+x/NO5GWgCI8jRJQ+V2mxjN4HpmbOozFo+8
hcIGbpV+Ho1Mp9OM/O+5a9saLvDUNAmQE693vlpggR5RIbx6NmVXSXCSEPoeSVDrUr7SKyrMt5Bq
zwDVshbHHWeVDGBwgwLHHXfyVkLsC/EZ7ANUUnMkRx1pOp5WGYQXojl2T+zNRu9GYcnOW+nJCO1R
DzQtHEAUZCq5sYLYpb5NS5LwYkN1wRitpWscvKrzdQRYek4Ff+gPmhMig+XuNkQFFHjSRwTLfPSK
suZ++gQVz9m2mQaMPC4J5N11drh5CjXmcb3S71/Ov30WQ48QSZf1VXl6TMdlo/76fCsgy3cdsXsK
yaG/h9iKgtGMennyD7KquFbsAcok+DRjbt8xLXEcz4AUuzko98wIMJO8vdQMbqbxZNX2MIzz/OY9
Q5OG5yv5MGn8wzo8z+3meM/3A4hV32Qa6dQw7FJXohaaLp2Mp6dE4aAQU5hWgIwAkQW8+ItTo0Yo
T0r5xzVdQUQRw0tR/3sA+bZd1OVdldte7lci3h8Bs38+8P3HEbWo9gJiOrbFjz3obkTvGrQjrCMz
xeQhDeUT3t1vlfC0Lxvmj2MpSsoDyoo/6VNrRxu7KwUtjYwCe9TC+8JsyEvG2hWi9J6vAYmQVZL5
qAo+lhdv+wfZ/hnJJxFWC/sHMuwZF8UOepvDrdag1+iX3/34AhqAG9Duim2Z0vSay1uJPWc+lF5u
ZRZa6iIfvuZntqtw9ZpbawqEXDE4OVeo+tyYqflY8blZ8IVmX054QIiWH2Ee4KaOJRHTABxYE/h1
BkFMnUixLN/7cKiKBD5lWnPZzORselnJHYFjVJ/Mb+N4Q0bBWpK2ZhPJJAk9X3+1/r/J3j2JA9h6
JzlICMYIWKVL0e4HQaogSzpecF1gpde5+5FIoIWx+x9hEThASQAezQZ4MOt1OU8y44Gam1qhyDj0
8h6e9EHXan6MJS0V/QS9gf303MNAc8ogh5SGPEdLxe9oXskOxlGCtgXYg7hPUxWGmkT4+9L/jFLZ
kvbVw/kMfwIIpvznSLc6n467B9g/6bdx8aWoBOyy/vxB1Ds2Dz8+cx5JPkFSalaKMLHGPF361uM2
E+7NwkXR5t6JSnl98nglF9vtPrAuMdYZZSXPf86SJW8MHGpRp5004v5xsSCySjUw5BrYGvNtqZA9
5TpzfMFRi8BU+Cmz++OYAkHlD0IaBEzicw8njsYOEHg/EwoYMUrhyqd1yMSFlwgQS2Fec94eXquX
6AxMcgZgjB6DVHKIVef1W4uy3X4MzI1FcCWd1XMHp4n6jRjc7nAj6ty669t1HY01awk5AQTRdQhb
OyYcFQM/eY/ST721TNHzr/Ye8pHdj1v+gbeoYxg++ZFino9+eaEhS4KASjsmKSr1/WCMz6wvSy2k
iEb9kGdVRX+gzLXiRKNJ+9xmZTBvQUHHEZFUlcYg1eBOxb4Y8Kliy+p1gRodudHeutZ+vqHs3bzQ
olrxUsY2lQAY97U/3EgskOAuFnHrzX1CKUwdn1qZHHSCysOrpThRDzBMAhMHkU6Ktk1THQBDInof
pCVd/3nwc0hL18c0j5r0LG2URvLT+19yS1bNeSaZIrbLktHUJVvBGZxNnH6oCXBUKocrdyx4VTDN
lQUOxZZ6TINitEIsKLpgk2doWjywFR+GBxOpkN68AOi3zyJ3mp41cuGm9IKmiuQph9jtAO5Hw8oT
GU7NqGtYfrQb2Im33a9cNlxjD6WJcDjXQ+Fqk136Y3kqkf0swHWofi4XbLEXYV5BjOvu5tsbZBQ4
+HECZR4rwX8CUjbb13Vl0uX5Z0C395pEwV2zb3vvogTFa9BCoqro2eIVIc5LL3W7TemnjQQqj/Br
PXIU0jo85zbP/R4gC2IkFAmqnzIEOW5ouUs1aHzbJxtONmWHHrCzDWO/1hH1rEF8nV7jYvQ7O1Jr
qM7rLnl+9McomHf7M+Fu8dCN+WiiR11PdWiSCKvxNm6Gbgap4O6JFM+Dj5XDdQJQtzkrAldVGsYA
Dpfr4SCWBUq69rws3vn9FZu6vS4Qhd1hqMDlAgMWwDQEObnIxL6XqdO0USmSl5XFHX/FtNC7lnZF
qb8pqXRgDRfZ80PPrd8RtmKcmm+EB8bK4wWvFBf2qniJqmuSgiKlW3b9j3+RsE+IRBLrYbhN6iPi
N7WsCnLbOo57g+64tXIWXDCIB+aC1oHlHoytB9OzP65nIAAX6qKcMtqERohfL81QXCSmUVeaHZkX
Vigm3CeqZil7U9n23rJXMx84afJHLXTnzsQhD1E/aaiohdhFFZhWulI2Jw0ItU7/O0RaEykZ+5AY
/id2pIJAJdDzzgAExJTpVCLS4Y+MSTxXtHv64LUQ7Xwe/2xaf/R8d7gw+zzes6i3Jh9xWZ5cjy/Q
Ac4Ig77/Rmrb2NRjCJ4qhdonib1CBeQv+BiGlzmOmi4/LaHZFoZKnkSgD0CaNZUlWWXkZct3m0mb
2Eh2NQN9Qzv+N1vKlvkbh925L4keFhCztsbFTfCGlJRMjAX5KtQppNU7M84oufhRGqLNvRm3mQyS
gdQ+JjBWBs4NydhR8yLooWJ5D5XLIdZYltGej6LqF+xwdd1cnLZY7I5BaR8LWiI+axNgtNEHhwbG
N1/xRt3IIisdmXc5vKlVRsMET7vRa90TGchFAIk/+MHcki69Taixl9FcMI90DxlLxUQedd/VNvBM
2saiRm+cNY8nR6n0sKflDcQNdDjFqjLxLcmF/8OPzpM3UxkgOSojnpO/wPH4eHz3qsPKFU3VmV5o
60RtXgDU1W6MHBW+Q7YHy6e7oxkTMNaqm6hIdYwLM4x0NbonNe4Nii2GlulbhkSQ8zrnXvIMu/QI
TtCtz6JR8WoxD+IeNbkyjVzSH/dUO1F8Wx8TXam5B+fVd9u8VCQ0CuIkFVe3MRcPPB1euWLuYRB0
IYklY8Sw2IBM4d/F4S61DDdqFF8mPqTvKregroktBNQTy1mBnF7UonA8/0xZXZeiktM3vZWZJZ6p
LLDu5a4P6azTJsj609IkrzrGsl9WP6rrx5rUuSvvhbYFQJcbq+oa3Gl0PZ5/y/dkwqUzEvAvxMdK
cVJvYs18SQhrrybbYNfW5dv6w+YW5Jx/Nh7f3L7SMcRpOWQJWpn6wy7e9i2H9P5xkV0vVmX/hQ9g
tZzflIZ84uTR48GzuWLK77ds/h16zx15fNOEUc9qrmB8Vn2Xa7/UFSCZSKK5DJfy0TWiBxKxEwFJ
3pc97EaHNVrJyv+DzmuIEJ3qyPu1L11sDnwG69aW9+OQQH251fSDzQCOA240an4iQuvTqn/28Jmz
or1ttVKxcWpjy8fn2T6DKcj+fifRFvk8HnjQ5dqIrWX9Uug+zk++XZf1Kutqspjdzn2g+AuX92QN
gVqffprlN9CSg8Nx1/gyWjikhnj8QTh8sDFg2Pnbl4x3XPB4Y+/woMehxcK3uVvv+rjG0ENx3Qjv
gu3DiptMpYxqgRumi3SwuSLh324ygcMBfHqMePqhvDB8FHHX0luGLBhi8rQtdpB0tTbvfL7agiBU
biK79HxQ27pATNoAxLjVZtUVyDvoA66PT/ejdRV8qeAV+bsmbBY9pvFnl9pAO0knmitzlmRf+Aba
R2X0ucMop/GWV+bOrByxPjv6mWJbCkNPbldBtuRpH64jWRiSAWM6oOrGiaWq5T7CqtKHPwnsW8Tc
4aDStxZxhhzvmwJ+SYUm/yqknEO8Kfwv9mI3ug1x09S+p+nj7/SL0cy65m0Ol62D+we0CR7uDb8N
i8X3/Iqs9y+hFwdzpshp6Yp8MC91HDJLulpb0nm50RB0QAO2fkOhNsE6fH9/4oO86cSY8ATtQung
FicA26lhhoJRuVcFbcftg9LatnYPcLhSc0B+dAYQjSUW1rurMTgHFJsiLyKpeJ/BB6LXtj3lkb0t
2JjJ/7xADVSQcBLBO8J2nl2HT4ini8HzRAjvmtS5oRWIagbTTvlIA6oY1bWp0FDp4YBMVQIFC7+v
Wi48jarb8Wlm/3bwBfM1rkyJgM0ZF07by9KkVkAuN5VfTZRNKS/9xWlrmxwXdY1VllU0hPxcUluY
HPbVRnCXRJMtooP2mhxH6lyC7j3PN+m/FJHK5faAYf2npYf5LntROwZ+btkP/8ZnVqQzAWBsvqLF
vRy0z+GvFVJ6PX1ykywxMQ8VHXzexLhPEe4Clm2SIFrWiaNKns3EOkqeBPa5ePROBlPEgBzpuceD
QW9ylnDrfrvOGpsiEw7HnlvUK7sM+OirN3av8Pp0Z3S0EXYbMl1NNuTV92/Gde3CRLizQJLRbQ/e
oG2ASTKO4dTQC6ujj78Y2vJNevh45H+5npwt3Y1sGG6jbd6kA13SEApSD9fjIxYoLt0w77ye3mqW
GLAoWGdCqKX2FT8P5exb9+JIGvaV+qHTx+iWaMiXONmoK98Nj/tHLCFlG5KBNBp4yVH+Y5hYAQHC
85diEDr7YdZNd2Un1YSybxKkpMwlc2iYj5zz5KzUDcVKl2MnMdvyPQirxtOb3E3wzzFRzvhH/pas
jcIi1ZObos/8O48gczEItofkFEUIiZPWgDlWWsLpFwxW3QYBJr6K5qIPx+E9rT6W8FSPs6A/4yLJ
t9gV9II1LeyblUCfnPtEppy7IZEiFRB1UvRhNVUWgFcgDioL9vT2Ks04GqGyDo4MdReUzHJxGmma
1Pm5rLWGASAk8hqb/QPEyUBIOQtZpFB0zGXVxtO+H+PadvaYu7uEezI9QWA+B6CN5zOH7YwGtbQl
s5Lj8AoM+0HCHhY3rU3iL94f9+Np5X5catIDvEpCSRJwtO42rpIBByEZUKngLtpjdtQbKRCZ8OxN
iKqA1GvVMsaiCmwJamoSKSRrAAn5GjvFXJMZLuOHKZjAFDd9rv0eLOcYWW1GFnhQ6AlEwLc1ULuh
ahkhCmtXBDdBIkddAPtGmdrk8rqMKwDASnxaM0L9FVMQjOXh6KwfPISuWVCGjhoNtVmjn2akT8io
RvlEjOCbeO4H15++8OSF08iuXBwsEFm0WcL5SheJH2Xc9FZwQrW8Q96dcv1SxvnyDj9i0EHkNrd9
tIgYH0ZEk/us3ENV5OI9sEOe3tOVmdISfeSY39te+z8/22NqrfPx6D+3pf9NxBBlaaJAm5ht1Hxr
lbQEWqJnJoeLJ+lvcZp8gPIxBoY3MgYcBfvv3QkK0DNlh0JrdtFr8q/vp6U8V5rB87V2/NJhYfo9
qwtpOA14Pn5vlxJMv8XpAr84vvWyR2PXCip0UPI+72IOf//VXpU8v8pOcHVouSMaLTXTnrojTmIx
qRPKZlM3O3uRol1FlgU7vdalUh4K3RnO6zjJ/qUCHQQzxcnP4mTR/FDq/GQAJFfFwPEXZ4uabfoF
+tF5XhZKIMCydIXuOIQjrQ4EytXDajTCWucmZAHQVb2RhT61RB7oftnqAk4jbT5P3FBQuK1DvM07
7FfnIt0a5mdkKm+mLIlZBjEzkLdYTSpFLejQ12Qa8PmVCk68PM5Jhxj43coTnAl0LJ2dSYqoJ77s
v53y3cUH8InG4s87X1ZgPJfCqCxBx+jCKoUyowPyt0TxDg4n3TOHNxQF97lRpN1evAoua3qD2rEx
nnsEbVbwTW7uSA6q1Vl0eXJ04dwauFCjH48UfKgxOjPqcK+Pf7SLuRn2JWzmPDr1Zc80SGMjL66n
1NF2AfLaYNjn1lUb9EhrdOl+tuSyJSW9jMSYmQUI1jDSrEaHpVcMX+gPhUk8qeG6ng0fULh7+NlV
Mr65FdG440Rm1dnGZr4tMpYqclLCzj77N2BFXJwtiIOnU89lIe2igPuFYBI404mw0JTff/WDWsac
CCmP8ZvNdPlNA8lJguX6ePHO4UhmO/qGIQec/gFkuRSlBo1djaP7+GCQKktsDz9H96LryS9tjbrx
gMz4JZKLaSoLgru3B0Hu8OySZHpuHG/EVt5rGLXO153kOckU1KuKXVNj+MWKhVinbgQmbHLBGmnl
8ZJyO9wQChogBjHlusRBexq11dJvnDNZsIhOiaw82e/sg4nu6e2v8mMnyOSOedic3bAWBhe88B+z
y7QJCNRc69z0sqwJRVMEg6kS6cPbsWreaiaWBN3ZXlaZg1K3GZw46qpZEe8EAIw4rpih+0aUayZn
ZkSU4CehdFp2rPqfJggUyipGnwR5iQMClWZoMmKotTJg9Ti3XL+WtUJLqwsKQ1hLikEq5tWs9Ii7
RoikUkRzgrfGt5nakA5LonPmtx2zNzqKJT12wqhzsHpsxGQi5cr3K7nR3eIpf1empsUMymucXcHK
C94gx2KgsoyCUgaGGq+w0lcfEkSeCkbzHeO8MzzIGaFMD5bSAD/wq5gg2mcz+NDyp/EW4S+Rcwtp
u5fbUoyZG+VT9uNtT7JRq/QoH/A26x/+d1WLv6YpfIZPO9dxpuLKYrtMQ4eW2Hnk7aHywa7T61LT
nHMnDWsyrkw1iQe3TZ+x/aiLhccJ/WSX9Mfaki18rYJIXruOBrH0okmjSpHmuSBccjjhpKs7u7BP
Q9pcTZ3mqI5ZnYkqyP4V62mLbf6+YpUf5uUcHXEcjVTYUo+VvZEfS//WFqvK0L0T/ErbU7gYGaSR
ime5HnI56l0kBjNDTtXa1juCfsi5kiSPTmIoso0apBfsQ5i96xdyJwHl1I9giHjJ54yFunNoUmkt
EaAnCStlH5VmurWmCOr79conhT6SwdU8kJj2xOGLNM2nz+SRKpNVQYGrRG7t8AUIUhlf9zkEY/Sy
fIS6yWVHC7IxKx6JdeGnBRmeb6ZvPzHJLrPRMuXWh79bDNG/XJCEy/Br/eq4qkX0fya1JxlHOpGc
44Bvj3tP9bLKXjlgmDmWPRfeBkajZFEOrqzeDORn6YcH5HUrElqBZ5YDUfnAELUUhAa/bMSmk+Ne
Qk9rjncH6iRjoA0c4EC5cAEHRv1s2K6BdXF+vrzGuh8OJ5vhUwVXooXvdikYd6uvCaD0RJWR+nf3
uSczMVh57xMYaIKbT4IKeZ8YYrYvB58XsLD7g0JIq3BwHin9hY0CjbD6LgS/149S/c5fYEBeN9OZ
qPBd8MqQ0asRXnp4Jf7BKP5OW2Jj6u0H7Wv/sGWpfKbdY2P+Grd/mQQ7eTFXr6lRTufe591U3VTr
9bZaLug/WzJC8T0QnMDU+d00KoUVcarYXj4wYljwvNPpDaOQttEBzOCBG/1MXxocN0m93elYE7vY
qtPW4TLZ0eSo3924wJyGREuirfQeHCiVXY60uxn8NtaKNFoSRsNDCxopFlZC41jF1kfVq34aI7sf
Dx4GbU5iXYofxlY0CeHfMfZJnC1mc8RZMW5tqEN64SujBGjaqidum1XAfVbr++1aV3Sg6eL41vZq
ANmaHrV8K5EP21LGGO4CZFGMPCyg0gkAQAzoXC70FytQXORnVmnRu5LTkGfX9ao7FiJfZeFnnXHq
pnXGEPc0Sl1SVmNlVoQBEOnLjXnhb219vdNZ4ehyHiljd9aS+l4paiWI6RvJWOyOLO8Rb0q/03hL
4V5+oVVfJKwCj+yEmIAO0UrbT9mnCDE8qxus6z2vi2Iv86QCdL6z2M5OSslqf6Oi9wq6dj+W2gIJ
LDKRyhXZ/MYakyd+gyeYJKLtzdILEUrVmEg3eRBQEjIBGqFeG2Zut4XDhtpwiE0K2sRl6cBsjomv
/fUQI9ERSbjp6FuxQw1FK572HQauAnVLlLCub0Ynl5k+Nv9ALDm+Ry9+kyeTpz3fTfUlXwn+68ad
rjEsJG7WYhgAEm9ZtwzorulhGfm+ofMJLW22aoAp/hAaRXkiJJvjY8BAkWLOrBbQjbz9zsLBx7LD
a9Wi/+++KgsWZKvW+fOqVfoQI+nVDB7Rg9GjJKUmB6+1XMkuEfN6OG0QH4e/Rc4fGWyZ58UDsY8O
DHaanYJOiV1C2ealFSwvZIDCo3+nK5oDrIU3n2G8kAOdIqzGxAQS3+YKfciQCFFkJidRnPYXYg5A
cNolUlV8dKmrlGLj9AiSo0OseMMEtGibrlx+DI+JMMX3U40KHpFVODkXRWvhydJWNt4u+9oDW6Th
eNp2QvLhnxWMQ4C+ybFakI6ijCJRfjyn+JWrQ/cXxyI3ewoRd/YOV/5gz8KvzZ2zIf/mwDwP01YA
bTcg9rNCzsD/3DjwHvYMU1u5Z1hmV34BcD0LPsDFgWvoPNDGpxXmxcmQhuVQ7ah2/Bms6h2pGfEC
dgwJMUuBV2WoVvvEH62AjUtNktEgGiMT+9o4AUaDQg8brnnadB6KSyBE54OfRQUjzDyFszONJsy5
bnmNceODfWCOBiRBwGxJ0RAdwKFSb/6u7XMUzMi/IVIQ5gz6+w4kX0lQqysybbUFO3V/vVoJ9cec
r9hvfeBhDQoqLyKCJJ9Xh0yM9dksnkY+Je1iujqaUsEbl1lcKXtV3xo9JFNkEp8oFh2JJwh03yuO
AvNJyCAQTmPkMUB435MvAu6r7QnLJlS5EA4TNAL4D34PYV9Rv9bwbsa5iG+rZetm5gX95+Wq9x2u
Jl8PPfygX0Ybn0KIEA0vsjn5G/7bCDE6fFcePp0ixZQsGNha0Su8FgWb1dGfDdQi+ObSIwiU1l0W
dTmMGz0FrSKh8LjOtadYT3naQZwrXO3f6Utitz1umfhGdFJsWAcBEMrgqpRJ7tpeTr05gD+N5loB
EOw6n+catM1vto8Lpd7uIKhhYV1Ezxpw4NnI923LZBqnpngPPe5RF47K6C/EdoyjRXxF7UYjM7Pv
XnRuvNPPt/14DGFolGbH2sdpLG8zMVxZy+0yfJezYBVfFMi5GBVY1FOxwMNz6zOa+0TL6aorbKGU
+D6kVtr9mDv2YpyCdPF9Y8QUM3x8mYDjkgbEEbUXx9HMpXM7Ja8g0mipCSod5AoGZ2Hx+ZGmCbKJ
q+Pwr3/cPhkWGMfCleU7Q9z/A2Tu5WpZSm19eEzn29pUBn27kXvhn1GdC1rDOtfdyPnBOL8Dapvw
Lhxz2oegP816eOEyfax1828zdEEG51DXicEr1uPUdZQe9ojezcG3eYkm8h0YaqK00PvU2VJyItZ8
Bo3r4C3x9greO896HU5tZvMYUeQlf///SNkCgtBhdq6iT35jTOC5bDF56qxzke+jZYLtaeJJ5yAR
VhdCWJnkqbwajhfqjZK6ZRUlymLOEnGKLAmf3GOBSWxqY3LTgJYD21UUueRTsZPRuUvMD52x+BIs
D/yapMDnY5OBPshbdGSqeaDG6U3EBCsMe8ZOk1fbxeQdoD5CWXMrRKwC+ZhGOjUjMXoy3/8LDpSa
3bubSFKsAsZIDMMs/fuEIcwsAAIThNREFBl3Ks1/WjpTIzcW8CNlcpn1NgBSznw0y+amGiEOVLJO
GgpJmR/AXvuc/RNomc5DqUj9E3Lz4hwFczUusfAgkPYhrwp9d39uf0ScB8vkEdJgNMhvBprvdLNh
pN9uZWgvHF9Jipe+ZBdnhgM0te7nptiTCzGWGrN8ETUxvQqv1rYaRBQcYdRCWCGukcpgy5i7aRgK
o5opC+LBf6yme7vgNbPcNgAwEOhlSLr3qakbxlK0aRnUW7qq0esCOF4mrX1rwWiWYFoMeMUW3Q1j
an5//e0ueaTNHTK356FTZRPoqixrU0hj/XDLvBeJuKYt5J9mEznSNv8oLEkiJ/EG3i8s155aH+Go
+wehiDxqWExkB5lOdWkKLHpa8rCkfdhxSlo+cQQuBSEb0Ts319EUdbPPvpvW269wpzkFyTC7YRqz
MyHIZ0XuIlSlB+KrvVQmlr/KiEJzY5ghN2T9fPckIHtQS54mmAtvkv3WRGKXuF/JE3Q7e7aOao6g
MN274wkl5Kie0wZqtxBeAyr9vbO+RyVKorE+0G7IwA/Ezgl+ONSr+L4noDCYGicqaUO3WjgRDRoU
Az8LeWDSjUWKL0f1Cc4qSIadGzxD4YvYPCmSHvy6cANj3nvttKk8I0bjzDmYPnm2WUeAvrKJJgFF
vAUqmkvO7bhvxSYqBEzd5I7eyScwSTnaYpZFsyYOcYihn5vTFfevXRE074VOzzZNZ8jhzEBtNaKp
9bXTrstzxWC8GFfx9PDDB1hokBHYzCwf7GDOmWKDIwpXgS4uCQkfRjoYN4y3wwmDMlxH3jJ4mt/I
qj1xSMVr6HF/JIzbdv0yhD3Y7PyITLc0zyOLiOETC6oVB8VBDC/5kJX3JIPIdZdWJAqxKJFcfTEH
UFOAErab6qdeJ7GvPwbm8G3UFxBja7TStnA5+Joocs7ElYIbnRdJh3euVbdoHtz+jtNvLSYx/9yw
5XQByuBhsjAYV2Hbv/E98lN6CtAKbAatR6N8LRYfL7+7RudkVUdFnjsrlivXvb+J8qvcYgDagCF4
p0FMkhvkXWDmg5TNg668xHTyTZEncZ0mc1aPpBtQ1Us3/VETjVe6PybLbhTnvTx81UlvwFoM25E/
B9ElI27Is4qZ4zUMRugURkVv2Zl6rDPMWghiEE38iSYCNNjhLsaffegeJAsv5mbmsrlRNktRx/CG
Wbo5n47COpqRPydt8cZNNubaSd+02jp/By22G2woyzVF3zNOcerP7ZElpAtqONcIbBuI9yNqCH/b
azb12gmxDOTlXSTXZ3n4Lggv+J8bffnPg0OmCUz68a52mItOt/1sMOfxbJPLSSp+b3Difd/I2QM6
2CJ2mhDkvuIQcZ6OsZ501MZcE+1kUso1giZJlBTbguWDbcSSbO+V5kKP5weR8uwhCxsWLFJN6wb3
w8jyxtpQbF/ToaUXtJdCplG06+f+0ls/rb/UhSkZuJNQzlhKzl+xamLVa2Go7HfsbEWWgtr9+E0/
LF0Nn2uTn5O3Fkd596Khd9MqwarMUQrPPPc7nmIK3zMIptD+6Tf5o/0ko+m69Y1sNSFULs9ENFHM
T90UgvtwtAimvtUXdkUHpuMNx+oPhEjk6RtvNKjBj2sBpNcR4bm9lbKe+gvWjh7/jI4yVD5QUXTi
iOvIJbWgcUZ+ZIiab+iPR1CdpVwbstm3YivubRSuSDwPEYqmNLHLIszrapqaCQpZK7soSXrrRaKp
n1DkeYafSXMQEDBkhVOpG1dFo4N7bz44NVX7OYD3TAeawGeX8rj0vDYYnsc/paoRebujkXxAKBUj
j4ZQ5RPibQQesgns7gVf6bqJHwakbEVMxJW0Hr4IMTrW0GAraUQMAFTeOyEkm4BJV4E6Ta05d2Ff
YwRVsA03pe8EHiAk8TxcNqaDkXZh3JgftWBiiZKqExHRZYwR6sRtrD/o0J+It9GCjLOTwGZX1A6n
840yhK8vgldJuBqtm/L0R99TfgPMiJDqS9AEm4T0n8V7ifm2swuX70EYRA/YQmENMzKQ+EJ9lWEK
nzr7xajnOdWoOkIPl+qXALr9KcbSdTCJrYTzM4eiyftMIUBCbuS1m1NY4mY6NbvIDBsFN8xT+2ch
Kv38NnvxrfmFBePbDLag5Gb003x1ZX1+yTVyzxNQjov3VVFuvYxVyZHSgmu5kQw72Kvb7gKwZI0u
QY/KN40Bu5I50uecVWQj0guDwTuyMiFBdiADChzvB32l9JCIKZA5iClSRkv+oq6keP+YayOU7ic0
fYsTbj2pglKkKI2uv4bUdYfdmo8gHuloVFXPS9bJhxQIY74de/rnM9iWyzAuhyah89fVIr0abeH7
/RVBskmMkF5mEFvUfDCp2guNLtvnqSI49JQvNczmVV6o56xk+y50jEqw1Ut2xEI29UqTKtpB4Xqx
W2bUXuFq7f2UX79F5mx5s0PayhnFdbt2thFDdRunVdQzeHjhYyCViDa+Jd189pnnWdWQDox5z1Lu
o2JcOIEHxXjXmxC78ui6tZDEGQwDOLOJWWKXIgpz8T8CR+fsK2Bx0R//JIq6bN591adhOJw8csjv
PkD7L1ObGKONYLgSsdvrhIi8recbG9lbhLqPtpMzJves8ntJXaQWFDpniITf+AaWwdRu33l48wXd
xvjIChqXhV/qan2ndirWB+syYfC5fxvhWrUUImIRrjuBMeTUBCgBEkpX6ZHKMYS44KcsBdPsoGPb
01VCL+70soIhhE1IJn1WnJAPQJMqKs0xb2WXAEGIiYTbuy3J9eQx08m4gIyab4ComwD6GtI/gs8g
VsvS2NtrneDXDWkRgxln0yzN8ROdQlBL6eTlAJt8BQQM+apWE5WJNZdxY9+W9Xud1RrqOzxyjH48
YlkdhEotxdTO32rEiKoyxsnQRBR2LlRf6NhZ/HEWVfriu3thP7Hp53Xlv0rqKnbaDvQGr9xPJZxa
2iwuGBCTwnM0N3zC9kjQOzvA01/bVco0vgiERPQ7SPWILSxBUvCENYLMkgCyhTmixgoVV6aTtHRZ
5WqGuPD5YoYLNX5pe49XkJ+99W6jTzIF6XUfbGJK/j3KYPx5RuGzlEYfZb8Mgx3V6ncmYL5HE5lL
hI8VOD5imuo8JcHc9LPbzdMaw+IsQmM5jPsgTst0FvDNIQmuN2RUxSYIAKoEaYLVLPsydbcSemnB
eZwydhxHnbtrcASOYW+hGlxI/IxPfhSfhesT1EbJgPAxEJPJ7nOc+BJt1+eWYGyUoW/xGjmJWGoJ
hX+a8ic3NXxFOWn3veZAyTHStUq8ic3511wklEJVjpWLS6/J7pq3WSNZhV9Zq/GQpp7bTQlm4Kjy
GvEDHd9pxrfAGfs4SCEq1dBauQTVtdjPys0eTQr/ZOGSrjUUR7KpABF+cuvj4EGBBVFMZZD5bhAH
LZHricqzo5S75m8H9TqYtd69CNBdKJDgXMP4cT2k15PgxFVZEhWi1z8IXsYDdCy6MrgligHrxgvV
yDyuSUMqFygaq5EaIKp7Oxk07sFxiiWXLDcN5meQ/JGST5S88hMa6/YpKbwkwta8UxaiY9bU3eOX
1Ad7wD8w04aZPfy12FSIFdK+FBKJmtj/47lwPfD6jbPFq+m2Ti0Yqx0Bks+Q0Chkjl4djr3o2x6H
EgBoVNn25e4VrrO9EUMf4wSG1xrMj7ym5XpzHGmuYwxlqBgpB7du4mGwEjnnxCLjQIkGKdiHF8GW
KJsfT4gN7Saa9eJBwx7TRiZkkUZBKpqEhTozkzO0qHGUUznorV/3ZCQlsg2zo6NukcU95GcqVQNJ
Fs/7Ik2Qh8WlWUy1fshswABIzJ0qPATn1xM8/E3CkJiXUmEYN/prSjKtSdY/+uIzchn2xM9swa1j
7FYAyJRM/0slYnb6wsobSU8g7KXHN1lYNhe33LhjmMc3DxFT8DUKyXPR+QTO3+I967/q4swtypNz
jRw+OAYNGsOHxgk1aNSqGBaKDlNVsnj2XBlBQCp1Tzd2fFUqOKY52vpda4mi4AtBFZfVAoviwKA6
4nA/LXyZdxpGj46ayf55q3FwU3KOfafJ/PlckV5rOzTaemMsS0SRtHNHUU1QYFXy3543QY1vbosY
kjAYBMkhyByR7wCK2FI6g67iewOUS86CLyG5j30dP3J2NL9tF0gTcWltAt694x2G5tbX37YNeSgA
MgA9A8xCOyjNBPWHEstyMHfFYl1HNAJ7QdtbJKCR283h8Ou4DRNkpa1KQ8IkKNrrs5T3Cp1Zm+m3
rnmyUXDxpd3aunXrh0hE66lSgljN+kRWQpl3EMqAy6lXOZ9ato8KJBNOtiY1QbcGvvOWqemIraAA
cI44xC3F6gE9qCXrix3FqeYCFmijcWiWYFXMsk9uF46FqN/r6R9KAq1Le26+eOWqIAmKZBIa4BLq
5wEuzIRQL7/y1ZWybHToaAWgdzC1waro/PKyjBxmgbwYkFhArGcXgJQMJB9XSnVL3/uXG7u0daeX
3dEPyEAUanM+vPSnaSYXXaBmdNzuHnb7Ip9qQoTUKGcu1boqYhmJoEHgs9PyF/5xnDa58ZdaKyu5
iK46gEs7aPa+B8v7Le1oRXVaZuC1ex/0LY+/rYbcX/s5zCqlg8/L3545PUiEUFEfxcWx0zaQqZCX
2KH+ReHozzibRJ/eKhKUQiXQQFr//yxaiTNe8McFUNLMiAblUeOOSlnetVtTzzsg70g1PdCEamV7
8J9dpIlHJ0vsNwl60YLofTR5G1wyEK1WsdAXCUng66vMTGNxZn0Ms4GZrGBlag9BCIYK2ExmI8YW
bPg4SnRXu6jbNU/nm2tbl+6g8sSdv8iMImtQ6+M2IQXIo8QG3rhZE7WEAtpLNd4p2akkFxLtuSr3
lMAmPQLYG72ZfkBNMcY8DgzxPUu8Raj/r3OqDA2i5yDNZDFmI5U36iwEsaOsXF4wcSb4nrBhh8qa
IRDbWHVYgHho0ZF9aeXUEFtXrkAYinATiFHIqLHZqeBDdIV16RFY+aHJn2B3//7V0LtpeyRZSX1W
MhmhkbXP73LDJRD8fsilE0htUbhxr1Jd9DvVO10KNm7pLDKapgcafyLRehcJcsh2MbHFCLlo8J+k
jYDL8vXP66WPtX7+S9VFXe7s5fSw1uQysyvSTSQ7JanlsV7fBJmSxMkcC/0cWYFHQYxvKAXOOKly
KXgC1Se/wMURIy4lS9Pk3xgPtLQV6W9zKMwYRGCbBAajbw1iPyfu+oqXr3dR1GhJ7LXvalhxtnA8
N22BwrtoP/ix0qxGD/KAm5OgZWg6OJ1lpuZL3M7ILlk3lmy31VOAS8Gq4EDE1P4DAgaB59thioCr
oe7KUtnWjJ5l48cJtr5NwSERa8szKh80fAze6Qnz7wFICZxVW1cnebvXM1IkvHqkui/+5AgjBOTs
uPD67+/RSXjOySTlD7nbeFkH7zRZX1XgJuqfKaeoyPTueXjTyOKRcnYinHobUMv84qJoP9dwQn0i
R6iZCNuDbIC8fkkmvcnCL6qBPELh++0V4zeZryM1oCcNKBdn2mSRjAY3y9CImsuermK55Z6QTA72
urPp+q/TfYuMhRScZgPO99YZ1ffEjb/uTpbJaSJVH6rS4Ow5BLXi/kXfWetQF/Zcjxvr2OL41s1z
7x2duuGfhIWqEU1eDcIF5Vmwc/6ciQF1t9/4YCh3agLphAJIeLe5CQN8hxSSE7l7U6u7K+ykw0PR
HzSpEQFpyMrx0Ucyel8znEc0ool9WgqE7QOwdNp4znNSTmMRGzQJAgDllwanZ0vl0/uDN3OVQ+aZ
PFeYxbThA3teuCdVB/SP/VSVuUwkgD7j9JZirLtxoTCZoARAhNrqFfAId1YzzzO0nWbWlKs/o+81
IBDMQVpsB8fNYCrkLxDFOu+NQg4ufeu6rTgLKWpGRb3F7tRD8iI3G6AQlw1XF8LJYte1MkWNz3Xg
/XFIEY2j0Q5Le8Hx3Zr0NF5UPtyGrj6C9vqrpFYg59SJ4GLGlhcGzxZ4hjUAu4ecZqzTYJDSppT3
x0rOEXnEJYzHtUqxvWPIWjP0gu8qYDjGs8W95psdhQmui0OIVoFwGb738cEcQ47TJCyMPGZtL5//
NJ4fKR49Ri5J3pWaXXGlFe3cy8vM/Eys2i+N/OWz00kiaJWRNrtsO1RjP7EjjpO45F7te9Bj93+F
W/DuJQFbG2btpl2iRNY568gXojJ+XXCC7vggPW9KOfeFFD+JsKYnZ+Fh1QxmhHyVj+dVxyg0ZlLN
Op1wjd2YEgsyNaX4TQzvqXaTPMyCZuyF/Pw9js5yUPW5PEAFqgbhgUfCJgrcGEPxjiALF9nvz638
yXQe09hJEvh2NbmWHXUxRwpa0SgDwGg6ixceGLkT+1nwl2xvhIUAwt3weJpdB0JimxQKOchf72s/
KXC2h7WTllwFYKR/WQ8Pp4cKjRPxSO88d3drp5mcIpGq1oZMTQVe+W0IFGEYrgTLEA+6QTYCMlfl
YOhhYbrMAccVVmuvWci7vR6u7DcD2p6Y9pz7bpEijgSBjRa99xjg3B8w4iCWxASW3wbMao2n1TTv
uOzBK2QEPQo/LLZc7tQl20zqgjcPvGHbMVcJ5TeQp5F6QQ4S/IKq+lvkblchK6jTWgL6RCJ705Os
wAFcFhbyro/OJfSSODzIIms4KqCyyQJXRJb7qmqPkInHmrK95KA1AQYzZXxY7leRrR4FdY2uMy2W
IFF8Guy+VlnnqK8H4Ils79jDE5tcRxFaNxVawvY6ztF7meKSA4s9G8iXF+51mr1JS5R1URkUg7Bc
B8FjkO0aYcnHEjQ5WNO4dDyh6eW2PQnRe45Xsr8NWYV+dti0Nj5lyL46Mo6oLbwxXwST56wf1Ppa
N0E6aIPuMaDuGoT7GrNVeFFL8lnJ2pZuwuysTgwU7d45zJOeOCfHvYD2m47DU0Una8mPFjKvksQ3
0SpbS2mv1kC9VacTmt0iKNFa25tP5BCmV0d8+mEQhR+YSqJSTum1ZmlrBxAhesw7Kj/RYE5I23E5
VnOMPei+Sw9xOjnwENaHxdCe8HiPmXEImeQTB+3eWrjmoSVb/ODH2NUTQyQRQQpwrilNAiWOloPr
of52f3LUPot91gIbMEtmAB6W8Gu1l5SXw7qaP/Z/PKqKcVa9a7D+qAuhj7UGIzcC0eRlRmUfAyTb
2JXIcFGjaSGycAIO6I0ew4tUjOdeALUpzGQce9J+wn8faCgl710cL8k13Q1/oI4F8R+maNj4IB1p
jKlhU/eunzUMQh19aeAJYmsHG8F/5ji5TNhMbmkdWvbKavNBi4davifG5IdIQaHmRw+0MoJhObGR
N70xX8Ekn4JcGwCJtK2RtnTfwQBKDyOlNPRL92v8O5HfpUsdC8Sw+SPh76e13i365QNAQCKUyAXQ
i4CLNJF/u5cQS99BnBSQJqatu3TSl4XxLaRc12r9bXmBpfBIeE1fq72OeSLpviPzKrV0qAe1b8q8
ZS3Jg4Ke0wkUumUZS/8zDfVd4jye12IO+nvzVlRQrsuF7yXw+Kd504qaiiE3i9/f6xr0poBrikW5
oyaxt2DRXI5g4h94A0nrrBQOoLos2qvSEUvmUImRFiwwIi8dYEqb0DM8CUr4AESlwyCmBzPzMw0c
OHTOwYGcFI8F8nIRhhOcEacjrA8wzrK2c7SCOEdzC7mAzd9mKiq5lqo9p4MWXsby63lj03v59h9Q
bisCsMU6lgZbNHsJlTb767ConoxqIzsU2yaE/w3ghjGVuXKkabOjtcG4KocQiN1xhDiDuG2kt8Lm
KCU9Qht7R32YS+OFJ7FEqhpnUbTou97Ufn+l4a2ahCzhYNOvULH9D8jkSp6Jn0emiVP7ZkJ9zNfi
Ebk7CTyQw+nthyNDFX25brN4GJX6J1V4xi6CwENSgRVxzjIHPADYj5HXPPAsJhvU46Yhld/VDQj3
CpI+W/BxtUa9ph+I++B3LpjE054dLA3Vz+Zl1vHv4fKstCeVyOskRHC+b7OoJ6nqUwB4dlJIJQRv
B+c3zOMcVA0y9bJoAhoNymSEXyM/+kvF/JVaJLAk4zJ8jI8bJk4OLhE5EtFV5pcuTPXgkju7HFqw
S6i5T/BIhG7fDjQsvnOMaSXKG9WvrY3n+gQ5DcaiuipDJU4fbW6i5sPAP1rVwrexkaIG2DePhwaT
d24ST69AOkBZ/mshJ6+iSYlRdmYNzCf0S6AQOCv1N/bGnZ18IoYn7n8mQ25KusMwykFE3z+tLbnT
mTqlzK1iPvI9XLsby3PtnqRUdx2zhhQkdWS3t3NRQ4sJ7BcY63Ye8+iB/erHyIrQVwr3twhO83lT
6NlLqBnZbizKIdweGQvjVbcr0kaNofq/Y/oG8vhzoNgBiiU4P/76BcjBsDBx94YSwgQ/Pm/oUu5p
ft9wXo5Oiwu8jbK2Dtd0Wzsb6khiQ5uK9ILq0PY/C2OOBx3HkrMTyQXWoCNFIVqWvKyciy23ywCr
MDGVS1lwfHIFjf1uDEVwkVGRZb5hpJrQuj4QEdrxUipNbGqDCCz9kGu0fpJ3hg69B7BdDh6G2TO+
i8AHdKNc7HXRO8yDW1Z6qprO3g1W8dkbDO7BuJ38WEybEeV2Wi0GHKapoi9QZ8/jhnV6AGk9XDj3
6ETJVp3M+lENOJTGdEmM0K4q+FO0mwe+br3oDTsgDyp8kDsUjBnIzH8AeYbdVZHTKiK3S6uB81DI
fcS2FCndgeoLsvR7UCTbJoFKUoeMLIjyU9J/EnCNn5yuCVY7r+6nNB890ewzDvdjH9m3VyU2nwLB
En/itw6Z5KBRW/lv6ipEcisk/miu5ejOu7SmcMJvcxFNVeanFgrJVtchbRYhN4e291fK4XYno/ok
kxHUcQH7TMBHfYP8z92Fn+5VKyCO+j2L7UU8VD1mmAlgeLgBKgVz07IvpFAspWZV1itRFtmn+FRm
mhozl8IG9Mce+tQ8grcMVL2kNldLaUwNQE+rac0ipInXmFewJ7zD39ONYZDxJx6hLIBKtbmwAT4T
QT6y2pwpyZ918v3ipwshgCgn8XKtDDuz7gen4iBOLtNjsrBfvrq+r7hz/RxyZeH1FcIYxwue73U7
aMFdHzo5yGLhq3KSdmmB/9YocDLErlCuOnYFMQDzZvWmJfVyBQCi3Roay62P3L5ZIWuVMoX88vOQ
9ALodT2Xt11FMX2PX1Y6vQz3DeIXO0wvx6HsnEjqf6C0L4kD3vW7tOCudmwBLXV3iDtDqtcdZLrE
ZSaoevq09Q4/ufkm3Q+se6We7CogZfYV18cwlgDviJDe5GwCxH8n+h8YudW/5auE4TdBR7nYQ16d
rmow2odcUB8tGKFzsrOG4x7i2T7RiWCAQGvEFMNIl+wnt/LKtT/vhL0m77OoOiTi7mCF90uJpmHX
f3SG4miVOhCBpWRDhE9M2s6pE+hx63uEdxF2NpGcmH6WECwnYr4zdXEIVtmY7cJFufBa1JlMxZXK
UnFYHW0oGCYpQq4BQQvrlS1DaCd9pnAahfB9+OcR44qM7PUo9OorFAyfFqUMKKJZNkrUjBe8+OYv
2zNJ2RXDmHpRLiAjqIAYbxBzUSKaPHgdB35kOHgs1HRQeeaAqgAX5m9SzNx0f4RiWqFbV7+nNPr7
cbfIfuhLOOhd4wU+aK+FzTMO6gX3ZvQPqB9aIjdNA/FfCgLQeRXoisj5nU7ZN+QPoqaa3D3EG3gp
6aRAIMndz1FPjfZhAd7vp/ndAFVrxpbEXOYGBNOkyehbkygKZnMFQ+kwD5Uf1qZe6A53PXdfBUqc
n2PVgVVlA/csQ/p1iTf9fw6jMR6zuSxQmUArMYSVKtG+s/HKsOD/031jwp83xN1u6QE5S+Coqrqb
4TVmjAmu3IMt9uOat1Y7KpdsDb4OVjd6NVuU0U/62hEWgO/Xa3keSL7tY3vCG22PBvPey5lp2iyE
GUxfFQxbUEKUzDcw+diOsvueKcpTa9gaUzMcdt5iTQJSdTrpdVR4YN/Tx9S7z7HYsedUMRTLq9hy
oJh2Wn0SxT3zA9eSJZWR1YxQTB6CAed7Jpzaia6mnifyIenPK0BSzhz8oPyX/yaGDdXtcEM6YWQ2
jViGbnO1VK0Jb2Ogpb+jYSHHrFxqktQPCFn40zepP5r8bydY9X3KSfkajEN/4fsMFaZi2GyFhH2n
dKTEYRIV8JV0UoCf6k0V2lmsrGyT3ZMZRhoIUo5/KimaxYz+1vnInjhqymIAYPRzv1nDSIG0HCLE
clevcFrQmocO0aMkSjP3HU1vsMMwFi3YLGE21iZ37XcjftXHurN/0gVEx5VEEQ3BntMbTCrPDjv4
WjhXbeBolCr6dOZlD6Oz+dgX4XGHGbPOyNirdZ+o7ofjQdlhT0CGeEGN08m4ZhYWR/hNOdJByzMI
XcUUTcuO4WZtSYBHO5+UnQs+9rv39fKKlxen81kMzAtIriAe0L5QR9+QDLKpaJBv5+32GCEBwXmv
tAkG9bvNd0OAXK2J4ung1EUAQKL8Lk7E1IG5aKkuk9y0tEkno1ltpubHv3LCeFTmNXH3Fv8Zuynh
11RO6XOH72/6vd3IDodp+QYSjWTA5RqE2GHl9mBulRhlC56AklWh5j2ATBhce+ZmQRFnoO9hb5u8
dsTtHftsqyBUCS3ijsxhN/PwRXuvMafcHrRitfkmjrT/bwjO/DYkqZCSTr9rtE0Lcv0h9OLCK+vY
Mck/gUlye8IFRsRHGRZlMLKRSUgWOC4iFJWQE5CBJUUnfK1JP8rSsS+8MSwFAVQmBGMQbUMAkwv6
ra1Og6H/peEx3yJl/bt9yLaFGnd2cdHuIXwCQccyZocajvGphx30DAaC1qu4IM7eqzT7ZSgQ7uPa
9hQ1EQ/+TqZMF1K1fQy+id4TP1fTqWbv4+znjhfjgHGQtBhfCOpm0VCVN6KAe/Pi1lVBP8kVD6ZH
DZqod0lslxv+AfJ00Pq5LYYMTrWdjLZ74gpNmMQOEL73lR9T7IFttvTMfU8IxepXgT6RWuiTcaHo
JhBat9x+AS+kbkCxN0bEwm4jhEsCBOsZzABLPdMrhvbKzceU1W66BffHkozSwTLGSvduIT1DJZTv
VT6kx0ZBHci6b80NJgh0lKL/PstdMaKfXPtd2PWDALhLCT/eVFx628PuUgrWaYCUMFiUwySVXeVU
LcQhIUCY6ZsUCFqlIvLSy86mN9Pgj0UuK3B/lxPoy5mEBnfHLDOoStzBgRgNi/iCG+KA8aHHZDSx
pJXprr1S1qQ9A2fB/P7b1yYljB2FoiO+wJDKjXaE5HtSesTiPSw9Oey6z0TJ7ORUWyNSPBVTC+d+
ZbVF8KkXLf3gM27EE75y8eAhh6iOg0a/Is4pZLLvGqpL4wWJZ2PLbg09Mbsh4YVoXkvy+gFFhPUd
WO0KHdyID5CKsCuuVkjLWiSWQiNn6bbTfCopmu6oPYlZGuDs5AWFljydGTevYNS2hTGC7uo7M0nx
ZgYkVvPO6/ULapH2zSnTNAYFK32GTmvNw+4fqLIuxtIm6rstqf29l3CmtF7nhy0EKHxyGU6GSQlY
kV/VeO1IiytXLPM3WAJkMM2fblYH8+O9O0uYMBbcCHcMUZ/pCOIL5HfFxaXBGxzd7gII+QtgbovZ
HE/UM31kSjjE5fHmiF9xiEkm8Xg/aymYvM9tRamA/YgyWsO6lLieIEZW5xcw0SlIDuxX7xvWOQ4y
HdoYltHR/R6SUF5oJh8qUlODnQgeHKg7Yqh+XkxQiSFmbk9PL88P8cn82vH5oEG0PbFEbNJu7RSR
d1102pcgqpMoi8+LFKAivzFlwRQgYxcxGyXY1OjGwFdpIEqkKmMCjEvV1zVlPMP6yOePtJl7pRa9
zqGHclFGS9vg2H7A5o07Z8TMCmrZNUz8asbOXVq4scq21lpN9RP29xKz+n6bDqHMETS8RuDSFpMo
eC3WpQpbhrHBOGXHr+ixxB+rFUetfyQyrohtkEZF01WH+tl1skM9hdlRDw/hzH1oWYrhORiuw31j
WnhNa4tXqwEFjzPwVqHD2jFQTsSsTZkOxDdn1ODnFdcvMDzXJHvNrnMXw7n7UF6/8O0sGJVqbHvQ
qsTzJr0xXQ39rZCuW45gapuV1t/uSg4yc2TulNO1j44i8IlBWIZW6hmw/2KTCAOpy42QK2+McN86
9YTlOhm0a2de8VL2zKgXVB7fQiAdvF6W4XSF9DeUsJbXwvsOb8UolYd6QqDeCRVpaLqIW0wQhvtm
ArHCQ8NAGAJN4e+wPIUqr+9yvCrvqJv5pBLzUdgTgbzD/P/iq+rY9EP0mhCOQPcX/Wi4Qh1102IC
O6ABvVRTem2/QHz6jK1utqRSLRO0DmJGyXf9QNXhHFYy/wAELBFpAiosLgwY9DBu8NX06W2Ro4cS
oN2OzGScHbgbk+nrSndZu6PaiSXCMNgCT6h+O+w6M+Jbs0wgOTmFtA6vVk5LsoF/mUN2hyvtgZ7K
59qQX+Qwf+FIvHoseDL22u+ZmQy3BsBosdUU5rdeOADrwYXcGLCy4BAmvN24fNpKiMI+YuzX47e7
DUN17in52x4bQcSQG1+dX/iV42RtlO/bNrefqo6UoV7ijd7DPp6IYPa9Tmqep/MGKNvInfuzmelz
oEOGCuciImojvwPEWf0iTRWEHokLC1JX9VfThqYGvMe7VDg2dtpbAcMdydhbryQC116bqtuLlVoj
Gujl5D/LIv9RTTMX3ttd9XbFnPxGp8SwJ+LFdDnWSkt2NXTKGbqBub/af4GHBSoipjT7jCFedrFj
PelOyoKJ35Gh+BpmmRO1i2p75AHAKwfONCE3bwvVdLJNKqbeOmYWPQRCoHahxsNDhRloy54/7t/k
tDjZcZqJiL9GBnGxFSk4IbUysjGfZU1t09Nf7KcvdzKhP/mIT24mSPNMw3i4KfAPet+btnrLgxVS
nI+e9fMXa8k1b2xnDJ/r1LVT2Db6afcOaDgzrbBYX/GA+qVVa8NMFqLyJA3Pl89fpvMXaKrUlK+j
bD4JIUn7oIQhpmV714BzcZ/FCPg0E8t8kM4GMyhfXyRgq8MjUPYwerseGJubWSPvZaO8+CPpj8Kv
zbMHHXMvdbB3a/7ghUDppptoVsRyx7CMqaP68x2OQJASoRpvFSBCWUSjxw6PAo5QwmFXt5scZJ+l
C0iAh9HjXy6V65SCvaiDHPxqAMwlRf4nd8Onp0Ris1Df+95HuPp/rC88ITEyRu24drvs8GsXX3/z
Q40x++E6Eo8AH96WSYsNsJd39lLDxgEnaHClQ8FgRBx+hnJheO15B6khMysHWqPU/D6cxL30Dhxo
sxJDTv3E4ubHIApMBVkk8sOLb8Vp/J11NnOLCwwcxVMaX2LyIAyltJO9JIAAsCjJU8Pzekq9H9k4
fZ/wm2jOBkFhP2mgDi3XCMqg/Y/NwuPydCJssIM/dqxbpl82hs1kXm424JAX2luRGbKAUfzzU3lI
sik4+xk7aANZqBi/SZivEeEq1P8XG/bYY0gDDN+50lycYu0gnEbyPcJ7+DFXtuI9Ypc173waVnsC
mZnie54huFl7BnQ112QpLfZOMtWsEu4vYwwaVcH/d4TCmvyrDXCMchlEH6XoLkK04sMyc6jvf0CQ
WfbqXb3c1UJ5p6Axe7/jrrEOP0niiuJ4PvxGR6+rtbto6diKcKy1akP+s1F8GxdU0YtDcvK03Mk4
mn12ADU0LVP+6lNZ5ltFCAYj3CUv0lsrVkphZuOzC6/BbgYA1zs9EBXk1UxOdxwIMae4rXWcwB/E
J0Dl3sLMhX4Zo84AECs6Dw2m+2/LmzYREZLAVWvMPRxvuIcg4kE1hEW1uKFqQhBV+mqhoYhExKKm
7Wa8a/TMfKQRdCPNZKT9wZT36iAdq4bP7jTcvbt+JZ5I1g0sRImCZ52ppXkyvUKome+bDstXz+p9
c2MrDGsXzGX8qlF0YgP7u9JKSroTHvBOi4zmd2rJy9X8TwEyj2i7Ty8yjWhMzjFeMkapV2/+Sf0H
mXZvZYfh96kFZ74aAm+gsy6PH4XHUnmqipixd2oU82xVOmmY9GbqlGRJ85hKIKr5/74ZGy1G2ZUm
+Q0YWF/2uXJLGYcSqo1NZ6uj8bWdcj3QeBxnxt/sVA0PsmSjV6doUV0Z5Pi9abIUTLql1beOFD4Z
9mORHlfCqo87fhfoXHzCFiIzeeLY01XtJro97jZazRnZIEOpLWK62npMlLCROxL8HLFPT+byyoiu
uF8faBb9ruSYquRZai4My5oOLFirrb/C6YdQ6mmGl+3SNwN2wFvlMibhXVcGg1IS1883SlGJmrkS
biH3N2v/963RhDLX9gjYWTYYjLKjIlxA8jFLYvXYx2Cv7rblVGH2ClK7qBWRub4xbLl1PJjhGpsZ
wWK99AGEoZrVt4TTaPAUCflmiC5e8HvK4yW2ITN2IB0IwMVUBY65HCvHi+1ScsSGIQcS8gwe7jYr
vJNWzFC00rK157SCFZPZGnyl2U6fDGGr0I7EE4L1RSNGBcTcpXo9jPqPHL1vUbyrJoBUZdijmZRR
4a3G/YWBNtP/PjfLhgrVqRfrf6aqk5mDZ7MZSZPh+pyZ9pRPRwyzdYCe0vB8hbKabCJkqzHZsK1k
fjGQoabrAZHxIL2Fk4Ma8aOS28tHyqjq4X1dTvgsIwPF/M/3ui4CwnltEFrzuDGgdWYPKZMMuRG4
DZGWolnPKH2niSkXV+HiIne0JNvvrOYY+2+w32kWnzcnYjfL9eLMhLA5M6bXnGjLe3AoDfuY5SRF
r+a58lb8YMc/Av8Xk8bNEz0lgSbYx99GN/f1NXp2F/TyfCgntDdq1/ftjFcglG6pBbNnO1+nfMrO
rNPcSh7pOu0iBIyI7Ev3Nv3iZh3x6qzbbjI+NkuJFjb7dmz091pvm9ANqa6uE6KGzwlMY2pteXLt
RDYJxMHe3TDNi+WObwOShWYi/oTY3uYhWihpHSzI6DnDaqdw48UaS9OKXoe31uLZOYPjk5oGnNuN
uq7aM1Tv0WKdOhzAJSKUPqwzWsUJb0ONe1wvVjqLJ40mpcxHS7yGdp+KvcWaqT2IZ1OzktlohPhP
SLEMzAsDh+8f/wp+OkDO+WbbYH2g4md1rB86OQoSx28hKcZu6lL24GNWC0pmfSsXFOykpGxcYV7c
6dpL6z/Q6FQc7kP6Bb0FvqFyRBGUzsZxtAD8jM9oHzdj8rbRBvbziLKH0J+5gJNsdj+6LG0URTPu
nkkAjNp1v2snChMZXMAeJnN7+SnQKWy6QfEof9G+zgsLSoufPiXpZobXeOxXo1Qsq5TJUKCkCuqw
E+WVjg8PqPbvWNjuLhnMNw6RWnqzhlvRRSFRhmXN1/Wknx2OIXdHnTObzjJBFcdM5ynoDXGAeNnK
Qmj3Bmp5KQyPH0t29xOjEQqKjVEIRcLCUPLtgEAq/cfe36Qngjc6O7zZh5/BlF32xfcLjUu0zZHy
7+UL5xQK1HpHOTCasQa6/xBAiU70pBOcnQBiF8DvNqa5ugBMk07HC17SR8hza7ENYRwLQX+fLoxL
2pc0QEAHMRxXD5Q+Fr8wNSMpU4fmuF33mkaObVy8MyHtcn9Eho3eIxY0KhPgiNUUn5GqlMNmRrG8
JkmWTuhp+VPKWX4lZLgIUrXV/ozmKSdJVOPz9HjZMbvosUECOXoyrS04hFMTlbWZNwDX9KpZkD/B
g7Dw+CQrl+MGdOUoiGjGhRo39Vo1pCWYrugIPvv08h+y7FPvSlFkRRyFn5JSm3PkDUCtAMj1Vr9B
jhY0sawT/Ibd0rbkygqzW31do+xahExST2aVOuedKhgmT/kzQ1DBruucIdVJvvWtI2BmenOQvm+h
aEl05z114SosBi/RnzZPEnBrwz/Cm3oX1iGS5eWRDjY/99xFOZT77y1s+J1O6bvK1EabIKzJ/aQU
9I4GY5q0nj4xaBVeOd94TRyI8/VrcIsCp2bq3HdCoYphKkWBPwaXzhXDIGQHt8RJgaKrGfWv1fht
n/nUx397mn1VEMZfWKYDTvLmCGD6g+sCyCDygMbvuSaYnJydkODYRMzhSMz8YUeZbNETkgOlTEga
KnlibslkPD3C/SApqa5TWhn91zmN2QaLpLtaN8bQSQ12YT7S3pXoLou2tiLxaJZBB8Pl4yx5U26G
Yb91yB/XVjBVqE9jTcM7wv/B8oXPRXAFAoJxZMo6xuAGfCdEoSQsCHMJ1m7tzjOhhBTsf0xsDpN7
VndyehkVauEwWI56uidEgrY4P2QEKb8NsnUhU0Gh+pi4RR2DmFPGKC7KaKoNVvEXCM5rTYePbPnN
cHJ9hABlsnUrrg2A8w4M8w4/Sk4MKe86HUFiDm5m2uW9i3E8JSDVBjDQfzqXjIGIzhlt6LNMvN7B
r2JUZlv9wySyHnTnzkd/MHgaAyz6LPua7pDlGJExpoGaCQ4V8LmWQB68ENOktFz3oSYHE4drGUJN
otbH3uIxVBRJy82Aky0UDu3713ZLHrmxYkQzBjZITeMjC2XulZIKd2IjToFyeMk0NMoQ4h9sJQmi
wPZT/JAXkVgfmlD6fSUxyaqwPITgNNxId/iavjBL8FCZvHotSYyzbyYP0D/cKCZOvQJhCOD2eTHf
eUxAWN+saGVrPA05UNfxaiVHQe9TpB9ptp5j//2OESMYWDhyrtWXMxNkdtZ8h73FRNjywS6WFuES
dWXdJ4BUDYMPLB2/an6GTXZU1CkZREM8SwV49sjmZ65VYB1ERZGAmk1K2E6uyeOgCv2CDAFESDiM
R8L5LgO85zhSoaXFr3jhdcujtns/QiD13Hs1mHOhJUSr8yIkTPl+FSlZL4XIqkfVgfrjHnb1FqnW
/yI8h+XVb8DlsCf7LHMgTM2L9G9QRM7SRA9+JXPZ5r8NYnS6FTbJKt4R2Zlu+4ek7uRjhIAKwa2S
x/g8kXlXTRs+P9XDVKhsNwiD/x8odNyPAvNYwklHIv1xqRZvn/p/2PaBjprTivfeWITFH9jgdjIT
MYg3g4RUuxWd5DWwGH64zzQA95NjDUtyETxByl/s+cbLB1Jf7joEOEjBRjX4aIFxBl5EoFZJUUKI
YdSPJoeFAQLU4GtoEwrWyTv8LHm3JeO8QBV2lUmi1PYWlJxLRSFWhTj6Lz+GnhxW6nRbID7DczR6
n5UjmUOjgsRaWMrpqrTBw+pE+moV8XQ2gG7PG9b2a45I2ZBE/H18HCdh0AYEuRj3BEiELBLHikZe
ELGcCCqGb7fCPIWtPOpxEzXS1nCE2wiGYSA+7sR92t0uTmkIgkVcnATAN0/nSv4iepEQq+ErMkJn
NMXO7Y1Mbh2t4gh1rfluEFuCi/SObgt3sCX+Sq0YDwNDyD/fQYjmveeRxn9UpfnB7eKXByfSt3BL
QxojbKUa5KgSflPfP0UsQJmINCoh6psYLLHGRyxps2QFAg4Z8jzqkbA/W0dM7bHQNvo8C9qGux/9
S5yYAyv3vdgKZ7juafjc5Zmf/1hB4fPecfJWi9rzhPrhvkwRZbgj9VgA/EsYM3qkGV00+9yb7Ekm
YswwwOSMzTP7uKVpFKMWu1asgv7BR0M/MsMLI5G/Ht0l/ePvy6uignspHPfTPDiP7l3Ixp84tk3D
uPQH056S76h3gn431Ls1RSJUN0Jnd4Un5hwdJgORstsOryBZnuFNdK0L4jY3nOb5EWn9hgLURnpa
Rl0lv5Hv7jc+xFSgyVrzCpvFmZpolTAwUrBjUHKh4okxFPX5iVRCOuHRzRZh6QNK/LQKYSrQ4q1l
dPfkpsyk9mS83qO51EF99suCIzZobrhxxnafAU/I6j4fX5iBGoUEm5iaOYN8FXT+bzg4WGxyYaz6
AqvM7+1X8mi9+VIKRxvYe17pHL9Ix4Pe3iMJVjBFqXeuEbsCrPi1H9WXP8WO1LR+tOqlvWD9uB6D
SU0D9OMnd1s0sMovaqAuG6i6BHDI7me0tzrMI6ndPCJuTdVoWuLZWKzhQSPsssHzQEU2QbxYmMcY
LGG6ChM2Z224UO2Y+zmzySp99WuR8RaYqeNs1URYnb4QnhYiE8zzoDT5meedYYQe7zI5c5zFya3w
OFCuQnHg48w5rdmgYDkDsOgd9oSSvLvW1+C13dd5s0ljBdxnXzqlWCYfix1WXzwFelfXJFdMeRt6
Pa/5gUawZvUCdYROBkkGkig0LkcUlHfarK/QYY+iKWRrtuniFdC2SSonujGKNPXNYa2fT9GGaWLX
ONy4jnuEk4ksDb8gzdc3Qt9Vt4DSWIFoZZk3sDYlzeeOfDRMptPVP8AV2ejKT8x2MOLc1bW9Kefe
pos/RjOkqZ/v90v5vnaSaQCR6Uc0UkHJtio4VO/PoY0sPyjfEQj1HIavNd545xzYXW9ACJ2abT/k
3eqfqYHF9H70WKewNIREKpsTBaTwm08DWg9xlJRq5nACGpSD+MEV20k878qJE+gayS3lzNMS0VXd
IcsSRrr6KB7/ymQ6qtXKrmypVwQQHxqn/agt/nDMEoThx+0d73QjAoYz1TwCoTbw41OcW6ohNoAe
PqIH7D/t6ekr9Otg5aV3AlftmMQsxjBiqNbJqH/aaU0CK81Efg4ZrJs4K2KeN+rZjXdKb5QIGc0r
h5qN6rQs6b3G5jtw4MDO9yIfYLgKdM6eUAWE7VQS3JZoeE0FhJBUu/VBnwkykH35lr9PRr4a7Njl
hh5j7orWMZnQ9vBSmEh/yz8iCXg8aYGGwEfFYbXpqGUU+x/HodJn8u2l9lY0HXwVGVhM0R2rhNfC
Q7dihNYZ5dpDSVZDk4z28iZqCt/VfXkLnS1AFJw+C8pg+Lvw7d4q9rVbmQNQ3NEwdH4qQAoCACLW
cdM2ljywu19VzMcJNMNjRmooQPLVulcI856THEu0GVX+w5hp3sO3hMfyIxD7FIj1S/uCrwrRu7iR
L3P2ecKmxsK63ScGWK6yjq48LLjPbPLkBujChOSfhKuaujEpJ6O/q1SHaL9t0hTIxG1O2+hNUxgH
JOktyh2ymVWH4WBRJl2KhalKM21+eGQKGMHgLTaEWpNkpHDubjb4j9HZgniJvg3Wogw1QGjAXXJW
OT1ab9oFgVDQZLdUQokuVsPqtiXfQDVUhviXafXX/U036JEdwpukzagw0bDNK9oNHIfOSxNwKtY3
Q9ysPTv0W6qi3E2dvzhygp+uZsF+pHoqIaGGsGD1M1KTlDdZxl1NsePJYl5fNJhb0PeKjbZhZpUH
JPJ+cLboVoTgJx1/JC+rb+9UQx9yFWvTkdV86uWhASnV8l/461W+yj+FkLGkQ4+cqsoqYl3T25N0
S947tZFmD5Nj9YOtFuxFlTiUy8gLbDLF30ffaCmg9SHJN6wRmzQoCFupzU//RhXO0tE2mEq24EPQ
Wmy5lKlHyO4Lh7uqfrB/8fgII4es2dl/EIg6i7o5+/Q5ChziwVYOEDC8U7GnzBFek54/VS6Q8qP/
TSq9CY9lyGng2rtxXL+lwltBaE75zDRc4OyLs8DE15wtHI8t6VbSecBhD0U1/q95yMsyCnflfjoK
YMQ5lBa73rQ6CuL3Y+gDier+IA6NpB+DOXd5iDw5wxORYeuxsWpdxugCjYxWe/rX35GqGbX04epj
ta6rex3W7FGAyPWW1Jdtd6gCHFIonAiXOZ9LXr/aVgzdP5og8MppsPnWvt25G7Q45y/k5q7EWXuu
cWY6yomkWzptJUpxHyHuRs1QWBePPBujIXU5n140yScYZ7Eq/1cqv/6JPlBQVpmcrw7rbeI4p3oN
e0XybrcolbvTAYFoCKojMYGURGF2l8NdQfEsWLNysqoWSrSuWLc0SFrsK5T0yhigq9lyrt18J1pF
So1as5dtY1C2zEEHGHJo4JATVMlEZyRQpgjdtB45KVSWYhgy393OF61DpsNL6B2LcNl01JoGI8am
dz0GrNiBpiIVZsU6BLyQs1PDHAn1GcAdthHIYi0//PJX+nVQar0MpWWgurgPlGJEbGVC190PHuW8
awLN6WC9VCSNdfoHHDU9/eeB3PbtWnSdMxkxDBY9OnafbgmM2eGqnfs73jM4Om7323t8m9yUiDgU
W6oA6/dfGH6KPJONZEH7M2eU188sUfCMC8K07BCfuFprvAF7Rx7WBZF7sL4QTZUk3fM+1PCdd7q6
RZD/y/jMd46Lg6i2WCMlMS8rIKlKvrWC2TV9GXOqLDu3+u1PXEhFeB11LXICuDL0txxN3KxbacHj
0qlMsF67dhey8vSm7l7uL/9u1y0ieAE35gKIFzgv2Jj2OJ1GBAgeKrf2+bmBOGqPVkPpGWpWcYkc
X3bJJdNv92OBrl8IfLJuvWm86Zc/Bi98QHXw/HnfVkN+BxVDYJNUHMfLLFN0X6q8fMxcjnUw7Nls
51Ijt9nYNH07ofH8RWZsO/GZGnlD1hJAHeK4gbj0xW0/tbeN9EVYMH7o7sqmd2L4jlg7wujNWTNm
j/M4nRgQ8cPTx/FpFaCAiUbLwCIPHAeftB0C57PWG6zeEDoyonyByDLy2aP0zum6MTGj3snlYRQc
e8vOmieLFkZoDmXx6l2a4yAVJi6PCA1yUEgfPlqLnmo1Xwx1fWI+Tcc4BSSUVS5ORCu1NqM20yuS
aIVqz6UHW1ncNe6caI3NZhmhZi7T5sFOQdylWNMA58+vrWSAePF86uTphyllVUgtrg4BTLmRfQyG
x/+lpuWtb4HnH96/8OxbOoV3CMLWR+QNxEbYootwBt69hgOP7v4Y3OdAayCRksx9UITLIzbHf+MS
gu49XOlCsBQE8fQ3C56eT9jJx905/vXoLy0GaZCZNeGjg37kGlkVcGe932qHXX4YssTNvtm2tEZ8
Is3ODN2N7gvEsb2Cjf2tFNlFks4cAuljnausKUJZUsgZ/Sc/abM9XbaX43HtgPaSXzLz8LwNAcGx
WTu5llIYskiiVgYl6ZWGGvuBtd4P0bEQipKj3S3B2D+u/TDcjcTvpxvgyBXjV6LZxLuk9NW7asdw
EmVPzYAXanYLWDDRG4d1f037dJlNKRVQncXT0bHw+kMznNcI81oz4TNGzvNWmi36I7gey1JHx6ai
O5Y/WGQs30MZK1l32P/62AF7RJvnngJX7aZMD4qEhQJKfaBLuzulz6S8t624/GkkqsVZZQT8MRVM
n28Bzp8HOyjXCk7Z+fT1Ak2kkJrWx8M/BtcuFPM7zNy+fjhsPEyg/+csJQwJj42kJkxJSfMVCgKs
eEMDYN8zWZcHqOecljxUQbZBvbQye0P0Vsvb/k8V6V/vXFQlYIeS6kF/KD5eWPfGrVUgB2x0e9Ql
I1rNK0w7EYrRvyhPcJuWTvw3M5CnsbEOho6NqDb5ZHvx3IwrVfio1u/4stWIWuZsusMTgHy3mRz3
9bryCbV7JprDqe6Pw232M+tpl2NDplUM1o/O5OQUmJVkRRrkKHakKCNQGNOsFIT9prZshA+OrRQK
/YLVcFsNMWr/zJy68n2IP+YCw7l2EAqTzcrEjDoCC7OPBo1OUtFMmHJaHCUAT8BM5OAJS3U1dH9X
eruvidUfN9KniJmiO4lmeiqz7vth3h0VQq7T0JVav2KEq1kD9DFhGTI5ykQ2jcBzfediOML+tfSw
BW6uygg3s0eR7CwLZ/wAyVrayCjzY27WWOoiLtYE0lT/YhfD3o4Soe4g6uD4pfz6CmIbuRMlnANH
sFCJWL6APJZ9vsv2rQFnZ7sFel+4foyq/LsJYUFO5T38HK8KfRnpCBNBdMQ5qMeUCK0c6DX/Qvpg
mEXEqRtlfZMEp1oAju7tzUnnNEceJloNkcJX49mxXyVNVAaLDTr7zfEn3IFOTcLIQsvaLZOUF+Eq
/36kcmwlrAviyP189YmRNa6Oygou3li/1UpkP9lS0vMhamK23RruZGoGfhgRGFSa2aACwEoV5c+F
xsAGjvUstiGbAIdoygFWHzs7bqQapaFOtS4vSfiMMOKSLUi4iolB+/poi7W0UnQRKeXdyoaetgAm
bCJVxp6sHJjL1Z2LvgfVO4Rq8Hn9/32+05486EtSEZur7AzOwKmG08mQ6Hja3LDTeQByvYRjY3lb
9wyjf8iEdraEWWu9W+LIU1Uu83AojYc5wa+N8rG6A7g4YHg60UdftomUzcYR70O4A4SJFD0RBnoh
oH/OnFYsXsN6aWa6BkJNHt0KHIrqCy7fRj/AWOzfPUwlAgPjP69UyHX2x/huwpsEiNvimOmLOiDa
QJYpnC6jJrmMaYnreBgk2mZiP7CnTdOqdGZfLlqF0djv1g2NY6/XjB1tq3kb7eCMAUcOfOulnsk8
6AnMhabDW0zSsWUKLWdMcO/RtXTs+52THMEX5tNsH+P8mVqkLgAycGAsAgiZoCXTK91F7HXWi6pV
YOUr529IxB/WMW6nMYy7jXRdTAr3r5FedP2zfsG5MXA65mtFwRwB29SLrds/iEtQstTViOCZyeRR
eN3Vpgsk+T1UFYbked7p+OILxkQIKX8rgx4GKfj5v3FaFWmoRRGR0Ib9VWeszIKGdY8LttvxnP0C
R48qc6i3bhXeO6Uwt7q97vcB8DQjp+0kMClQCOt5FCLlE7iwQB/uXsJziLvmjdjH2/obcO2F8XJC
qXdhdYk2EdFt5lZK5iWiessNasukKdWGpLgbF1WE+qqvTCXIuUGmMR+vBdSKGtxvMEQT8NGULhna
eoYxT7M0LLXqchY4x1SWNKxEqPA8u/uB0RvmzQs0q0sNszC/Bv5uv4CfFOtz1VbcWxkqXDgGl2hY
bz1l3qIXoT6N80ZZY+Q0HVic/PgY8MFj78HTwDbu7P9zOeW8w85PN5DxgF7sExexIFxBJ1ECE7HB
CH9kcuwq58dc9w4OvKXE0BfHXLT4D695F19NKqNzSqev/wVAAHJjYlo21SUyPLz68kGdTVy1qYdq
VB5bV1c4sGaXw+k7LQ8Of0sTtBWXrLQv4lWtJBdIUWFMxWKhjMi9D/8dagi1Ek2zdeGqlH+5Mnb/
ZDbI73QR0jgwjPUtuFux+ZltPMvcsWgsxJaaMu35wBBjWtNwoUrdgyhXAjQq425mPRz4XbTcgOVl
KaUDJvpCGP4740O1kE0q+WL9cnQWk/dXYM0+5M/BmNIFAt0OGcmvsJXRGDdcdEW1R0UYH4EkK4UE
hyxdVMHaHsTh7Kauw8CJsHNR07J3LmH/FE+OQ2xJLGfAS9IaPVP72bo1TgM8OwDSxRyIkH1dWeGD
7KKz3tfQkhHPoj5UKlrDTpAIMTH1tluYJVBr693pQbqs3G8zDIlt1UXiOtYx88wQrdvAYI1PaBfP
asHuhV1X4x7G3LPVsJPentxH378M1S0izZ8o8lpxn53jWrzKt59t6RTgVHAxhsTy5eULotCgLZ+R
Vn0BCYv6d1sp9LMNz97wqdaZFosW21T/JJqEE7LJ+E6szIQz6zLt86qWC95r98MUfzKauyDmq7j/
HjDrM4ZKfYePtbwLp5Ggy1q1liSaEufCBpjCdVdOrTPHJaU6A/7sUmusX69xZ7ASQqtjnHCxIvV1
P5oh7zljbq6KdBaU5q8Ot0a1SOLgg0MxjitUzlKwk54I3TLUOUaEo9hLpMtkk0brK37g5BiywyQJ
RBHntsgD41FPl8yrlzRh2k28v5Jjm0RyAitfuXy97/BOvlvs55+YMDDKrLzNuIhm3RX2T0CqsgOj
Jk32eU60bxxUdGY1TOcPUfh7RHtLL+MUjWKOh5G37q9LWiLkN+HmYSuhaVGhcHZAisdEvuygF9r8
LwG6rfwFHOhAKXo9ps6siNjtOs0warCzgHdjxEen6YIp3IOLWbOrtZe4dO1X6qEmgR91s4rYBYSh
5TMRUXca+CqKQvz7niPJHTf3kC7waH34klZoQOVy6kH+R3whMM3/nnh/1mvWFQjI92x62b2UDVLf
bur5M/otByYLNUrznntOX0+DrZpzxNF98suIMUN194B8wqJaUWmJujPUZDiYnh4oniGRzvK0aLiO
F4BSsipLftMQTvA5rGafUW/HFUYDEz398ib2EHtCXvv3OC1w0uxmmASV1/lRfmgfqpk3saXqVCLT
TwvEhIA3Er+VYYDOByoF7EoI/oUHZiGywo3SAWmbk6Zwdjrz5eLf22k4/gSjHLwR0Hq5lzGM6CRv
uX4iH9l0MrY/04rz+dgvU815riQvlHG9ZalDY+80up4IAekJ45dEovXhKTc7xHRm+ha1xTLlxas4
/4WMFr9EpZiLrJ3ghFsZa0soZuk6ZJso1/S4HckAAZSAHn0u4IMZoIP8cYMlIN+3U+ntreGGX1mn
GvL9uElgMO0oqDiRyu5dkES8rM93EeJ7GV8vOr4E1UwShV4tJuYdo/x4pN2lxV7WDOylJjZJbTdw
pn+EQEraGdLSn76NOqAC0V7mpAAHBw7+e/oIpayZhW9r/TfXcEN7o/XXTgCx75ZyxvZJXIaVFNRn
I2c/lOGlwGA4wh3+gCsmHCk+SgqdeZcmzzHQSvTXLs6UoxUz22ZSFiUB1cMZmEKWTtrIRK09Wqjt
h889L6ODVPC60gYPB3neN9uv8gVOLiSb4XUc7M4GML3OOPz4mlSuzdt9CxBOmn9cTg0lqpSmce8y
cfnuRrInZEWgrafkZVGRsI8VQ6NiJp1NbwM7MP9vbY2MPLJ1ZFYBG7rNy5/lg4rE9apr1YNUEDJd
VNMJkE49Qw+OgO9FJqufXnqeegm9rR2KcmizQi1fmXGRKn/nyVB5sQFyPEVV/4y+aELin1Q+XY1C
HsC5ORIbj+FcGRHD9Cj4Wf0LgVDg1AudBP3lBf3gsIYc9NLOPDIyQrsPyRGmSXTXLhPotzrPiu/S
JDryXvgx5Fh0YyNthiYSEeQVmw3TtopFxG3m06lKWzwjS0ZI1WmjXU+yfT4dcb/F0ppa7sMgk+Ce
T9YQu+AjKm2YunSGCkT6zJVLZgLa/tP7i2FjzjOaYZynkxSlD5LTgDW343UyN81AhgFkRpaw2JR5
T7DbV9QP05LpUx9r0SpgEAsjCR+2mV4L0BpLG4/YHnZUnPc5rucYjTEo/GZ9ZCScLtA2/seVMTQM
jj64s+H7xQQm5vFoIw1HVOdveqiu9wJSaf42TeKFt7FU5BPYJSyWP2G9NnT3yAo9fQ6tFet1B85y
HynJEWQJBVMdhxAc3+E5dNSd9j6YjSzmbEd3+S4PWkv19iPway0ZyjzroqGqkYEApjrtoKCVFfKx
fNJTZ+nbU2AH4k1+F8t/UDZLTjBQWrn0cO+2OL//sqL0oBf09xRm3JfuWXaH3nkXsdFoXmQflGSg
PEYB0ied+4IuUlEvOAym0CLv6VEqoapEBH+dNcTV3P4WyEEEXS8fWlarRm/2foJuXDAIXet4f0XV
8AJ1XuCakRJwSoQ7Q9uNjFgBgy5Tzj1BjKtXUE2S8kUAG2h8rwJi6P+td2SKzgbEsjol2uFLObfs
YZWLHV3OFCZtrY21kr94W+uGglmUHzVt9OYJXkfGiANmUcObX19W4FADadoJJKAG00DInXVG6DWs
lWNw/upmcbuDGpCQas0DdXetOAhr6opDiTVpYNqUV0LlXvhUuV7kda+HjTmA7tJ64H9YOCWRRNov
lF/IlbQI6/tKSU3qoRW46XmmJBLnQWn9z0Dal94OQlsluqDDr9trSr1G3coJt8GSLQ3lvrBnraPY
akh4ejTP1XLq6eVVUL1SpNM9bucLqU4YkIP2sI0+S4YG2VLFzTU1h72f1csLl8l8L2nE+hgUI/OB
4OwMN4NbkmuqchUKCQl5lF0JSY+PxT7PXH8tl/cgNK6Gtrhu+gSefHn9pL7Muh26qfepsaULqclp
PhNtTR53NMMTJeiUql4fnpn+gWFJ4F/KEUjZgVD2rYOn7NW/lrEF9dSphaKyiNGj9nsK6nzsrAjR
EAE6QDCij3RAU2vPl9EeHTqaVrSy68OhXv/F1M6LeDo8hi5lm7r284iGsd56G5dFEgrlCD5277OW
iPpIsD1TxKXCdUjqs5w2to+yRvpdFPCbIcx1aRIPTSKH7hGn1lxDjQQrsFq9SuREtpxNU+KaRwld
NVkPzgD9GZh6zLfv6rrocjzIvoWmA2lwkDz56w/sOw/apxnOF6++ndlyDHDdVzxKhknmCf3+8wOw
CPmwXPMTm5MZ5ya/ZIYliXus6A9AiAXTK70hC1OZCW8MFDPePOLB2ZOQylXqPdObkgZEKCOJUWt8
L6zE+5FOFWK7zURt+g9+M4gcRIWRU5thB7iUkkkivHT9NfKyvO8X9D8r/GEAdaNs6Ux8v1rESf0x
5lxCSQRVNF7Vs8rwiEJWL1W5YIusZ2JNakkkhaHZSuvPpFUz2IGjzVPf6zTI4WpiEUtq81EBmuuW
6SZioQgtxIMnueGgWjFAFEL2zcfSQKsnDXFV0u91bYOEoP1jqgTAhvxig07fnvDWn0P/rvgaqsuJ
TEWboMxuYtWViXakFuCbhcBUpOGDnBXSx4SzXi5m3C5HhQoZDoeN18dMP/7vfz6h32DCy/3FMQOg
weW5F5+nPGgqMFf45PTBqPysbv1QlrLZMEH8jjdYi3uMRfchBz47ZSLnwoExLtKY3cogrcGJqB69
Vel3sHVPV/KdPXQF9Us8yOMYmjuSZp+Az58tRtC4NkfFkrKwk3waJA+3cfJ/bGpN5yBvVgH3go1l
JgbPs/oUc0zzIrLFmSrrMF3Pn+ryZQaGhSUFUKxQ4CD8bQYdfO2OHQUqMF+iiMYvB6Op+b5FrO9f
/fOhcm9VqItUzduhRU7AhTBbKttJCgm3lNHaFDfaUcA89SFWvFBMP5hvgy/k3Eg72NjvlXuIFqvt
wax6pat1gseE5Um1EtlqZ9QMrfnI7XouUTASCk1L94+F1VgBTSRiI9QoTKU0fSTP7R6CDMVc8osd
LLyiptU51UyMOovyo24WvLnetAMg8h7fkVg1iyuwVqIpxfjzdX7TWhamDPvqFIv6kcNV9esKgTbK
8D+d8zJot+wLXQQRKhmD0TKx6w5mJJVeKxph61MRmVLDohqb8IUG7sYXxFqHAxgIzaEJYwpjg5fJ
9zvBQ70lgfKl1WvpVxrz/xPtQBT8teUeLesJk6zHtgagNV2TpQkNrf79N7cnM+dzHvMU977BY9+K
MFZCuK8ErbY9YAFjTn+wpPPNUQ3nknEwfTf4ANiI6bDigKlzpe5UlPb2pvr4CRMTswIC48QnPcCe
pbCbsG36I/6GFJ+0FOdoFKaOPZyHuIOu/DY2lOvOhbXPjZumuDLFFBCNMUcuz26gy6rQB2XoZQG7
kFlR/gHhSu0tm7SMDCFEjP+owQf3GALnfu4oAAkakOZfcjBAbAEqOdFC3DCdW0L6SgMdJ171lq6F
y4Km8HJ6x+Rj3zk03j9kb1NzneODRbZss3QMQu4rhxvO880/qpNsesBB9o9w/qSxOt33RXHAw8B1
97NAu6exXVLmywNsQNXJeF1H1WGKBRGv9YwjfilSd31Kq+eX4hbqpKcz0a9p5j5TQvrtYaXvyaEN
+IrotV2Z7bhcA71+6o5RW4ivwrab02Z9hUEqeiQgPZBX3qpRRjYGbhqkwDKsuA1CIKwP78SBs0XK
gj+MkN4nt99TCcWQJsLSR61f3M8I36xbHr7+NiHmfeiAbmhd5yslhghOVtOshEL87FGS0bxLip1q
4qR5PtW2eHg8QKoIeLjVlN2S9R0Djx1fHHW485nKuwOiHZ5ETKSExe43faLLGMRA7byhdy8JFD7P
HgWGYQyPm/vEm/ZaGUSe+WfZMi06FYTivfa0KRGTMOg6u5hGmcN3kxpr0Nw7Fu73aEQOY1etfSNR
PFxkPsHbtDMsLOoL2/0hAouA/1cXPpJbi4VpQoY0bOCaonM7vpbOGO4s2D+WXeh2Twq3x5Ge1O9R
zczcHG6f+IxEE55o8pQ12lLDW/S4gbbsHuO7ABIj6R+iUJFSTftpsheOOr01Wf8/hfP8s6EbG2y9
PwlMg3TjOE6kIud1AZ0dU4pYiQi7EMsdeFy5jSgaQ7mzWTilt+BZup2CoS310WxsIv7c5Un8auFt
qX+KTQiKmtjY+fy+XVwSId/hMrKXSNzMxOu6lmUlpXsHxxJIgf9b0LCkib1yqY2iG35nN3MCAbj/
AX1J36PL+mWmEAva+5qXawRvNYWH4+pFxMg7vEhJ/xjNv+7L1Om4E+SPxGBak/xniUJNIMSOWK4x
IoQqD+PX3AlYmD9Rtj8jluOAGS6ji/Y6ZWe5OmGaJidSt4l1SwcxNUkVZYdxNuLViua4iBzuDSbI
6OTn2UGnJbq5yDadAgCJ7mZO0OMDCgRpyNWD6gdHYHGQlQLU9x+Da/ekpE+sfk1VdBVFQ/WlUD6C
u2FQRxX6vmvI9vsmr5o4+ZpSypCz8fYWzDxtuA5Uh6uR1lLOum7BkxHb4T2b9mQUQHBYSAM0/lt2
AS8e1hotNJMf2U4udTNhMix/iTfHNOCFdoPOOUzrw/soVQovJmxsmZzxE+yyI4ieejKW8lSSVyT9
4GIxeMITng6o5kJmfpTrIaa52FwqscIMWtxGucUVOWjx6Z/Gmt/fSJ/XUU/FVli8iVhvmpi2DybI
y26G39vgngdwk0u7XZooYb2C3gozaTIvJCitU69cX/ZdGoznZwmjLUkPBPVezpfZzFJfc71SZkno
K2l9V25Tibza1GpjhEqAN1/sLJkM5vh+158ZblPP82pv66EcRSXyFD3BrcnMF/MM8TF9hrg4US03
yipiNEYQdIrNBe4ymlqUyN082qtzXM+tr2ROR0v8xBXxpjVQ1H9M5rPMpAn85JU9p3M/O6ykfYKK
KWhbbgZqKRw1L0EEgvGD9n4AyC2WE8IZcW6G6xT8uKtO3ixsjpIzhEqzS8Ydg9FMXdk8x+sPfSqN
rIkQiNiGoipK3vhxC3En2T7lYfL7vCZglHMcB4h6Ly5gzsh24bRn8bicX9KUF3GGSzYPlMjiqjE+
txmov/bSJO9n1YkslH8mil9zZOUY3i7ad4kxXSR2J2HD/V0beZNg0aKCaWDum7ki47igjD+IFot8
Su7kmZMJYgjaAaexRkVD6ZXUlFSZZuCOcf2u55hnqYa2TZt1B17lhjA+XKPqFRZc/0NAdUJoyG1z
ULlzNvaOexaPVVMYTKu8PPrHfIp0DauaX8f/s5b0TJcIJw69ZjArDVRhFsTjqVqQdqXu5+RObZCv
jZMzqHzX7c/GOWlnT6Q7UfP8C72EZ2yKgINHkLEHdgT5g6dqwg6O9fw2OrvPS/a7AmkMuY4lkdlU
gkVvoDLohCHe/aXszVVfRq2vCtFqNfX/BZcg1Xs1uYVV45d8pQoB3g8KhtYddxNfdxiEGnu/wckQ
J2oe0VlcvlSlisKTYnMnD4Zh0ZbAcjqnLd8WMKXfvjnD/7C2xLyUl4OrUuGSvFuyjXGO4EFoXCqy
2Yemf43GOONg7n0Ofz3fNMFinCtB+YK9umf/Ifdh4DsszoJSYq3i/1ZMaaROegALxEnCPcSkZPXR
Ww0pURjzWl3EXolm4pRDUaJT5fzw4XJ75QKifAU3Pds426K0oR5X7zTx5+HUt/WQ1EuoVi813EOx
pPsxq6UHOI5fk+SVlYBldkAt+3lzizz4ScHjNdm0S40E4uX9eSzkOTpMsus6lERETWzbk2mtVDAE
IMfOm83ao36D3OuRtGDnuXrd2L5YODYrilmhJ4S03RdJ44Y/ll6fv6JMqt1xBRM38z7ysKXpymyU
JnfMJNG4MkjOamIvbqRNwVUAo7kSYeqkF96yCzQmv2NLJWcXINawQnQ+rD8D5tp/xRqG7CyUFfJo
Nx22smzY3axGe7ACBM8h+9rj4bIzF7l4SswgbZRGgcRCsyTd2OsCmGj1LFFIBEbShHeRdTG09fE2
ZbFXnUmK2W1ETHjgnaC3YnydttGFGC4UzahROTkpzyjiCiNsCbnWbl8SFtuoHkGNkVokPP0eRjG9
Q9txLmLT/vwnl5/65BBXrvk11PGLJQTQ+nNPFnDcVNFOH/rkHo1lhHmY5a8E3jyuLSlfUQF7ikJl
0Haekgs42Wl1AHjhqfZqiJOUAM/eCI/QXOzB8Qaf6vxbaPgz8UyXG7JqAI7S2dHzh7AOqSyDp3DQ
ZaPUT6rW3NUgppyJiNiGUOvwlfnpO/o+SEl+qatybMR7YJpQ7hT3uBQe1vBq+bN8XYTNT8OTVgsr
jBVVbJJgagR3p7GLkwjIaeRcwWUxcgfY+NOT2t9IL8HsZFH3FMMld66TQyCpSJmWFjJiNalkM0JV
Utjt9Dia5oFHIR/bv5/Z/Z1RyRCNfIPqFLaPGUzjyYbZc6fh0YQChhbZjfskONlZEvbXpPk0z3Rt
bgGuoA9LMrpVG84hs8i2yrnMuvhyqwDTwmS/REC0UQMTMZOOBlNRnn4mGswEHiwOZvJ6U+2dcP21
l6tm3tJ9c+FDpJjVjhsffmZLVdJdYFOod0usR4mz7BUCg8RTmmd+pu4zjEoOY1IAIdEAOWIHdZ/f
ISeBOJpZetvXbpQWR0Yso+dHFYYKTB0mZT0mfpEN97kWYB8U5kVkEt3nsuv+mNI9FVWObue6jnRu
LcHg7R3SUnVI1AAnpucC4YvnZiO6/ASZ+qNL4mLrKbtiHcWKmjDWwMCqJ/wqZDoArYFbeLHgWRxb
7oE0mnEfideX4KifdALlJCrXJqMad7pm4TzfAyvmqFxg+1B+kgvk6i2eKcKs2tpnMoxcag9u4Fx+
Yrh4kS1NJ3SS10UJSU/YrRj8r3QxpKacx1cZjPRKnIAS5GA63q9h3pbKlfb2mXl8Ba0bGC30Nssl
fTUe9ITDoBwr+ih0HfgEfejAZvcePvF22C6kdYP7JD/xqLMJeFeVFkfuG+yNM4LF1I3AXPadw/k2
guyRT8DCdp+Qw/zssckWRP7N5YWp6NFQaRFBz5Agu/VyTn2KAQvQlsXxM86pjHxATBL3vGzdqD46
bq5rXCP7vsD7NW9vUGDeCvpFwIr3aCGHROd/XQxuGvqwoCVtteJjRpvk7ZL7Q0v8A9oMdA1pu1To
YI+HxabuaUXzAvWxafWUsS3Vu1RxEaknptOI871wjp0CbjfoITQWJ+GQju7+CD2L7/b1sxpCukGN
JyBu7CLcaJieBE8L1/G+5b2T1ANmXGyOkZk11UEYdHmGv1N/dWFMNHZgiKe0xWRjcoL5vpMrKZv5
e802/FEoTb8cjGfkis0CTuyQC/ltXhfBFlu5z70naC/lySNAolOi4v6eHeTL3BunYZ4w3zmzUCfp
o74GlTTMosdyDyKYRPLwixWjqPChGzKe4aJ6oDUEWw4oY3CpRTYohbBaaw1DANkIieRApKg0Ze4a
+ea/2NPGoR+jfw7mFGuzlv6GBnnWltOBADEZkplCY2Iw5EIsOI8NOOydgCDAub5nlXVttieP96rX
8mxB2brM2MHSF2Rfti1kS0zNq757TguRQ3nXISwYK6CDHKPxdj3iakkeniIIhNZQXD5HSImNzA9V
r9DZJyVSEO826LyrxrutppPzkubK1eZ7pyTY8AEBHEY/yC+gEmDhzG9rAbmaLP3ASyQetj0S8Uk9
/3mEQV55P+FcnoQObIzMdVm67XvyznmOSVrZS6Xq6EJmMvgtj9g8022vWwMfU6UK8t3yYXfETWpn
Te/DENn8VrtEaaY8GaNiNxqtx77yb9noscNAHDVuPO/9UQdOVHxftbN4PYSCNO0QFQJMWNuYStrb
qXqsYJqz+XChL5tCOQmMN7DM3oSloMskpM2dGcE4yq8u+OPlPVovtgPKhOug03gZ/pHmLpLj5J/H
DCfQqHFK9I8ibx7MkXQro3+5S6url2EmtFf57zqfpNo611DTjLrZ67nhWL33rGt+CcJnBjR3RzYy
AOnWl61K/fau9aiSvS7V12bOVXo/h4dE8ZyphbrMgEbGUb58D+oGhmQbCRi8FfVthR13znfEWhN4
wsrqSfQTaFZNqxkmFFys8QTR5J3ZHKp1Swie3fp24+xyZYNL4gqGFMGsWzhEdpdzzU0DIvGF+p4V
wHBLUYFzBVl6SK6DSSWcKK7la7P7Pm8D6oPPayWXh/r7IB8w8ForW9zClXWwEF3QeLN38FDBksDU
yx9j9bvulygd+/x7hcqmT4+OOFeYxLUs8kqyIYAumQMM+sI1eMzAgkIJy/pHoxzPaQ7nR+HwVxhG
j5gtzrsDHEL5Vpt+wLFh7TpEKb1fekrCE9S856d8hTEzrnUkI7ekcQTUx73kkT5vCHaanaPF5mkN
MY5GqleREEoQzxbd8fJ4XGoJ+yL5Eflg/mmA1cEklVW11+7SCpWzVgGK2YliNcjO6fpj89MXOjsA
gH4TJEiQyVsZyorytv4RYuqJ8w6CLCad7HkyKLgxRTiMtUGgqL1YJ6mUvE7Aa7ebukETnm2RUfd2
kqdeJ7zJE7PpiEhGyF9dMuAtz5/lPBjoNpYfyZqmX7thZiHqzNhJh9CUTRObkEWpBMAQmEEoBRZ9
bN09KNOuSbZDC3R8I8QmW/qOUr8al561gZt8THYAz2Mz5dNJEy+Ofp25BfmJ81fTONenaHR+FZ0M
+hK1WrFQ55+m+M3dcpV45dxaJN7oIc/Zp+/nY1+E5NQIeB5K27fIj8CY5Jv5gJFgzlGtcwwlZFRG
3TR8K0ulpzVEnajuEzcI/3IGFpZ+iZFcSmprV+WiUWlRNz9+UhRnq+AYpGcghLW/B/bYXkAtfw3u
+lKxlk+i5yVRfBojqwDDT7IdGnyEBryEYZdNn5twnlT6uKsIXGacDTjd4F217WCjuMnPJjwBuu1M
qNJFaAZqQpV9bT6h8N4gkWpSD6gAi4q28GOC8w8TdAEzK3iXqiGWU3/IYXG2fgNeWM5f5kBXSyyo
K6QKzJzC3O4Q9QomOyk5SarDzDKS7rvuK1/KeMf7yk+GbgmTWQK8sqbQnR6ZkisWul8ejA+vGUCC
pLbvozwY4KY4p1mZitfFdZ5zg1j3r5n0N6zjvNDJA2lX9vKx0vrfGYL5qQhroezxF0QMvgFepm0w
Dve6bAP4GPusDPtFsdkwsua10Vi+PzjaAol5TMUpwj5a7l0YGLtNZE/oLRMHwJKjlU/M3gtMXPqP
mCcU27vWWGV2/A5taOjs80/1RIK+8iM9YkxexSbU36E5cOugdMZScAZiMhuYON9pBK29r6aBnYu8
Ln2l4kXtaV8H6Zos4lRTgY8eRwKxNkCw3Gga288EQbj8aSfKbkOC9wCY4DJLKrYbM2IzVJE6hWZf
C9YzrDvuHsiahNZto2hq2gF6hfGUhPTjem2m1VuVGFwxjTjOC4xnSXBAOqJHwWsTRXPRdW5r+3VN
b0qlVekglkfZes6804Y4XyVNJxrNKxooTaP1rlS693aW+zNf8wiaTYg208dwdEJx0CH4jBg6tCz2
bCrNP5WcUU2YOx+Z5WJy8UeXs91xXnaEtE+NhwfT6gRgvn8+f+4KxqLVDB4bxNNBV1j3zu4siw6x
x4bHvnufEUL7X2byjSXUhpVXjJbOiqrejiV/CBSkwgDfy5PsS8mIVoZu/WHGlNor+8tGjVXM3lZd
/+3c0oF2U39wT8xsHf3A4YtXr4sKioDscHVib2jVs474sQPviU2hHfGUZ0mbhA8Vl2hz/UQIR9aU
B/bsCWP06PrUaFCcbTQd9/uXPq2b0SLXD6pZgUiEyC2EiM7i+owjZrsxNhLcwmJdo7HAJWws2Hjd
Vy+agdoobj5cNqZJ70zzCkn69IqSKbEyLyfk2gSg4lwgrfgXF3DWplgvcT0b68FU2MjWXP9fLBuI
d39MtHicx7wdL4jmHdbAYdeK1KnwW/cyBHtbdRePbFDEUv6+ocgKLem6L/stvHJPjZY9OEl4hnNl
ufB2nQf7vUW19bgfdozProrPedf9KbvC1y9EKdUtWrNlymAPv6+KvlOz3tCV0Hubfl3Kdl/eqHqK
hQOPrOstgpWfOqCk05Qkw/es2OLM0gM6uL2JPHAutuU26x9Tl9Pl80pw6aBe6fqBli/dY8/v6LtS
An/Nwv5HdYo4KDYEIcTiv2UCfc9EUbR7Q7zcC6mVegNwGKDp7ji2E7vhmAryjpm8UIK4VcIXFuTg
V1j+PWN+mIe/YgCJetmcMG2VrouuRbdPIBycn0mVpSuFTF+Pd0yhc2Bvz0kNvNflvwgSesSlJ1mA
RXcKaa0gN1tvmWWPXdDBb8irD2x1aMy2QVw2TOZgM1nV6jsdL7utcYYBKMC2cUlW/gx3sh7siFgu
jFJQAP6ukWP9qDvqBm9pOWvBntCYc5jJOLTc2bgezVSXAuaIyprt3FELFw8D2QVRDzys4iOQ1AAX
gVkhOUGx5XfNg4iU7CU8g5Ijjw1B3CGzXwWv7UD3Wd1cY2WulbRuoxvZaJ2qqj3NbBXAvKvpyA5i
mW3uq+EnvhQUAfh1ixKK35a2qPOfWJRvyi20BSVYArCunwu19ZzrKeve3lrODl5QalGVFwSiy8/c
sGMz4JV6QnYGKK/mxK0MVw5To5xKk9fJW2WeuE9QgIXNC6qyZlxDWaM6fKSrhMANFbb3wZHpYIfP
qg+J2kVc1z7JlD5ozkmSQMo5i52noxuFIUVhZs8+HJ7frzhYqgFNCFU9N55R/CF7m0f/+ua4dEZH
/cSUeiu22wd8heDEDI1+g6p6xsp83iapG3dEUo7wQ91KFdKOqdeYxaevGU+PlBhfU8bEeP3uDXUz
ogwW6hdxTWyOAqtxMNJM8OcO1uI1dAqlooTu3UqkvT+wrMXrCNI+TCJ8D5FQvdWevvhjT7vFQ+bs
KfO0nmrjs9CHve8PBUDi2jZ8XlVQH/5B/6Mtg/jToxTJiv3kA5hN13v70pYA69DlQOQHLhRn4IVS
kiaztU5McSU3ShrGAjTEihMBHc+duQs+8vosct67DcjVtzbZVlnxqlClQGbnxuLW75rxvZmNmwhF
pLfXsJ/OaMB2bmjU4xcXwZBsnrHHNrUBmFhkbJnhwW6ZNQu0k4JiPNeG5OA2NExYBsklqyUsAKiT
Skb91Kuij9KuiYd+Lm96lkSrX+0fIW4vF9gaaq+nWgiHDX3tW6rYXYSG8naXkG/8DvaLYrVSB1br
+QKpNdfPDJCtOSH+7L1LFzKzEB2JkCdSQDl+POtsBtKeTvfcQwNQDW9nLfrNKn3qk+PoWpHL2JAD
4/h8uCl0Dy7znEw7xE+xdBwkL+oFnVVrFVI10lcpWS4xaRmfVzgUG2B72pTzkWrkpQPiRV+BfMcV
Gs5Eqj77eWgNjOWOrh3ZWZcoozNBrDzv4B+3lLkhE0eQOUWBq07t8+5kwKlaiSNJrCHyr/EKffK4
2IjvGX+jgskxFdQQwMz19iZa+JA8CMZrOWHJBhsAL3eiu9/8MhoEfVjvn06ZnW6aninN/sOB5nlC
7R/iomd9FACQdUokpu19DuF0mwOoi0KQua5rNw0+9c1jVCzKIYQ9nIPtitdljyzjUIFobH4+d3s4
BMZoQtlOlJdR6j1y5erLok/A/4oaNB4fYQQOmpdp9yNKemum5vJCaFdK8T7wkt3Fu5473nFJXucn
C7MmmurIXWfPdCWnHgmtxTMwUmJ1CJVte81mO9XBg3O2WIaOwJ5hb5q85VsPDtr4NhvZxEVVdkiq
I1gFOvntEyTiZ6/Bk5lJ3FUJX76LMrZne9lllYmg+gIN+2RZ3WyHP+M5zoP9WqKwgUNoD6EUHwpN
29/8VI3aVWgEAvPWcRxTcKT+elyEZ5jeAbsadi7c6LTXOvio07QjzPAoa5Rkda6KBFlfYKtjro9M
szF4PgB5pt/sJGD1LUNGHJ9eGvW6cd8Mpk4MWOEzV6updc/2TQXXlF5wjnWIGoDhGuNXnEHCDrkK
cKG3rw7DiXuvSFniuQw8x/Uj04AiKsCcK5vcIf8ukhA56rl46AdlQWt/SsgCGKYwOJraZuBlCntu
Mb1aSGFLvVhTFQim4o0h2uxMjuqe1jf8DpfI9cNdlXWsKoS2l9g8AYmCT4gTwbqvHSW33WTwn1pU
/8uVVV/hKtoPaS4RyEGCoPeEYwAkZ19l3Mw/UFd3OCv07BtIrMR8ydq64EYSOEZr2lHU2Aw48FrF
Gk9S0BebEHIQmUjBeVErzr0FjB3MZcIy+YIBPxEuL7ozlS5uZKbQ8qz7KE8THysEEqd6x+nD4ZyT
HAjQVb7arrGkZEdVmR+aVHgU3CrRkcIgTmML/6nwq+Hf+3AiUyd6xNl4FNeACFH0LJIuqd+rZRLK
4MsAIbokVL1oS4MaIlY2ReOV8kpzvxQAHwEj7TdUVBB+Fk60nTnlec4Pxryga6SBOVcgsQxufehM
9cCxoRBjfBTky50FNqf4hFyqE9Bv3YVf50g9RLEXBR8/VnOb3uEUDyiFfjjFM/WP8+ev3SaD64wC
IoJdXwMQ2XzCqO0Gezf8aIqzViXpBFMXzORXK+YT9rwUM4MhihcWsAENA8GpZIebf0XBsTSfU5Ta
HMUfpzW2VyGyJPLwL701eFcgQr+Zzn1H0WxrcvpEyzjR/7fpFSeljAygvqrg9WquFY6Xa/XJKfAg
vKBo6LDFnQQCCZhNplz5/0sCAKgEB9V2Y3nwQHwO5Bni9OfAt3t/CZtZr4QQb+2DLbks52V3lppQ
YHIO5opPRXqZvr3YSuvzPFEwp58HxJiujiXDeaa/ALQZgwum9QAxEufMAmf2YD8pJXbMarcW7yl0
DhQJk5sN/NEXkNOKAWZ95IlNEVmN+mO8UO2BQRV47iRp4Cg4M7eUG98yVy0gOEDz45W2spGqn7VV
S+UArLaWZQ0wK8l4xAYsUXIuwG6qHHqpNSM5bNJdTC8yTaKHovXjFMgs8iMqhVfxDvQuelq5kxd+
J0zJ7FSv54EhpqMVjSaEjS1ee3iIV3cVnOGfg7MEDY+IDSCezB8Yk+bHOrp1UEdgVlh+7wuqpRyV
wFsQa7l+/fCiKCRKDoLwE1js0NuGTozi03rRqp5qLsmrmNjIZhoicFWY7WFOlRDNJHQjtoFZey3B
E11RMFYgicQNflWQ/QY+xBoPK5H91z4zfbmXU7CKKox/zgxZdOI/efJC2WXj1zoT7AfToGzW1T3H
Oydzb4hzVlH4c8xVwQwgZ+PjzBYuCV/OTY6dU6VTkCuWdk2tOIMfiarf53eTElkZ3PlF/M2bimF/
thf9G0z43wlk6gWndRlznru9GlLFvU6sFJB0KSVjmoB6Jgv2u7agPSaW+0+JQW7sqb9TQanwsE39
q2Je61FeaaN5c1fiPc56swfUv1jdFdhb7u8dKTrVc4cti+Xh27+aTqcSLltL7c8w05+KQBaCqzct
U+yXApcOo4fCtLzUtEgx8RalhsO/1lS3pLd45ofin9po89cWXIwmz8Jak+U1anxMwffqiALP0Bfp
J0s9MtQrL7gGa6Pmh/HEcmIRQTeXlmPK00tbfYscL5mLXTNqoFsnva4NHSYOz9Q7M1CjiNS/VLVD
zjDScenzAtkpZeUvQbw79NGCM3V/LtAFVjMmA0iyZwGSsvD5sToMfihWg2+dSjicnFxEzHItEOuV
mRT7c8Au8xZ9NrpV0NkhBbtY7GSqZ1cMNweeg/lHuwI2d9I/FzNgDp6E3QkZGJN6Xx8yTKIrboQW
EEVFPenK04xOtjdCwwC77TwfS8rWQz6Y8FOnkwyskKlDeml1A+F34wcl4JG1bZWL30zFIdf29aE6
RLqWybKBeNMUDsYHt5Sl5ndbp33/t/xTv/4kLxOVckHtm+cJhuvazCVY74eK5Wbreoa9y1mnT7y8
MqLQA0s2UhrTmcp6MvUM6zfmRVQ+88RthnVEscK2/W3GsLg80s7Li6T1o2lT2AXecLIgBYZ70keF
U33yljXqN3/MVJAwsQVjGhmG5kfLF6g2KtCTSiGVeluMhj9/csY6ZsYr/j2O4mbadqq8vd4EPg7q
Sz91Daw28vyBrwiSbVDpTJ9ZrHQPMQtq3BfV78PalXBcWhYkVfzwakEPr8Nk/enMriqn2jaTCRcb
W0dN2R0db+OUF6nUncMVXpu/x+BYy798KV8YSRxwLvIW+j8wXanr6yaQcEYL5UQ7PC5OlX7XzDWZ
j8DiuLtKJNe7fJ2DNf5CpGbU8TZsQ+CW+h2juFWvZQk4FuaVgySOhj53lzxMVgmglhFRvY/9jEJh
jTkEjDcHNepoRjIipCuB0zOc4Dp/4hf1e43Rf1A8WlMSwtd01NcOrUELJZniKRv9dG/4IbVQ0aN+
xWN7vxNDiTqwgjE7+2u0SQIdwrExCqXiheY4NEupG7Ofr9SrzFNEY1wZO253sf/HjbuA2ZYZ01P4
ygEXmKIxqbh7IMCao4P3ToNCwAs2GBP8fTVxVhZn0I3uYfiD2/l//n+SEMFNAchYEN+4d/VaISuW
udJFr4WdVYtWdEIAf+zc9uXxpheVCWUatidvSBiUHqkeeMnlee2JcAZyQK5zONVgkfexo60a+e5d
LdL4lwit/v1++TudX/eA9tXryA1gYjgJtXXR1rfxdbOte1epjn4TFHjSDD4qAQaeKVzsGDZJfNpb
QDO/qUCIGNYSmVoNywIhC9I6BoZ88dfqQUjd7C08QKpVSG1fCKGUwfVOv6TMI59tlM5GpOWuijG6
P+qQlenPvNZfeSGw5g81bamnTLSu+VYJ62UXhldIGdIaUQojobQOx2D3gn9ul5hPcQRh8Fv20t+R
ShkLbUchuTYsdhL5HCL+oHHtwWnj929iNd48llIqN7bdOeemqAZQBfQengrInwbHz7HKBEoGinGD
zEZBzn/MgsT5GwG7PrK253+ADGYy8H3JAo5cAck/2PNkC+Kf40DobsU4ALvJ7rXV77YGVZ33eXKe
ANtfMTsJBF//9bUi1ilMp3pCop6UgnMi2ywh07ZueytPIseEHxkpXvRXXg+yv6HltXysOFZx3SjW
HTdWdKVQAuatjgPgCkWwxeMb+R6s10kLfAbJB88SnS4gXp4tf2m67eVeGx4wKi739zTGzbyPdO4c
wW5bC9sLBM10Qhy3nVDeidHxpz0Dl7HgOxsb11Mm/vuYx8rtR/Xb0U5xcCpDyHqhsUE7VaO6HdlG
JukqH1GE4tHj7TKniCOPCHRNULp+TQ4i5dTWGGQm9S5ZomTDzla69Rxyg2/Zfelv62O4V0wfmSyd
f4uxSKF9bI0/r8TY+hBmjjUtoB4PZFnMuEBM0bZPxAFyWjEY4l4pr30RoA4uX93jTSSy7KSEob5W
jFtsecnD2R7sQzf76l/taBhILvse0hPlEEwsoWriVQC309hUL/a2KWyk4dzl82rLjN0VQiQqV7QJ
SvGRn9dXMRBHbpj5BSSdGYM6bkwMQGKxvSMfwPsgt5zDmIJRbWx+8TYY3pZLb0unQ8fFjU2vi4Pj
K7IS82HZD0XNtAAc4WufLD2tGV6k3nsVmP8gO2EK2CSMxi4qYd/ljjbU/YNzTb/I3YD7KL4HJadm
JIUo2n+qizvKDOT246nFvmcrIOXO1BY+PLNstbBPUmg7nmN2OYys1cNaETyQ57LzOubPOhvnHbbk
gt3FuPit9iLWgz4CmhFpzcX63QuxhoGa7u9iAT/6jov6sacR5ZuuHD4IpOJPfX8CLCdw59s8GGZt
XisPYhW6XyDR9pbeJ3COcyZR/GhOinItx0uYQkalt3w6G7F33JWO6rm/XeUN+oieq0OMGiTadbn3
jW9piWE5qzREyLXdSsuERbNQwq1mF7GP/DLL1DI/A1i2QiS3eG8q99WtkCFp9vlp5EJIC2Ux5B5I
hfXxOjudad7vWHDT4VHIC+7L1acnzKSaUAcOy6ND4GaiHIbVmDKPjICfatWdz7wcQew1wBXdTRYY
i8Pqny5PXTGnZW0B428aoCLKPeeFV/I6gL4MRHoDIjvPTs5XD3d9NM08r2X+DL9hRZeF05jm4KOZ
Nqc3jgZxLF8frN+e5Y2YIxa0w5gN1O8dLne0qmx2CA0yPjQCffNh6POyviGLQP9IL23P/UcbPcXZ
h58cQ210IF7E492u3UQ1CEPh77iZ+68VYrik3xx1Z8J1oiLrE8EPJ/HBHEV8aR3UDlwgTpW/nLBR
2pbLAvZNzQf9adZ/V8OSzIyDJk//a2Zk6ZaR/KEVJTtoea+EjEDDvaUAGFACK9pIGmWM5d8CEtua
ZkU9d2PrxB/I4UVow2OKjj+/Rh1uUil0GY+uoQihNQVvh7m5ZSNVpqeZb7TTQ6akqZeAyD4QmAlu
ttQKw4jxrbHZ95nfh6z34/UJPl+VcIkL09NpCa2xtydhlg5n2TbwtbpnMuXOp7j1zQ5GEk0GTEck
e48bbgBhPcj/qifZXOG24axjP3hNzvFtdnn1aylbHib1E5v5ztzCAbf8b+S+rrBqVDRVoB5t7Y7r
90rKf1itdrS4gPYwCr0cjosy0gAwBVHXSMM3kemEFR/zdl+TGwm5JJSYiLB+VHO8Am0xTnY0As6K
HSUGRZM2O3AB3wKdNh7Bnj44v8La4lJoTqimrGiCRoSuQCB0SXxcUNaWIrBrGgdjSEwTSGNx+p28
pEjFg/TGXvTE+Gos+ANSSXQr6TU2zACQFECDfe4kBajLs5ZlnaNP8g/PIxMGasj2ixZBJ0t14Rz9
aY5I71jRtRhB3ou4aLSBIMS+YuUX2Nuog995g3s9CxItru14/KQ2usruP9lSt5iC52uEK5f2Xmbc
8GIOwXtE7bpnOWSNNMB7zO2s6BWL/Ah1jmmhuH/pzyxKeZlVzUGp05D1FChW9GXk5SyrZOEG1RR3
u+R90WrGPxD8baJtDOdbWkZ4SIoldG2m4Ja19/+aLnYqNsb/F6i+Y/oExJFyQn3BjAW1rEqj6e/v
ZPkf8ZgkV5NKE8CABr9Q0POoBBYbln0xSsIiYJ1qo9aMPnatHCmsj8cMDaFvRrkiqA77SMSIcoVR
AhxPPnK+OAeLGE8PZgXfzhymtHWOxQh8I3NJLXkgawHnYjVTPcZQ/IDjnEBcbko4jWJOfGfTC5k2
PLlyTe3Cc4CoYGe2LnxlIPMjbXmyaC32VZvlVUwux1qEq1Gc1oWBbiuETD4wuELqCkVVofvzuHGp
bj6s8CshGpCf3so/8R6tuDWJHxWSVZ1RZ/y9WBti+QxLHCVrUpZ3z44CdjpCf+aw5DhFg5qM/eTU
gmfvSbMh9M+D+EpFU9M/MvsVFEzn3zj2h0nf5lHPkrAMRoNsnrHBd/jyAqfaTl6eHfbB6xeUei3W
lOLQieRD/wvUQNEnj4cXBZ1tzCyrLtF33KI11BJdx7PKOWeMBteYeicpmsNkkOiwavl53mCGr9cU
JlQMvKYKk6ejAVQo2JR/jg72JP7Y4tl/b70l63rTKxqIFUXo4iJvi3apL9PXb1ekRaDkW9VCi99R
0VklJlfOOsDkgJS50Pvtg/1omziYxtEM4Mj4mQ6NLDxSC97hqxb2UEWJ36y5Yz6bv+1Ws4Xl92kc
jpU82kDJaXmLTM8AJO8Z9dxPZ7jNIWl1iUg/u45lYAW8AXGuFnrADW4nKVsFcIC2PD84YnxsYbS6
wIIUV7y0IU3i2clQXcNsBHlR/Qi06mOJrWs09D7VkOykvTtvc8Kk0IPKYKlHaXr5G8vRqymaGrGD
0qvs+EirpKIxvOYaVZcS1aiFyOa8bZRyVQwiy9rGwixb8g5uJaCZ/hZTa1TTEcRpoTWF6uIpGvZC
Vec/k2mwLfv1SOIlrETO9Xaqy8ooG6BmoGkqx46igosXvG7QO1Ru3VwUttLXoACeKTnmk+rIC6dz
7JWX0H7MaGZeOB+TVbPLha64jN7ypmgZ1FsFgEkp3dA89I2I6XOUfQo7eBSlOboFB/5jCEG5bZlA
Vwj2iI5d8Plb2oalYnaIWa/eWWSK5YpoiIJmQFtfG7SQQXksQhdoEaQXParvHQpO/zL2lB21cPaE
viLmKjgj4reBFcOPL+R42tEjN3qpYpo20QYhXNbGkU5lTUPnWhacfNyrv0oT8UIgVWxB3wVDMnWR
CvFxqLKlHdlHBGrnQYwcVbDDJOgqncSUhdelstJ4uIFqgHISFaFIDnI7FEGEBe5t7AaGozf7r7eJ
r2qB33auIlpONouXG/4XFYVlAL1lOMaqUGkXTsal1i22mK8LzYXHXWjgLJl1wZHWhMo1rO3shBdb
1k/ZDoFZWPr/hwYRU1W80Tgmjgn2ll3yfEaenfd/aUw6iyCoQP6tTl7BYvAsEnsboiQURkogBC9t
+1d7UanM/kDENR2QH1akLQI0Cj0uKdX/swiBmXRpCBsTaG1febapKH2Yv5617Kqv2L6ri5q/u9bY
7VqzgCZ9KM1wWtF8X5woL2fw/MUAxuv04Dw618JpDbOaNepdxXFpdfjWSyUbKyl4lwfnlQKdR+lM
HjWm+K6g1+hYsyP6G4XMVEieKwcaT3/cRE/NVVoVR2FRhJpxVyZcY+ncX7lj3E5ccJE1/sGrZxrz
pl3FTSLD+L0fo+M8jP01h3qWYyhsarsOHa/tuGO76+9ZXZjoLyjxn7/FkT4PNh2Nf1+auoWNq702
1jMpiPnSEwfWuhUWY1tJaHxd7b/f0xOIL5IsiTbszt2LHXX6KhhcDYhvhcQhqn3hbUT3uocCnSYJ
BDwoAut/ltUPR4KToOs027cBet76/djoPVmh2xflEa9mafLHdhR8bL1qUS5LqeUbUpFT7DJHPqXe
iuMzh6VeqmRWNeNv6ebkQLOfbLNJONRBNrPy6w+xn18gRIca/Y0BE/gsWNRSsFpLnMqCSBpKIaYc
/ee3LNjvy108U8u2YRU4CipCfYT2s558AS79GHuNR3coYf7jPFh2b7Hc4L5p/K9JowkMsrYCUA+A
iCjEcNBmuIX+5B/9O0FKCDGLNQSqhqHaQ539Sc9wACvNJnglTnXgBqCXEsiotdIFJZTEsTmdJMN8
Chgjr6hvXMTih99v0Y89RohJgTMZhFy/1E5EgH3Ka27umq52lwXhPWjFRtn+y2VbGgMo4Z6YUUnK
y9Cs7SPKmNGqjzoKqw3jxduH5zUQRkx8Mmbi0tSOZSgMDqL6Js5ZOQ7kp41oEwF/f4iwhUTLtFsF
mImexqOGWVy73W4uEgf0IQPuJeII+nfNQLM4dLufsz63nilc1wimrNltj4rioPfL1oB7fngzq9v2
7zGyVkyUgqRx0PvLQnE4Y7Af8/xzuF+A+gPPPXSRe7iiqnN62d4COJKcZee+zQWbqj2doQiWiDbp
Fkrl0LEaQUPiELo1+SzPy6+bkwghhBBXoWUZuW59/QO8jrhQ49ifFtbmRPEFjvcTmLA+nZZNuvkP
lv8yYVIc20C13vX7DN3BA2Lp5upG8dvbbuzlBLKRxUpYVu11Ju7LGY6D6/3eAo+GwjMa2Wrw7Vt6
LB/7GtaEmQ4K/QleYip1LV+REKuRNqhn6PxnrJLxz0sAK8ws0TXaY5HATCfHgCFwg+wHQYYBs80p
PCZepUMEeil0MCUcWnNBmrvMatQloY8J0ngm4Wfu79w2bWt5Y8jFhIKtHFkNVsksmAC+WqMcbS/f
/yhzQA9lgGItRpcde+T/O6kUFj3hMKk0qYKB4nFCwnmwUP+f78lzUPCm8jFLq9vSNTh9Tw4HrSzk
akEwWf++DhbrGGO8ioNZgqKb1FxJCxOulbUM0M7NLA4z5bYet5vDEA4+Cwszg1Le3O0Dj2gonyQz
K2Hfd4Ehj04Sl5BqbjJgpI9FoSYFpej7DKh2fOA2tq35NJafHSALnRKXAKdSg8jFBVGc6WQO46rk
ap9DfzVSfe4k92yscTp3XbPRNTHyX5CsCeJMeNgdR5JWPjZP6pnFYNfL4WzE381PWHp/myEmVOgP
8ZJqTsUeYdywStzDwVCqAdJNrbi2EkUYo5YtSXKvzN2qHWeTjgkV1BI3RIisukwvdzB3F/jpVS5S
A+tsywOgPzi1LtC5TgdXQGYh5AHM2ynmIQho/vhV94tH7f0HEeLWguNDi8ykPZ7F0oxgUFsZBz9V
pGwYtnDdTfAA1GtfTIbmVYGidcCU90jmwy3res+YoAUSxFyu6eluGUVVUzIMa0HWPjoj/jVfKj3e
wpsy9cu3rikMmxZxMpax0M+2BTMABWGyb0DwtZ7DbBe6MB6TBHvB1H8GriNpvgNxETHoBbwfWiPp
sfAbwPGf5Twzz/44Ew4odC6PasNFyxhp05HSCToBM9m/TF2fEi1WLzZcA7rQsZLuATuINgNYWN/w
n8shz/P9bcupD3sQBrKynSguWmJIWKWiRzuAJhgZyp++yKz9S3DgXSwa6slEzZAlkDcND8TlIQ6v
H0vcyWVOqpE+dJr3d0kvCOR5c4j/Hgz2sUCXzfgfKy9sozYBKHNuUl5+lLa/VpSyKQR63GTv22au
acvv0SP2zPElR0wjhqbGxxaLtbk2No2JpJ6Hj01j8cldXxiFUtzcAY+ijLyUg89mzli8nbcW75fJ
ijqds6ncLsoIGZf5d9SYHGdFrZGnZX7ne55U/Nrjy+sp/4yK3oFYKSneCZM/qJxI8wCZr+vfwF9G
IeKV/9tJkzL/eQ/tZ7RD9kABH/TIDrppPfBi7iwNPvVmc9RtXSNUGomvivNG8Sk5juj0hdxxCz6b
bNMjoKYnNCQkp/GfDzUYSgDk8zeXZKSF4wEXOoKDJcIXOlWVW88WiQhGQzdGrBOyzSQCq2eYCRIb
N0Ia4Km1ifbZYwn+tFggp04mzcPmmYjX9nnnWiElu1xuxHX49K+VAdbhf5KP36TO/3JXG+Jpt6eq
cEpX9efhy+CVZtuxrYCZ1pmioO2WrzadxUwUogtQRwlY2jBN9HlFVfzugUz4GUdnO1ziAsmXV+Zt
zyX5CbBDRglFJWEOgJ0GVE4nxRqWLoaWlyMSxHgMoj/d9dkPYpT6T96x6URDxYAwwOZU3mD5l1C2
gghssAHP2mioLpBvW77OgPRd8p6KKQshFX+5I6EPeXt/KGv9xBJRu1763O4nbQy7NX1Kl+DKPZOD
XSNPBLJbPqZehJvP4lJbnrvbrve5J0qeenFyW22sOwk/igC+hGspkPyCSHiRyT9rgEVFddzE6Rbd
YqDT+6d6HsP/IzKoLxKLLREXLGN7RWQZWkMcSRJyMmqF1DXj39NYbrHQKSt0jB5ixXtIxCDxnam6
LItPHvfiGtc6b3n/H0s/11dz2IZsx09LaFO+4+f/5Xk/JhDIsLnS8Dn0+/7LFzMDjAmi/eqtmR1L
sx1j9P3wfpaItc5J+phGuaxKvu8jMLbZTEBuKsg6oy6Du0L0IbeSgt0gq9dnBLpCRI8L9JYijzYh
jatbkl0V4uhfYZmQsx5Xssk5WOPlPef2htnFdh5xa6b3nQJaZ1cSYKMP5CRM6nH1NCe/8iLRtHMQ
YkL1AVZIpURRZPArQs2+ibEdGp5ibI3e5dRMKyUpjBgGs5cDMh2Fjavhc09GP4HmVa7Pc9FUCWMV
DbcSPHluolTgonX5ag69qjNoCnTlZXjC4/aVHkjbNrMUbxRgqJrhWzYPCd2krRVTjLNenX2XAhKG
ekopITbUBwXHrKyt0g7N5/epjONF/DP2Wg5f8dqQ4Q2I5x1i+qIboXoD2kQC7EJuKD4TVJg5G5Nc
nAunagOVISmbop1QAQ24oxZz8zHzZ11tyGkjry4hUkJdxPlkB/M+kuw2KMRZ0Qc59qfW0vcXhDDy
YtmYoCtt0+RvfxPV2cLnG7bufsckvL5OtebELQSq02GQaKK7uLmddyBEIsyI/3jqCfxRHj0OzlS3
+dJPo2NhqpAPAfYnuqSwob5nCZHXd7cVJR04mEFlfNqaf07MeocanrHeVM3mUnGBP3sE/uLMWI1J
3dEMwBNVnusyeQmEq99YK3ZyNLAFivFnkXP/ujqd/vaHxxqx53Y7CAdOL2+4YnuRThfqRMblV7la
qaxoQUOKWGugAW0nHInR+kPDIUcuc8HY4jwDc6Yd2j0XvUFI8VOsOvwi8vBKxGa8l1pgMRelcP0t
rh2YvoMRhEy69xfvb26WU4r+3JGRzcHKizfc0G3KfEMBnuH3q2Rb0w2kxZF3aeTbPFEZ0VNeCMXO
uC+8nHpFCodK4/K/F4YBGu7UTrW+ABuvSPhNfVurUuTMU+JaxU7ef1M81eyNGJfuSCUS4vY45Tc9
jjSeZd/6tB/UAIa7lpnDsBSkkrtCHiY5wObSpT/qiGzAfZGY70u1Is0Lywplhy9waFAI8tkBCl7j
Dz68Gy1uB7m5x3Bq7NOF3JMx/QJ7ypsXja3m9xHvOnd9yQ5ZOg/Y6sBsz8s515ak8BCBRAfI+dI+
KncEypE7ICNnUwQ/O4BpbT4mXw6Y3/WyqPnP8NwJlnzAR9m3/UZNgwP8wjDJ6UDZDGQwpbXzHCSE
sc9DdTtLaahY4m/LwJAEeH5GSizzx+JC8sjwyMTsSaTiMP82rOKHW2hXXppJkfDU/DaEST80MlVH
EYOKkbOeq0n/LF3fkFeEqGeDsZYGtByRG6/2zXZR/Er9TnG7QRSgJmeptA875mozBW0FzuvgJWxz
dfmZKYzMrFsP9jeawpzmS610B9GOpYradPQsIPxD9q9azRCF8g3UClxZHyss41X+f0iLmmzDbyrZ
tfCVlvKbkUmN4dkm1ENoWB3YEXzna8agels23yGMiEI33D/uYWqq/pQT8CUiJypCQpI7kZPNfmZ3
j6oMkQtFpYICPBxxQlvQf7psNWKbeUY/V4T/X+1L8LlOQklNodIOZmGikj2pbyBKp7wo7niR9G+l
UMCwZbWihYanHN2jB3qWBqsF+5bed+CsPQn5tZqz2dl4UaVxsLoqNtwEj1ujVZEE5x0i4h8Z8M7F
Ppe2jyvVB1LuNwzOjKGah7jkM96p9cY2jlFr5WCIYxlAIlrL1w++f25llt72dDNbB+etF4WaQPLR
2Y5vnXk7mkIDc4ZV5GhXqQkPCZpYPxstG3Hws/T4f0Ee+xBsw/lBx08/Pl7ZpoOX3Fd1/UlrO19z
Q+jz7o639ana5ix9qMmr+4atRuUzdG6kkZumq9DJKKRvdXj++ru25enI/VF9ivcXUl5ZUhRajLQU
BerXwyBrL8i8nwkKgsgYWcJmtt/xHmA8ymutBljsegtRKhri2Q23Xy4zQvWlWRbIZDBYm7+Zlo+5
0prTVM65o1zhigj5M57S6GiePbSXTumlRAVi2s9xH+5ixnikcJnfsPxCxf5Nj4XixXXrC+2zHaee
IbjXIDYOfr3mEtpZthavcSLU5pe0XIyVFjIaXnkpLEvbnBhR78xqBguW+Ues1OZuRISb0tzw0+tj
Eq3a1FXu9cCQzUw15f0jsDs4EnDVooc3HyO71A6fCmrgNnerthTcvXWEGAjghh3bVaeC7UAadLw/
PUGf+O6JIPSi/hL+Ew4NYG2MT5XFurTTLxu7dPZNNwd0j8ihFhLD3PYXSVkt61buFNNSfuLrXLgu
byF09IuVVl3KDn4EFzog51cMmfINMIaAazX/0Ur4NxO7QgfFHEdGZCkwj1hiuO1VA/7Prmo1hfrC
ZCLS/QRnmSrCNzqnyagj+h2Dhw9GtpGClE+M5XrDrWi5+re8ZDz2A0x3TAb0vnd4rXG6ovkq53Dd
fxphO1bxA4+cfn/mJpk/1Is+ygKXTGx3AhiCBZdIaTzBDPCAHWDyi4sG2aI1OJLWhi7dotXVvTTV
INpYuL1rq8pmU9yoGyWWyBR/olbMMXLryztfR+xwbwaj7eqEfIlDB1qk4Yu1T/S2u4ys0LS3o7Hq
h1XVHHHJHeoRuYSnNrltg7kVujRMz9dq2Qp/+Q4zRhh8Z/vjSeQKz3QNP+9ypQ0GQZ76uikT9dsk
p3t3ZOZMtM0Dr865fL0PItyihaotQDC7L/5jnLn+kZkoqEZPqPcS0eYfyghsMKikt4nFnjsaC7wF
VoihwWL5pnZ2GI2q1ZFLgiSaGU/XeROf31C3xgkHRZDdokdQZ82kJmDYvfQ9K/7w2GVi3KH3XvX5
1cn9ifno/7LmKTZr6lKAhVTtQX3wehtaXLQ+lKb1t4X6w9Nxksam2kCGrzI0NJY3bBtiEZ8VUmfG
PxaZm+CGaUcGh1en6uOPG4x05/pN7GhrJgdXLLzpLpKotFgh4HSRPCBdtKJ7G+3e2DW72KCcVufy
qb41bEjH+lPPVvwaCmYNErVLkfjqqKGeaRlFKxe5VfddFYYN+LaX+mNgQQa7WhW/CvZoQuyFOv6o
PvOUheSN8YziYkquz/Jdpx4tv/9rC6LotB7gQTcgIl1UjuPO/tKWgnHzlESPkseSTlIsbqV40Gam
eyfSS+VXVPFTIndLQ/LbhITleYO+u/BwOriEEXPSSsIv2m2qrjDbrXuTAnRE3Qt0fHm2lBHL+5vU
nzzDyxmA066E/Tcf98ybzypF5XKIL3QcjSZhw4SdB7XLh4EqsEx3672E1JtvdYpdvKlteYfd5P5P
FWqFqPbv9hg+GXZE4awUM0KxAMhk7Nq0hFY8gugfSltVGh+1rU622LbXQd5ZM9F3NCrX0M6j11Hx
0gFTQ7IymzKgxZhUiqONyn2WgJOap00jV9BLJAZ9Xuz/L5I6GWUNhB0zQVDliUd03qt6AAGmGv6D
UuMQj2q+oV6oaeg0wmdPfmnQQuh7Uk/u2mZriCBndA7QIolwToJ6j4uBWapUaaD8EmgYuEtFFD2Y
wdW7KOE1KCQYGgMFogKEVulfmgU2KOOuxbUqqFeeQKy33o0ak05ukXtHNre3gqQxZTbZ8HdS4GZQ
WcAWCDiY5tZYlTchSkxv9FbjzrlzT+6TtIJeTl/wHPW2A8oayjjbUwiaHZBML2S5Z24K9XIVWRiJ
OC73Qduc/H9tpUhtCEPMnHkQyS65cw3fUcNqdOeW40k7PXyQYhaFWq+aPDKtkUST6hK1jZArzoeE
O/atsGTCLneB71BiqDJXK/BhB/M2gTJTJeF99pxllcd7a5qyX/rKZi1BmtkGh5hclT4sGzLXr4o1
wAMzFnsxNDChoiGgXl3R9zOTsL25GIurTzc9CODxfybprBXZYfbMwYqypnmYBdYw4tLN4N1HN5zW
poNlGC0DkqjE0D1y0LxFfsrQ7pmaafgfTt9zRLoAbMChqJPukR9iVsIbF2FrQJhpQvjwjCX6q3Bn
uJ8/wvBmdAwYHIEoFQSvpld0zlJxJ7+p2J8z5kNOnUuI4k7relXb3nxEjT93L/QNhLI2IxPHgiqz
ZCA1dX/Ojkp1ByUBjfQyDvWXJfwU56ThGmpe9JjEjk51WbA59BDAFsX3HmTOrMzSJ243+x/RAfI3
/olBMwf2sGI5k7hScx4yFsFhj+Ki61gbzVhGvnP8yk5Asf/R+fPkdAkPU3ADHwjO2do+XlYLt3OI
+KAcue+zdXQxbwyyLEP/UHKGl90/nuZ300HG3h2b+X2rb2kEiuRrCq2ie/wk1S57TYDu+cIW9kQx
hwZnVzmLQg3Q0eYoY62T/48FyAco5/ffGAMSPPDRnEqlmkF3TmqA9kYoUrzXV59TEtUMhppjzpjW
tI3L/O13RbwoFBbKRKw+m3HQRYNrdQhLXtuHqXowhu+kJLIQpI8B++Ib++68DmE64dggN53nPFmI
5U9LG9OEuQ4QIaSw0oIv2QlOUHB/5COLyjRLMmk3PHeAwA4rBFpDD64GKR8Z48J1uEXVMNUFNy4G
7drtBKIJ1vjkd0+zNjnXBR4DDtm49e30z/QaAZXh2hlg9e9qEv21qndT+MBjfm8eMmg2DtsMUKC+
51QcjP7IXlD/BFUSLT7AF59t4zZsW8/x+CxiSb0Dig8sr6H0yrW3zuserKRzJ9/mC1hbBfcS3Uf9
39JDJkAwopVl1W2a/gxsHAmmGP/8swdg7MArl3Nm/2eu42OjRm/H2Hh/CFYLS2MALoiK5b8NJ+V5
k9vBli7nTVjsvloINGV1aQ3nKrfxyVpOLbiaH2HeIc0zc7QCK4Fgrc3TV0YmdYNc/Z9CAvmChk4j
z2gsK/wwE0XFWPk5+7fu+PVSbmpZ26eX4cc6eWSzRRM5HcqVlJVIBqfDl5UISiJDbEAyIwycmrdc
x5+qdmHLDEEe0Fa6WjlnXsPEa6CBDuo/LrEdl0YO/b00Kf7giVXiZ4nG+j0edBI5Jn5HIIb2deHJ
JM2AW5G3Y5z8tWUguz+w5z1L3dUv87GnlYU57QWrqbfIfr7z9CtpwdigPsFajQw5d/2vLb8QCoXV
mn7L1YQ1FXQLBI2/HTp+IafhUV8/YgPCnS004W2iv+fL+T4rgKoe44XggjMNQ2XKcREaa0s5CARw
T/TxIYjEX5iUy9SbEVz5YYnZksCyjsvcj+P+UopH4r73mJWgNPKMxVUpkirCCAiXQhQipcc8kI9q
0bDZl6D34T2/x6teIX/DQ+f1CjphhefoGAROi7fZ7mGjc+QjF1fC2+vEK3TC5ZLJhkCWaQbNedS0
/DxU2j2Tq0IgrqV0pyMunUYwqdCeQcYvS/NKc+z0UTl8q6KrXj+2Ch+mHUyHSqX/Gu3UsErECaKZ
pSpRyNBO0V7104FzjaBOh0TVuGjoWVd9Ayv4DJ/RcMCA/+8ZIaNwC0/ScqKXGnC/cHVoP5aMnjS5
RGULHfr9ziGqKc4Up5WmsErsAA6f90sy6caTC4ncRGdUQOMxh3D5xQlQbhxjm5HibZHtoBGYtU/u
p8CWmCjPy4a3xpKHxckMjNGa3ZnBrhezLSgOISZ6wStnPqr1cDrk4LERnXLWTNQ8Mr8APcia3k6r
Rlrg4VGDkdrmp5lGiG2cZxg3qMcc/A3KLA0/c5wzff9siVUMdKy4wlsvyuqZ4+7O9b4LjSFOB3AI
VXQxKE3hhkDfugPG+1Kr5E5b3YtTs9uH5MStD08ECdwuxsWNqEFiZVdBw0s6kWIm5iPBHDAq6qXa
rUDhBuBtqAQY/4te5Rp1qwJZb8ptA+xeJMDcAOPUd5BaWqfxn3NujRi6lEw0uUfREJ10QuD0MSFx
4WHc2uY9gG/j2HhCfz7zqt9R2DurN9lbHEV9z9LagcEkgTtaAfv5YYDu2cHXI5HHR2b62L7fAUWX
3WritHsHnv535GISqyXd3ITAI9jpNVmd2JNyj2SaxYecCXAgijJ8Vra/jYcnWViOpcZ6B1VbgdBI
FFGdfEuzwz+95sc8ALiu0uow4rCLZUmoldXtvVjNxn/csHagKtSVm/N869TpJLnLUgtcxTKlmagz
Wuj5RTOWWGMfUb6vH/AwPk+jc5wd2Xd8ewEkl+OOCLGQKk2j+dh9yPBWtftD7zxucD1cVJkDrkt8
+r31CrKoe//x4zobUctlrCQb6eYaxDhbfitg5L2JhOUUjppCDfExcPVR0GuQpHiQ8zO6hmaOTPiy
3xqCbCqDsgXI16MQcJgMmGXHHGES4AXXa45BkClpzgS6pa2H/0ftjXSUgLeYUXUp4INiCa6KfKfX
LinpPM02uu4M2dtv/KG3MqayIunbU5QPsAX+frkysB/JSGJ3vdkD7Lj3k2s3FiIbRmicEfZVEatW
JQRx6sp6uVyilf0tBujGcxqpf498bgAavcZlbpBT4ojpwIt19LCQ062V0FRFlmyElaPCxWGH7jEw
orqL4hDq4okHbW+9ExRB65HOM6nAmd4E32iDSdRBp2CPGeHF5Ubux3ZRBSXCEuOaxfbw3q2j+n3i
clLz5exI3peFGSEzmPQvfQZrHaMatazYajmqo38meDdoTON9Tt9XTNcQPJLFFFCtPPXHp/DPy4fF
JOU5QzQS83etDawm5bwlXlfsm5de0uT88SfOgi2Ll+loTC3VacojG8Q08/uZiNgMzl8dhG53F4FE
oFsI4dgLHyK3ZozWM/WEhRKq73yO4uJ2AkbEcLIfZAWYcOQXVA1r6tR8CfTMurtID8S4pvSu5JWS
J0cubvPn2XVsOW/AOedzNprW5NFndUViKUZlZrl+GxoIaVZuHKPN9beotaRrFVKQZ4ZUEN3an9/E
m637MmTMK4vgtKEhNyBPZ4+MW5H2F54wIXw8AaiMtEJhBKJaaF1Jk8Cr0DdlJETPX0HtaFu+TO/R
BN5Hry49VZXVM8GLTOq8ZlOaIyt1EEOUMQzltXpIj0EgN96OdKRIZIQ3mOyIJbOARLbssrYw4swG
RstrtPJkrOnt/uyw9nNplb3WwBtBV63IR5AM8sRCxsybIJlzJdl0KBqxH91SJvNvSL8o/JbTmxVP
e4YLuBt+d4KhwZzl4Kh8TOG42QGY8enD0YAaR+Yxa75JnpcMxvN4UjjvX1OTvrpdjPPxRJmXGFF2
ith4RDYLtWgL5jVb5qlWNbCMeMgkwphowRJar5AtoGe55UDlFjd6NcdYJ17uTQ0BO2SGgCx1es+f
wN3Q7+yXPIx7WPACThKgQdxeV91rPykN0D52BMfDe5IXXWtxS5ACyGMgNOJHT8Fq//0YT//70jJF
m3spfvYg1w+QZdCDCh/IqabbdSOOwgTc5jX66C97WnqDx7bsOLLvvpZlGlI5n0RKjPJfUOvp/kUm
VwbleperGHMOlTVsQXe+UmLDfbB6TYQZqzutwd1dTWmLxVAIdKK0v41LcsTnwjwtyyawtf4Cet1M
z9yORVuEIeD9+Hnq45YaAp+NOn2tWhIoQbCGTYUt6jVx3PIk9Q1Ct/yT8d9jNe5Z4VmtyUEapP/Q
hfdHbRHDp+LUkS3Rd1CSRJSg44eWbsBQrftlazXUtcrgMxDKetlTpjf8/oCNPS/qCl1jG4g4WIjF
RASa0rRvKwKQzH9WdrRaHxs4H+ShxJALPcmrYA827lqGQJsLeIWAIGJB6hbAeHt4/DNb4IQKLJ6D
N4mfJjdZ7a+tmq4i7PzN/Ld3WOAYtoiumbORDmNcZhvzbTPYd73ZFoEp9l/WnkqEBpigBH1Cxjgs
cu7o9IgGN71qohZuawJ2p+bj/q1st+yHZEgeJVnKSy6OMqMYXfq0LPGwNtN2/idEwDWrLisOq973
/hNwYVkOAQgJhudBMmNy1ebacGG1Ba6Yv+/FCQKRj3TulpulzNU5dlMcyUBouOo7Eh0cNnl4rcYN
d+MXyXnYuNdKMxSz7LtcPcv29jr2BwJH/7UffQPiMIU/jEfM2e06mHJ5bM/yOHoMglqI/9B4MUnE
rcf7hJxO58tl1g7pHUrnrqkQXMWpO5Vc7TdYIjOXnWviOlFJREIbwHaICWQ7aTFEfQGn3R54fs60
0WYv0Fb1FWInf7ZlGCnA1/oY/CSCqgbdzOOwinQC3eGMY/tvR2gLd1sgvLO3UYjxrh+h4wuSnatf
MmOdJRFtu2OnzE723YhFFm9UvhgjZPQbw12pyu7i0k0bmc2a/MgZrTbuNoAwrfS7yFUCGpEFGJIz
Tps/eKs1jh1aYUFMVnLcoDtKJhqolYAMP5fLL+1aSCt3J5wtEysHpB9MO68OhGLMLlzOv1y4DBcj
8E2t1QJNgzN03pti2I8se6c9bAsIl7Rqp3+gVSaFlX7eTQKtXvYhMWZbI/sWGAF+4OEyNRApv8BU
Ikyt1+GKsoYqRPxHIt80gGPxDGvpNzoI6Gf58nXDZjbepm2ee65YJqjkg6ZzFNhFQQsKHw/e1wOn
X8DyOJNDEaqceUgcINuz6rkBH4neSI4yKtMzNh1ew7+onLHwiR0yNnI8omNZTqWBSsvbai2peBDf
+5f/Ilxh+iU5cW1HrxtZlJx7x6lcZrl6q2EgCSFWyxdJ3/mHVRuO+OL2n/aqowhDeAkZZQ569brO
aSkIsaXt/Vgx/toO7+3Hr7kTcolWMM3XhERwI2RElzsPwE9dvAlX+k8K0nit7o5fIHnDsW1L0t3q
ifM5RWaNO6YIjMInrvZcJkg/II/rAe9ez3nj5jOlzg/DsxSaSeoJFC8gm8OwQTIXPEw40RDHTiF1
XEZnp3ZTNR9HtJM/3kVpuIhs4UlbRWLBRy8wBc30Tbs+1AedyIQmme9eZgHCjnrshWZUsP7rm3wZ
/hWRDw4Uwp1MLRQlvyD4DocxPN09O68xbxySiYQyvtBz3lTC20j7hLBc6Lp0yrm3C5lP89vsrC+D
kW2kUY/GYgecSZgf234RJ39qMYw1vf6jSwM+U4BP2axbRAG33w/QYxC36LO8a/t5xQ8JHXkTlYzU
UjOfYx3HtX0zhzBLBeSWvEHgjvAo/v401SZY6curCavKGPyvzAlNyUHpJZbyFVHyVpK0ZFCwkk0T
laTfnoU/HZRQ022LhZT799FyKGC4rMqDrtmhZqLnkyJl8r5k2oFmtdEPYh4dmva4WPqbRJfz0Ee4
tlyWdgwXBq+lEZjGkn4GdEmVUEI75InzbD6uRi74k7STqNwToVYj9W1hJZZ712nUL/9jOPSM4HIN
qeshxZ4BnijK622q6T2+RhrpiDFFyobh0gfgsS1ugKqamIbbpMjW0NqjCQQdQMusa0XipypLnupI
jTL6nJkuABDmPzaZpDMMDoH3Lfur5dZxkODQ8Masp5oXpoQeYtVp7yr5/pOuiZi5k8stEq91Kxvh
SE+a3qbLYOZXyDUbsSv+LDYDD1rmpxzpQWp/jHuIimVobfDpHJhJqg2kbtxLBHOc6+ezBMoqqxKg
qCnTqLtbG/oVTKPk2s+LTEgPWCw4W33svzcXoPpE5PbDPPGlZaF4F7fkRxFTFt+MVFGuZb+tUXxG
bJnbxYjIIwQVAwbG6WNpjBeEpQtrwwo5ZA/GiMpEEIXjhS7n8Tb9RM4p97ZyH8xGWrZaGcbM94p4
kX6yzGEBK5uHvyn5VR5OPqfrsxDoIORRezPOPSULpZYy7srYd9WACpaU8kTthQrUTMofhsficmI9
jhU4LO3D4ENHxew5VjYePdZf7LNW1lnuzd2iqcP3EGDUj3en86I9geRzN8JXiFswtvVSfP2nyMEw
A1nZJ1OBfy9YQXYpiRZ0jGJsCE97LugfqcEGS082N1G76/ku9jxyy4Qfs/wa+zC4/c47BXFuOKfc
3rb8j2FB1stfhfhRn1g8uvgYZVDKuwp9JLSAKDBH4zNmjjez1xHyS00MuMHQ/emXlyvEJW6jJEmr
FXxfRj2n4j9Jg4+LwKw454fzZFCQKpcWwn9/HyhLxcMR7nb92mD6e7ba5qGE1s/7NFbDYYWIQd3L
Q5a/SjNFG0Ez9hCVK9tD6LWx1wclAqjKl2IjyLvLdgsp/5zuaPThePV8vHj6dby5n8k/BaEUK4Rc
TQAjbg/MgTKOXpN/0nRv0www0ffj9vvPtiLJwiv2WnhFJ2hL/X1bHZzIDiKIAJus9cOuVIdXqQRX
k2D1/HORRgdeyvINzcrcrOF3NYDhWjNKQ9cc/lmgeRT+sE38v5BxzJPN+c8nEFeqbZdVDUJycdIF
oae4oCg7xzJL7yys2fpnyurAkXtFFRfyzijpqae/+oEHXm+nd1rVYDKjeOTmp5XqkiGI67ocGAra
zNftHafNRBqNa7ld62BiL99TBhf9oF7fjVFA+1+VWR4OTf02AOEXMtqlEgzLCdqfYafYWiLL3ri1
ZDkfomj1NvdtqO3lf5TUvsF9N/sRbeSA+L2e2QC2Z8OQjUwR1Xl69vPaEPTomA863jB2+My57rOr
7Ddc7ThmKcb2EBIl8yKyfzba0hH2EPy9c9662v/Xh5RzuA+wvfOx2A0UF1HMq5rJWEYQyrM/I9sp
ZUzSl5o/ttBTK8ZuOUTEn/wDwdp4rN7X6ezqnxI/F9P0q9/jR7xUDXC18JaiqIX8wCUU/RtMEnCg
EyUhrncSKuRwdGbqBhNeAWoza/5MOobhiI+SRpMCSg2+4IvPkFIop5e6cAJdi8O3iPIEBgVd4ypA
ehqrKgkO95I4f0VHTu1K5AguKn8pOO1g4SdpCx4q30ZdCjqETYh7uyor5uxjs1b1NwCuRw7TchwW
lMgX+qnP9pYQpVb1eLPpxBzRdkp/pNHL3pjYIpbmg1YayMlXPH0daIK2S53bRL0xaKpki1A4IX9B
rgdIDIrRQomtcmTwfsfu5oADkeCOmkYwFdxvoIykK02lLG8hpWbiVny+GJ9z7pRNUvpz37wh2YLp
a8opWJun/vHq+c3QWlT5F3aCy2rhCKL83JzKrCVhApYdePtf9Qdxs/crWTMu0z5FUbMampWjhZ//
F2TH0eZ4jXlpFVRamGb/Y34cqz61HWQ+XfGGvtjuqveVNg/CwdAxBvz5+P9r4eFfAlhLZBgHUD5S
nKqH2sielr7do2MZDlwKQamjDdNQACc9+VnzFy3lUNfsJe1gyxwD49JilllE0R0mSHpVygSjxLkY
0nZT5CwuJxqoIWvNDDRB2nIFh6jlT/mY6QBIOHlRJ7bCnYbVz7bj/h8rebZLdpURcD1Y0KUNFgV6
dp/MaIa7eNppIENrZR401ADu1DNetUqqgQLbGozladakiAgQA27Zcwbqp4BkzSyq70hxXlr24I9m
VfiHiCV0qVtojp5IOWuR8tkRD1xgj1WQU17A8GxugO7awxm84s157eXHoQ9GfoX7T5U5o5WczO35
KIE8yXIXhsoTBGk2NnZ2CVISmSkxLD7E/tButlUaNWvI8SZLxAC9qwdPq7Yu7dUyuJuMeufbXjLf
aWfif3vC9BDnERqjxtucHg83ijsJyuE9/hr5rQX0v4bs+wW6IhcziD00ldvJZ9LkUZKec0LypqWW
QYR7yVqxX2PPmKqu3qsLdd+nZGibzVYmi3IGxettm+FOFdp0lEQpk7qH+k2C19149OTC5bnPnDS0
a5r/LTpqqxkkVzj+aMd2JRmfQv+HJNfUnXOC/z9eT951NitlKBL6oLnPm8yyQ47GlBBGUF2ID5FO
YP8QgmefWg9Der0Zmhvrc35g0xmIPNmveMN3jJ84JFe7+h3P0Kmm/Ak03hUex9tnDlOBbGMM0Ay6
Bc3wUweP2fQMnKSTDJDe2/RHjdtEa6XnSN8SNXX6ZtTPLpqdHdpcI+VZRA7ajuXWJ43e37s4uOpf
FFTDMXQqepeoiJ2/7u1kk9FUnwPLId8A6POgdW5XJG2Qc2J/iUcG+76NzPED8Z24ZR7DKj6kJlDb
O+F2Eqo8rlcW/mMlmEbWzKlUl2Yj1jNnEn7ocxILv8qLOTrnhlJD4AY+DHCfr42ii4aPZaM0Ett/
lDRkWzT3VXeW7rtyMdqeRxCFSJaXYEJk4to9pqUtzdDFb/tteSm7FvSfcoV0nsEhPveSo27jjmdy
Le2QzKlulyKp8ihdbfFcCyMqbzGvWi6QNbic6ZfCGxY0k+CBwLX3a1pXGPVLOjBp0HFe6BFcyfzl
p+RJcMYnJ6GUgqgGrctQ3ENXGwP2a2Ko3rdrv98RrD4ts/5rcCS7snWtb0SwNeLeo8p5KmE4JtjC
SXI//33o59h3OxxIKTEzr4VEDgIOGnqOeJmT6wS/NGtPTw08IQObnXJD9aldce67w+hxg/L4nZ6P
5QlHVuTavNwB0SP7Ho2t9dq230I1/1pAoBl/CiO0yc5WTGPZf32ss4nMZXe5bI6xMcQy7UwxD17a
F9gGE/GOXPKyYEXzN10R4KIlzAU0nADoAnhe/nJbj+clXN9O3KZ53fgfBn0ioxnqeDOZjbAiRURn
nRt5oTg7IvnEli9JUqKKJ3G3CcSlwfehwvAM30GHtpA4Gz4mNhIJI5Fng0Cyz2OHckRzHZFBBuaq
01PrawDVfIqDotD43DPbp70ge/ufVkpRdXcukBNoPi6zEu5kjr01UXgGGFCDwPQcOmMgevnH+eeE
QlHf2hTWGXcT97gR+RHvGRdz3mDxiTPKHOZYhwVyCf2fjQa1RhSV1Ik4MxQVqC3sQrjXuR+0g5gD
E56dS65VINJ8bf0yGjj+71loZQHK59nPOCzA5suYPSkPIpFI9nwnXDB2Ro309mNSvwwAiss4bDJk
PkY5rmuUHUCmBMD5jF9W3+oIa5kBlSv2/waqYIUTnIiH9LOq11SQ+YQEvztuvfr1fsTA9HQrE+21
C0r5vtdfFLo3dtZjyDU+hDfNi+EiNP7QqpK9sy3c9l91Bh2FhlYgs7Sug3PR1ZeKJHm3diytwsJJ
uK3VTT6yPT2ijYL7sY1xNaT+TkycZL8zIgmIQMAqB3DdEABL6DVVEHqE5rrbh8kZNJeJ2EgkpZae
voCpC8K9lM6oeJquLxQ8Uh59op6kGiHWwygVBQ+dzceopc6q2GDxG4jzoHg/SdVyjwFOJ2b25Lxx
kyquaci7n11E8Kr1KBs+0HcXM8/I8+ZX6h34/j6Hc6aTrhPxiCQzCkQZehvyqoW3OdjUJkTzBm+v
shnP9GFVR+SnyVSFNL7lPwg93eTMbRl91VEFA558E4uMK6JPLrNqSMtBJyOvUGucAy6aG4ClAaHi
RvUCtxgbce++2PMYwfe26vJHw1gRfggE/P4d+q4RrTZEDePcm9q7Nuuun6dZwF9MTgiW91+8vU6Y
0MoG8QHNM6zbuk46ueJPVR67HoB88n3/lpYNTV45t0fPHHU3XV0H/iEbw3uGQQzAK0B9tDUymKWI
iflSiKw32Y5LdCV9FRFyIBhNJOpld1/JDKoOXMb++KDmPxki3C4LKp1NScW51vhupXzFq2FHVr9e
j2jvvDCt+mdOSP8+1CJL9plS5KJFnRnLS9NHPo07OmPiZrSS3wO+SH+Rqp9Pac8i77VuHkCO0z7B
GkxjkuIZv4cHdtt2jB0tMjlzZXFp39a5++EYA55rltXYswPAl5hZmurDGdahZcpQH6Wm9tuAtAMz
2pKlnuNjkXqT46JJECUj+ZNovEDP4yzd75Fa6FGtVVdQEmrx7aDqCdwHK8hw7zkDXiu7y4fXgsFT
89+G8TztEFkcCJJZ7AheIFB0BDxyzKlHxrm2AEzZQmHef9lZCpV6bcfw8+vLE0x7/hMyg+BdF6fJ
iKlJm+iTeiVxXZ/EnWDWg2wQMV7cnW25nzJ1tnrqIPiNp+0VTkelxhV8tM482aM9uB/yC8IfOd6p
5amP8ivvG3VZd4HZGOVtj5JUzcyLZCTvniuix4nQHXinBvJSqPbbBUPcZuMROAuPPdvvLCo1u1YJ
JsVAsV0O4sisWF8xrXSl5OOrzkv0KHfMqVaGhgrE98ng241kCzDSyqXKSuKPsaz/hXUDjaKi1YGH
1QwaqgX2aBWZX4ohRCzjuOSuoLVkrZEaw7NjNNfmRZK0S/3754mNEPqSIjAUr3C7mrdlTD7dZaNR
SPf7/2f3z4gO7Ge2zZOAGleBDR0n0/5+0CwjpREKT4XjEz1P226FojtPOnPqvVJzFgdhfIV/BCHV
Z//gUetvBOdJszoT8ZJT/LT3Fpcmf/Yj57jOwTJlZAmCnIUD/LBIU4TA12f/tP9jYJPZVlP0r8Wt
7BquJdrc6m+7sdADNb3ZhkFKXEu48j3WlQwmB2RblXpZcGBvWFT0EiK9wwz0qT+8nvrMii2Rf3Vb
JyaCG35ALFovz73Hg1asBjCrpoZmoXTuFJqB/Bvnv2pUSG3172V73xzS3DSRsjt1/3vFLCumfRuT
UpJcCB+6jMgXqcBoqbBM4AcmcFb/hFY/SxagUcdt1QAiwKvnJ06eybIUF5vT5fFlrBB7NLI+nLNT
cRB5O5Vt7kxE08STpM9AtzbyjKcTOuILKxdzUqLv5XMRGnLRg2tNbl0jUiEgkTwAf+YZsHIVol4I
+dnV6cHEasd76bvyAyOpzh0SQgK2gdH2Cd3bzTAXBk467isZf+s7AxuvduUQ/eO5ZhQAcspIPdSb
QV1hxd02MYVipg2X+tev/m/yg4BoeuzL2aEwtPAQPRFYM8CFpf/G5Y0ZhJyaHww+ANdlbfI27OIN
butY6ylH0YJt5F2yQeO7mBw0hjnffUIvzJhszIsoLCQ3uLTVPdSmhZmCLzqgQ9OdUI64SrH1QrxF
VHEXliOc2KT8tmBrEdIpVzMkonfyu7belSj3nnQA1ddcgvGQz4GyvUTn2YD8LaZSF2xfLRzzryEL
BSreqjuE8Ll6Iiju/eiJrlObwIN7HmNVit6UGZmeOaEBTK/62608an5jhjM1QgwIu6dRV27AvUqn
3fn54oXefeVrtD93XqQGYPT+vxeWln/aOWxbOkxnWT3BngGo60zaHRmRk5KMz5GJJpLFKcWfHWcx
stK7dxuqwkeqfZeq3P8Z9FMLSFznlSjOyu5WODDP4JH1JmNjCDDDs0YXwb+sp6x+HqXl6K+qTosR
bNhpfludrjas6SqJUrwP3Mq/nB/7ptyuNvwjnpYWySWxAfMPMky4C029h3fLb2TUu3/eqY1scwTS
mqlwTS2L7yYSUV+Gs5J6rkoI9sbWKvY3OR9a8I7jNiNu8YJmT4HqdgYp1+eBdWG72cGVZyAfoo+S
rp9e41wZZpo5mrAIj35SMy9l5ilI+dn+9kTCQDAv1A4bkVGumOjcoQVu94//jyyvj5FVemCHbNA0
PY5eRlCyD3TivauYxH9v0mUz8XS9xoNOiVOGycF6mgzjqxLNF+778tqrG+IrgCu16d+JG8sKu1tx
0Huu95jBy3keTAYJh1Is1ln9z9S82Fs6fHE135y3mj+4XaamU7kmaoQiBcEAjdBiAySME6+lHiTP
ip+sf8wnalwHaS27Vn+0jjr3c0Tn8HLp4yNL1px/e01J8e2qgtsavHDX5XHwuVyU8jGwAjbRTBOp
pJk2jdtJ8QcWhJ6dJy6L5hJIB8AUbqdpsxVBLrCX1HJn2IS0GgxL0Ndn4gQZkAk6WrqnAVrBYe0L
DUJeFIJDSl2Uinkadjdq6WNtUv7jNjy6Gtw48DmSbWwl6VhofIlYf8ydRv154qb8RaCNZ20b7ybh
ju043YyUG2ImHER49fYNyNylPYffVTXxMz/WkWJiNzYrnRa9jNO5V2kmyzwcvdir5b5tPl138qvR
NL+n6RU2D97DdDiog8KkOyBo5Nqa4F4VCznvg0/FWhXNciASBQc/npwGruzXr28PlLFD6ykuTH/G
GQALZxshIM0RTt66rg5CcI/eM2fnEwuSewquuY4x5UlL03GQ3uHYR1qVVuGnJ/F3yZguJ1cVc+ct
C4xOjMLIaPTX8mabRKCJt6A1GMKlyriZ7DYmYh3G4gcCs1hYqbzHKZy6eFq6SwCIMxfWE4+OUW8X
SWWb9ZMS0EZXjXFBflGswIaeIFQCWj3/XMl386UIEFbqzqROV5mlQatnwvpL9XzKAtsGpGJHBFtS
UxmwJrNKU7WV2qcnUkML62WazUyc+cx7dVrLgt+bjQtBKddJXPbJsqmGZjTc3eA8IyEVZdG7Ajme
gf+bOY+IcnQoxTFD+XbH/4ME3i/cS9SgkvURLSHWpLO2/ya+EdUGt/RXQLKD0bTUPZVMIraJY8uG
ovgyQn3uJ/pLa8a0tWeZGNq5pOd7EZkWCT9OhVL0jJUh5UlgxswCgQ1Pc8T2Ok/kk/12E7u8ml7X
m3cOREgKwmEBfuOsWsbvO510GEOT3e0Yc7Fy1mgUZ/LI/ghTp9RsfefNAanYrywv6ZhBzIyELGRh
jYGvdf0LssypnofI8xPBjyBN07ZCm9rry5LAx99bnUuT+umdT820UaHSFj7rouRqHsNvXuke5KeC
wI/zj67xsR1gjKawVOsHW/Jp2fSHE4QrtBsclB3w0qs1MiBBL7i6QOSmBPBJg72Bm1CaWW8qD1Os
AURvhSoycTvocXK2Hzt2BW7loW+GZfyAdk+3mA9iREFz2z63vKtU08mU/R4d6geVdnUy7rBnnF08
q3B/4RCCVI6jaWjzx4hmNqxPwdNOy2p8ESYBf+6dzi7pyJGfwkYdGIevDyaYq1LPI0Vgk8DX57Ms
qcozt0Cr9M1DPRNn1KR8nttBaXM1zJz43jS0rUvpEuZwwryqsJc4ZtMdvueKjx63cy9/jyzG48jL
vNqETYoupc98FqMDVUCm2peNQTyTts8v7f0A+BdY0I87QAmOykIy46ZMiAMenFZIoTlQiRTf3ESy
Lh5KQAigEnA+ZmrlWUsQ5l3Bpp7vu/QRgQDHpfoeIvuQFscDk7IOHzp1SL2LRh2RBp8LgXcV4ZTU
kqC1Vx9ldXZjWoYUaB2E20+CKkDUpZQ0kLTA02ITOir2GtFPnAUKVtnjTTvkcy5DInCYqKHzlL1E
fEnVwxLM2EfpSohJ4vh2eenQxpfnE1TksIShdYkCVtsUelmrFQeA6mVh1mvxhq3xXYNUotkMaPjb
wx4h5O7r29APbwFUBszdU+XiTFG+tTpWfxQdVe/A33mB1/yF9FekXFY6BfehhoKVCu/gRZs0f7+J
QZ0zHIb1wBGcvn6gn6kydIoHxS4QU8b0iqff+a+Q+iOLvMo2Pcao5+lCD1Ax11+J3QGZ1GKAEkqs
w+QBrKEyo3w1339c0Z+3V0+BwkFLMsAtHHukSOMWjZHBNzVUn5/SQkgDYPcROmQOjCBProu2xV35
M5vFkqgK0OtB0phWeXzjOVie1GPIX0bcK40c13wMYWaZQLwBBmS/XpEAU6XK1NfrYtursMplw7YF
0LoJj8X+Ld5L4WKTRBcqLvjBgkjr/dhVEQ1BLI9x1gB+sekkrpB8vRDtmJbnp5llOK3d3nuKInhk
HA+wluLJgMrTGFEpxlkV1yFxBQySrCge/1zhs8GK0XRrrNtLSWP4WAPTIN2V1fGpzyTYtUvZ+pyE
rHoIkBMX6ynoTi7lju/NFNvo2xxeMRT8bAqo7c97dI0XOxgIsav7jDSekykltnZMTx0uVonXjXpg
aqsgUznvxTo97Ac5mRgtfwLR/dKcndwxjxuJiYb3pfqhSwMVV++/RbN4IW7cay9S16a98/dHZnsy
z5/gJmBrOwrdKIoPd4bEyhirnqs7jvBEOTf4vQQya3KFQRE5M4UFM37c8seXiMOxambMwQcZHh7H
T6qQ2w6FkdJeb6tF0llC9IJKqEDiT6nKcH3OnQtRmgP+toUfQHcShQPMBIkWNiHiQml6t6w4AWEl
13Vi7STeizLqtitnkzEILtjscNlwA09tKMAqJdGXtWJ5IAwZ9ysLgerH2ADqp3lURdMOJIENOele
lGmax7j/1r+3bhjrUAvK8+dH9/cY96/VBjSTKXbeshqxCNlbW5krFqQp9w6z/9GKlmG9Jbrx/JKt
3E+RZNNuYK/sx7ravUg0HCowbkRmEkVJukiAJ3FJJFaYJOwXO+BGmYo6xWAX8Cc8oTEyZbC9TyAo
QsK4lM87NHxn9dvoXKs3NGjGmZn/hoDIwfk/iZcQ8wwpH1SVPCp6XbM/jR+Ta/x2SNYLkR3QJPVC
GbyPqbTnqzN/Ny/27/mXeZ0wO/zO0GEkInTzds0LdN5tp2kD95HjfJvEryCFu2wbU7liceiyJE70
ZDV2JDQXdT6AOP0mvo/e9Xz28Oqq74NHsixtv33/T82N1CirOeUiQWC3W5GBcMk71bZQVxcTdZ/x
4V900T7dY/EejSzls2SUqQyNBGmDy804YxjAkuF7MlS1jKR8wmUAnAefxL5pa4ZZ1xk8W2ljatJj
7iPJB6HXqQjNWINqXl3wa1llEz5+A1Ok7FYG20BrbIGS/CrDmf94jsm0cnPvfVWzvmgEkkd9kifv
KGNt1zE39+QAOqwcUPfNJdrRLG1tlWGtnZg6/eK4uJkqRbcSiA7QoVQoi4M2mTE1kL021Sbbih5A
ippq/IgXkiTdKjKl3QIr4Jq4l2TzxmBzzEXEsboRWk0hdyURrHazCtBRTWwbP+P5SPN6SpQvKTAZ
sBOGmcfbPnh+Rgfv4YWhFz0mQ4upaTXfW0/XF8E8aTaONvcPX839XeNmZDgRuutvaDEn8ojS2Hhk
cPSSMVSYVOecI4bW8Zaz4HUdMdBOt6iWLbu19X2kOBFPUbW2RDVU+a/M3YQm7/eKKT/shAAso3Lx
mcRbITpOSa7waWLNyIbWbC4Aabi/vohbfwLmXZrzGg8aynCTiKGaY8XJ3Xx3WrmTtJmPSjoJiUyT
x63/YbGLBzJFeQbr/GoL/ShlSlNpKPYlKE6pX/q56gHgI0oUYvWmtWm5r+pdMxcPP6+ePI5KW333
r2IZYHG+BY9sKHvsnCz0fagQQyT/9O1IjzD4lMIKxmNJYqTHlJqy4KQyOt+lEulu8w/M1/qT/m+U
pEqz2MDd5nlJ2WG2EXy6GDs+EeLwmq9CSNsUv6zyQXGVBLuyr8GhZ3m8RraaP8BEOHGdasB6x6pD
fLtsiYlA8HTRC1VTVrhiBtPay2d88KCTF7iiAupEjdSSWjXRxNgd53ido+w2ov+2j/lZlOYg7aG6
u+9zlxsJOWCBJvEtdCmveQFAmL39CQWawzqSlEAnGevoG7DVeIJhvzC49CdjqWSzb3QG7Pp5xX7j
zZwmiLH1b4/+01gLMWHyNWZawIQr6rzsBJEbXajiNpAfwiSSkuLwFs+zQDUHD5KofWVsUPxhvHZ3
6UWjDlPEJwdjSRLd1DPlu9p2KPsaBuhggavpSAh1PnAo43/bG24jIHMmeDMOmqH1kiOcRlOd5kRz
Vygmwz3YkNmYCOf+NEwx3xuUqJIH+QZsgcPl6LTWDqziPrJWH1CNmTWzMhdzaf7s2EVjTjTSGnwv
GcENn23u44hlvm5zXX9kqoH5/6010iBYy25qHThKXhc+CwCtCTRHVK8Wgi+YjRHmjyf1YGsY6/d2
D8Gvby9xDOfp2/M7M7lJjHa9CP0CGL4oMCs0nuII275hoBzVJnUwER9QTYJZ3I7vHlGaPrey69VU
25d5Wz79XCpaimBo7G9mQZ6W7yOmloV9bVFwTQ5Wvnqz9+bLbFvhvLJv5AUDRLwKpim2/8j/aR9w
2IJViIpC5aIM23K2RbjiH+CX+g9wFwqj4w72eRENkfoCOrB5LCeLeWqrxq6SPq23r5FOwjC6rPCq
XksORXfbeXln/uEbozqNK73UNqEU9K3T6ErUdFqgvRQ0IVNcpOjGxQ+eRBMB5q916wEEvY2ETZnO
AUENIncaGC5poVlx4QyfKhppVrY4xwI3ryEX09O+FpVgczCCvdpaZr30DMKljiLbg1RL1b+oW07V
WFMvQefVSOyQsbXX3Jqtr/Y544WITBxnV7bOtsXn1qWzEuVNZaU+Urr1J8bRGK1QK4mUNAmHLuM4
CRPte2EW0ojQ6Gxv3l3fCNC/8LBseQZoCoz5iumFWS4dgVnF71MujaPUpwfoaM8s+OhC4DRlJfCJ
hm8fUkthNZqJw7sw8a/5KrOdn7TA95cCCVkeBDKZ+5s3nzLqF+chfghparDmPPqjps+MkQxXqpE7
4mXZj/29wWYoP3LcWTOg7/yOg+U198ru4XymC2ndWLFyk5EcpbHWkNT7qSudAxrmVpTL+73qRa3f
uLmYHbIbW4Y+l9jlc4U/8c+msp9Ltf2yPBv9RDS/O2hlJnG73W588Go8IOtB68lSsjovXQeNgcvL
R2ep3ihgIF53sUXRtk1HuOW2zENdSxn045RaGPew+xuRcdAX8wTJD1xaLmo0CF3TT0r8HHI/cOcO
38iycgm83LrvsWVDBLL7vSJr3AzulwmziUrmlJ8knnt8TNnFFS1qw/pC7CC6VmJ/P1OwmnqqXYpo
W+se9jmK2rDbwsdK8p1n0Fre6VN6WbGNMkGV0auaQymBijrdoDFRR1YvNOxzL6DMrr003Gp0VxVA
JjKylizVIeCF1pROXOb7lSpBinyMySTXVwbGs0sEWgDOrP3H7w6NeHJxrnclwBYfuDsXKsrDtg0z
MHDGFVX+/PkZRXHZ+0KspPdowfTQNJP8x5miS+RguQgL529HnhrsO0vySa9a1GbnXZd+AFDRJggg
JxvQ6j9yDCsyPD0C2qNPL1+/5F7Mna9/l8yt7cK6dOIqqVMCO8DnZCSGKu6yG5xNP7S6P2232waJ
KdJd891XGYWSVWDg+tAXXCnPK55pJGQTGdXZVD1ZsT0e6zhTb3XfFGHSRVj4iwRI/Nj3vptlQNxI
XwttUOJnx6TSNtuP8pp/Dy0VWJQsZPWpflW8v+IYFcaG/RFOfEI7OJuEdluUdD/JMwSRR+EFJX93
OLi79hcRKswPIJQQClCFWXpqsitXIhxQclB1Ho/GE3upHHe2igb5RCqFjMmwow73pa0V5c6LNMNC
efiH3M4XNzJUXWI3BvWoU8b09BAhSzvlqa/KE8folA9w8SvNGgzhrcSgdok+eEp/0UKV7KOjFFXV
l9j34NGMzgjXsG2idmEv8WtowwdWeqNMt9yYogTXK/g2zbXSmVAhQ81HDatP8bVb8lV8MHgRgw4w
+TCTAYJHFK2IsjQth7l7tkIflNkZJDIDwhJFtVJGPVuyVDVUReOlNeaL0u2EeDxExftjo+H9WU+H
Gvjxqa6WojAHQSQpQaGS1encJd/cS4BuuNZk1WCPaNtUceVqUoi0WK23DdRqFj2IIqAUK+BNQk1v
Q9747RUcW425trFb/DoM/TSl2k9GHRrxY1iWU/tx12DWuXj4xaROeRa2m8r1y96ySKvjhZ+vnPXm
XAX1q3DR0ztnPiHKYxGtgmDvvzeqNN1ygrQWZc8lx9minLbXT0GtEkqTn+wuQweuU7fc1zb/oVf6
a/NoKKf0WGowtXqkBFFWyKecyPh4ZgRrYz5YpMdUWZtY61e39kLRJJQyQfrRVWSHABuPuhkkveZw
9Lnmdh4LH/N/s4l9ubNxMOskHr5tgJavUBWKczicisFwCgt8HZYHxWLT1uSKzhEPLBPK8p5xNiYN
87pRlf2rbrrpxgHaWQvQj+tkbRjTj/9HTlCOfBcXdxr7Ek8THRy6cS64O1p6Mk0WgJNhPxpfpXNi
mar7Z+hkmgpRnssrbusChVfS8FVaZXO1PttOW+MBblNTZdPl5ii/fIlsgFrhQ4xtbFCeN7QWMAWI
9bklbv5rDat2qvAHL6uzOM3UKyYqNzbbXcb9d+BmuVD+8ynIhr2OY93RJfQ46rjmeinyGDSE2f4y
vQcwlNyTlIdflPlI92rw+bFhYXcMw71hjJMPFdS+D43V+YJXYHhOMLPDWgfcxsxZPBESfm87jPQP
uOSl7VK+8xLSve+JJyu114PD7CO8v2DVhF0luMPOXbEUFYdMJyW0vlfXbegNxy369kBcgrmjrxNI
cafnxSsqKZ5yC4lXO4WS2vVIutU1Sx2Ysfn/63hVdcDA01oz0/6pD+HjgxywcNz2L1Maor/GFiHP
bNu4uwynVMGzhyfwKEm9Kk+aq31l0Od3mLu36UKHJ6nK4BSyjRqzHaFIkr1qVjz8IcAN+5G2CB/3
QO7CuvZ1by00nQ3nXav8ItZ/UGD6Z0Wq8NBz5Sk5SWgx13P1h4e784oGlcRErDYR7gJhRSOB9PLZ
l/VDSKx6oRSruodyTKV+TJWe1lpGDGBdf8GwvihxW2CZUi5uogali2YL07ZlEqBiHQyqRQ9M6gxQ
MzK4WF7BwUWvQd6/uYN6KLFC9lF+ZpX6dtXyW+KZSnyxgRaLNb8K2agZ3xxt2sz92+8VKoETZAxD
7kXPxzusnzTQ3oPvZa64nLeybuCcy6MbJhYJnBn3d+ydz2F3VLh32JNPfJgOgd+zeXS2FE9iNrw0
vTLCHZt9rGGv5LSLSd2MFsWvt9X6/PBivmHKccwhGVeJTrsKUtKiLX6RcJifYo7lJwEjoNSvqKxy
OU1S0K6HyilQwvKER3C3KzY0QrI798Hfg8u5Ua8css0XTz1DUMUh0YheiwcbOTHECtZ0QV2qKXTl
Q0HBYXYozr2jhxpfLN57edhiCMOJwCl3NVOHIO8k7el9W13XYUKJ20xbgB6ebIfOPkATduW0rO5g
dMcKR+31ucVRYHoDVGeFy0aS8kr1NX7tBa1mJZJbYCZG+aMd+nV+ZjNdg3vgQDGAW92pdAQsmZBH
ClukCWlCSTDGKwr95KYckbyAPRO2USzrSPtFYpxjGQsHyMoCsAaazWCXipB2LxWu1dLdH1xAMXsf
aYb7yCaSGz7ZQFRIJItiNvZoZzDqwtHOqRf87qDroAtd8eE8ST0+8x7s1ob/toDyQmqsegfDkwsF
OqBCydzXFGpzvGHx2UIE3AW0TDgeMekb4yY/9oCNkIolzQJjIiVAVGLgUyhpl1rRgnno5+wMyrLo
HBUE2d1SMkoMSFeqD51+tuZXt4YQcDG0ZX+F7q/wracE/tGBuvXyHw3nIwiQ6mDh9qUD3mw1sTCf
kWSK8KOfU5Ctkdd7umVs8RuGu8ncANWWEtP0S7Sa5fFfLm6fmNamuOfUPrfYBu6ktKhWjAKnHleq
zoinLaDdwZPQ8IxYy5F8kRaEY0Pw4jaV0aoHOeSxR/q66c/vavlTjWNUr5SQg3/bE0JGFvYbFEbq
1CoSj6NZUh5YLJauyapTQezokNNUoUXP9lLiE6BsnrM/Xt7+yI1igurK41eJXs9C0afLH/IR+0Tc
koS3Dw31bag5xZ/fglPSE/YWZH7FpI45LmaxOCNVn7sfrP/Q/XwTlTnmNJOQliMHFBKWII0ZNoaW
jzchVX1oq58ywlDu+FHnhvJpVSF0QosNttJkeD6pEfDF9snTWBuhA/EIPWlcapS0lsIuUXS1Y04z
NEmKMrgeEkM3O4Yia8DkaAqiHQ8sqtHrtWzCoT6VfDxNqehjVBMmCwOfy5cmLc5KkL8ndmun6P0n
idVATdvJZwbAmTni77WJpLiLRKOU5LJ3MsuIhPZEI4FS5MF1QG0j6bbp1bqWn38abjNkKYiJuWka
55BTKgmLwFMSys7P5SZhrucY8mORlZno9+xcpqV+vo65c6+Q3Yas+r9lNTSly8u+5bQ5iTWiizqb
Mv31sFThxdg4ES0Ix8dVKTzlUqzUoN/LahdnPIMso5m7LYIW+8xgY4o9T1yu/Bq9eaLGXJGswyFl
X9fs2g7bjxoUhxrCHKrGQ1axaOv0jVbgd+3Tzy+monEVrb6fUO5EByVpQrMpAUp1knQ9+nErSPoI
y9WUzIOKJJPw1y/4Pzva+2xY3Z0A12rrcm0JS/PoeqL/6V7IS9TmtyK5hyKt6hciauPLabyDO1mJ
fD6JFI+wFgPnn8qkrDdftTs5TIRSqcS93BxNG2+1pgsIpgL4KdajrpW4DzFfZid6lACkxj0QGbU+
aMp+JAg8ebYeYwSAqWGuJpx6U1YLQqpmDQE3egUZCJn5N8zi1JbAFazDTtm8BxXF1ws7hNHcUF9D
RyUYKP7/8hUYorg2+nTnw51oFIlBe9RXeP0wWgbak+QU15dUCr83oUPNb1PAECb0nQALLiJMoIpI
W+MPXVYlx6vUUxL62kAGsiNfu75DOM+8z+T5VcJSRD4vb6vSvsTLbMDWXcWViGCZzqZX9qO8qs9H
DOTImMdi/6jEWCcBhrhKaXPqZrXhpnR8OshltKHuI/eVBQP2NbXqZa0Imp5OXjccUzKV0rohmYE0
Ht6KvpoPQNC5FE+2W4vP+c2WFIUcemqK7HLVThuF8TRWWJgKvzSiErhDGMbRs/Jq/4xUhdE++Liw
8c2a+o5/mbGk1nGq0gYWJAS5d4r10EH5EznZExIJJ5/Ckl9q0l0s0dOJxX55TjFtuoVLBX9W6wC7
dXqj3wVJn9YVkeh3Xk3ndfE1h4JCzWijS9B8qrGoOIbqcmty99LKIJL7lL4CSYj4lLGhyrcGfZOc
AehjUcOzky2bY8ZKHixGfhGE7qBqeXE3yaORqWrLCJD2EnKjLBUL8UPBgd3FJECzTbu6bMaEmQ8J
i4zgmEDPm06PEDhENROSg1GpK5GeiAe3afKPMg6imU4QNiyod9snbbgKCdhApNZjXEIqifjBZ5r8
+vtWkCSe2RaKm3JPUchFdhtggdlvhZliXhkaVArmqkycsjdTL3TXbLMo/nSry9i8znLC9SI5XHPr
S3VIX0EszedKJ+tx1Fs6s/fd1BnR0EHcnpJfjPvthe9pDonu46YNBsyku9/SWKJFwkBnAR8BZIWg
S+s0rrtNerj2Pzk87uijrvOwmc3HboUi+FN8zqYPAJ0sIdFZazss+oTCZZfzvOCB1AQH91Kr2MHt
gNyIJJlej8ACQiShE2PvUsjLQrTrD3BAV6A3L3MhnYml3GfWa4pniq1RpDICge9aleY6Kixu0q4V
nTB0PS8kjzQsLD34HKVBYouRhgOf7NJ7sLpd6Kua+rxcKdO9ETL2ia6OBTgbcga+gAK+YgBpFjqi
Dd2lL4xObotMGOVymzkadQvy6Hi/ZTQxIrzEtUadbRrxwdKy3e+5z+urrDD7lBw+f8agG4UP22CW
XEXwLeCx8kxh9Ol+TnD2gsw/EQfUD0x5PgmccQ0z/hXZUIRiWkUcQ4MQdyiyNL5uJqQE15V0wHjw
+f13Cw7C3YUAVd3LhvViY+cgYuSVsbhDDO26mtvUHnuVmtIpvhdB6TDlp197hGUNsXPVpBW9r2Wv
jTOm2wGw8EKtA5MkA4cmD3bMvJEmSjbxfDj9a8N3PUN/hS5s4I6CHAvfewv+lfNbSwC8+SnaQ4HH
EHISO8EMDe+2crun4qBs5qY+WVG1rN9gd4GFmW2P9yCTrW7P96cLQ7a/O4bRd62JjrjPoalSpve4
a9ktKohG+ngq9ROFmpqZJycDc1jsHn2auoogQdi+aZJ6obslDd9+ZukbvsYrWLef3uY3M3x9nJpa
K44HLqDCqDCXZ6Abj0+ZcE2gx7qfCImUG8RrwrIm/g2p/tjpf+jfiC7x1lU49jR5SiTfqoPKUYt8
c0GtkACHCXSPnM74keF20zdhlcd4PZaESb8XbIwEFm4QVTfuwKswRb0dEcf3pxB017eEibn32y7S
X3aafoZ/VBhQatCPhXM7Rp3edqDHTfEbRx+fX8nyWBDouXqozMeo/ZrOrNYB6DXxUvJSqWHh8f0D
Bo0GabcypZK367LROFAw1C9wKAtV3EbSrOCHSgtdp+qysnCk9JwMwmEj5Q4t20F6kaOYu3be6jzR
C1SuzEW6q1QucmMdR/t655AGCeia7PUjsHUyJ+viVrFKOWEMK2v0f5evStO0Uh4pICd4SGF0m07F
TjgqQ1EKJ4v0B+huY+/825K1SKPfnWzCuDx+Bv9QkwpJeSCRL4piujzXdzLibZ0D8uhjBMhj28gV
wjTPT5pv4RUX1oMj7HFXJihg+nUG5ZZS7oRrFh2I8+0MmY8b/49C9pVsNU0VFvkVAKRNCFHVb24Z
l+N78gUprgjn9hHkjBbnZcg1BMlDilJhQ3x02hGK0UW7AdzF+i6hfS9FSCjvS/jPduX87+VejVh6
07ckdIN5GlrRw9p5CzEQPfIsMPyN/1r1EnVZ7L7Ku+pHHfuYoLfNU1K6XtJom+6ytOz2w/gR9WPY
egxfd9a8kyv5QSzCyS/136Br93AWm4B3cnSSI8NB4W5OD6YSbhLo7STNfFvIOLtMBqos8L9eKHjC
FMpm7G744yp0lIx7rFtAA8RpdeWKypGvbk5eh5q4yu2G/r6Mqiw7mvbD3Pn3HWewe6MfKPDMyXaP
LYqWEtMxDcysKOB4tATA98YmQma2ZuxMzS7Tr2vg12vlgtXk8AwU20LjdR3nOc2hdE6jNXOem8O7
VrKgY+1kp5cm6YWkmZkFmpf0VQEOVeoNmHhmas+Va7SuEFkMYDxnStSqVcf1cviLCEy0x65gGOer
CNM+FrtvDLfTWRQuY/zZDEXgrqbmDGiAj8oRbA0eXHH34DUx5+BJ9v2llKjUMUnPRq70h00rJMcu
QpG0mKxxqT96Hv7dEcEv34iCMDC4XY7m144sxIzlOV50bPDnQEmn5/JVp1LbASxu0zTwm73cxwyC
CTdCTGTi+eH/6Irb0P9rnRjYe5J2QcRDAAArxkddyr8bsDIEjf3uya3+DI4N75AZuV6LmnLiGRIk
46wqnvtxEpkyBXW/RqzkB3jBsAHroIi5gSPYZMWla/9Y8FaMUr+u/rT0SYGM3hsQMWgPJmJHuQx2
7HUv7vu1kUMr9GB5Gy5SFTSwV2rTAh/Xb2fkq8h6fXMgoPeU8qOtpTjSWlFKjkZ3mrzyHw+ivZIV
yi2vNfjSfjOnGFr6Au5zEUX+Ka26ub5CmGDKHvTDI/5BxTxy5Q8p5Wx7cQKG0Md/AcjvXaLPiD1S
lz7vtf0Xhk35Rv+ThZzTZGSOdsEQ/rKsNyZ8LnpfC7a/07/pt+jo90KAtB1Sd4XAZiYdDFdUBEGy
yJLGHcRUiPuJcnzBUhrYpp9z2ZitRMMKZKsxS9WdgiEyfTiJmRny4DdRlQvujPDrWUSF2c1OLOas
b015+i70nUYwv0nKVTIGX7mGrpUm9gRf7KsJGW0EHIE2PQbTyCIWa4N/SpzL6xm/ya2rTf+g7N9s
T6f9BMpA3zBORN610/u4S6jvvjFjp7Vi3clRmuk3LvAvIinvJiM1WcA3P/OcLBoz3tX7+s5Dz3w/
qX1427Cb0c5zRAt1d4Wvt/yFVEbDlbRbCb+7+ZH2AUuIMdK1Ic4OkMbzW9GMrM4QlVlvPr7KvRPi
wZpe1B4Nqw+V1eUX6jviMSNnrVCnZEbpaIe8DGV62rhM4hEabiMxMjyNSyChpz88ib9T8145CKEB
sRqRBZgT2TmpxqyRqNt98W05YJzkWQ+uScJL+4I2tKT9FWjSutuS9McBfhSRQCLx3fbENm5cTT1g
kI0vbpFwI4sZ/wJQ9lk6qSNy8iZmhYWC8EJqhx54hM+WF634QeJmR8rvXt67xL8KK7FtlTOuieTw
dp/A+dtsIQOYBaoPUUEz2RmbnkxB6QjX2EezGHDHkQZFhlrgxpNlJfnJX1gjie3Ldy9LLXyFN3Up
IlimhZXcfN+PVTn4VjVB4J4iYs57w5v6UU0a01+ms3f3RCbFI/W1a0ILxwnR6hFv8pd9TWZex8EN
iRYdfc5zlrols7y9CKEedd93kuKTjIpjunVoMfmvvVTC/Uhulv5yV5YXBOs46MsHk86sjxccfSu+
FmqxbEiExX1ZR9aNrXOg5cTjiynLctpSfM1u0+ZapN5NyQGoQVtWk7brGRFucXqbhiAoZJbCy/19
w4KrY495l/6fpgjiZMU+n/85z8v3elfkXHYngQ7zje49/O21CPJhpGLQnzXR1a3OEkGLwUEyzRjj
qmHBeWYZoQb4WVB+AtrW2RjvUqO7MekFUX9mwkqFNTnFpsUw9Q7gGM+ko9CQlG54Up61aBmlkIRD
V4ATGZjLMhd88Xs2URLQkYKvvXPyFBrMYRfbH60CHMRFCDjsiLNkQFSZWANw3BobrZkrjox0cFWI
4iltXw8veCK7QT5OApGCCZ7aV6JwMK+FYSTX2GHADGppU4c/X5TGmX1rEeb8o7tOCFyPe/lBgTEd
6F+2UZn/RLqeONlwT9ZJN0RCkJrgfHz6hc8xvgiaNh6GosN3SQYCIdr6ssdO0MQR92X+Csp9IJwb
SR4A7KrLKCrRW9ITGd7jRV1tBC9fIDgdSi2/17MJHG9HaAe+c0h8NXOfiv0dgG91A5UV035eXrGb
ZvqpB7p+Yl1+9tdvOmy3fmFLh0qosk6bTD5EFO1axla4AG3PFEqiCYI1qDLrfj6kbPfCIFQTBEXQ
nGNLx9y5y3kOtjwWy6llX/HA82Uqf79qkYRTBXbJZOOYNYOpLqJbZ1MoG0AfEnRW8bt5awyK4STL
AtGHVmxU09HQmKHuNXVTcWxRuOrRa7rWDcIE81Maqk4weh2FAfK5BluRLP5odoKORY5C0a/4inoI
ZBPaD8w5t4biv/wkP/LtovbtpibuZ8wboQ+VodFb3NK5qqkuB/GCDTP3SKM0NyybxlUN1KHGZGVR
RJ6/uKnU4A1UypK0ID2QQgfRsc9lhfkmFGQx6CUWpi0JpiRFOanPDRzZYDpzJZ9DgBKy1m3nSaN8
zIc5ZSZ/mDldkXM0xdQhSMvJvLtlzi5y8frHSa1if4cbNq0aK/8kZu0jNSu1XQwltJpNnpAYkUgd
Tcm3WjmwIJqPSSFgCmHOKdQk+Vdklp4ERswueWqLRq6+1v0r1DJBnkI77lkb1tCBavGHvSf0HHZU
zW5sbZpKiGntIAMINe6SijHwV4ov7SvQ2JT7Xa8z3JlQ0qfll7XJZ3ZkZaRrDT1pU9XWr8pymNxm
5AfKGKxZuiPQZv8bv8q5iJeV77wDMjRAbRR6w3A6JD5qjcFUNJUcUYmv+txRR6he8K5RzbGlCJMl
0Q4R+yNzCf73Gx8OWq5Eh7C+eIZm2d1VQ5S3iwkuIcftxtlF+R4OF5luZJV59mm3S6KDIUZRrGY0
177DIAn0/Pw/yXtLDuWjYCqK1U3XD0FIuI0mGgV/MbQx8N+5xM/kwG8G5TUVzt1v53HWgEKqj9Mt
Y4+Mzqlf7dq7dbYsvVHV0I3uLIcDb4w+2m4iuYwqT6GUwfR1hIYLADkb6uuimeNMmJYm+ND7yWu/
jgLI1VkWwg8Mv/ezjYDP40NTBo8/mG45jNB8lJ+aDIWWFUP59aHKvt8LXVdd3g/1Bas51lSf2MTk
X9LgiZVy8Lasv/cHerDkiFbrZOirjzUEprekpaZa9APHNkV4zbOBnnTqy9vKnLR39758/3W11mX5
bG0gNJjdtOjiOzXQ9zeJfjgZDrtK55hcl8hW4RG7yqmW8Q3M9xvvz9bCIjS9+yS3hIv0NzilUZzY
3r19C5oSqn2pBgEFilwZnVvI9be1UTGxHPozeuAHl9qjOkqaaGRynD0ibswcIAyR8BJvSkk4HL1K
MLxFU9DIlROmFJbGkCKYX1ubG4g45czqB8bsnuNIWtJFfI6VcBPy+Oe6YMq5aq1fGrNr8kHFgELC
ybnQFENWxOGrk8NzLzhYq1m2yp4bCekMdXwKr5sGz3NYvAflwYUwsxO6MXTbkHbDak40g03Alhp3
J4yy7688xf5bZA5azzRWlBzI8z+QO3f4HRfXH9erZXprs0b4r2N9KTDOZpzlWqfMJqBUVKUD8dIG
8nb020kLF9C3BO4U18gl3ukfRZw86zDieTBo1nGQc3ZaAa6TXTtMIu5UZKXCyeQLXHHid++ILCCX
43pjlE3RpD41/PxVM8CHVhCJtLm04vXjgFjz3Vd3aCezfLogRhcFFSyZXQCSGESj2E8Fgih5iYgq
5ZBMc1VshpdLQI2reTjobJaVVaz0NvrPV1IY5C2Q5Pxf14rWELPh6HSVxiB+kjSSXL19qQ2jgQ7L
Dcc1Nzp0XOkxj1/GVPe1CBFUKQFwY7Ggcm13pMckw4ppzOqVQp67fM81XerW3XtLqhu5cUnJynUR
wmRas1aLj4Ll46sKS3UKcA17N3UcJTcQzoRQyKLNX0HNsZI9HZ4jyxhgot+mwSzVX/uzHjZqfNVo
lG2zccsd2s1n4vxYM6GlPhAZq6772rPoGZyJEMtJpeTpH2ljx+dd4nLVVGBhj83WkRscoUlUSpnq
o2lXjhf72aRN7ZMms+iwos9dFpi5l5S/87YVSo2CzYAbJFOpJO5KpA0D0xLYNzFjLXaoFKRt0aZH
kRUyzL1Ti5fHlvRCO+5EJbB7q8q1cMi7C/Fw1eMz5kHM93+MeNOFmyY3dT9mmtPfZyCVq5tkbp28
m1aSWxeEFm6fV8Hs5d8tzpwe+YUJ+jlyuhduTRq53MkDCa+mGq/MBj/nvbdw+rvMSO4xtTEx/rGC
EgtayTXxBL0ft06/IzgppGFEVqTwPcL2JzBpLoA5SYgoro7Vt77AILTzSJbB1KZ8eDBnLmx/Sej4
L3XSUnhBXc8JZsNqAuledY8Y4i91fMdTGHFAAAXBwg5lQF28WoyFJzJY305A56Bl8nyB+JNQjRVr
5BGbDmjvhUWzRnO7/GRUEjzdN1F0sGGzWOPTXLBfWJvS/Xuqf3UUbzEjlEZ/sneHq0RNsjU7JvWV
fkueEOUm6ovNoWLCaX9ZSgjOIAsmQCyKvZLBqheBk6b8A1sEwjEy5iuHSsbGwKc56e8Xxd8WzEHg
VvSooXMTMnS08IPdYWXyvHbQtvdOmxRQNUitT3vnuwIv7lSuIadkSyASHfWAVM1fFjnI71urV4xm
Tj+S432ANvb/oAWzetsy7024zNOafkaax9+Uq8zeRTBF3A8FPa0rcP+fPFV3173XhmpzWujspLQx
LiZCWp6d0nPLM2+gyTtuqULyRDHDVbaO+fk7PYPWAJOGJwYHHQOIyLO5pBDi2S1BgNTv4g5lQOqc
XcrVWTde1B589e6LlcK0nSiCGb0A2vpfxdAxoBH1v8W7CPBhlJaZhXg0QPC9mDP8vzxuFXEcnUBH
QAZ2axklrZwUR00Y1lWrxEQPcqifww0CiryfIF35ONZozSxy9WUW8oLJaNHdfC29HSoLGJ67MAMB
9dtuWHDDpn272RFZUGY74HhIggfpXI0sEBog0BpMlGLUutkM4AHbOGEyINYH2PyPAaIn6WQpuQ+x
VWBnJ5IPDyBpPUlWXpQcSt9nfy20TWnLFfJNtVF7hW9pRFW1Xs4R2DsnOnTyOZ5mo3YGwZAkmmki
c5Xzs/Puejy38nTFdzBNrA+GNLsRCHj3h0dZoPKdwl0sr7Th1Vbuho99KM03TBigd15YCyoa8Lvx
Z3NonO1O6T+plAXeEKKZHxMeY6Ys7JBGf2FiEE6MLcx6qdI/63jJS8XpqFNciOkR3Cd9mn2oWJ5G
EPFRw7bI1A1FgCV8kAqoWI8LEsvaocToZ9pxU4WC09NvM1AVcW1n79GTFLUcU6ob7dNqcN2LOOC3
Vl8JCNN4JPc034k+TLzzmgImWiYMgKrvcZsoS0p/9c+dtzevYcxwBsm1EjHB0WZUDenXXL9z4k8X
1AIKJGkyYPQCMVNJ5D8V5wtA2jIFvA13jSYJdpiGe/vNqN0anWLWDoGtIEXA+NiC7asIiUvTb8Og
TlsiJLwc0IH+4zDnqhF1NhVYkrZ8+R9O5uFQKGlfEuEMUGFt2JZm5qpLDaKJxZFpi6QHDo90968Q
SwHNk5c+f84ikG7EAzx8noJjaqUgoHWTLCuQbxXLOnmlZScXnB++30fHio79CSUxE6QAX4Mf+ihM
O0ar5shIDF8Z3MujpYUfOrJCRDz2xXj4oUj944qdODEgPv9PWRwIn1ccY598dFBLP1D2eHLhd5BC
H9hXMxJAkFTrQxzTTEPGn9F6t2jpwTTPuhUL0e+XAZvQyFynPllyuJl5MseBA2A7SToMZSfk3xig
TGKE/E+j+HIXRL9c1MrxP/xJZ50ezmsuX+/voJWvmvRXi0K/0SsN7f7CuuCi9f1iD0fJ1eqt1Gjd
LzXi98P/uh1jsEG6+w+2AF0C7uK2uw5pt7Ek69FcMYUmUJlzvDz9mfzNTcGd2YssJqkM3H2dO4pF
XS4C86znCvYmGQdPhUIkwItCV2oXTpgL3pcZwRwSCjBI+/6Y+nnfwJ1CTCtXMyLFFd7qTedXpVsx
fbk1DXe4zUhk5B+zDgn62Pnwu//y/1it7QZGIcQW+CWHZpMzmpoMJwP0kfu4mPJAa0/BLU5XW6VM
pflks/ODXLHRW65OyhYKNPs85X0MsHTLFOH+UVvaRkDrfkQ1y4m1GQiigOu5j/+lPcD3etL5y2fm
g7fv5/MwxMuECLSMoZvqTU21scgIir/Ejvy9SVcEHYb61WoCg6sjjR6mWqy9iAdR1O0pgixtKncI
nm4nmx0r1XCsEMphcX3DUZiVWss02v5ITqeO9+2YYxkniX4mRYhe5x3zIoyaRa2VBsMLtLLw4ohg
RIBXBvnJs8UicbKjWMVez2Cm4nBUi3eAesRMLuEHIVzUGGkqZhaUUaDjZaDM8Y63hoT+gd6r+kIR
HaYoCFcgc3d20ZNiHYK9ZBdK9/ehJvIgLG1+RAu2gPpj90bYJqUkPEBn9700cufxCE/nT45b1tlF
5m9UmbO3xaLzRALwxqfr6gxKB1AmL42byG9wE/vlb/NZN2gce5Li+gs1iH8cTc1jA6cvoLoCifPY
yLjIbHq8vM1vTijzGDaO5hFvBDO0RjDGlOAG/rSxn2xZ9tlo6wA6jRghYDzdHjsgSboKKvB+YgUt
5ZKrY+nwlNAY/Y0A6g2zk0ho01qPpUezscGNrCb5YCbxqxtTPbIQ6B+43S2H/HmGud11rjYhIeDu
5FMLVMswUlXWgAJmgEyAA0lz1ctKyV17VktO9CVNKI+Jl6lZ8TDVDq8nbXP+VEUb3GlBxKJxrv98
9QnJcJbXvQ5x9psgxMiACHWC6W8VOXinO5NGpQEX80NbgV/+tQ6XQSxqweBwoywJeGFCKC9jmJYf
Ouv/WePBlOZSDY/jTWPYjXbZ0/QWkXNjaHfFI7ZIDz9q/GCM83A1UvbWg0xl8eUmmzgaJOxoMC6/
M6gwFywgAsI5u5b3/n5iHqb+4nxS0DkhnFxfAkTqjRsijhGON2F3W/oLrXuN75P0sbSoytGyo3Np
jGzrvqAZ4AoHjz/z+ilZYS7O+qPuGF3ZICHMi50+kl55EFP05NlaKu+5M1GoZQURkXak3ZWpvi6G
zlj+86akv4f6MujsJ0VICCiZGXfar4wiUKnKRp+pX2KWZm66ypXvAzOj9T37lYZWf/BrHbcoISAZ
VZEt9PHJWyVZhTs5Csd0dwz1vgQcuoeymwSlfgTPbOgGNtEukrS/KLfVRjSTAGdPRxgdboMXW6IH
0FZErMOrgaqfQWlyeG2eFmacy5e0O7tpgo+yDqKSjEgGQzA5CL7U34Xxz6RwwEzZN2gU8UGo+IZm
yuBYTV2vnWScj9aExtQbi+Uo3jPM4qmjwTDvbPkKEt0s1qxWxTPT0zCPI/lWbafBRwrY0rJhjt1n
cob+UYOuQmN6GFQjNgZaFS/TCPAGqQGQibRP6MisNrLv/VRuVyXuTApUoWKHENSqjMgoGvoQyDaR
S0TQUUlDRYA7TkHF7kUOawN0kFfZP0KAKfkTs2ggMvZRt1JicfnwPtwKNlQ9wWuR2UKh0Cp2l7fm
kRDoeTQX7nOeCKyUuxdVLs6DVV4vqwpCpTjHtVM4sX5fAPwRAnmgc6U/fPiXlinofDJYS9mQFirO
KHYi7iLWbMneN6+CQN6SX+UvNG1nFoQTuqVuCn/4ADKi2DEf2kCRX8VEHFEb7NuVKaZeHH/nYWke
sKvEjmwsVPmn/kOhQ6TnfBI/9m1+25FYMKxWBgEQ2L+FhJ+5RZHQ9EbeSIFAdSCgrGH1+XECqMf0
cDpOqJkd9H+cn9TR8+Rw+wi9MiLR4cw8ffKerS3oQ+8rQpfkoRQuopnk+8LkYCA8eo2vXBuh1mzC
AiERrVF00oOXsv2yVqai0L/qinF64HtevBbms7yO2fqq+ISM3AGM4Nruab5QrY0yclHQSr8mPp75
YGhhc1yMFkPT5FeSxvvD/oSTFLCKJES76do5D4bfnKGQ7+YJhgw3RV9ZU8uF4T1h7LIfko2JYLYf
Gh90fjOrC7xys1fL1ivU0MwFLxyYG3oPsC1QQYeFTHwHg08Gt3cMqknjTgWMkYFEWCsKR+WQe6ck
/7ghZILIys1+OIZj75Or5DfD7xtSWGqS48P0cluDfx1v4TI/9TGgwQ7S2PaikznW33MfWhhe8Ufy
xRRHPhcyuLtDkIyI/Ascx9X6RUPD2ZloCLFp1im/wW9+8NUVdu6DYjQWv79ksGnF1uZXWYaZeNKJ
JYovUl+3lMwv2t8/C9qjxKuIhCoRcsXyhVwlsDthvgQjWDrXJvBOaC31BKqp0hAbZmUXEiCv+4z7
N+redF/kqJghzl4G7JkpBVIS73vnD3L48dvBOwjipeqV+/CoMl7EkYOncBNru+aQzxDmsXj4sOpl
B96VtmVvgabrnu9jwpR02oH/BTBlA0FoYPsyN64dL1G7UYFlhRLUPZYbZ1eT+rNV+VRHv4ZGmCSy
q6qxZCC8PQ4Pu2lAYkYmSAwcPFPMGHwMy+qKQsnVR6HfvpBRrJ4Pnqi5rpoE5cVZmYazYnJ9CGiy
VCzrI8LDui6T8jkQO2cTsqEWE0Qn+zPSF+KCyDE7CgPjZZDOJSbqJp4FdTxmVJ5g8ccCeJJ7SmXm
RL9dvxlHiLE3HecqyjU/szvF9EdssXbmGRLB+WAXNrMwc2N8YFSmwPZWGyTHHfjw/QbUSNFTA8FP
Rfv9qtRWKOiPUbSPtED0zHVmW1oliDrs9FNLDcwzbbz5tx8rhmzZbLjW1v+ruJ4VOAQ4PkUdQpjA
pEj5cVVN2m9luHghljYrC10aMykP/uQfrX33G7KRP8cqCeUqTuIrURxeLqthMsKk36pRchcmU4gz
dt/eyzpuHT/QljeLhblHvi3UyiTaSSOaRkikfNTLUj+Th3jGZDu+Mhk4q3JTUbVsessSZlyaZ7Xm
kxpG4hSh8muDvPbRAhz83oHLhkHk5nRx53kHl0EF372rYYM+rTcI61iiBFNgK6tu80xgslZWApBO
ZdXw+4Ph85v3IqQ4SJQQOuk7n9fWDxaXBCbnvy4t8fehftmXI+1O2h7ZAlhlwk8Is417/jAabcZm
imWH966Fqm2AnFWTEZ0cYQO8Hw6AA3yvl6z1oR7rHO+tD2k8yqcwWam2DKx+kMGtKNjC3Hl2ydCL
Nezs+IKaqxWf0CbIe40PkI/fqoEs33touR7fASGC8a5O7nb3NdK1q7/HLlfqexNxv0Dinc61nGIE
WgGGV5xRHY25V62Zb8bxf1golupqIkugkEolR9VdU3FKAOj5+YPnGuaBiBOUuXY8zmebH5fy0uZA
RNT5zEvEAmlEDiA/1K0yPTgYfTv7bRftWr5aQcQYEm3W1XPFEs7ohATdcIn05y47GvNdBUFsEEvp
syFFBPS4/AhSrQRXtKn9yWkEuEFRLkFDGMESkwgzDs324oOv3m0mD+lTTtIxzvZtPrEkgbYmIuxU
Zek7j0Qebx9Nb8+gY7AKPIGu4MMi+RX1/FEmCyJge7YpkCh1aI1sbSELOfAkQGKDsI5wYKkN3iPd
SZxnRIrFtYZBLHFQfEfTZyuoToiTZ5fgW930BghvLZUMS9ylbmTy8w3Ofg16aA94xYh6LsUriLG1
dLGiTMyXTDIbw8Ex4JPzEzkLXgCbELzwB/q1+keeR0TxF08m5N2Pr4g5yDvjsH4FifOyCUfn3vPc
A4mzGc8mmlA3TET4jyJNstbf/FpBJ/LLq1UUrgR7nWSHuWyhQfIey3At0kQZbX2xjIkfA3cN3YZZ
hHAmNOlKzpZepRvifcety0R067Kmix35ii3JxFOCDSPAobcGqBb4+2idSbQ+8gqFYX1lOnj5/AFC
VcR17s/fi8+VKnZktZnvEcWpXdpo485d7nOhppsreKmTn+0PFqzOdxybt6leZeGcHRPY38EGrXGD
yneN5p71FsQAn1rERGTKZXLnpRdAkrjFR0JuM6H4lNJajOWQsiPJAFMjwXk+lxi+bJFHgWCHwQuk
x8AgEixW3a3x6niSdGFS/XKTwQP1O0iNHdVd8hYT+YdAm/XaC1O7LOrKBJNkTYHKwFVDJoijD6ZE
yF4qik4utiDorQfSIYmzB5ui9tn/SBgmJVs8w7zwcRZqeK8hcx9/AFTkQjlMRwVIeGwYGYoqCedB
DwtXT04rmaEKqOjqcetgqzZBI//gj6vFHrI67frnIuvIx6GMl0GZrNc6QvdxwQxvxhEw48BK8C80
z8DLRcpweLLaDRyJA0l3QeUO3dJJCY1b9JeMuP/gykSY5mDxHTUPbswmCD3zxaw/HPpkNcxI3G31
z9eZS1WPpxSClNaVXpn/cMci1xfFecPQ7TTm+s9ASAtu1IMtva13pHwEuq7mjcmNQa73m46R8VTR
fO8iyc+T9ntHBms0PbRu9K4+YMzsE2ZJ3gWdTzboGKCCVMIAUYjsWlv8pULxqMY71N2iOKsB9OdJ
vzBRDXwpbsptaIqsUlf1C+81PjXokSFdMkZo5S4fkQpTwb00eJ59MlgTSShaDFGmOx6IHhgBeBHK
J6HkgKnLV2l/m9PTvGIIjpc7OAuMqXOWbU39KTW6NvroxCW3bmvJPsLyLVUSiw72zO3To92rD3KC
tl3e/RR4qvtG/oT5lZaHgKOSUZ66exzkBGPdeG0x4eFC2k+fG3zLhJd7Mr2cNm6Ni2Yqf1bo2cE+
f1865TczuuZc+lM5d0iF1JdtGQJfsFpe2rHTGMxM1HmRuQAjsQ49ZnOgZBApe0qLL0zcK5G2vXjr
C7SnMN6giJd1vfp+mDard1lfOH1PWY8l0SyBhUuii9JyuoHwd9rpsNIpLjHdi8V7aI7+yY9Olury
FGQwx+YbwfH/M/FPPsCVRjAcTnip5KTUSUlXhTZuxM57W8MJRuTeOXhQ9FvZc6LoI7OJ/yadf4Jv
IBvQCZrBd8CrhR6d20Z9aaeo09SucgF/j/uXn1HwzqtB5DM8+QcZIYQfSxqVG6p5f6i2GEQ/I0yj
9Ffjg8OQOWdEQwGUjSknZqoaF6voCFOAqX30om2YKSFKSuo4OuEDvP3PWLlQz0w8n8pilORW5W7n
bmNcg1F29FMZFKV8jIIN8yZfmxXcn74mu/yMGtDNTjpWzDEXvvyUHycUgZyuqf3yT+DTHgbWLV9h
GGjbOAKXYdoacLbZbyFHYtjPSUsqluvG33U0S8MrZChTgKVOIkLISXysO5p/p77/s8Dip0KFj9gb
oLC/OA9dUaxv301YH9BTwhVcYFE5JVY4j2mXgXQDMIYcMWdJgPPZlhYb7CJpde90Twe8PJfx1LOe
JYt0GzlQMDgyHoctoGeibnlKFeGzwjLKHEueU4UgSMjUAFaNnkcKvBc/X5kaTBTcIDyrbfsaRLp6
3C7VL3IHaUdVFqJGyih76RhcsmRw4NiLpyQy+5cHPB18TbfR6HUmyFaFr+WVJmR1baKUml8X44Q1
9tqKvRtW1M8CuyvIGnEfFssj2dkNCgin00ZJyLjwUKS5Ucc3YMhAnkTZ6B2o8Te1Ro02wfiDFnlj
1mfJ8czDHYUVBIxrB5Ue7N1x/vnwKM/8V2dXKes9UYMOg5XvoAodsQ1JKRafTL09BQ9DKet9AfS1
W95Bhqu8UtQufWUoTgUGTvAs3NR93kaLti6zwUIBk3OU49UjOHjBSUM1cGTn3IJnZ5V62ZvLessP
jEjtSn3UIfIH1f/UEOpjh1ldnzxd++1HrqP5csz66jAb2uouEh4cVLyizl00hG6G1Wo5dquwzg/K
mjkH3oEyITwxLBrIpRx9elFFgSMIIMGK/AVTzrYwgzZBxT5ZfSUVNwPMxbZ5TZZ4zDQX1IU5qds1
+KAk9W2NOu1f6YTkhCYqiBN5d5DghUvpsYN95rm5Yzac27Ijv1NT6gtaDnHlA7uldG1hkYKB4HaK
rRGj8Of9dFD+B5JE8bdtvpS1N/35Je8SU1h9aoS30iz1RlyUK/kbR+4OuYG9Oect5PtyuuZjbsru
qk+D2AwPOPNxY0kk3YtS9Hqi8J+9CB26f9cL89AJFXySFILIEfW/as0qcGwzhctY+Gd5d8C2P8UK
wWMJmCzR0wPoczTsdyddm4qgJCcrwHucFj6f9zrpfX/zm0awiVLLM5Xwm3xgId+arnCe1FzD6Q4a
lZzrHto0ZfGGu+szE9rB6ImrYqbrQxIxtpJy5y7VM5gpmmX9MLT4pM7gtRycdzCrxzM80q0P2rj8
w/uXA/9dvtdvQvt+4fSmCY3d4RhqT281yHMfvJ7nhaWXgX1UKVClzVxH7LKLfBptP1HQYl/8rbEu
sStescwdcR7OQZxSHWIEyxCnBdf8bEaJ8ns8vQhHIBDIhNJ6eZnbjmi0fbsRAEw7hl0Bz2zdVebh
rB5k9L6pdcOTlakZWNx21fSK4IOqvvEuoRMwzsqJeGcd4NnSVK08LMWKi/jB/mfG/LeyhHlrKMaH
BsowFdm6CBf6B1KL0+ACAaL1T6LG8smUK9LyfelF1Ii5evUoUb3DovDDxiNCQbRrYHVpFyNytWUS
J8kDTgfV7NCo30/cL6QHcopRiyJd28LAimiQVmg08BFm2SSJW/b9C4Uja1zgPXwrdWAVWqd9itCL
luuqBIcnHeajhhhDz30he8CLyLfyqSAAQEysvg53h4cwCADHeFwjSGeaecJi+FsdVM+5NzDVPSjT
lKQ6atljpPeZLvy2K8zx/BBlRtwblkpgts6YW+1dXp6VOjNcegbvEdHXlc0oEJotni1oHKHNunmg
H9QpVlFPqo/0sXeI/JKtcWc+vx21uhZ/dTMx+tnaO9On5JrW7Wqa3na3tWP9Pq2UahHwwWNT6kOP
gQqyD4Y6IlJ9Tjpg8AwlT0o4zQePw+tWiDxMJYz2upXpY/9S4bgcGIPtbwqkU2c8sZweytvSu2M5
nw9/wedq/dEndhqKEbVc2pePGmtaLIH3pPsaRDuKz4FMcsiTNAyP2lNEZbaEY+D8oKqDcFmW7CIX
W+jMd0bFYazOe1sgfe2hpkiqGI+UFkGId3uAb6CFtanCmAJDhJ18nVd2zMAUhCeABrW1tBogC6KU
sshLvCGMlnZlW0i8amdRHfXUCdbpy/7oQzGWK2MEVNrJhvzrIYQjNsxp6gUKZx5yG5XGU3+DaI9H
jJoBo+xdycOhu0zssjCYZFrDxRbDC8woFNZnj/NKiuHxPAe8zSuEwiK6X3IbK9Ng25f6ZuUPajZ/
+UmO2TSVVjH7C3qO9t+w1CKytYE30XihhMt6D4ax/4L2M7qmRdYSFD4JojmzTdNmRdszZRJ8vuh3
orCY5Y1syJLWkYOqQoD5dvrg+CfH16bTde+Q19EuXVADCB7Gh0Ll0vKxKp+GOM6I9Q10gA+cZ8sS
o2b2E/lkeFML4PmO0/5KoLVdxbEtXeWsg7O1GIdFQ/NywK26yCByCRpyiY+QGf8ifNvhvx7OrCDY
YNuiKcG4X3mcPn8LnJRUXgB9mMC1rQc6yZ2WNIScrjZAbvSGr/UxStliEwaAzlWzKHCizsqV6vaM
vLYKiy1yLWPTv6KS8cByxVSaXH29OpQFM3DF80ijDkIj/ZV3wXNZTRDTpY0PCD1I+o94LNaxC7iK
BdoAxZtLLjuD6CQzbY/eFjhx6hWqMCcBZnFFams3cwfVk6yzpCMCfl2rSywIEfrhTKfw1Kes2+n0
iFiRm9jMy2GufV4nSyatZYxfUgRi0KJ5ePPBe8xakeT3aZwga3cTEE6BV1PWtvvD68bnbn7Cte/9
V0BJiP8iJCGVUdTFAuqomq+EEphU60zJZYdNYd66fiyIkOgQQvk8SL9NzD+brzvhI1t8b/x8nbHL
/XKh4QB70ReuLssw6LyBzAsLPrkHeB5BgSX++nyzi3LNCsMrQj4ov2fpmi8q1bRYqoJVExhjiQRb
hcTAt7KfI2rMSJKTPdEs/SN6gGX/JCPjwh0P/nrqqdGUVLONm1VagmAANeQZ5Op4Ll71xyG9hwbT
s54RkQRO+flxsTLLi6eZyW3wo4JjG3cA/0Kq4/8osEPURKbx/Lzxmscmq3znb2QSIcihMvuMZXed
M8XEUWHIUbOg13FbSCzEcLZL3Ua0pr+IOFYbT5BkRPi0ESvsMhIQkaxScw2CYSQ3iWNCEjOr0fJv
2N9NLa9HqOIvEbbAiFSOTQ+ArOww0YuBviBxCyt4YeXYvwFZ136Nt8fTo37MFNyMuHs4ghSb6OLm
Ki8UufyYpmEIM4FW+cxpbC4wnst1oASUeVcT7f+36s9UHIbxKl11sqfy+skYPmvOjdv2KXJhhGPd
/m8ijpb5/SHCwpdVbPbMOIr0pWkilQD9HDMNtas7NK8nF84oXlfv/m5nNDZv+chwE4pPbRQPU54z
NHrWSjX/DuByczxyHCxN1UoKRts81uFC9uIi4G3pAecWcGY6Oszki7ngibuB4gEq0yqiivnNgzA3
ZCLPRM+8WdndtS51Hx3632H5TuHMqs7oYHc+jIFnSSnGpAAR/w4Kr1CS0hettF0k5HQPiMMpBLGE
fppCQUJJhFhsTOyMXsJGtMs5e6o4yDtVkf1/k+om5DSeWSqlei4vJAspxuuJaP9bowcE+ethVlsg
XMsb/dSev16hIeH+/zo3hM8sRHS4Zpk1yVCQHLK0AOwvECGlVi8+m4h/g1TW5Yb2Q52fB3Ee8l2o
cccl1WT7t9lo2tsXJsgv/3Ya0QjiC4q5GoSJLJ8fkfv/caK3iCy9y92soIzYR0DnUgwvrJzG3dcL
cEHPDeCW3h/hbD7HMzMKlAo65tID1TjHX7e7L3NFm1w6nvTEWYP81Vk1cusxclQ3mVIiVFcFpAGl
iKpDWYhRwSfCPj/3ZAUhal90uX8bp838cu1A1Po333ARL87Kc9Ci9k4vePARVeRMz46PoLBUlx9n
ITuKybdxgB/e5jzIV8jbtaNfhRU+2b4GOVMfh3xR76fZkyrmH0iDB3Ac1OSM29oOD1kcUe5iPCCE
/wHaE0oKTsW95X83wQylbRNtTEZNmy5hEShHnVUX7YKX9oi2b8gMnI5cpG1XcBMJO8BhzLr6By9i
mLcsGa7Yj+ftQ9S/cl5L8Bt5MvURSvTgJ9tzb1x+6h/L+hUlRTYX1884293gm/7ufDiemUZpi1pr
GhZxe+TVzUN8CLZWW0t8cPrgueqtINp4iZOSMZq1YBK+nyRYHx6Kw6vEnt2EdRqw+K/mEqrJM0vL
A/B0cJ977GHgRRVtNb6wWCjZU7AtJtJ2V5L25cGt3nIidVmwZjZGWq5Fn4ZkgNx1DjZ9FCQlMpBT
tYa7NdFVZzE3+iutwz25zEHwLoetnm2E3yK/aK1UyoKEYskfdLI77oY5kJC0HEIPP/4ub/WGTZsR
nlJ7GIMg6QDCsgdi1IR7a9AEqusOvjjA7LlCcTicJ2HOC7FwdCLNq4RD4DLzn/PKXAvofqpmcHIC
Mk2znP3WJoW+RS4tPCJoMq9hBJEDsZt6T3iJR2mDMHefUs3UtyAs/Y3ol7biiYvcFz69cz7Q8mPI
CV0XSRaNrYRy8amJA+/k10vM0mYRMwv/gY7lSuW7cpZIBsmUROEGuLe0NafyjXcDIi16uHwRCWcz
FuSJiqoJF2XX86181JYS0+OfY/e5uFd00FCHZO/yk25GcUcdRk/yVfmwN/2tKZAH9m9VyFxlyS/L
pPV9JYZ3GS6WvYOhV04GJSRa21GZe63UykqIPY78WMNyFlfchuTalRajlvuDeqwpB1pHomQ3dGgt
AtSapPfEJWdz+H6i3DNiBjqtp+LrnneEOL7Pvq99C0wKhtQr9Kc5iiZ4DS0bd5JSCf4ykp1XteRx
FeDCGL0KAFuxM0xAasZTjM937VIpOnFZfnJte5SUkv7H6jVHZwPnPbS1rk/5tZieLyxBdIZjiQsa
hNp3LxSpeDrvlfDu/yffe0K1p6ok5Da04Ut7JFp91S/kBgMbGKwjjlrsDzYAlajiWoqAErIL6Ewj
kN74RgcZ+lcNua9aDJRWMQmSoPRzox9dDhGX8OTbCMyUlw/Ns83OPoM9L9uoGYSEjk4Sj1tNIGNm
wWygNUrNjWpER8rOlYHbXEjN+Mzt98Uofk6qDUfpSx7v5+bDucuKFCqcPsflRrPg1GaZkf5sR9hB
I8jEVc26aQqEslp4d8k2tjMP+qRmwk5GAKcpN+UALI3FClQnhGtnZJ3tWW7Aoyx6pSxXZwFzCCLV
Nm2jJNhUbrO99yyZkYLtTFB/+T0m3RXffbmEcsMAYRUI+02ltd+MaJtN7CwXCaiQneoIwlZsn+yz
nv42kqx/Q5d/cT9MD3tp4gCsnBFV0XaxHotQGILr2roTIvU3uS1zC7hxTZSVZx1iMoq0W1A+N7M7
j9BxaQR+REmxhcII4KdbfWrROZeu9nFkilXMcnTc1jHVCW/LNFwfvpEm4RWi5E1lf/JOm5EB+BRo
hzVwll9xl/f6FdKGFfnnZUynpRaTzBGy4B9tpf5x4HvTLkIqr8Ne/uMN34U8JPelWB1DhRfrsfQD
Tu/GwhYePQH4vRoV3K9SxL9egmCK180qfMQIHtBw6YVep37cct4uTmGKocvRPG3p3YQxh8RDNb0A
LfWQfym+aXC1IcgY/Lmb8bcqPc1gdC5N2kgrRrzIp75qM7k2rvNgwv2DWN7K8U7WnUG3L3dBIW0Z
MMWe42MkD46g8zjRoapRQXblBUn6JN7wvMrl5+2nV6yCZnPyUNCcESvx7gR1i01bBwHuFAsKuf8w
e35VLdnE8ZFzCujUNqNDIoRObNRSy7Tcr2XOwAaRHOBBP5Uw14Ii8uDaHB1Cvxr8IfxIZruYqO1C
BLVXpUpHkwRA6TjeELBkH54P1+zq8rFBji99IqTfWCTdzb63/NWtFBzlZxlFUQqnOgZ6BuHUd2be
ghquNJE6Q2v1hmhoTlOp4rwLcH1K2S3Mk2+z32nhWgxNtjARMWqW5wtcDUo9RallVU3R4gdF8uF2
vNlpiEgKcEKAdeRczR3yLdOZreN8Tki3cpbWgBdGP4BpeXIW2CFLJ6VWjx1PURr8zbhLcNHb+3Jl
/0X36aBDjZjWjLLrYcdjtEODL7DU997n9JvSqx+dY1CwpbtOvxqTwqKGslrdW2SXLCqC0tM3sIle
4TcaEfAV9N3w/uS2aI5bYZQ9RiGOSM0MBHozgW9eZbWrvhjVlD4ch4s9cI6s7VWQmluuOkF1Zm0M
oqx0ksPjOaNr2MAOUMciA02UBO++SJrp0gA6KubiV9mD8cTnFRH/C4iVpEyZmFx0kFbbCec7cMi2
CdYQfRpVJXl/7cjdvase5nfhwZnPogG3ad27iI0v1AOymW1fkMwNcLv+itAWaXg5+Jn1vlM5Hw2/
jHRojewrrvI9SBY+f3ZV1UVOBxBjZK3b+IsvZZ8n7GJ12ln8Sat3dmORcvsvH5xgA/bqyisHf7Ux
OgdI3MZoaHvzW3Jm/tvHrCwm7ki0ChSdWjDY5yah2RIj70vd/7x9PN5I7cudIvROhnMkKYcm9wSK
Jr2GbLgW9lIazaP47f1BlYudxstWPjgNTPjh/Kk5P+Il5i5/5015KEXOW4eEzsr22yxmHHbw1aSO
+Ri+fAUIaAh4hVMvnR/JkezOwQDNwSLsE8Gva40xmWX9WnLnyKks4YEZNDA2iSIgJZWuwCW1/MDS
a2eX/k2sSHgAVzg+fQLX6pxTPJ5kezTcaN3Ki77orl604m2GtIjbyNDmKhzWfauCf165Q1qo64rA
GDoU1jjvhPm6qJcRK5vdQ0aK+qxaJxXS31At2dHJdKTyxqEkwEtWcucIkcjOI1u8RdLVh1DrCh+g
shL4nhzC0VzzAZ+3jAtba7FkSf0cOJrdpZ5NjcMJjMgE86jxMZIMRI0XcBqhzRfqJE/6O06rJccv
23U1tRreiKT4j7Mj3uEAiblpF3625MQBByhY2bFGr9jI2RTRC8dXR0tP6HTQwFMXeeznAggg4HZo
PPv7F2tId5xZkzfpgJdMQ/vzBUrNYzmcydV4sRPNpHmvvNkLwmslhG6Fuo3LmTF00QKN4t89l8hT
s10Og338TXtBnx+ARZDruABVAgR/KeRRICvckwWjqC0hkU8EMQa7nOY0RgnQhFhLOM6MwDVgXOnj
MbHkmPEvMjfycgbwKAVzXwuOE74TZ13lmg2RTDoAVdPusUZA/Tx5oBEB0LH9N2fKtNNXSDCnxm2n
TDYxt8z9te9EtXncztjfI7F4Rbi26w0ZVNXBYv7jhortnz2vsobLN3O+dK6267k3+FRR+1pS0vMg
540euBNVtAzXMX7OIYTAQGAreSBUN3TFEd7lpUBUqI/0w0w38Zl+A0ZudQ0n7grdyXX44mNymGWE
QOVNrr6rnrVBGu5ACh6KAlvxqgWuyQDUvEq6EeL3ejg40AaXDXwlF9PYeVFKA0dYpJHBcAeJLyAc
h2OZLDyulq611/JdiMgtoq2r8u3so1sx23MImBhw5rFBQiizwZpO81KjsmCTe1tsvYpgSX8oOxOc
3gBwR2OOtzFiTLc41vIspwaQ1V3lMBUToWSZ5laWORhrmMjzRLbklNRzhZDPJ733WNtIWwfNUB9p
Rozz9ZOSBTBMh4IMMw0uJeSp5hcjGfo+Aa6oTJwnohBFEw5ZFU1Z/vNelaK+VbwmMcOQcXistnBi
c72BAmm1cZWBe7qmaX15FNe+Co6MJlJa6hBG/QNRwlo26CevuC8j/l8WXjt/Fg0LSce6o7LBOdky
vyseX2WxNgoa/rKxoPWIAkhPujC6M3RoSKJZb3mfbtj2sg7KMY6EtWY6xR/QCrDDM/BAOqPxVOgf
7V/arUix1OsZnUX+EavLwqDgObm6F9am96TWMpCD9UP+MSVoGTD0KdaYpBgxx0Tq8LcQkqcEm4Pl
ACQDo5Shn1WkpBGzMoVAjE8pKnDMquY4SK/aXO3Ym67VIxr9VIFyy4QHZya5q0YKxTvpZpo52MSs
sFLKggGfLuBFuLWpo6awvfVoUi8nOQoiJrD/c4iwaS7FBFDa0bUnQ16k3GpthA8UQlRLZxjq8TMv
PSSlEHZdytbJpnEP/WfDtRgFL8lEJS1QFeoiS5GI0kA58ABHWHireJEAxBQ3g4pHsIiWFPqp+K80
7mKbovzvs4URKhPwa4p2UDBYDMTeEeyKR3wPaBuGEeAWgCWmQI6xtX/Scq2BFd5edTN9AhXs0apk
KW2Do5sPkVw7bYiQegAG0013msys+oPoOtu+qEpCrE7c9RC1xemlIjS49y6/CYmFEvmzlLCN1X3p
Y/n+riO/fGXdGU1u0a5TmAjfi99LyddLPHco0KHkp15CyGO1+32n21UkeZJvCvhckG6IFAZMEpU2
AizctZL5K18asD6tR1kMW+6GDFnzjlVG2Uy1ZqSv3/7sBKUhKn1CLE+wvuVwD6judDmnhsFGguIO
ybds8qRq91wqog44tsVKl6PsIAOKdTzkciIsWc1BMofgx2QWP4J0JBOdPAbr9AeCQiWCMWsbJlhY
igwtLs0ZrKWgmt5SuNRjkTBtjvalUBvPa7s8duu5syxTiVvIYGnuBqlOVoK8e/q1qdUe7cAspK7A
mFXyxtlAq2X8BoGx9rJjlVwnOcrO2kOSFul7EAZ33DmI7yMb6sO56BvHtRpkXnmMF7fTekPPy3/5
t5SIhOY5yrWiJdvCmFsXcvVWEdu9tOnLc8ZF33r8Y+HmpEjdcyzfHcnG8iBQLqoMqTAfJc9l2Q7y
ukoO1w5cUdEJpcFIQ0LA/InVNqX4ndh0z2Cyu7khEmULElLa57x/mzDu1OKAPqo6HH+sW5gpr2lU
4R11EatIuhKZ+EkJ0+p+1G0QcjKYyLEujP/S4lOlKynAia3QcgGvijxWmjF68rtLe1HrrO/X1T6d
1WssTuhAH5HpTkMcV56MAyp/CSD54plIWww0XShQnsDTTe73PY21AXvMDbj668y93eVyOkgv1AL9
O6PAj/FbQcKFp6HuvH5kDt0xpkslv+LvF5Mxz1fJn9N10PZRyFJdDtBnRDVQ0o/1wwsIHmIBp1x6
JITTh0GNh3z7TrROLRcodRedIfN48eIDVImP05MY97cumI30Mxt6AH1yx+fvGLwncZhg6c1XMeQ9
CLXO1IzZc1HC3gDveCR+YegQil4SQcrvI14L4Xg4rIYvMlljbVx4XnRaT50xO9OwUCoDjS0bIcUa
7Spn5q+4Okv2ejO4qf+AVHGbI0hcihsraP45tW/22e2sRaOU7Z12q1PTH+J4fW2wzvvk7dPNF586
jeIQ8I53Ssq+URBU5TADlSjGvuotQ3h1CGxKGWaAnH3Zt/ZSht6u8xP958XP8hpNEQGelWchIhj0
ERwKbwNrJr9jPOFtoB5kiaPum9DEpIyxe8Gq337X+L7d+f4onfdWv9CkW818OwihDUO/YjARAuWl
Jbicn0O3xVSl/OHXlXT+dGpgYuRu/v7lwEZIhPpIc1ozSYqhDaeSoTPj6/6qXhDAfZX9YBHRfbsZ
9SprhjAyEOoIXB8qDcaN12RIPSEgoZmu3dDLWYTNlstEXbifqBjubX/iriuutXm9fwc9KG/Hukt9
oEyqbcEnOWKU0aMQtpkeccpinEy5QdkoGttaMEeGNfiLzoDeT6dl/H0VySL9OBQSN/0yZXcrGNci
JYVkwEiILAxw453IMdysIa/rIHlR6GvLnJp/APA5Pa41N/fc3oeHheXTCm7HDRp81PLxjmGsy/pf
H/s2iE7GHAF2CqYqHIYyuJOfamd2dXLBa5J57iinqiGqdI+Ur55A0OY7fia+5Jap6QvxgD6sP3dk
m1NgFkJzpGNC9LFOE9CbTlCW3quZqbP2Omg4417nrDjyDPTETuADLJ5QVKPbhAlBOW8/in5tOFJF
d5YktyPA+zPYhRBlpEvk3yBhwUDIFIU5WuaI3W3g3kcx91hOs6zYrWgXrnhK41hfP69IRFDegDWM
8w4tSajZh/xOp2Dd/alWT8rR3e76Iw0bLSiUcXZTcvXOVefhIyuWQ1W3I3v0bDCFHqo+5Lz7I6Z2
ZwnW8xsSmndtkhLBYl3fDfGFt5YymxBlVf6979u4LTMTyttGFc5dL/r2ZmfmVMnHXXHkD6+/p6sX
gp/z0EmP4z63Fky9jPPerK7r9TjX0Qjn9wm/2bbE5aAC+w3xB0o60GllNh7gipZ/o4nTojV8KMCO
9qKZUcUa32UtFaOWTyoU7fh2CuX6O+l9lxNFMtCztySKjRWiz8/vl+3FrraCie/konjlRZego2k2
kZSDDLLSxP3YY3ymWiTk0odBBbrw3UfUYx5Zuvsz7zZXUkQsgzHyiyqHyzknyk1jsEX3ke5NBQ5d
tkt50qkex4vVjHVc/F3oyYLaVvQTKRPVNgorN0Vo+qw+fQVANEeGsqw+uz17jnswCe19cepjR7Vu
XSaClhs1nqieTuT36IzC2o6kXwitJxUYyzDJWKYQwFdXM+Cuj97/4litxX91ykdJtlX781GiqH51
61kqkdMzXIRindo4gqxytH0x0CaZnDh6Edx/Y0fgOW82v9/dVJ9w2Xlc04/3KGzeA+uxF2AA1k+u
xeVzw0Lvoyen9UvEMgRbOZPRl0W+FoYtR/3s4cy67eWOCbuCNNKycQTUhzzH3Aa/x4r6D177EoxZ
/Z5QEUjzRti7Jw7hw3jttCgw0KHlQC+HAbCgO9qE5aPMRXOS7+n1eJh9cAq8pP/5yYACJ7quZ2cC
Zpv2MSGuoryk2rAmsmnA1TmFSgyTVbXGqg6bN9cDygKSTsJRiW/oMFiLfmC1EvNQMQrzNxPHahhV
uR1q3WxDzNno3PR3JTY6GhCVjAtPGLO0F1vS1zxlVW8F/3e7MO9BiRXu4ivmRCHVeJEJyGPrdBFw
Hm6h7mxW8HvZuKyYYAPmOKHUY3FadAb8c041At588GBPwpv339/26tbOjoZ1rfitFqTeZtFaYNaB
mtRAWdNEdZlKYawTujQFGLGEty7Nr1fpU/DrFtNAPPtW8Pd/9Utq8p5r2eN0aHIfgrHS2g1OM6zT
LUaBcQbSaEWhavXiP3kLtbHXV11uBrr/w6oUOOOBkGJteKmPsCE3OirpmZqQk+vXmdR9Rx+8EsTF
914ihBLmqEiVfmZc3Dy1zS39CiDUBsf/OxRuFNwhddyTDzjjzjexfqpr5zfE/t5iVtToRIUSEwP3
whHBgtrfK2vPE7e4NC65MqTFbWGfcnjzj3x7BbBUBvT6yPW1ktPppdct1dv+n3Q7vuB6v6O/R7KX
pCO1wDgtdt2GNDWFg0W+4FVILh7aFc7gjORPAEahSPvnEhqOyUrsc6I3yqeC13uFH4EKyfVXsvmj
uh3SSBdCz5h0BsOJmF/tR6ScOdj7wtJftM/b4FRrcGhqP5nswnbDpS2GTbueVF/60eIAN2hueP5E
kwza28gY41wA9Doh2LhpBSCT+Pzv3RSuIR8TMdnlD/TIDj9s/BKuvZcGWMbeL9KuNgyXIl8HY28s
OitZIDE7odss9fog28V12KY4ilXGW2sujgyVWCeS6pLSVY8o5OqmxFziFYcNJq6uln0DFuraZI2r
h8XUBcxJFGsMh+8XDAj9JR6NQk++BQ0BXXhBghux0ueWCn7NrT5v/wwz7/oHB3LTCVAcP7VRQvDN
qK6Ss4S4Vb9E7NNy2C4ncEtyNuw0lhQ9ORkcnHVwHipmGYuq0L//DuhVxZVxd4YIPOB9lsVwI8Ra
6An+MojvGsUBZj19JJuVztnJZhpXPTEXnsof/6LaqHw0UbZvkh4Kqs3ScUv8Ev/SRK0bY0XWhmMU
0oqqc6sFEmkqqdNjzXZ26J/oa/QyTXZVx6krQfudpXLt9TDEUUJTlcM84SVZtuI17U55ytKxs4uU
Llht1ShgFC+Oy66LC9rFOoFeqQPEJb7xp6jqIE2gMxmwJaxVqxdEwVTOYWzDNv/Bb8Ybc1O427YT
tBjueCluZCG7iP3GgT1VQTesID/uD/iA9AR5ZYBoP9GYpGT7P5dpZo1dQXv4z6HjkfaOjgwALxqe
DzPZjo5Hgrs+2EZKUhDOnZzoU/DrZufLO7dp4Dl2MEM33/7rqV2Nau8Z//T0tzOr+LbS70/HRM23
cwOTbgxP7hn2b9oWYO0W/Wi4878rxxrsn74MiyyCj8LrEMFnoxf5f+kIbzRWHG/roVqjDJPQ0UXm
bS/8R8/JBr2EwrpOYAc6TXsiKU7JaznHfsnk4W471usvTY3lhL7x5FMx1Ocj5Bs8OKS/Dcu/9sdm
OyPmkBgex2jzarjOaJa2uAFeyEMC30m656P8wUsOOLjtBY63X6+HCAw6cyo8Cf79VzodQWATaImv
8nGyhamuhjTAQkDPE8BPYMoPRwFPshJ3Tyo5o0Q0e8vd///ztr3+qhQAn2U2vbuJJSda4288XKOJ
Akej+PavA/vDx8B2JAc8TkpUBxK1jHgqh0cRu91Tls+n6fapikpYMybyCdxacryjMrn7v8Dm9zxw
2RqwtJl4aDC1uqcdCfQcZ5BeiQYkib2adVHZ4qyKItyw2AvUsT+IY5brgOg3nWb9mt8+Ttr6r2Qz
FbHDnDsZ0f7KhxqeQmRN73w7uR5yyfygzxbHxpNSxjmli7pJ0qFcf407Zg+YWPU/RkQgwEwQAzgU
tOHXm0TU1h6ewCD8U5J2BUg7PUIiM2evKN7jvUqRk+y4lKZr0JKnC7/k8x5gnLP+ZAafHbOM6Api
Rg8HNzePA+tGgk8NbyFuBskz7/FSgyT9JfcwPTwfvwQkV/ZeUPV+Tm9Agg0A9bQITBOCaLQmNt+o
MSCww8bARlVDg42DKtPJ5oo+j9u6pCHQ6g6Y+zHGoOd1XEN9T2gbT1M8pwUjPf+RlnY5D1+z6TPj
d6QcruNEFjzTTOKjneLmB4Ctd+8uI2MyhFGIiRSgwKpEjrddAkdHsGBevKSoUb8z15v4NUO1SpiU
jNLVwWSRV1h5ztQjgwZiIe6/uBbUKxmbMwMdtZ6yDMLRNHkBB/YVK8ENEBJWIyAkBNg/x1rTSv8L
TWoeY7070hw9WqU1xx03LQZOckHV1zC/YBa1JBwlLRDyRWpOgbrvW5TQ4icBvwdu5B+DqZtja/2b
uj5KR1Jgwav4IvCdeKD5UNk55lJnqo0YaqHvL0MykZtNupDYy6CtmyCjr98sGDM43cM/scT9QMjU
RQ5pqsOhP0IWed/3mLrtgVoyoJL3G0kvx8QUGC9mHM5G59/mF/TsdMXKsmEqJb0Iep2ypKE4+d5z
N5ifUdKLWbSMhIMcaxGQjPE1UYm97M6/j5J/zDwfDRI+Vkf6+npHUrq+D9XrMPLMGcsq1oz5+IlG
zGrRDCBARp+ra+q0to5Tt43OIad1eBz22iw2QgWATeWD7/L+ZTnLpE9b1VBuKHzFA6fhdmWVOd/x
2/YnlkzNLb9qs/EDbbO+FsD0SPBYSDfBEyOWIEGfQf1hnH8B+PjJzXuOKmvfJp3XG19Um7FXS5ZI
CiFGGN1vtqaZmsg7taFTPqYk+Lg9wo3/5jvECOa4aowRune/ATxT9nqGyqKlEJ5AR7Aw6hb0Kwi4
ZxSXYsxHMnEmZ3D85/La0Sb4wk90uthKv0NsyqI1Sag7R5EB4GlApaJRE40BSTl+VxINBxK6Xr5f
RdPjk9cdqHaBKrNOHtoLjwy6hWDR65oSbqQv2ugdWkF1gmWmNT066x3gOLNxbwl8P89gGviqd8GL
cQepLYnxiSw/EMP5O0RJAp+TLmKAltvoNDsEWSpEHZqBoh+JitLymoIEMK0At+cp/ac59wOcZZiC
DpJXY72G/tCt89ppX24mmTwZLCdNWIwkgLV+jdwWsR8hbBppjx+lumbEGYEh24RkQeOnIoW3CY/t
G7RzNVsVt3W4V8BT6MKQEAj8IcAGnmlYfN+36jyRBPAj7ZHodQxNbrA/bK+fQJxiufQ3yEaYRbUg
1jXd/lvsKw+YPHlVGQhSgqbBaaferaCKXQBpnzeOfwzFm5FmecbJT9sBwq5MjuWVdQ3h1eI39y/7
f37YxOZV6j2B8xVnSc4ZpGdKI36neIS/dWahKR/jyB1MDSuw2Ue/B10RcYWpRlY7AoWKmke4vT5i
Hg7FcyYSKYoLXb7lRmCVhYBqP5y1OGgjS1yFHf/X/ema3iH3s/BnahyGW7U6auCMiK/4ipLrPEg1
w4EaKlBCIK0ODBertzJzNMMeJAhOJb/Yqegyzt94Xi7mjBa0nmEZWIUecsVVz8/zLCgV5zM8HraC
R8Ttyr4Lt0pxVTH+wEiHkM9TUlz4MV49kzQR1sLeAt1nSonajlJAo8OIyDxE0z5O0mms/OUGBxkg
pYIS2iq0KfghB8VuM70rgbsovwMNJ37LwJfDQGXsGiAGEO6h5qpPtP9L8n46Fz/XAkXHbSPVXSAZ
TfwkiZsxzJSXgcVJ1zT2MxJKr0pclZYdmDCy7tj/keFz7WISgtKWNKQtJ17IZru9m8dDeRMSYkGH
LKU8smJ4BTuJUVW1aJfQerOU3ibA7+wuU8oPCJB30kAGppONtjsI1GqJGgeWDyJ8TPrQV1WU7TeY
i3zGr2KzV5A9BrEetXR9TzZID+2c2+rWpZvfj6wjirhknzuf9wyMFDOk+/zuFUsoW/dlRrabExi7
gHwIRFEalRXZBl+WKRQXxryJOBND364QyVjNzcwU+vBBbfpMSdjoyvGV8Kxlu07hBqkmrzjUnLWr
3oiXbxjswkGF6fvVZDH6TfVRseoIXBIe9aKPxqPlGuHSHcMTdJpOIt9Xj03FY+xo04vyKR9j7qkC
0xFBhCOxwa9ycUDPOW+wAgC5tN2Ap8vnIYOsR7pOxkKaonC8uz48Tu2sei0upPFqyEn3CVGvcxlz
yFZ6EDN1HBNREnN0zMllTXs7WKs66s3vnZVAYqmlR3lUPw8/3S0CXhKMS17GKseszrxGYuuVt7wf
acqwPC9v4CKql7XzgAi8iwcX2HnSVQP0i9XfGR+ikM936Ju4ihcW45z7AYYTakLMGuuqgYDfi6Jz
M0vKOTjtmGb6AO/WsDQfvG43oePYrXSQE/PcjcCPJlY/RfPZx6PXVkbV/RpJ5ldch5r6O7mzlkbn
2lTGotW9uaHkKJC9NCGpYGPJgiky1+FLDpT08SogbNfkKa7A+aGdlmGaGqRvr4s5xziSICWjkxiB
fmg+au6LBp296Lifi66V2sgBI/WZzVIB0b6YuX2cQ9gniL4VdkNCw3onF9gVQux0FzCVKZbR9/yZ
W4gKYv9k+fXVpI7jCCZiYvyJ+47DswEz38b9Q3fKnsJ1USvlHUkSQ5KIU2lw+hH4bxNhJsR18jNy
O47oL1lgOzjF1Yl8JWa8Hcbs+Ur/J0tiXIngb6/YzCMZC6Y9aY+qg9dptTnQ63dNdS9BWNZacoZ4
XYsWUOi4nPeXFnq649AYyC2uvi8AJQOA6lRFdwxdbLXy4PGfpMHDkHIgVdOolOPYcJyN0vL+4MgM
i9aTlW4OezY8T6jzwxBgX8708qGZ8CQHCjmM3xgtJzrf+uzkLV2V45llK4TkPZhrfRLAbWLLh9Nj
1jNopAvUDLvVyPOP62NFewSgn9RQg9pyGrPavRO4GFl/sm75Jxqk4BZ68jBN1p63r0QPl5JdjAdl
Uo+yktfZ7sW6RXkAAtkl9gjLR2tTk2a8FJO0Gnq/NVmKVix49H5jVy++hs+2sqMiMYV+pji6rmK0
Lbf9GvhxtOLAzQAITlQteU5yhB5cGQthSiBONSvX3UB8lsGHmG1+JwZmCsMFK61B9Te/WB/Jl46d
FYyC8lGlP3CfpmbPDkwAyKCvLT4B9LEZtE5SzNJd96AYJrOXnYvxVffQ7cffcCAwUXoha7pqAqQl
NjGhosYKhdx4ckHFcE+b1Cx/3hsMm4XZR7HGwIzYJLP5ZxEgZAuDkFs2PyrUH7JH5jAuIptBbN5p
1WabZ/j/PPxcYKZRRtYVhgjC5ipPVwTzlAklb04ycPGNnZPpGzrL+vPv9Tzvn3zHPjzPRQBf8NFG
k/ocebRRlNV5GZ+AIqaXb0Jtb/4lsFjngsoe/h47K2AJimHJnaagIQ53huT6+YIHx1o3h7ixW1gb
gcBuhBpsYgeyxZ0R15t6EUGVV1QgDJ6Q+jZZevGPCwEiuRoqpBiTUiiB12/nlZFozGnVSUPwNw5s
Bty7qNx3SNqBcxHX/s8hMI7TRqDNoIkOwbXmP8I0KLJoG+E7BEeGJF7BLOD8O+ps6eT7kSLGAUGD
7UGQZwVPZc4b4/98mlibIYkGTr+NrBdaYMH13fxVS+z/F/9hmYrg5Ly4pEg9zKZ3261CBLuRTrwY
4HY2HKQNuKkB9WTFxJawAPnS31s1qX8QYV2sjomBRd69YuAkMEF4g2mfCjtupIQ6n2cVQzfpyKnn
VNDnGtT9XiE3+AYQmQFYFVRJBzxiH/Mli1NS9HPy5PzhcBiz/wG4Esj+YSZQYpo3M2hui/qfJq4r
JDOPubaaeJP8V7UL6O7bsgJTUj2ewjeV+OtxphqwTJa4iiqHByfzILa1+iqspvIYLEARPh4pgjN4
wE6jJCIuizWUzGHKOp0nTvwsHPq4Q8AaVUQ3mbQHTyiU+DZ6qMWygWULfuIB4Hfpiqh2IeBTt774
ZIuodRliG9ibfeis+cS9dUjHzEB0cL0BKoBVF7DJNquDfP3hpKnEq+rPryaexmBkkrjJOYmI+AjK
o6IRcGHHI1jJMOOYf//IWssd1P51Si1v8vmRwT5hQinBk/9vIn0r9yTuw6wG/LaeNXkt+98MdMo8
gBjLMRTRjPljaMqcwcqpiIlyPQ8RD8o5JLkqcOyYz5r4XrYzJuAOOSMJnC1S5Po/nh2FDIt6UhhS
gnn0N4onymFip3hCXbFRAzYNbe/fKqLiDo1hNNEvDUdKUC2rtIHjk20zlRrzPZQRVIb3gaN/kvWJ
Z6ldITfRNOFJnQZAmSy6bpPUaeSd2OIjNM+B23QJujwthwODxjvX1WGALivqxQXukNsxuyfYcjNv
bauNeCynmEugpxCOWdtBbCD7nBfYLsc5rhxLb1M8jQf3HunZPlTDoJjlcfygUsyqKBQO92FYtiSx
D6LmmLpM486qdVyePxSFTiz/rwauiS8/e5Axsj87C2KKNwSa/0QYH85YpF4XYrDnHzbxq4byIWmx
Uo2awS9ffnH/1q92nUIFyrXre0Db29jTnC6je6k3tqgmHqxnZbUvORXVsovLmTP/WtSaGL+Z6o94
HTAOXjzS9+YE68R8QK+sPrYMbpuUqK4aUQdksfanL0jUBKqu5oZD/QI03JV6ceyXl0KdyPRa/ZqF
ryiKRD9gosd8Sod6q4I6PQ4nw6WzuxGoGFPGKmI4NODF2vUysK1oRrjfCWsXl3vr5+4JRArfd6pA
azfYRffguBdv818Jwt+03dNO3BR+j22X+Fp6SqXHLMyMmEWshoQg9EeSmvz3RPNocbyUjnqUVWIq
TXo/JWUhbEhHp1Qs6klfRZg9qHhIKQaxq+HMZbnaf8TLy7ssTnyhHV6okhMoQB6Mq1JOeRmzeV/+
OP0z2J0JQ2RAGvOfHgxpGMLGn8eecyeq71mXHw9iq1HcyW6iyYln6atJtnCmvVTU6kGG+ScU26wQ
9scJMqTWJEx/EDEA2t5tYJh/9EovM6iuTcJppqEQ6eeUpSojeUGXJuYwSHQ/wPerrmLFGiJnm0q4
MEADPV2KPf59AhXsg2Ny+NsHhNbkwtnTY804NnQcOVGzRwC0Q/PZSf0ozQ4f/TOPpcyqq9s1d8oT
ZttL7Nj5daweeAjQBMAgPsGykuKRzqJdcdNotIesStfhlv/A9dHkst7NtOycl7201jc6dXvoyrJz
JYIEA4HQsiIH9w+c5NtiDUCdEkUUpBop5W0w7pEsiwTtGWg7Qlryzwub+gZCK7JQMPMBUo7P9wOo
AO7SF3M+EQbjDIw7nDlJ3hzQfMq8wsWDe1oW8H7BD3dotscwghLvvec1k62QFLU6Ia/Oc9telsLx
EGkm8f+olwrN1BPvc2sa6e3IOWHhfGKrWtYeI+R4wCvfRssIy28/wDKUzoFpklIsF/zQ1mQ/qza1
qrzUkJT6NB25hTXPu3b4Niqcw5YIe60rVJXDEgYBSFPXLulC0lt+JWuVIRSMjzIpqkMXAC8qmFob
f3olMiMiQB0km4Sz8Yvw8fen8FpFn4W9yi75J0qHoc8RShLC8dRu4nwkyVWXnlB8SAs5KjOFt7FL
1KAez8beAzJ37WrUNI+s28oZSJ+mS9UymjqxVEWmT3cS8P99bsV5skkkUMSCww0rroL0s1D2Ca8O
zuUFV2lgFAWspo8AZiT81p95CbDyVKtBbCpg6S4Ngny3RVQNpzv0w0Hw5fHkyO0VvIFGoNU69Dy8
1IgJpgf5va4ZpOARQLjVDe+tz9WxCdOphqZz6IYpo8qsQxkBILricvMZpx2L/dLtF5x2HJlCd4+V
waHK67JQM9aSSVksI4Ymm5HBaMUJgZ2kUEcdM72MmsXkKmJpvcPPF/pCrIOBniUu2HeR2Y2QCT9I
iXx3qoo22oDjxe7XnDkprMdYVx3k/DKLnmEXxh3uegWx/lpxGixoz5X50EO/MRXevk18AT24bg5j
0lG0LXmCMuWGts1sPdkJ3a+sUEkn3W9/Tll9t1zGr4iLutx3yAld2mWb08fAvlWsGLKWhuS6rCWp
PCXD9QBh0zE+6f1oLGx3t1lN5OBaC9XvttpocJoRIfikYotikYVZU4SzwAFAY4xAnRTea9bYfOXs
xPzcgYc3n7fOQpnYecA+WaZUGk8n51tkioPwlq5D5h/IbW30p8EV27B+rGoUCf3FO6pq9/ly+4wC
krhWiE12YkhBZHisyIcdIo1A5qFUWF2b4RQU3LTVBjAfbmSSsEt/8c97cSdUuuZSOePx6xZUl/ql
c4Fojhq2nZsNSdFGGSlt46oRI/XuRI22838JEo9hzLXRy4yMT0Iu2YauXt2YSHY9GugU6rJwPOXi
VRj/jaolsS6QLLitlkF+yrmV+BtrdVRD5Kjlxt5pk52WpZYRO9WYFCIZL0bNSZicxP5KNX3dQl2g
BC7aJYZdSMhoeQMUZEBhJnJnGlQS6z+TQ7dsJE7PYyEZCbBmCdQ57xscQN6kCtCZIynUfXaA/anT
ndvrN5keSNplNvzLjWYGbT/qNuE+QBmfoI6/TFgIy9LQPoF1NvhQjHNarbdCk/an8l6Khih49AEz
9/EfVoqucTsdDYU7yovtWhPYZIGgKUSTbGHM9bCjRlND7EANfRhbgBz+7Y86ENk1yeb4AJv0YFNb
yYwATiOtr2jCqRQSjaFD7ovH4qtpIq8BTXLKf7nke7zn7nqQRNqqoKFemcq4IHS+235l/3AwGBXM
LXrmvDqmhU/dTX4S18fiEvCZGEmjYM1UhItEYcy3QUcNwsKE6pwS6dWK3zVCjscs11pUM8NxCK9p
+vQZbhCy5Vr5kWZuO+7Rw6L2X7BuHOaTrupfZDAvVWrDmIXPpkICDvqFks1o5HwMHxUi/lBNrQ3m
1qqCKyYlw3zZ+C6VP1rBrge4FP9oklJpcIlm5vA8PmWHZpXzfHBvMiXcuzI+7JbgP3XmLLCgMANj
scGwW+RN7TcTJbyEwGClRpv3KgsAOOBoXFb1hjxWSsFDuTjK7U2X4VlkYYKgsrNqKTo7JRMjdWAI
hcA63b2wgaJpAm6Lp+bWth2dnJ523qDEhG3Denx+oFhqQxaYJ6rhpOjv4/elsNBEGbnxl37ycE8s
Ruibsg8gyvS10ZGYm3/jWuGULaW8yr/QkjdeyVVYcgW7JzflF0OUlUpA4f/RDY58Qq6JIY0bbY6k
NlklepRPNeqdSZmF5Cxbhv997jYOCZDbnhbbz169P1ILkml/sbfIYqibqz2h+kAbcmFelHgceEqb
UzLoB2k9yqzTCL+tLm8cAP/Wgns9hcHygOOv8gRg+GLwVsGfW2Z9Vj27BLwTP72b/CDxSF0zScaK
f7WWTLCccbiNmjAZ7cihn35IRL5Ri/abtVQ17qgpMbhLu/ZA76f4wqhLWA4jIu6QIcikCpaAB6fN
91c2YTw8m94j8I7aZHENJMELhdMkX8e7Gq7sSY9+K9urnAm4+8HYElyeQvaR09vY1NqVKxi1jJPR
V5nUChv3bXfsdv8/1zK5cXXM5dchvL/F6/+YanOJq43zwxKW9egG4JZT6fQ/Av/tg7pfO645/lUr
b92dGQPAFfezAcL2+FnLJhAtoJlmZ/idQniJytduKeCPDzYdD+BLbkc15s2rATlxV5WzSYXMDPAY
MFzfBgmvCI5cTAquOAS4zIyZT9OMlT7U0RxTSfPyESCj6m3DgujevuBdo5IDmsVXnvwUevDI96Fn
LYfLCSHaXeBCE5MEFRnW42auYV8Upt19WcXJyJBitRcw7kylJd1mo3u9kIjSkz24/LGaNvGawhO2
JQ+EYCNiOmcwY0lC6J7LrMKDovA8SGonRcTUSSpA/QYwON6NROQ4ZlYkLLbDkDZxiZAkY8NhGkaJ
rK2R2hMWENcjf6h3xe6ZYpO51Ky/960CflHxr92TF4reaYac4F3c4g2vCziAASIbXT/L294JX1xb
dxOKbho0a7ChmrR8JMxXu4BXiU+Z0SAgmz7wq7X1uc69cJKt1GhHuk7W5ChkLDvlUvN3Oy+JKXeW
T68V9a05MouAz7u3FldvGickALqgduZazf5SA7MuPHIXlsVZyiPtD6fEbHifT17UupPNSZNnrkjc
/9hKbCyH4gXZkbGZ+YgP7mKK/9T4xoFRD2vJSsjTAM/6KMbB8RgZlJBKcs2UwqPHaUdupAqUqBmB
/9YtGQkUcWYSGYVKdYxxf1HKdB8oe75RDHdMw7GZqyAJu+1tDB8awxQgB7Hg2rNZG/O3CaZBxfyC
enS1IMxdwMeRY3vCd2e4RZtBJYg7ggg8lXelOkFr5Mvv7ADqk7t1QkLdYK1jT6X9o/o2K+kpsEdC
29pwEbV2+dFvl24FYAaXN9OTFgRxDOtLX6NFCokp1rh3EjidcZ++FYmVl4QC5uboqpzArNO7Ei35
+Xv1oBHRFcMKoTeOe43v/riY3SdWAzCdy6sSjZJD7B42DqXSh7WLeosPiwMt4uHQo7d3VKyHeO1e
THeWEGQwJzRZ5r0bN/anOiQafCfNpuGi3MWYjucuDdLbkmS7jFRLSbtxvY1S6YKPKizkwHEwf/Bm
WbzhH3z+1+ci21c6xtlD4jEC8+LLL4s9iQv5SW8fW+GzIBbuvmck3XAWjIWHYAdZ/1pzGO2Nij7c
VfB1Vfu/7n5kDf2N++3EtSQ1a9Tx3niD9+ZyXmeOGd3GIT0rapY1N6NUjcsL+VBzTwO2zU0ntBoK
LXKTaiKAnRQDX+jOhSypzZzg8WEhOaxStjDk8WbV+sKhqYBnqkGh7Y1xMWWlSZMMiv8dd7MERYMW
KSWPn8dXIoNHYUIPxSXwKtWntjAH0jJzaecvLv846HfNoT4RqDXgerU3TxLFRoYXSgO3yzE0GlkO
maUxqBgInk3tQAFDofnmpDSGinkANC+X9UuGl8zvXjRDaKJaVOCUrvQhqfrhAhhwsEnA5lc9fjJA
CgvO9FRtLMXVUvxpl/+OaWXMkT9GXksoA6g0t8Y1RcQJyynJ1Cmy4BVWIHAIuwVplU5cwxVQiJJ+
68FW/W2NGwCY4QoTvooqCPUVsfgTTtzN4PZ0iNysGbS5nLoKvcYsz46vMDhMbsSANtTNKuiQzvJn
IyDBMKNvrF9Q0X803dUbabLbSbBqtUPnAGTet/0k81AZKQdaMFK9WQ6ul04v9vG8O0JmZZM2AAgE
gTOfBUHZBZLb7GMe9VDbsKenpjIFLSI43kL3ADjyO8+MeX/bIYCEIX2d6RNZWhaEywNjIYc0VmHn
zokDShyycJu3KIk8kayRHpOWWWiu63T4NT12do9SwSMP8f8vWTGcZbLyT+lVNxIHQLP8mFDfx2ym
MFNnFZqDNRYnhtrVkkwGnfbObCcA4UHjLbr9KpNCOPBBSe9W0pLOZlgeZAiFbL1qpz0zmEAYSbrl
qiNLdcNfMgM9dxCdD4GuiSXS9ydUl59wivopmIxtq80YH4zGAFJifvAX0dEopqERwC3ZIN76PZ7+
ILFfA4ThH4sBCDWq7r8OSG2uvxi1Pl4M4GADNQNWyCIGzPrD/1YqcEquUdEC+dp1P8+RiT0ShSS5
PA01bTFWCOy00UykRNyP/B9nuFYybBEqzCsd0qQDXsmUaUHojN7hh95zQV+yuymXk9nRVvwTXE+p
ROu7eEcYZR9+rV7EAQpphSo69DkSWxE9tcb0hP0wOqYMtxbcV2UkfK0lIaYzzmmwP7UM37tw9+a3
V50G4PkDSAJTMiw2Cpy9ne+YaM34wa1MfwKmVfCAhrSWkSOpV0hOVOOuYOArbWp0WqlclWxxi3X2
QGFfKBxvEClj8Yl5UYGXNFO7JFpyox6kUraoqqiQM9HD2btNC6j9ESl0WTrIHm8mob2JaCTA/BfD
iQtpOlKQwQw7HWC0s1O+avf4cpdWqbQ2oaOvnSAfoeSkzpHlug4W4WQZOnqpPGtppQTMZEVjkbGf
CHkKSw8yCCZsQawnDSkPgoWqs6B1p1A5qgCA4c4urRFcE0jJxOYZXezF4udXmvLDaBHPPLEMSgXV
yG4OyOkWP0AhAw9zDmx//TDY2+YtGEK1eLBgTN/CJCsScX5zI0nwAWpc5axnG+jtjRbDgBBOtcpf
HtrsAmB73kBpnLzHV+53x+75w5VMJCcsSEiL09ep3iPr50QCqQ0HWq6PCP28Jrm+QpI7BwSF0kGy
427lOQN49S81ABzaLiIVZampFjPWBbn7bvr+sdqbCmogwa848rX0Drtp9c5wxtFLioX6Q+8Ftton
zGJbClGde0piTX8w/Sg9Xfx99/VTEvSmwvhbS4M/syIGb6K6sv+3WelA1AhOJ9olDuVZIdI3DF6S
ePXw3Ak7DY78Vdo4niZ8iCiMySv2KxsfFFprEgvoyQHqH4Oi4iq1EGZB2ANe3ltWozXMRdy2uz0t
AttI+hYBdttE2ffBdaPi9/GDWtpKKHv6/oT6B0cA1fI/iDxw4OS6j3Qz5QpwCOlt8Ie/XhoCtlQO
7c1egXWTFr0NOQKIdVKrzyMkKHoIWjeT4kG8oIRDyRF6egJmt9eYF3bMAgMQhjJSSrjV0HV92dz6
xt5Eu74F9Hx2f4V7+Ew7QYvcHzjelFfuQL9dRZEySJ3HT/iUwcbYGzT86ubQuS1MTcpsGOtjoyZZ
JgVpy6qPiqLFYEs90hg8x+UhwM4gpdYNecIomyU47AscARFENYIw64wrD9atdNWKSZhLco/AQKqH
BmpViIBVT8d4nIY1KlOz8B7MUHyKQ0hQySq/s5ZKcTYObir3vqsE/HUHfsNexD9i2Mn1CQ5lCf3R
z2WMEl7WmpgHyYiZb3Yg+jFhE0mlZnFo4FoLZmblXqi3bXQS013mPGG7AjlrkgT+pgxZsEtAnSrP
3/5lbOzH2GwUlC0avEQ3Lg5x8Cl9NOUmWMAO0V6e8i7M6qZw0ms2sVa+Xl8WgqHIedV2C4k6ScyC
CfYgLc5IfphxqBn0oMMDWggPmyzJ6J3ePTtWfk8GyqHgd+R7LwNFs5CbkbW6Z4m3OSvzmATKbbVe
UGtVRY6OHWA478a5LJ+tLwPHo86HLfIqvNsrI295MdH8bBRs0RIRKBkpyrOs+u6zXO6i8dB/xniz
n6optsCtrU0NqlJUyic+mt9PbbTSvWXDkIpfZlIsrPqE+ibpIu4YJEt9nQ3Q269CsNbdoqdXYX4X
LbGzQTDtQmiP/PiU7cJskZR+0bkRATnTSrutAptwa14UK1lbITcKPoGm0ZiJzAC7NpEuVKImEZxM
Nkl3sIAQRumpF+5G7pdAANEKBTM8T9JNqY130NRjLUgRU04qf6U9vrqOQwctEapU0ifa5VAAsjYJ
fM5AQjA7VnsdWCa84flyv2bc/ICQqbuFjuCxVD7kFDD36vxSk6b+ySArh9ngttA6Lh5XcDagofrZ
uzGU1a+xXNYiIC2aWDQqxOhYMw7Bgk+Xch816GaVP8tZ4TLVKgOsyKbNQS8kZyMg42i6pn8cSn47
1FVwoLhvJygFNy9/V9Hnu9m1DVVtNuWM+y+O4EyTLkjqhNyvkxUI3b+D+N6wFcoTY98WA1fsNAHQ
s4vZIx6KRCZ/xxxKMYIn/M6MgH0JGuSId/ZmNjg87pRDevmcksJNzRNsh/uEkTDqrEnOkV4XD0/q
gNJFXZgBSCO3uJoSdcMSFQMZLytDzErm/0PTHkw9tPoPYxQ+gaJvRfjT3+0uN2Y7W2ImuoBJOHrC
Th+7CwWQMmMxpkmdknwX2OcZU6QmFlmp8+QnrkyJ5foxQ7KX71AC/ZE4U0hovVWE8cr6kPMMUEZ3
LOM5SzQNzh+7rYfVkUnMRj1V/SZ7BmDu0+xgJSQjPgWI2mwfii72VPsP2jPD4cfC7ktGWQjj21Nf
bTj3UkJNlv16itvCbL0vaEcHsUq30J1Xgif3C3eVarv0smJIoRzZ4MxfnEN/pd97NnVhK4cCjOtr
ay6iAPaowdetDKxgzqL6nGkzYsXdX9axdkBCL19qldo2PuosVXq+dpbzIbevZfWiG839pf+tfBjS
j/yBhOLaoUkuwRcMv/P/6D0tExL/Uuq6JV3vtoZyTuuwMOa/P4ZSEEhyp/3CdjwfgYhXTjr2v4Jd
rBJADlLo5E2bO/uFxcnWplLgm2DUWThT1l1mP7UUGOSLxHyv52KdTMERwNMM5fk9LeYbuJm9YGtd
GGIOQ+0gsmlS0Nta7m6a+UhMkvCYohkNUZKaFQrw7jUB2/oYxC0huVCWX5NvYj1Lxc8N/7wRsuEf
lUt7hTCVD+5xPQrBwNchdqs+G8vHlaoAO2vxFrLMuNy96DTOuskYb/WqCaRCkKsIgafFPDRTdlUA
FG5a+ofIWjjYempA7Thr8iLWlr8yvsvxmknhXgxMl37Fcf6dmN7hsFbizzMvBeLxHTmfkygXuUjS
WgFplAWvGHSl2t6M/90ixYjm10BAihkP3uHuoEFfW6guV7jlZ6xitAFTT4GqBj7MWz5kpyOdEIGI
XJtUKrL5XqAsObjJ8TGfmwZOtOOMr8AXglz3xeDRb9eO8cDvqNMveU2b2MY710tofqqfL473TVQ4
4/cFAb6hui+wi4AER1MfGwPBONvDKLpV/oVePvkc27uzyvEFC9y2+A9vA+SPEeDJ145izWu2bpaq
siLWe88Qz4O9PftLxeM7FMjHgalZjt/MpZZlxB0WjmtfWFz1V4+qBLdxk8rywShkrC4z/pk7Sh7+
ZMaY48FuGkFi8MpwpHZRotPLPxUlBUjLOwHQLJuERKUd9KaXfUal+dbc/9ydM1z5SKh/rBzu2kW/
ScoPpQAfQypOwuWpTTmZTKJLW7bJ+uDJtqQu5w3bTKWhOfw4xOiBA+0GoGN3CNwBrbN+1dbEEWet
Ok5shnwp0Y3n1pURtuR9nebIxTh82Wc6N0PwSgOc2lZrF2czghzsK5R2y2muofA2g/h9GTDkND9d
v517nHzhqc2uQ/OJKsqn0DG5+OfpOTSVF6/oZ5qI1XoTbc3aYMw5COZSU4+MhFnOOHT6IzztyqMV
IZxAUAMW7Ig/JKrF2MMG96STx5P9G9WVQqvlUqqpN6pgx3A/rLDkoLhprUpG2t0jn7pdv0uzv3+Q
GqOjVzlbG3mSh1WCiScdqwY1FcT4ftJY2Vw629GES/Q3tRnX0XRc0wT6/hxxfrTDU8Erzpd7cR0H
lNkACIaVSYBX8PCJcGsodcIWZNHvG79GMqvVTkdWuFlMahxI+5GhQnLUlhYPSUOJFwOq/Hd7u0ON
55R0wT5rOn/VrIF//VzDvLQ5YXCY1d3olNpJpo/cd3pP/t4gaLCa+AsmZUsS8My8Ec1r/J7yXRsp
+HTF8gv4YqDdnwbCu3bjSCWC+v+n6RTTukLTdV3bqAoQQ7iEYfft6rqLjr4QVxCHm2zEb8NQuh+I
Nov0MjVhlGGUD+KvfKxBmXqbJoLOFfomWozMMxHyAkHe6OxZoUuD7wQKXzfjLmtRPGM0L5q+N+bP
xKUCZl/otVG2YYkB1DSKEPIZmxsr19tpR+ci3OVJEp/ltXjalKUva8zsiIttfQ5eAE28j2jZ34r5
OuXMeRsveI0CuEOJd/AU0JZd6p1Ltp9oLVBzZIVVzoRUwDEOSwiHspRFXHBqHND07rXQhDE1/Y8k
kBaNgllhKS2mXBJq3yFx80pPIwGOtFBrqpC6i7VZR6sahYc+HUrtgpAcg6G9W25E64xAEGAWafXb
CgDchxqxDKSM+aYUQIsP71kvDuRxHb3Ce/I7ux55a2Y5y4cIR9oMQmCY9fXD8aOM0s9WZ2XpPNAS
ajLJImCrmOap0c29ox6ITE5kVkqXsibYNMptVWxZyQPtLikiEC5CgDgqf7ARGm2NMZOn7SkD/plg
04vAxRSXlrdaRN720cKRNzpxUDVj65KZv1Pl0qrJiB/vD60ZG6fxmilISi4x1MHncYS2NuY/NVe2
+pNEo4KCfiapLoywBxK/k1wSriZN8TyBjtG7744AC5TnuSfaLddcUNb1VnULUUEVLPDErxPGMfSr
nu7+d6AtThP0nfHetoV+sITzVMS3UT49/HRdlv9Pl/LjXV7IsVqfWg5mcDVwGOZJjg2hH571dL0Z
X5yx49g9T//WrBp6iLoTZzQxwaebEkTofnLIwzSxTGymNMML2+RVmFMjGo3uzSySBzaojPOuWJXG
SY6YmJlD7frflbBnvvPFTGASSAqmr1/DXzhS6GS4x45mu0GrVBt45hsonq0DEZAqejV4cih+BVoQ
C9yBuai4xKkYpozz7pGmOGCpMiJDP7zGRpRrCqj74xVcTHkeBOwk4WdYnkOl4LXhA+jgrcsrYct8
LBcfjUCxxByYI2MNsun4R3UFAx454Hk1KzC8TO2MKg+JhTQxcynyvLEW7lew7T0wzWJ9n/N9uj6N
a9y6Qnhv+WdNi+c1X+680+r3z1egRR1+Kbm/hqxOftehnZN4hu8I9Ti9PL1FqGX+r9lPv0hjUxXp
HmYi6MJrRxvyVP5LGeECjzGncNXNCKtJlutYUuguQLq9lnpBlpJdIxlMyL66Y8yoN4NxMD+ug1uT
WSsoKPvk1sxyJm4TVm2Nw7BgVv4RE9XlyVb9A37uFRI6pLjJxGR5q/MzR0G7cPu5gyFTvEquFMmc
9MPre4HzJUf9WRyh/HU4j+Svl13vPAcXZqevdVr6w9kVIa1FYAB8gdx0meA69pB6Yh8iPxhnoZKl
8fHlYDODSsMefshmhbKs2LEWaBiFJUTK5Sp4H02lLyzKt98/2P4TMdGrOcmYDathBZZyPKFufhIq
VXJXwxt0hbFrFWL0dptTTjC05PSOl9uT3aQluYeW3yh4WBpoFefg98lbBYwssR3lyIQ2s6sRgUGl
wrH0NWwb4pQlboPMTKgikhiicQEOkTMHscMZoFSYySOC4gWs8UjkOhq1yP0DDSi8olNRvDASeJx9
NcmSgucJUcd6bKuv5brKHOuMUCbJS56IqPK3RbVF8mplk0sc49W4DBgt96/+pzMV3ehpX8lvWhPO
t1hawa+KI74h5kyUAkUonM6nxbfetaJoJjMOODBDmjylM8pZqiSXDIsVUWyPCwf7cJjySEL3pAa1
XV781b+fgU3Rr7t1SVqZXvxFEE1VV/qBRDJYXBHsI7OBwmAPdG0ha9lF/xccdFcO9h4qW7VMkA3t
VF++XXj+xiIdi6A+jDjm+Spm2KAY0KZyb4YQ6YErK8Sm02vCGoqIMbCIG2X/nDkKjvpv4ZD80Pz8
JGpxRF3j431GTKqRAfUuTdBAJqimnkf3rJdN59nrSt+CHFjZC4NmHmc1pzuXz1fpAaxvuSXe0+IZ
I1LI0861E/KOHQdYnqVRJlQE7Qt9eaiXtoNcSi/sExvlTLBno16RV9fWGzNZlnexu56kTuFs2/NQ
szkDyeNR8bZ5p8wr0DMBdgxARca9FimKZGO+JmcQgNqsEZ1Z7bQsPxZdBONmv0+tbBbgdCiOgCfd
rJ+Z74TJkwnWXOrIGEGA/sFPR5uoAdYwIOMs/3GBy/9LaTnesH8s9ORt/719Xq8W+9MDWcyEIdo+
szNfGwlaQCmQKYG97NFPzU2EoMeFE2j1EALWXxvzxJcNieW6DYYZYEMMWvXn4kQ9aKbJ0WMePNgw
UQ41iYQGIpn+YuBEByDg8/oryltOdAZnwKFATcJ1t7s4nEqU+iStBQeXkvzyZ7YaPTRflXJQVKOT
2TDHK751UdnbtMYehBlVqiYS3mFftRA7YE0e01WHOEVX76C/rssPborPnK9b8yH3CpBX7Zh3jJ6G
fVLOvhZFbHGteg+pDwa82WAsE7iILvi3prlBwE6m98EKgHQVflpATXlqGeKtbEN7HHnHpeCheHOW
3lf0cxqFRqNwFf8RJwfSwPqFg/wYx7kmKzRqtpKf2VauS9nXi6JnzN1O7ji1iUa5HR4FaJOFkMJF
VZ9MMvvupmMlMP12DpiEQyY0lry0ORkEUSKO8l0i1fkDLfqTCBDBoJ4aOvlADnh/W20G/wcp8sde
4/Qd7VjLxlVmB2F9rP2iWBGFwavm13AQR/QSN9lNMOv/j6VvmPm9E+25RjXOqKP/OBwTCPvNtRPN
KnBETskG6Uph0d0mLj6Gmau7YmWiMjCrTiGAuEVWfn63kwv4Qq1g0A1IxJtKjoxxG/9rwzovfDp2
L/OnVZhrkybOJdOX7+j7/8yU/Zvq3QFNc0D2H4/Medx1Bpcc/VWJ89Pd740UovFF0euoLb6oHcWZ
dNsu+ry0gmgdpaS7PJOKkdujfQ4yY8JYE599qQ26dxW6lar/EIIpvYEhwED0s0X079JNVO/aIhjc
4v8hwsD4drVP+Q5AFiop8QsW9t4CuAfTtxUzEeKZikSQiLU5ijCYnHlaorX1BiQUZS1YTqfVJnQo
aqj6x5W1IytrsawL/MoopicwTMIORS1Mrmy5In/tfA50BzrtQzy0jCT036f8+ApTmiaVO5tcqWR7
L9pt/s7Int/r5Sl7dL5oP0kK4f2W2qvXqyyMlGn83b3rf1krMh+pa5/+BT4RKOwr5HIQKhngIA8+
Ai9IdoQoK+GRs/YpaLKsFec+ni+vpmvUsu48eT/pYNF0Pj1OXe2kXyetGS2X2BJ06fKuSWDV/CJw
INXwpbUyC0SzZrZYT8oahWdHgfQxuLLy2s2YSd58zuLmajsA/r/dkUBuwImaGfsFv5HTje0R6n4Q
2jZFoDQm0E/uKP041KvrATotLpfzjVeyOLV0ve7tDwKEQ+Du5psr+4wfWEIU9A3ovNMVhASlhGCs
YtUoBgTREbd3pQRlS38su3Gc6/i6cb+zqNrKufNyfOpiDd+k0YLldG4GXcFxDlj6bO9nRkFcKB0D
rLEFNIeIkoxBgMKzOXgSifTsrD0LGeLk2BY8tl4odZXUQJCJMtqpVpc14z+3jO1Q9F0D1S/1nFDd
HeAkNQPO3X34SbrlvKnVIUMoL6sl8vsrypvHdWB56tL/fiCNSbEedOnNM9ZsgldHj8cpj5WKpWoE
0TcPSr1TTH+EPVGidzJqnbBNPuW8SvGjhJ/VP9uNkXOx7JU2YknP3zH8uLO8L63/9zNM/IcM0GIm
QOcPR44LN9ofjApVjJNYyqgmWxDTsTRug13WiRJBSLVoOXXGf8B9mo19iWT2vg1nuKTZUnAc9wV4
7F8T0V8455P4jbrUcmuuj8CYWAq3cBpf8Omzgj1AH6O3As71oj51cmZbBWp/fR2J3Y/afuFqUhRA
D2KVdNfmRufXFpISDAaL/nJTxH/f22PcminEgB8I/qPIHmI/SHtwuLIZn0GJWzbG+gvUhhogUyRk
Yn4K/FIDnFldj7J6xwmUpSTc9jKWEhK6KzTxzyAVVx/h+QKvee+Yj0BHKqX2A67Gvu3n7INsedJ7
h6y4iemv9Jj/S2leOxy1mkyQvs3J2uhOpH87K0E2Wu5oZ84wYEukPhBc3PtTpcbT/vlRBdSqJrFU
Es99h4+ekFovwSbnjCBFmj2P+yMY7wVyAtnJFf50P2HlNdhEq9V/X7xMjk0th/0sXUvDNA3/UM/i
586NLR0S0K4bpAOexQs5GVN/o3H4/NbeKzvXweeksH7DvHPdGm9UbbRkmdNGgPal9/h+z4pVeHrU
Q2B96zdxdOeEHPDZkk3xBLEulwoRlOE6FwOK1twWUHAtJaAS88ZRUs+SRyHT0y92egOPmUwz2hjt
tKKOLSDTQGMz5ZQTWiXRDBw66e1+FHv5LN8+Waofe5lub/R0ay/KnqcXZR7PkcaoaTWrsUXW8+CJ
/dq9ikc6qQrtsYfnYi6iYX+uj7KnmwfNP2RMXlyrcXkifNzvHeqTgsHhV08vJ8hEg9ABegtqoUCf
+kK0JxYXZ3DtjRQT/voN+OHUJ+awSXGwxRJTrweBQ7AUunKtmn8zJqd4Rj2Mo2+g82lCVfpUe1wn
4phLFMNI7U1VFBFq8dIzlgsCD6CNyqomUM2yn8wtOMS+B/66rwmT7IbHB4bKR57dijcVifbFEgSO
LBw20LeOA4c3Xfd53yqCKuPA8pP6oXC8FZlyJg8OCk4CgIdSeSPpnUwN7dImXeKEeFk6uFbpVJy7
vnL34um8Z7qDMFIlyN/WKVERGVN9ZvO0ktgtnCtU70yZUtDNaCtfFjZwujrjK2URQumcxjAKlfFT
gVYQgAE/DK96AHebwV3xtnQmIJj9VmcjNjnWVY1H85xmZTEuIyb5bhWjPFI7/d6gohkXCLiglSvM
yf/kDZho+2ca6Hncz91ENv4vysgkPOE5Vb717V/OmrWou1g+2jkG2QL3fCy3YXMkKugHwFaQuDJY
dOthdo2sV+CVEgGUITBP39h7nbA/ddPBwFhC9TT5VrgYRF0DhAg/bafGU/QrYvCKzyJDJsQIJKjR
9LjuBknqwOOheO8Qua/KnNLjdIswcNlCQHjJ2XFeea9zw0u+AWSjl5BxcSSWYq9amd9dOKKqVe5V
28VDrON8k87e5AK7bMKUQIxkZvUNpd8awsIDtHQoNEopqEsriySsl86+gofIsFMqxpfVx7VwSczN
mJ+8RT/55YCfAya21jvGLfU8U1Rq3jYp34w5tz5OdrmW+jwD6YiuW/ZwybDkHizxJRY364BuBD9C
Hs5wC4jkl+sgD5cW6nd3pnXL9I2goiydDAK8Vz7JaLxWSdzVkYzaby934XxuZpw/b9E+703XOWSD
TFo6zwg9Kva5+Mp7HCKbguMPXAIoYlAVFENdDCpNLKpjKJCH5R1dM3dItFIiyENZL0YbFn9WXQrN
1v7V46rTJ37EUeTxUXygPP8xbXiAbu22pSRyzGzBq3v7h+wLFa6ADfHdo2HvjFn7c9M4K6U0iQ8w
1m2TTh46XUt9o6kdVpWZaT9neywEJTn/lJGbd0Q2EpZ14+4wE9ld6frroBF1QZFF6a80lNiTJ+S6
mtCR88TcjH706YVeoZCzbXnk3Q/kQ2uCuA6mQ27s67rpL7ekSnzcs14Qe9zTaMzFTrDNW2MUKwxU
8KZtJY72ad8U9LPkHNYNGj25RxwFNwo3rXK4M2I+ifu0wgmRDhZrluUIMxLfUrXUDNhlUiTVxENH
yljmMrlsPlmJVDqPF+e2/IP6v6+0PGACwQSfSQk7jUFcpHBzq3qTV2kI46M0fBCM4V6YoxnZSeMz
wBQo5Jt8r3gTHMhl4/Qp9TYRowG4bun3gqoVM/pMYh1oOEFmA1SR8XpFhhQkqrqVHqY+CQ+i16WZ
oUJUCosrg3EiTJOE7YxYML5mL7yZNCwDLoQDu9qhNQXJKIbBdu0DTJ39wLq3rkD3+ykOa0ZBT3qj
rA6dazggavylVTo9SE49DHMzmIclllgvz+L+NkFWg3BHveTAIdvbQOkaZKdC+g6FibGpeg6OncMx
vvkNSDdWAA+9UXAKA5lvR5xxvOiY/G+i8ZdOsU7IfFIq+dP7xgrbjj+5+hd3ASPHCY8uECu3h7kQ
eiwq7JLlS47RKC/tTgIeyTioulSp+LQ64XAtjfhF0yjkfY6NprYIigceNQqUTSCcYxMn1HZvdh2p
oqky3qrx0J+fSRPhomSJnBGBAqckfehvq/CA2VuaL5WnwWoT3ecOFpJgtGHsEvf86kSRKin3IS5G
ZLekr+Qk/yDIeXwp7XHQ5nO3BnYuuvHuT8ooN40q0K3OONIpazrslPJ7PVnTXz1vTQbzMXMB+ic2
Tj129yKIyESpz0LlxtfOneYOYPHHsR7yLRClY8GFaCqxT5579YD5nKtw0W394ELB3CUpxd/XHOe/
VsGkfUU7n7XBqtyPPlIkYMBoxn1OGZsb/W1Yq7xufAT58NsRNBspXyvNoYlbZdSd7nmnKJPStDEI
sbYzfA6Kznp+gZ/ULsnUCbufcnwBg9LY3cwIOOkGxuF6lw4QY4zuc7r3DRX7PbopXBKb3v/FgG+A
tTsq2H9HF18AGACAA0zdSj3HW1VQKolgFLoMizgIk6fTrP5E78ORCh6o++JXdsCeL1mD+2HwOLOR
Yrdwf/7NHMyvhnutru0a826X3OiAnu9T0rJmXlQc7JrKm9HOM6HWTm6pBRn+7z6ZR3B+t0HpIQm7
ae/Qbc11ap2U0Om1hvWpOX70ca8Gk6Hj3fMKj668WpTo8/Ra/bgvJ4P2kUaDq1sgryKhMsLvn6ch
7oVWYlT8jNCFpz6TVVV/Ef7hlowwV1yznHOwwg9tEBsctl2rgm/mZuWMKirNU9JznPzuYuLdHtbm
yN7yoULxVqkCFMnhvpgGc52nuV3pFKM71DycLUYM1jkZgzf+kZ5AnZP19acWROYJua10DE1EHG97
U9SSrm0+PK76XZdY4JVc3twgqlFz3Ux3U/y63p5GmHjYL6myvnw6dkcy0E5mYt3xrC+u8SiPjiKn
K6Y2Kk52WEFMVMPerBNSu4oaQwUBhsZuDIxLCWOWplDCUKanEn4ChADzHj5FwQT5eX9gOH5fm7ci
nZfZQgjYM9M4JcSD3CO7IffbxFKeMb2u0g8qAjpMA3qQ7Mah1l/T0MgfHfGHLWJ2i4FhxzYpLIaq
jU192PDmtZrUAMN8E1dkuKHQpzgi2pt/vsWlKOtdTzuVDS1/ujTNsAYDgzfWqxc/VpjNH6rK+JNh
4D0jUU2NeqdHnxw1ELruJml4IodDS5McDglebkr34+kHJG7GTEuGEnjs+RdXz5wQb7t2Aik/UrkD
oAuycso+5tklT7O2Iy7mRjKm2Ntabpf/HQeinHFRhmu3agMYwjQ+mWkbV70Mbjez+bHIsYMPOuy3
Ucm0QlB8jUSVWKKRwK/IFI0XeXQDDjCsOuUW/huGoKbG9RVB/+VuZQ8Z65erZgBtTov0UopWAsjO
cUlNxcxNd32Oi1QbZ5ieqXiKeuzVwn3C/NwhHhtbOuFLl+w0vbM86l1V1rEviaBrdAGimBXy/Dm0
463T/bz/SlsPFcfNfKyHUAX1GukNTiZHpTZi+bSm+xNpx8WYGX8e/Z+Nu2EmIBMoHO7jbOU2QNZ4
Wwgk1mH5fkfm4Rus7cS7XoN/l4Zdnync8VEXH08VdBRAlkKDHyTFxjjeyQnZtlBRGh/AnwTU+dR9
2zw0UEkYoQwf2Pn9kGYXH4vHW3Ymh6Gk2zkaHgAGQ2u/JvPYF0y2oN+4ceigFsi26AQROATkINPi
ipBLJDbUtLoBnJ2wsEpiDkNf7i/gRkEGP9Fz3vKQZ55D6raoDTHQruZk4rl6CtcTrjXmn5Yjg9/g
uavndvM4KkqrtIEwXGZAofu4jo7afFhoPoQ0KmFqTnc2E+8prCXKJUBaxp7Dhvdn2+adAsNSkNk0
j6ALQdsfUD8hDqgamyjOZniTqWW6uVETSEdtXxcjGll8FuVBvEafBdYypDhPwOuVK9MiNonQb9sY
TxoCQVfdWyaa+cKrO/99IF7S3vNh3H0op/W13jm+F4TKU0K2g3tkOfgshHDV86PV6JkGE9+Fx1x7
L4DKT6AYpNvysqNSAesjHSuIAI9JzHi5NBHfkZKp4UKon9LCr2sLlhThgd4R5Pteuwjy874CuiNR
3gRORsmgDfASDr+Qrt2iJZiR0toeIEJEJHkLMtcZl2nT75+osFvr2BqWdZrRU9Ka5zhFsq5SaThC
VX7XeJEXumX2SuRJwdPTsAlqza8sBnpODrmWp0uURqgZb0RzG8RI5PtI+0B5xQHW+f3ls20iC1Wr
plipEC+9iJR7vUJgHsF5gx7MKcFgT8HBVJUkrGxMvQ4ORAN9RuBbAkv0J3G6/gKfVZE1VLzhfWY+
Rzy+foC6Mjw42qYRHw+TFscyb3dkySE3ssG6bgABNuiMNLIg5MkPKn06NSMpifiRnXARIrjO5O27
XqnniuVfrftRzRCQifxAVKSHlOMlGF7g3nzUXuM+QttOwZK7eCDXpgWD5PhZAR+y1M4xQdNmr73D
cf+Yq1eVhcXHW1YeF2YU6S/k8Isj0tdP/DRtVf9IQLWF2biCWUngr65g/dZzj2xO4jLaMyLfFyyc
hm5dAQPFRzsMMIeYatuilpvC1oolEIvuIWLuoJpnYliY3qDU9hhu7HjfpoxQFIuTyjHFaNErJqeo
Frkcnn8OYRtpcYokC6lDRiRJbvvhv7lZW/AG8wVXM+0EwyNf9YS18TTb0Xv8c2zZOrbqgxbzR9kH
vvmWWW4+JyRdi1965okn17Ivl3ujXPVAkyCJzE5pPsPNsIpEiXA5N4kpwUikf09LFcNSYgb6LVQY
ozYjxA3gxAG9WNbYryHbXMTmBtKhrGaI+57tGDnmff5BXCTwlSwqAEwOAgSHCblfZ91+zYvaGBfg
VziqCnbrmcvJloDBizztgrFfxuqK44ftd7g3omDUf1kiYvoOBM3k5V6/1MA6jtcexUDodH+kqiTq
OJpmbL4ZbfZh2Siq9S/BscJa+Njsxh3qlI563AIk5g4LjD+o1Wsqb1H7WZGcOXOvdE/a4Pd3UvqD
dYTksQKSryrQfDIFnuc3VqTLiVSJnO6M6olaK+uKDQcPii4Iq9F2GZojOYO2peH1dRdSOFHgMnbs
PhKh4bPlI0uKXXiEdspj+nUEgN2LnVAyRtVseT5DFMrh+c1QOmHApz2jKY6vBCfRiSN+PskQ/D8m
q9pFKX6DAeUmbdp9AvxGUsoLnjtoTHbddq9mY3/dTe2ZyGExRc7ydzI9wmkCWOPJXQmu7h52xcKt
mnYMriUSfyOf/g8VksqUm5wpEmM9oxGoB9B0CLvc6SOcasV++32gFlVjcMdVpLMxZ7W1H7YCF6O3
LHz+BcAggNZPAu8XuEYOFal2bXHhk979q6Z4QtHFJ7A2QpIkcV172tYkJ8WALAgTGwIoXga14iLH
YZWbkLma5KyVtIgiqq4bNVvew8OkWlQyzfUVuPqZdw4+A94roecr2OwM7Fvle7yMD5O5Ze7Yg4AP
bs6dEQeB7IFT2AEqHXDoXhf+47pT015LBmsiGR+XVLVEoAytr342siAUGoS9PDANV9Np4DVQXYSt
rz6J8jQio7+xqKvrstJ8Xkwzqw8YRyVZxdfUD5kO+dd7uIzbgkZ8B9yBd++3sZLiZnXnqJCiTSRf
CDrN+6TM5v4E3JVcTgSMl+TegM+1j3TvMNRpWxR+yU1TfsnN51rwEmcmWokrzGgSTg9YZ77kCBEQ
rADUu0GpZWsX3k+C9o/DbyORTuUm3g2uYmFZVZ+9LbNkFwV01VlMTKOqDiD0rPDvnkqhmL05wqs3
bkknGOJec60Y13Uyxd5Qo6gfEczLCJQYZLcU53GplcaOOsCW+p3ti7Q+z/Y7iyl0aofcOb7bqQm8
YGVgpB2Emb+IgTvGaGUuc24Uo3aa4HVYApbIffwmZKHSE1sm5ZefekUnW+M81QqdAScaZ0j2a3ge
n+v8TIKvqfN5o+/dg2loiN+N/Oai9Gs9ohYbEbHqrWzWEhBOOqyb2Jwt7rL0UOspg8uFK9xc5mze
UetZFQIyyUjRISL/ZiU2XCycNGj7GGcdq1ypdQHZ4GL2PHGKLHU+rjglIOo392zuBcxHQ7ZYf+p+
HDlmy2N45/8DDdNkIzfBovXaRzuN5Zz/R3UHo6tINtL1scXAKIB+CJElX+OU+VMt60xmXBXXCApe
k4y9c5NuNqe3qaTxpxuVb5kZU7d5zHJXtYqARwqHCFzOMZlgLSVQ2jdqaO9mwu3jjPYLhoi1nA2v
Uq3CaF5SvjycFBlXsUtCMeF6viSr4QSwrcnNODVj/8cNmsj4h1w5kCz83bgidCEnCO4p39krgGEk
2fLExRZJ12wxyD+Hac0UZo8DVaO1Tsn5qJT6Yp6V05umMeb6s67jwQvAwSYUlxISwWvV8i4Bm5gQ
qMBzyevUoTF7nEC9gugoXSXJvHNdzZjJSUn1VWZa837BKXVkSNhA7urG/k4mdY4hUfD90L3kO/Mz
g4jk0Yz8RTQuMD4KTFWYel5FRmqx0HepE2hcDQxvcD7n01p3mASM+7YLnB0KxvbGBiIFKQk1p3qp
5FrnBuP2/8yLjBLxYCvD6Kj5kvki7ayNRXUvCvRHsDJdPCsoDI6a0WtNFZWSkQSiX6QdgnUpL8qA
D5UpD8g32/IyKuVvv97TGK08WVg2LxSlzkJPlN3FC9LXcNInkfnlf7Pt3Xs9myvEhqeXVhUE8cVu
1D9XSOBJzCaN3guEcQ6APPq03GLdenGPxSJEn82fkZOe1MGhHtK6l7QAmBGZ0rfwTvpnf05WDGmU
4wXJchOkhGV0kKq/q3lO78idpFkSDoIOqMbOIuEaziUnS4yWfQfRLPlgfcl2+TiOmyjihh0ZfdWX
Tblz5jaGigHNwcscptrbm2I9w/36sogEKT1dMfH/o+ys8ddgE0XIFlnyAzbt8ObDaMGADoqYPsL1
ewpRbUR0HDu8H5tQgJMKTrkpgF6cUWftMWAcGAsOmTO0feJntfIK0r9KVQ9Fhs3W8J2J00DNe78S
eduRcSvnMQwvz2iCJB/Dh0XtlmUMpUdglE07ChqSOTHUyvBQhysSGMPqN1tM3M0tTJr4gFNmKtof
BIYMweXA6sT7eQ75MQF/y+LDMie9yME92RCWntwhiCTGiDcNfrVSM839W9VxSPDCXJ4MGj6UwKXo
TTsBSDgmsSu/XAXsaOM1i6UhsXCmlXcv7GVCmkG8ucP+OTUgrH8nPjH5zzEhZck3HLked4nNc6dn
LnX82xeF1h/f+yjw9cQ+0N1EsRqKlSVLCalRMJDgLi/XG+sdLlBkljEjQBKUzHLg0KhYnXFPuWCC
n7fAyqP7XxCBZ4FJ4lGxREyIFiV+WfwzPbgtSLwBXuh6YW5sEIp+4s0MynK82PEs7nTNwhuw0KS8
a9NOh22ou6GYSH+YysunetYCmegxIujJSS/dIA2NfwNpIV4E8JDYxHJv1XF1xLdkqejWoLZGccZS
nq4QE1obm1M64dRCCfn57gO7c4K2glrjrO5iUtJl4RGj1VapXJNAhuN+/GH1zXcueHYZu2V9rJTM
3+wonORimh+TLCusNV/IRQXsyJqjPdrtCWcwY/FuxIMilzH5L3vl4Gwqroirxttby3la8UCc8bLB
dzhwO1MjtAHYY/m+99kXR/ZPd+z0pm2VJNyO1XxczJwk4vDnLXH6igHA7ZBtL9ep7VzI4WvrPPAc
xx3I11rbUcHhnWrFOfUgru75k02rUmI3oVCglf35l81YBbQ2pslVFxOcl4iKZjZpG8dX75Wjy5kE
1znGnjlLgVGl0SAyJK9oqGCpQjoenDOKFGTsJd2/ksXolLg6QZaPGLZOx5gZDEVlpKx8cctI7AKs
KZHbMYaVUJZWYVfO9ANOMz28DAFrjEK54jEIA+fqzFMgo/DrhsYRrfTNyumaJYwT3NpXThz9wWgr
JpAKDk/6+gv9OcECji3DsJMJwOHN40JYfVO1ixDqQl1bPlwIHbV7fTr217PJU3I1hjL8pOST5/aG
0ezQ6J3w3ItcKf5eeT0cWj1K+heRepmwk5rxDVg0k2qusZZIjF5ZXfnvv84hm/eASqiUrDX/Jo3I
5HunL4b9W2TEkyoAS2MA9iuPZn9eT19VSQfvap3Zh2q2CtfguIFDl7foPfFi2gmPP/tEeNdc9NkK
wEeYQmv8glfJBiMb27bQ+uFA98ObpAZh67fZLaehutpJKybhAwVx7UQDCCgD/gD3xdLectntiLKA
xm/nfXbBOGQZtQuzu0WNCx6be46jAxJUdO9CnCnOtkvO7ZWm3T8GNl5YCSPTYRuqGtPb6o2HMbeg
Zpl5bCchYtJ/aIhq0ghO8mDPnuaXLREDhhDotlSaG2fMg1DU1BrUOXeUnWVy9ahD993zFgM0kQWC
nRnR1jcChoTA3t5HUyxM9ytsMEiZjKQo0DqywjJ5rZp+IXQJDatknwmcnc4iYwtWiPqfsYBPwyv0
TmycZ+qMDRQKopC37j23J2mfCvcqbjqZRsCZIWZYzKQbeoJcgWru8uqcn1g8znf4pbmS6m5Sr4Ta
BKdierTKKaUdXw/ctDJ1UruMVYAwYiUqRRq2x/veYEI3OIfCkEQxRn63V+wWW5MCJ+U2YiZbuBOU
uTq9sBW6Hmcx3gp4y246yDahFYsSyBm3H9RloMQIIZbJTpXKmmpgE+oqwRPw85ygV58Y0gg6Jyaq
WuLPy/MnVb5hOaE4843jSdSW/OmoPIzqFmMptvWnxaQxOfEc9BRUnoa7DXQmuATWWOAvi/4XsbJg
haPRAfK6vpTopyOkSdUAlqgU2+Zjh85Q6pKYbGNapkpVgakb8XC18T2Qa8mo52QmHfU8PYl/4Gty
eCtMSnl7+5esptKSoZnBqLk5QC4dyTQUmtRvh21qX9AuO9TavBDwgZxXxbJcdrzwA7POq4ARp5xk
a2yKEs/DiFgd0Qb+dbzTNdnOAocY1SVmnU++8Dr6Z1eUyooHEQU6g0lf+vneQ+k2CYo0RqLso7qT
/buH7sjxO6e8blSIPEcrWKber+UWZR90l6/IJR+P32ma+3bx3QPTqOgy6tnztK0G95/FNrZOM6hL
9RclG1THsPeCNqsHFeaKr0SiTwmtEySO7zKhtOG/yQXwSPad8Q77ZxdH7JlTBXvfPtqOeiJjH2H0
t4cETufCH90Vr0gcytMRyp2ndijsMqAHSS7vpmYF877Mhqg5dyi5xqFIi3HhWsFS54GNy6SgOVwt
0lprGjD08u3ikRFy9gfySHzgSdXXUmvzJ4KFOFadWOxNfIp5aIZfeF8OmtyY2D3jJtld9NCeY0kg
WNgaWXAjDdgF+Po4VHb2RMGB0lGtte4JaxrUguYG47zNyosR7DZNb9HTU+z5A2Q6s624ROvlxgaA
b4YxCGBFhGVu3BIcy7qZ2N/dhaYBL0xGLxkerLd9M4Xcwovnxv+ci62Qw+VGOF8EBKUSOtiuRCj/
hcncDp+3H/KHJZhecwGU/2MR1HVXKQEyIZkmSXx0dUM69l9bl7NbbCTAxDQXXEtl1eSffUob0yZk
KDz9C9XAa9kNjv71Hjk6aahZPR6JGzFHCUyfJqG5OcvJGuAZDSMRmFn9WlRqCpsMENDdby/JjD0q
kMNsFBXEG0B/3s4Mx1tu+Km7QAYlg69knokiPCs6iGwzveUU61gzEtLk4IGlHSnDCGCXNH+aHS3N
0yFW01XeuUyQ7308Cn+sYhMmEPVccSIM2u/LPyBV5g8TXZ3tgu7+8mfK0fdJGzSBII4mMsX/K3YZ
VeCLq7zGlwWOsbJzM2re0fVuibeZlx/gAGZVa06cp40S0fGMOybxH9g/MTYoMad5G+pe/xoBVL3b
CUpp72oj9MSgN0ABL5UGX9s9aurbNVKzXGX9F39HgjzVsIG7+AyzX0b+5TlVf0VnaVXqQGcM4ZQ6
ylKXOfQnVWE8m8pbV6XoSWMjhSiubfeiEoXEhl3yKKeJE4kcOZXcXv++muyKs2qdJ8C3qtYGptzS
dSZf0gIhfd6+KS2cINWjQDSTVxNJwUr243yvQevW7kNUaEYYHSdUD6d6RkLk351lNhamY/LhdSTq
JijpdRAeTV6w4mshRMwAZuBcXDghL8RM4y59qf52gO6qy8e3nZAQLTdNRPIufiejaJerbqsjPgnk
GkWt+QZN3ukD8XvQxxV/ihe9gcYOM6aQdEEN6ZBkoamb8zPFjI9eK1JCpDmzAtbvGtUg5CWCN9lc
lzXQNJZ9cmeFgpdRySAkGW0Fj5V4rOifX2Qx++zXST+kYYDH7svZIYTVGfqHoLM+JF3TN0J84NBx
RsNJ8ElXlNnVqquUK64gc2yewmbsNguLg/NsPNsfODKFG9ygorinQ6zbZgE1mj5Sb8xuoLySQZs3
cPlokQ1C1HSuheqZnuHiqe0J9EyQpyEYok4QpAIhFCbGPhSmgywFZTCZ+0ZEoGmbMPw185PXR1BC
9i4z2E15/clZpZjVWL10h/UXmuIz0TNfYVD/1oRpjQpRUAXwDrUIvJ+BVFmN96v29LgC1oYjyECF
xFzx4gPkN4pXJOO8mk2X+f7/f0hB29EKbH8Durr+su97n2cL7XvpKOC7E6jgcvh6JnUddJx73lBa
7gkawLBb06o3BwPB07chWezc1QKWWX4FihfvyC08B6e9gnVmS0lmFKKfOMsPL9mrjBP5XkDBxolA
gugZaPtqSR5rnwa19Z2P5k3eaXusNBHqFv9k1tmKnzXZIbibp2VmcTaCWvPXkNkW62ayaCSD9Bk4
1qvGicNCAl4uSB/kiWFajB8XPAthgJcPWGuraM/6KGiIj8Z4Wk746YIJilUgVqtdAi43W8kP3Gt0
V19Q1ypDwwdI8ieNpIyrx8kpxAWKt0UZs2SfTKVwYhh5lVN1Dq6sUAH6BKKDr4/4LVbjcvpSIPcI
cnjVIgktfGsOQ5Gm1CkTDNnlE6uLGmG/8LraFzyoED9LCmGSqGCDRlumxgumiedx4VFsU3GUnRMc
4XsVCN2JKoSdqGry9ZwQpBwQRp07ETioExqNtybmDH4+TkPu5cuZIX5ATqkP/FQBusz+tOmzwQ1b
tWaeqh4C2CGQtVxGPf6rhkzGf9hgwxBEXnkxDjUgCuR8MrvIMW0hwb7ka7FfXk2Hx6XsdJnY0gjz
8+bDbhkiJWjgKB6Cngwkpg0E+KVK3DbfjPjFpfZrJBCttDhJPq6Vtxfl9FgWTMLKVH6W/VAT7nuH
hAC4uQCWj3xpKsB2TBfowzJNCfFhZXUAomlU3EgkbzocaV7/2ZFaJTPgP679bRqcO7JOOn8wVxhB
GEpOYfeULN8E4zZW8qtWab0XVy/veTe5P8mXVkGU3QZbbcQGv5nUq3sggN3aGGhY4Sj4ar3pVSNn
BNO9jwNLnp0BvyhkgNEfMgQRl2mwdJKpsM4Ul7V1SeXTOw8324sdCKsTqlgPoq/W0whhmXKoIGVm
5BHA/BqVrQxvm0cHUCNFHlL5OwBXssK4A2ygTiUWjV5P8p0PztcDAlH6dXYs04+YwnqtemLiPly3
vE/QCikU8BCt8TkikVSP1flLPsJu6w3/1YrmDIhJl20uvlH0PosKgcBKMKFbgUcinjjOr/0JNs6w
FORSXLjJZZyAnNjtUP6pbpk+2nNn5pbp7G4fUM+bBW7ZfWdcjPSF0YQHnbZrR9Tf0MdncMBEXbiB
1ePREnMPaoE/IQIrt6c8+7bg/uCnFCkR57lmP7WyS7EcOgj6YUHDeaPrWl8LyArB58aMVhud/6I2
tOXSoROiZPqtiwrTUeCw4slbEqxLf/g4g5QQ/YHB0g1iHLuVFND29476d67Cn/nVdSN5BAHtoujV
XDkTzibmfD0sR/+mP0vSMxMNe3wmI0ZPQ42PEsDxxxOQZgrxSahUAWavn1gdEt16VD0UIIdjoLMG
ohizwO0ONjgqDA/jLt9gyW9XnOAGAWjBIFyK2cNFcf6l9y6WqixmaUoXkQzIL9rf9GfJyqnrthvk
nb5ZsvXumzmWY7jtIs7qSYvY9G3VkdCk66mcMSBt8NMy90pNaxIazhaBKsypRqlpBQc4vj58BP6P
RG3BYQdcOzG8lmpI0l7ut3M14+3t24qg4sEqgiQw6QHfEAajsya7ci39Rane9O4LhBKz1fVSAFAj
l3HZ5eWkNOuwAyZ/ilIRDDiI8sOz365bY3DWVXVG4Km6j/NYUqtXAe/Hv7WPVUJ3FQjVHcmS/KQl
augGT4upyCz0ZsuunUhvj8FBXMRK4t0KF9GThI5PZJAY6lXVXAjfTT46LWfOJ/FLrp1+yKL7BptU
btcVn/fGj0gfdK2FcdLu9zJTvTRj8W8iUnW4Zt7uIDk1mo4JlzwopzN41bdJ+PabnQwAiiBMc+Bw
Vlzn9BdDmL0lT4gFTjrqy7sVjz/iroNl7ishqY+I75DLTbak7VBPGntIZ9BAqEoaZcQhSt3uvgZr
riV6yd2huonnW5YwkJhF/wwWQDpDr7JSyfdZI8lw8+9SQnr2zUHcy2u39fROueSw8TnMkg1uZ7Ho
riZppUUmDtjca1v8JfnYsCr2VXE6AM4q0RqAfdJBMdwQ0NKgT4B1jDnGugJu8WYQogvdoCLjf4Vf
OUW2IOr3TU5DUeEnKan69VJU5iFnw44hj3GwDlV0LXFZAVZs8RKEEEKguv1NgI5GcgkdQvA/8BkU
eo5j67ff33fnZN3Nn9f/TkiipnV9U3z0AKVDecNldb7SpOlHUwJSegUBKRbSE8sG8T4bVlhGJr1M
xgjNPLMttIHtvfmJUTWDn5IKcMxuTmxFt0ng2ak+voc04vlmv/SLJXf4wgsCaNzHtM5C9uZSQyY6
ZzvsZz6Cl4gDJhCX60ScCO8MBXDvGhnZI+F/K/FMdXZe7vG1gPGJqqZ2LbvTwqRorwEIX/RqmyAk
Ak102hBiEA1nRziC+jW0010/qtLnUJzgyxe9zORG0pOb/ZXtDAL6qClTpQgJavdcVkTUdEqhv8U7
nlYbFtRWtBA2uAJB2JMqfscI8SZikYqTWK1jDk0PCsy+3oQJsK/jYCf1epzFOQ1B2rv12S/o/Izl
V8WJxEML1kl+B4Hi8C7gKg9Lou5M9EzqsIucmK8SLo8BbT3j3bp9XwtklbmszHiV3/qJLXy+Z49f
RMOekYEeflmui1HBsh/OMN+hqwB7oa6CzssuxoSOguw4BCLBLLf4IQb3SVhAFDaoSf0hP4BJT9tM
Qz0g6chl82co0Gp0TrjCnnv/2ko6N0kW9KwX82tbEIa24wpEqeFXULr6eyWgYHM+Mi8psj649fxt
89zvpKkmHKT/01XbytvTqf26MFTx3d8Ys++bfDce26FCUrvbtzCEZzUcwLe9FKdGGwObPOOljGv0
jxRhlw6+gUVIUkyYXsvtiL29VOTHXc+OyGAfc4SLJE18GCq+4tQXp+KWmKGtLpJfvZmYyqddSNvl
1A73WFpRICT9LO5nigl8uV6esfwxzdhYnacCG/2LXKFcm7n8/l4nxvqUaniYGH5Wdyoil1Lx1r8a
oK9AhGc2I9df5ghIqcujpXskKtuFArTMi5tSw9LYUnbtkB9nDenicajXy4HrOTF6VHgoIGRYo5Dp
zUQK1lKB8zjvW/SaRMPFsmZLK6pprFoswFowL/0fPmSYyN+0ZfwxYzOenjJc+SA1cZ4MFx/ZromH
CdXF2ktXjScCwMDWzQ14TbSnmywLcTdcuQJdExWN8T0fpezRWzfqb6AlMTwAio3cyXfwzn6UtxKl
BIisz/EU1WA+Oi1FoPswEHVXmdi5y6/cNElk9wHTWO4ZrVwkWQ7maErKM6GJWrwsE3YtnHqkALbF
l479w7kZPlgqf9vpcAm9Z94pXlNvkd4tDGiWPcvUxpu1dWQbmujhZamTrUpy7OK/tSQKc2gUUB4T
zuCpL6/zEHwLSKSeX3Tw6Xy+EcXslvD6+0sJYZKJ2d/6hZwErxQy0oiaO2RzIPCT6r3lcAjORpJn
vJHWS36N12a7cbaPVak=
`pragma protect end_protected
