��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����Ղ�@��G�(!w:tt�M:��VA}$�zȗ����e�uT]i;g��`�\Q~� �k��D|�����7L׹
�#6�J}����н��Ա���IL�Hl]�Y�ȬFE�r NUN}�\hS�,�[�Bp���O �b����ɊK3�&��=�B��U$�&m!5��F#�k�VZ웮�����i�^RB\�-Ϲ��F������l�+�ǻ�{�H��%�O�RG��;��-~v�C1S���K?ԙq@���hc��T-�G綳��>/l±C[GVi6,A�����_�?U�A�A�%u:Zf��5����7q So۳�&ܾ��߁��?��^&�[<�S�D|��-��
A��L1�H�OdyGc�9	{�㑗�z��R�h<9�>�������� [�p*o��M!�ː�/�&;������oYZg��W=R�A�<���Е�*$�Iæ],69$�vEv����blq�&��'C�IQ�,��{�=ь��F��ɓ���'�q<d�)GB;�A���W�k��T�lv�922+���N�p"z���T����sg��c���lR3�9����g�h�v�Zf�5���Qe���F�=w�~s5�s��E!����N����O1�ou���V��7���܀����^	�	\́��ear\{����5����F� v3=�WM�0����p�f¼M��~������	����a��R�	3�}��&��AsN�r�����wOYSm"��f&��X�M�u%xj��T�6�Dy�lg0��ں�D�=���d����5�mO�TB�b���/�J�����KBe��Ze�˨7���>R�>�����ޝ�y�,��d��JQ��7��(� �����~���[C ��Я��"�Q�q���o��˲~g�a�8��#�N$9�.*�Xx-g���wS0p�aG&ϕX�m���Հe����6B&w5	�)�9;��I���"V��-�~x����8�����ñ��߈$�Hqޅ_�1Vp��D<$�rQx��v[���zԕ�2>�)e�mᚲ�v���"���p�rOѓ��g��B����4�<1am� l0�����pd���7`fW2S�����81��o~�� l�Ŏ��;5PdbR7�:�
�찱�8��]7�Pܳ�̏U57!����7�MO���1�3�`WqL�K[s��(C��dq�#7��)f�~��� �*��t0f<�9�e��E�ކ^�'(����j�!�e6�׊\|���	�����9m�+��:�ֲ6$4Y�5\>�
={ؾ���A����@�(�U5�z��w}�?�n�@Z�X2�*�=/i���ʸԹlIc ���t��d"4��W0]��2GD�S@��cV�JP������+X7S}�f��z]�ΫY�K�t/��YQd���B����kR�:���ग �56S������dH�t߼� �Ur�M���o��eG��H�>r=Yl��5���uI��ޯ�`�����A�F�8T��Q�D@l�,�0��HU�3n�����Y$���.o�������@���O�$������]�'�>30�X�,���7�
$gjb�n�(_��hQp+eXѐH����DB'I��"J�Y��7����1�Nա�;��g���.�϶��^��fId�B&���d��e� �eU���-qO�֯6�B#��w9����-��v/���f�n���;��}h�,Et�;��(��,K������̢];����6�W{����� )OF^�����x�g���%�\�i�o�MD�>���"��Ա��Kd�8*�ГX:�@����A�=P�_S��M��*���D�rj�z�Nl�y�D��`+�xY�"�|A�OA�Y2�))?D	��Z�JT�żo��_7�#�쐂���di�:<�����6�}�	6K+p)�o
��|N�+�y��\��x��M�*�h��j�D��Q��.&���k[@Pp
ܻ�q�Bs���~)���^�bv��Ũ���5��#���/�K��}�;��B����b�^��r�čUO������&r��k��M���A	i.ys|���y�˳HT&�t�JF��Sty�w<c^��0���M,��� 5�w���96zl��ł�����ڌ��o��G���=$��D[*&��h]����	.��ڃ���,U�lSTs�@'���]��P��P�1�k7�M@���2��|({�Pb�{S�U���ǀКB렠)��H��)�0�?:���+��f�����<L(O��=-����G�(WA>�'�܁� ��k9�eh���I-G��7nƊOڲ���e��]�zq^�[/
�*x�+-H6�=��3oi�,�*B�lRy�9�{m0�{���U/��Y�V��n���Aj5�hx#��YWh����+ ԇ�������oe Hw�Z�ɋȪ�f`���.h�N��c��4$M�5-�K�I)�dʈ��m��i���D��F��塚��ECy�-��Ɩ�us���LZ0Iwr�hl-t�ӽ�A�e�9�H��"2�Î�y����-�ca��w����q����3�>�N��S�
U����R���(����Q�2��\ƭ~T�)��9�Ϣ�~���?c	Za0�g����#0���fw8�5�S������,�c�6�݋�(��`�&��h��q�`e����~`K�9� I��A�>ᩏ��	�)���&��|�gA�p�>%Z	�:�t9b�����,G<�k��딍1	I���B$�6�>�W덬��+ѣ��E���4҆�}��_h��J��Xy�.:���!E���} ,����-��2�KX�%���2���8��mn��21�x��W�fR�l?��c���-Eer�[!(���N�n�T��vG�[,�7ЮHD7B�)��L�gO�0�+���v�N�E��y�g|�]׽*��M����cEK��</;������� ٸT&� ��9���Qp��t(�s͒vV�sR���������&)��R�8|%[����Mn�v$uc>��O����8��~��ǌ���o�G��5Mk������ˑ{+i���D|t�t��f��w^9��T��m�:��=-H�����|^�~������q�s�d�w$�³֣�!j	W��VW|F�@!{�:�`$���?�ϼb$*���ƈ����Kbڠ�m}��cw�s�ֶ���
�@�J�ĽXzXj(;���#�n]S�7�:6��S�ѩ����M)�

U>;@�8� �[����8�P �I,���Y䁰W)�8r�\���
g@�D�����"��Jy�o&��<�	�c�s3�ǭ7[�"��i0���f�϶�YȎ�_�
{��"�\ftx���}Lo�~�"�'d���i\�_?Q���723 f���-��A��್�Gع{��Z��uH�w�d��R��	����O:�X��~�0s^[$P��,1}�fy�x=�jz����,Y<�&���A�?܉��u�<t_��1�$�-�B��F�]�u[�j`��T�]ʦQɐ8i���,�������Ƀ�����4u/i��������@Qo^��.w��rU0N��<�
wxtY��t��=�":az3�����Ț�]�cI����7%��a�lދtSu��z��#� �oA&�R
E�3�
��$>Y�DV�$Qi	6EA�C����
��W��%� ��x��/E'�;�e��Б��o����@���_�� 9���(�	� [\�P��yMw�V��Gh������6�T?#�����jy��1K-��'�������6�\���ok��R���M������mu����AEv4ַ��j?� �'�^w=,"1hbUɬV�n�l��\W�ҡ�5��b&(}%�v��>b\��UX�$ʻ	d�B�[�>'��ڵ K�7���c�����7 ə&���.h��Y� �DSm����E[���U�� ���܊Y��T�ڢ�7ilvw�(����0�+�o��#q��ȪY�1�o�g7�µ)A�\vD���ͤ�vx!�?�ݿ5B�s��}����r�XU�l�zp����*&�H�Y\.��}�����(b\�����݈Ϸ�Ӊ��P��M��)@�[^c�c�qڸ�ƀ%v�Hl��(���h�k�����e�E\��<�b@D6ИI��0��n���D�d
��'�����T׍H����-�I�s��w`���/�˴F�%�
X'>�������D�fs��t���6�:�tDq�����H =��T0��ms3x�-�`7SMu�����E����\���t�D&9w�rup�I>�Kh��t/���X}AǷ���n=I4�ZKs�^� }]�a�)��^
��H��d��g-�߻j�4�ᇬ�F����Q���[���f5Ƨ�'��k=���)<��t͹��:�u��d�͔���P&�f2��\�;=tSt�?ki�<9�gP(�5l	�H�pTZ�R�/7D��`[���ա�Sy]�S)۳Pf$��"T���Aw	u@����Uf�0@@�`!��iFNT���O!�<6O��"��H�E	Tw{qm��sɫf�-��V18��C�b�Ox�Xf�[yIp�i���ͼ^`�����=��?/��e�è焵�dK��R��<�Bs
���e*TVeЉ�K�tY���u� @WS�a�z۪.�#�W��NH��K�-����GB	���l��.�! ���$@Z*��g�J:���g��.�(���{�#��Q�Q�B�e���Dk�w���h���A�D+/����`���輆�o�~�o���s�e���:q&��w\�|�xO��-'Yu*pwØWÚF
8Y8�hh&^Z��1NR��(�>�|�4�?"'��V��u�Elc�=�
XA����q�c�01��*��G��o�QB�N4��85�Ma��t_���t=��e�mnJ`	Q,s����$Bũ`.�	�! ��	9�-����
ʨ���nu�r	A=�ǺgmE���/��N����D��-�,K%ՓP���$��
{]^0-|D�>�2�y�
��K������
��a���I�}i���;�l��m���A
!C���0B��5	%jZ�$���Ou�]�������#C%ٍ6��.�曦��NzO��"�8P��/��e7,<�G滎���CD�Ş�No|_xBZ-�ë%a�"���$�IVv�Z�x���8g��;�Cn;���5l�oz�����7�� �|� '^���&����C򚒳�H&�s�PN�uj7�r��a�C�6?~͓,c$�J]fp�h[LO��R, �o�|�8'|�@�͢�	����@V#_n���Hl��:��h��r����7���V���i;7׹�[e�WJ���ިL�J���U����rjdd���i��RXD�j;<��p,�צa�F56N����z�x�S�~[7�o�텍�7O4�rB���3��E��[�+���{24"�U���b�E��A�6���n��P�;2i�iG4]<ĺ��J�	���ǫi�ޣ[n���>�q-���d~jf���Qh��mN)�nz��	xkT��ѧ�;�ؼ���oδ?2�M��W}͂�u��}����9ݶ����KG���.�yY�f�`,v��������{y҂���\�
�&����,�LZ=d�nl.D��l��H��G}zfY�!E��Y���e��-�" <{��˵���\%�޸�����?��__�~�Ƙ�=j��3�e���,�.��߼A���+h�MҲ���þ����C��|�i�'҆�y��#��[:zG෰*|��,#*5�W3��ʢQc��#������d�35��QS�5��n�[1Y��e_�}�}׋Jo;9j��qA�	�e��g���_�Qt7�ߞ���������F�a�Z�p1��9����$��d�J1�m�Q6Y��/���YS4�n>T��R�pI7�1:0����/�A��Gպ��'�X�u�T�2����4�2N���>���@�RGx��y{8|�}�APLa�� \b���>�Ahg"�_�e��h0�>q;n�W��M�W �Z��b}��3,�C��kLaR6�VD&R�u�Gu�(��@\*ȘBmQ�O�w����>���`�5���oz�T���������0�<|�|������
"1Up:H��0� ,�%L�/,:sv`��	��>���}���#��?}Yn����o��r���']	�b��3W���e�YvI�Q�5�u�Gb1�0͹�����5% ��'*c1�Tjw��ܒڿ��fT_���� �90}��z%j^�8����{��I�Bf� &!w��%�%�cHH��������zf��!��o�C��3'��s]���+�F��>���e���I��+zT3�b�#E���w�֕"��]{\,����M�%I5�3����]R?7s�fYr݂���F�b��~���� �R���L��F�pG�L��_`	(�	��;�)��p�Q��K�m7�F��/��)�>�ͫT6��:���y���G�����������cu9���`]l�SX��*v߃��)}H$��m>����ޭ`EJ������o��� 뺳y�Ц��!Ԕ�L�-��4�����>ӎ]И���qR�r�$��Yo^C��O���z�o�����F=ᛩ3��uJj+T8�W���*!?u�j���c9�m8��J��($QeQk5_\�ҨnqV)�}'j�n���V��IYs�����k��%��}H�Nؼ�
��
��QGA�{b�ӂ�e��&-C�v����8�ȡ��ͬ_{���#+�4i�}R_�6ׅQ�_3�΃�����I�L��%i�������V=#H��Y&���W�\"�߮/��$��w.��h>T���h@���72U�%�k��g������3x�Q3�h�!��"~8W㒃��7_#|1q��{�Z��c! ��TI�9wR�7�!]�DB��+�d7C�_xK �0j����W���tt�L6���ekN�s�M���,��x�Nr�w�bM𿄥�Q�X-�M����) u�i8.Y�n�u�?�4#�,��D��B���D����B��&$���X�D��k5o�����'x&7
�b.�Y��ӈ5R�ǮY/L�ބ�(��\����~�����.Fq�VS�ď��ua{�:��<גּ5A����G�n"�Fp��j�X<Ɲ��h�s=�D?�MV���J1;���>���9�Eu��$�Q �{]<df�ꞟ����*U%�����@�$�����k��i��V�%c�����u[〃�v���b���Z��q&�>�r�z~������,��W[���m��O7���zc~?���Q!��c@_�J�;n��w԰�a2(�ɝ��oƋ�Q����M�a��t��ٶ`v?���:}���t�� ��5>�E�lt�vܺ�i�|��"l�m�a���\��->�AJ�̋'��?	}��e}�޼�������n�9!�+���ޒ믶�b���m��,�Պ@��H�_���̢<�0��%�0O��U.��x�KC��D!�P4G?�6�B|v�=/L�\��+?�$:���{ͨ����>��i�ҭ�h�����ϊNG*.�Oxr�\��7�k!y�.}��橥F"�R���2�J��c[`�тN��p
�ȤSu"�N�&��>��i6@(���w��n?R~��h��G�l�_ϐ����j��f'�>0e��M��=#���W��~q4�i��.YW&M�#;خ��VnbqR����+���4�r�ɟ<rgϐ��Я��S��Sd|S�=l��x;̳�a��;�7�^�ᝮ��J����m�����ܵ!f֕��@����9��80C����o)�ց�M<��>%gI<�ތᓈ����i�HC��M�5��,��2����$q���3u�)Mm����q"S�3�<���?,�r�[��]���LF���[s)1*W̌�j��U)*N�}���7�_�ϙԘ�Gw��W_�(���1��A�V3����9������\���������� �%�(��]L���h��39�T�')���g3�t�i��(ߔ��Q�bY�\���J�w�d]k�	}!�U(kQW3�<M� m�	3�Ov�D�$����sM�ɲ��X��W�Pb���I5�*/PMg���Q,�M�9�J�xK=q[$.^�5�u�gt�����3A+�*y(F���|��JWT��܇�'�{��ހ�]�k��:� ��й�>+���C?X�S�>�)�[���6��כ|6�]���:)�D��@���͆�&X�d` �����8y3kBL�������|O��;�~�?�$�0�D�Fp�h�a����,�P׼b���n���Q�@��Y�쫽��� �OF�OfL�@����
����j�)�������x�(%��5�LW�2��{��tzz^���"X�b�d
!yrX��v��X@L>s!�V�'�zw2�M��K@���3=�@��d�J�tN��e���:d�o(dA����sm*� ��v���\5c���,~E��v�NO��*➒�2~bk��q���0d�-p:([@��Kx�_�I�o��^l�0�������u+ �y�g�����Y�� ��)��Bȳ�)�Σ��?�A��ڿ����'COU�����y$�hkG��_N�5�79矩ܝ堋����p�2�`��Y#���KS1�{��!'88�D*�,p�$�@�ppCdc9�]��YBo?����
��j�^$ҽ��l��XBs�Ғ��Yu1DL����
Bڠ�CZf���N#�0��z�q�ڟQ�c̶Z���wly���|�jv]�������]/���m��Ii��6�1t�[��:�o��b��^B���~�8���X�|��X�ס��a����o�SJ�]*��G�� �!�_d��T(i^pi�Ϫ���
���S̎�7B�be�aN�Lx�fB�TwY�y�y�{i�r�X������,w롃r�%�D�2����3ѫx��|�ddR�W�D�z$p'����4K����iN��#�bFDW��]��'w�/��t(�wX��^cB%J��g%��]�L̯wc���ǟ�b���ݦxt�d"3s��{hL&1�Y�H��4�{�m1b
�����#sKH;!�/.��5E���P`�`}��J�� /,%��'-�"�.�A��+��L��QE�H7bn��[UdM��"�^al�'����y>�ޗ���-�E�B���-��%�*���R-����W���/�6N���I����
X�	@Y�+
��W~�Ӈue�$�%LQ6��9/:���s�m�K_�!�3�ː����CFp$Ɔ��Ay5��)]�C�����
c��4i�GOCW�;>?YD�{>\�D;���(�>���O�� �ų:@�V��Nz�!o�C6��t��^s���]]�蟴�P���6�*�AIA}/��P�a��L�6[  �X�6I5'�y���2)��9C�GӂA�-@'���� L�:p�W����F�u�|Vm��,�0M�d=BG���俨�"���M�w#�0B܋�F�%T���b�E��wJ���ރ�6�lPm�l��%Ek:
��������c6X�/��jۓzy|���2W����n�R����
�+B;�*�}i�ks��Q�y!� �b��ǩ{i���G��n���h�+A1�ѸO��M`�����JN�K��6#���eqE�h�<s.�N��`!��y2I�m�aF7�����4G�ӊ�B^7����t5%3t���9����<@Ѧ�
��`�,���ѥ9㌘�ؐ�Ju����`�g��TxV���o���_���#����[Q�_$r�,won��o�X䄺���=G���0�50T��/��>����x�}��2Z1ba��F�������ʍ���d}��\#���0�V���ˣ�	w��!����T������/�/��
��w�S��¨
��La�:�j�n�DM5�}�m�9��̙��`i]��L��a�Q;���E?��&��Ӎ_a�s��%ݜ{�sѤ��'/s3l\�X�t�M�Ц^n��	ɷA �����y���TV�/+����������(mZVV�1���9��We� ::ܜF3�����􏅁+��ţ=)Y#�ƬK��J���+ʎ�x�@h؀��:R)����W �F�y�8'���k�����2$ҤB��	�Vװb�~ �آ��F+�)uN�A�U4�8P���\e��x3I�^:�D~���lb��wG5s��L�JK�1�j�B	�c�=VT8�P��/���v�q����՘��Ha��_�AI��Q��A�]f~[�qJ�%ªծ�Kh%X;_�X��;�<�H~�v��cP�,񉘦�LԬ�#�ؐ x:&��S�2��*�͡d@�0��K�E�ݴ\�uA�n��q����oAۭ��|���pwB8*���+q+N�۷c��!R�&9��]��V�KR��e�j�{������M�yuk����7�Mt�.Fe�fi
W�m9��䵌��yr�:~�xӼhYό�|�\�C�w��I�9�I����`\�e������t\���I5Y�t8�)�ߵnhd�D}O�J��=�T:��wF�����ڞv_F0y�	%�%87q��i$��d���CR|�vB]+��A��:	�[ĥ��^4�>��O.������G�%�S�B�Ǭ꣬���$�rH���E����9���p2�^�;:;.�#��g��%��Y4�ϰ����adF^!Qfw�y��χ����~�	9��"�|\������^�����y�����5t6TI^�^)�U/#����G�M"��4��N��i����\�_�.���x������P:O�Y�e�z�%�8o*��H��|��6p&CX?��/�k�M��.f��S�@�� �+�=̋(�Z�FO������W�ŭ)پ��Ζ�l�36��a�:jyڄ��:�V:Y�@�g��l��|RЅM�ց$W*���P"�-��{�Uy z��k�k�X|��*i0�"W���B�*��6%��4:9�'�C5ʘ�WۓG��K!�eZxBvH ߢHڷ�x�-Y�b�(�];����Pc?Sj��B��}���{��-B\&]��"�ۄX��ӄ�r;,�j�=@<��z"��!���PL=��vw�(�b�0ys�Y2��u��U�yJ�ٺ����ށ�]�{�s���09��f��+LsH+�ݹ��iޘ��t��R�_s��W�r1�}A!�\��|�Űx�,�.�m�=��Z�Ǿ"�=��y�WO��y��nUb�&�_>�x(k.mxa=�"_�z,�7�|�_Z��JˀٜJ`ŗ���;|w��Q1��x��_�pe�Z'#%���({n�Ʈ)� N5���GJ��rQs�:����U�7�B���e�<�ZC����2�EZ�ۨ{��P�μ��v!�������ׁTЈ!�k`͠O�o�$��^H�x����'�@�r��E=v[�|��:�r2Xi+y�1���ľЙ`��V��5�h̳�dRm�V��L�!���@��8��+l�?�>dfBh�U7�
��8� �w$�;B��=s�2�w,��f�����ю�B�5T�m�P�x멡S/�i'a���ߢ>+n��C�h����<��Qى���i� ���A*�GC���"#����i[Z��`�_�N���<������wh#�aV�5���AVc�E����s��i�c=�<��ԍ��6 ����廽D�3��7lc�:��c?�k�����@��-i�Y�hN�:�I��0��\�W���m�}�_�?0vţ����jK�;ek��v�acyc/�,�l���mҬ��t���`H�;68�@�D�?;c��C��I�Z�RE8���4��%��A��Y1_�Q�6D�1�4�K$���ݺ�(�Yק�;�ӏkB�Fk�<�'�A��XYI�u��ᮉ���rDc���TK���"w�����*1@c�]�����V���{S֤D�g�����JC3*3Х�v3N=��3b���h�*R�,8��3��F��R�\�W��G�gV���o��7�g*&C����(���o�LI�J��*��4`�X)1v@{R�D�~�	�i�{02�P8Աϝ�7.�i��;���߰P�r�����H������h#�۬ga�AA���g��
ެ�`5�n��c�J��h��B��&Ӱ7'դqb����P��sr#9�����p2WI�v�3��r;�͗�rj�3��Ii��\Lwt����6�ZO�	��'v� _���0���8p���(`U���jԶJVᖤ����W^���v���(���	.j�#W! s�������vh�7z 5in"{G2y'���\p���*�`:�d�}�x�*�w�d�}�/-}>�6Q�
@$�b��@.��ձ���K�1|j��Z�o��/�x�G��� s��`tuq#A��M!�N��Jx����,/�KԺUl��/0>�!�&�e��/=ޣש����a[��%2$˔�FUyeF���^K����i>�eu
����ag���Z�ZJ�W+Hi��k�RѶ붂g�@�HAm<S ������jP��YL���n-Ā��K��ll�G�'�vIa	��/����8�O<@s��5�2��/^����S�X�E��@�$���]�:�)��2�r$0��� �V�]S$_n��0v�eb.���
1��@���v �#/6�csb}�9�F+��1�M���0ϝ�����W˦ʱ��� >sMM�$�M�K��Y�kF:�"Î!��;�*0���Ɠ���}���:��e���0�!�iO�#��b>����E�f�-Ӱq^�n�[��PT}]�;"��e��zT��x�2�r3{��1[�6���
1\��9"��aX��c� U�x��-���z��W#�>�V=}��Ȇ=/�_���:� �f(���um.��.���>ǖ�ٮ��e��y���ձ�F^�珁�n���췣�R��+Ɔ�/"/ʱl��������9]�BBvyo1�H2�_gu���4JȖ͵�����k;ʬ+�/��9`c�g-��#{0��j���l���080,����1���b��dL�4�*�X��e��݄$J��v�X�dN)3d�4�(���#R�/���X�����4�"H�g����9��.��7�j͏�
�d���$��x�/{�[#d7�Y��(XL�(���0�����G��x�U��9�n%�����v��O&t 蒔8���0^��˨�� w�w�����B��+��عt�;��ǒ�r�����YV�㉍��-O4��®�x,}�Cl��t+��Gҏ�̑P%'��y�z<�ƾ�R���V��oAG�e-ӳ\���|�Ƽ03�L�ӗ�%�)?�.ID��A��bU�-(�
��WT�xoTyf��'�GvC�A1��jo�~h�y��blۋ��,��=;./z5�������FAN���(Q�B��2_��6pr��40( ��"�B�G|���Z(�+�˕�F���؝��w;�XI��[��31�j䤉��i�߹,L6ܥM�Wn:D�Em���<a�@���9�T
e��׷'&���I���0 2�+��-a!�������it�C잁�^j/K�ѕ}=�p���I3�� b�
ݲF�c��Ӕ�2�R,���Z�k�+�=h�Q`���\4�=ߺ���#�0�ܻPp*>7�j��ˣ��Z����(�έ�X	oV���G������4Z��DrZp*�u�k1?l���%������	.H���n�T �9�򡛧�f�7rBj6�re_d�}<�P��>�i��wn����Q��ݡ�jBÐ@=�f	ۜq��n����d�A�v�̓�`����v�΀N�ou�,��B-"_%<��:�+�H5�\�	��x/�gj��8�z�Hf��Gt�c�~��d��c���Z� �Д�2��=_���p���S�A�72ܫ��ieM�oZ,�7����F#*���?�|�x����d�Hw��B�����/?��@��Wd$Cs!��>�cZ����B>�����}�V�v�R��33������[�+���-e0�D�i��ͫ��$�yK��_T8�O)�mߏQ\g*��p�K��n1L.�w�k�6�_��)�W�e�˒���o�t���j���Q>�ƙ���µό/������%�����fyee*XS���ȉ̭�G�m�h0�M�Ĵ�Lp�%;+�u�mC;�ózG,=��B�Uk'�(D��W�x	/@첾ь�n����;.��f����5��/��k�0t1�Z.nUߑ�p'�$ׂӺ�l��;��.4���>b<����Et��Q�'�L��������m��t.�y���LZP-i����Fz��'�5��x-#����QV	�4��pE���	����w҇����zy�+}< �U{��*e�B�G{ęG����(��!.������R�1jO,9��u�b��$����Nѡc�N 9��;l�_5Y~�Z��h�������8���8q�L`��fگW�̽��85���Ʃ�1 �3�T�
�5��F

�G��V�Έ~k�֟���j�aΊ24O�7&c���_���P���zQ��A�o��Ԟ�¼RK�o�&{�iB`4e�	y�13b�B_2̜�w��Dzv�}K�{�w ��D��Y�Kؗ��M����L�������B����.��U�ă��͠	Byc�FhU��Õ�X��-��\�[�3ᠢPD\�k+91��s�_J�%�{�a��h$�	�S>QoT�:�nFn��@��y�-'���D�Hb�����ֆPR�~Q���d�C<�xz���ڏ&�tx����ŏ	�O�ӱ��N��jw����ts��R��>K�(W��C���E5�d~��+��_A�^����ϛ�|��d��L�������Ĭ��%�..9��m����/�����m$��pR�IW�u���v:�:��Z��y&�Һ�͛^BZ�p�˕w*�����W������)�N��X�/c���7g����r�� }�{������ʭ��h��?��k�R��s�Zs�a7�G�k�����!����Ϻ��� �:��!N?1U;�i^�&j,&�;U�zw��F�)u���fm�� �i[�+����y�ߠ��lD}|��ُHΐ���-��Q��pn�ۘ0V�=i;��RXXP��hUF�W��š�[Զ�<���"���g��eRQqcb50�9�,�M�a*d�:�1�l��1�s�b(B獚���&�AB��@��Q�=*�!�^��А;�H.�h�sy���|�1�K�@�ai\
�j����ԨF,+�r�����}�X
>[���v�%��v�����!���j˥q��������}L,/�#z^�����n1["����!b�r�"�a���3O���/_�뾣g9���:UF祈חh`��pbS	��
q�[_d�n��X��ck�\�V�H�|�_D5z�Ȍ����ꅡ�&b��Z0 �{��@�?TwJ�)��fN�ߴ.
�Q47݄4Ίh꿉f���4T���l���J[�5~X͏�x3�� 
��zcNI���\v���Ĺ��Ԗ�L����e��^�Ө�$oY�\2���a�j��o�W3Ҧ�{[�I����b���O
V�ic�8g��Z�T�Cpݍ�0��8�78�.������B�g�V��]������g����^֏7fp$�^OӒ���/�qC,d֢���)�"�򔠷�CG.~%��-J�o5�����`��X����&�=-�Q�=��!�sT��{�wJ4�*�AܐPwE�W]6�m�5����GO�l�5��v��Dυ���-��g�l���^(k�#�W�fQ���4��bv1'Aa�3��}M��Ҷ�Ё\�m���� ��A�ür�ВD��F���e�1#�˱�);tʞr�-����v`k[ʱ��`=���^��Naco���ޯ;���hNe�$�k3Y�G��c\�̿�2P���+�T�1la�{����&��L_+�d>�������l�Xy�'��p]�p�Kl*�|1_S�7`̂�ԟ��>�gC�Ƚ|�[�y��!��A�U�z�X��&�_`Qln�v�vV���j��.m�	�e���8����rӐuQ���� N��_����Ł���"����H�X�G;�O��%n��U�����I�!�cxď��� =
ǫ�5�$�l>Y���{y$���ب�+�Wr��aK`u�q0���Hm��|�ξvA�Y�k5������-ѯ�8��wU�$�$46��)��
������_�fE�I���/�F�&��,̬;Kd�����;��}���Q'����3�,�T)�K����mV�o���ɼ���G��E�ng�*x=�a�B��w8�` ;؊��;Y8�C��Tr{ Q@gg��h)���&����~��:�}� d�,�M���L�N�p����_c�U��c�Kxg�?� j��!Xߖ���fg��2�5q���;�f�\lZ��j�M�'��ĝ�ҡ�_=|�*E+��,�4~���:�ɸ�ӘF,eU�x뒘#�u@��t�P��Կ�^H	�޲r$v	�~��j~��^*3!�w޸��� H�HMBYS��Li%�,���=uNvT��d,���T�×�x�i��j�\ژ�{(���yD�)Dӧ���`��u�i���R��%�YZd�}���c���C���$�Ly��yo\�8�(�h)EJ�<D�y�9��~.�usS:6�f��q$�ɮ���`5џ����_-�=�p�V��J�/~:�怔'ma��FP )��|+S$�-����Z@�R�?j�<��2dȇԿ-`+G֘����lF}��u��z�Լ�� 2=���/��u�Y����D�ϴ��'�~���X�yߠct�F��I& ��ZցAT�7��dO�6�Ic�������kh�c��J�b�Ō�@!Οx�>�И!Pg���uj�G~BF#�X�~D	S�̹�.�dj��?�"a��:�ov׎<nT����zv�j��wp[�]��D�r�yŧ��D�5��-}?�/���˂���f�~6��7�=�O�Ƒa�RԾ��S�Ԥ!}6Ǣ�˷a��'n��5���	��TE�����T`/ʹ�n��P%�!K?A4��L���Q=l�m����[�Sq�$�aa�x���q������� �fk�;XG����釄� ��҃'N`.^�<ҏ+���}�J��&:��P��o��J�.��~��,���"u�>�L���t�fSs����Z�[��w�bp�J�y���❾}q��k+���ԉA>�`{��OW��?�>���L�]3c���`4�P��>�d�-W���}��H�3��|�x���'u~��%kѸ�oI���Hrn1��$t����v���i���	qՕ��V���7w�D�b�?g-Xy���W|@��B������#b�U�ٝ�z��#n�6�+�;J�UZÒ�ܯk�(=��Q.���������+��Æ�6���D�p�*A�t8�ϱ�G
f"O�	o��N�����4�=��q-P�P0�f���j{��?=�t�&�PEpԴ���}��ω��u���M��=�*�f�?G�N�ns�Ms���w��\���
V'8I����M�Ν� "�	�g`Y6+z��V2�eB]�t�%�^���ڙ�h�f�_�@����(�������9Xz���1�q����F�.�x��P_;�����JyO`��u��Y`p]��o���*�a��T6�N�t�?a�d<E��7U�%>�_�JTL'��یČQOY<���Ĳ㋀��T|��i-P�k��DA�9�"��+{T陆~�8�뿧j���R�-+˔7�� ��� �O�2���2�9���ѣBQ��<�.%��d���f��8>���e�8���K��dR����^��`k�+nߜ�Vg�㻠@Yn����xf�i�i�#lu��;������Th��[�P������E8����WJ-�D>VaZ�A}���g9��xxhZ�v[�$w)i�6��pg]ڐ�P�f^ D��K�G9�������G݊�^DH��L�j�DE�]�;��вRA+t͆t=cX�v��"����9��>�>4Eo�A�mZ z!���|�9���n�g>^�z�s��9X]���%�<�B�<0S3@�q\6�yݍ6��Z+?Ҫ*�Im�'��QNӝh꥚L�Gc�H�w_�3�h����������qԲVT'�ﯯ®3cÉ��p��g<et2�aw���܈�Pv`�f@��:C^̰�xʉ��]4i>s83�Č��	����.�������8���X�4��t��U1�)h&��/7sR��uz +n�C	F_�1g+���'�l��;�opJ���cr�iʌ�wQ�V%��HU\��TA4A_F�����s���B���Q�C�,th��%�9U��ؑ-�/Ѓ��FSڙ��������lfP�,��)�͓�~�g*J.d�
�[�����S;��kO���"��Ҧ�}1E/��:��o0#[�S!{;���$m���UA,�K�Dlt�~�6�����V�;)���S?M��z�I#A��$��R.N=����8�o�hDJ{�_w�-y�{ɬ�
��F��J@()��Ya[%��"{�FȠ?�/��_8XN��u�+��m"{7��[	J?��=�t�wjf����������L�a}��dO��S=�6��-�8��r��vi }��x�=��iٮ �N�� 
"q��H�����D���"���ö�=-����P�o�>+P�/2eq~wq�CMT�>��O���\��u��Q��
�X�
ٷj�&�YH���������jT8�k=㷆�.��O��)l�7p@z���rȠB�'L�����m��PıƮ�y��PΤS�
���&�����F���+-��e|��Ldo/��7y�)7� �=�[��.�P�!�=��Xŷ�ؼJ����0fC��>��A�`H���P�^��$�I�5_�U�߆?�Ax�)�y.�}+Qy0Y(��A\���v{G擑� CRE^j�7�E���6Ӵ�:	����P�л\C����)|+b�6�=?r�j_��C%\�:�+���|}!�ex����m�^��5���u:��b��o��+G�i �{d�38MFv������$n4���}�j턽
��W�^��j�^Js��GE��\���`�W��[���<o������7(�jS��r���}�Ƽ���E�a��X�d1���[�KiS"�(4���;I4MظW�_,�-�SI����?�3��k�(���e�0%/u$���3N�KP�8p��?�{��S�A� �Z��H�I�/�z���hob�I&�9��Ɨ4�x�̶٣Dq,׾�;�9\~��y�pQb5�y�-bOO�Q�9��ˉU|C�H�$�>���0�wU�*&�Yk_<������u�8IQw�������Q"JR������̆�{�dbN�}4�t�\��Z8��ژ��������B,�ew���h�89$d7@��637~�th1j��ZdQ.�|����Mo@�Aw`	����u^��Z%��*16�K����[h��J4	���CV�J�Dw��`G����O�a�Mge�M�o�Km���6'J��m��V��}a��a���|�LZJ�Ē����!I^'��
%p�T��>E-��l���5�W�������)d9�ARf��&Ƈ(��p �vk�Zg�Tu�N���0���yB�1��V�|E�"a$Ғ~yj�3��q�������=B�̖;��f]~j�X=❁��q����t�D='B����?sF�K�v�0�1I'���-�v��Gϓ�ǃ���'ٮ,[&O�M]�_2ɗ�Oc�aRL5��ݡ���.��T#������{j-�qi�6�\��gb�C��uW�؋"��z�/����>���fn�6��8�r AK�4�x +?Լ�|&�Ț
2�����.���7�r	M�b�0�]~�Rf���]�0a4CHw����2����'������g+��yݥ'��K�v��j�1�������<\��T� ������`���҅�ń]Ǜ�R�앻�"��0���OSdn�8��F�=�:s�,V�8�N2�_S�yK�3,�v��������� ��Ė�$#;fi`�kt'�sM�n6%�&��"�̽W xH��c �W �f���-[�Х�Y�J<�q���D�u��ݚl�4��[]��b DWrK��}��l���=���Έ���N@6���C\�άԮ��ȐF��6�� �O����`�d�p(E�uԖ�Yw�& �����β���AQ@&�K��Fa���*y!N6"T�l��#��[���x�t����q�,���T�sa���i��F��V�(1�P��ǽ�9Z��yH�頭O�Ѹ�O�&f��`�"5 ;o��uOoa�'.ߧ�U&R��M5�,��g��ҕq<j�a�	�ģt���#��Ln���'�M/JԿ�_�g���`Cu����K����:�=��߀�+��Y��͞�x�9�C~�Q�S�=/@	�1���G��CTT'��
�6H�'عY�*z�{6c�8
���4�R��TW�C�(Ǥ-�*��L-XPtj��Ʀ줎�.Χ�p�LYS���f�Iz�W!�l�jU�x�E1�C�����:Db�:�)���Z�̌-W@�>l������EY���,�f��D����Eig�����V�����ϥNm��	�l%iua�
�U�.n<�����[�� ��@+\���!j)0]K�fpQv"���|'L����������YYb�W;�Y�L%��E#c&��h]�
�}}\(��p`�p&N�ӯ���M����ee^���Q��D�u]~�'���eIe�=ph�?��*� ���������)~�T���+{�3�0�j9G?���v�~�޸4[��ϓ�� č��5R�d�rY�"#��GN���1�f�b�Â�hT ���A���	������X=�y�J>[�Þ�Z�e�V�,?@����*��g�މ�"��P�d���2�02���~���Xy�Hf@�nz@ ��p15�B��\�&�%��D��)X�`�7iD�!�e���<@ZL�oaZ�"?���|P+���h`t�.�}�OQ��]��\���p�N�h��ׯE�e�'qE�gԂr�H��U<M!!r��� �#��"P-[b�1|�*��!��ce��FS�'�vҨ��r�5ڴd�����mN˗�w4͐�j�+
+V���٧<Z�۠>t}��?�3I�����Ӏ�q�s�Р�m"���-zT���A�����f�v�^k���-�>�������b ���'�Sm����Ƣy}s� �hsF�Oʍ��7#��b4`ގ��H�-g�(aG�����)튈�jn��s���F������_V3��e�f��|�nb�}�_�2c �
��Ƚs�,�mn��_����c���I.w���q�b+n�{�2�
���.pW)�x��`�
�"ài�d4NT�5�o*&�\�<��$�����S��gG���xfP�x1AO.A4MG�P��3����|Ć_ٶ�4\���7r̕ο���e����H����kv����ŝT��:���K- ��� �]��Ml1��.E+&�MV��
e��xH%�{�<�þ��c�
���n�Փ/��r`�eDU}�as�=eϤ�&�099��&�!���ۛ�%1H:�D �=��Ϧ4��S2
߾��0�jr�ija��r�h�Ov�ӂjQ�X�K;��-iL�*�:1>FX����2o�<-��l���׍1r�z��)��ӫ�"P��[{h��T����X5�*T��C��lsg^�`#Y��6��DUN���zr�����Iw4 W%�xдG���#��]N���M�k�h,#���1�Ь�&|�<��{��{^CA����èv�%����<����W7�l�8��T�sK��BS��
�Jn��wβ��Dܠ�ڴ�����X m�a��<a/3�0_�c��-��9_��N^����Ji�9�ky��.չRJ�Va7{v�E4��ިf��:�z��]�%��ځP|rI�gG]�{Y���EE�A+�)R�����T�'X�	֣E��5B}n|;$8����L��w(������U.�4)�?�5�jד^v�
����|��΂ٳ��k&���7n����ܙ����:�h�(,N�L���7LI��,�zU���lC޸?��՛����G�ى�|��XP?2:������S.�0׽�>9m>T�&�ʦ³J}� 1�����嫏DʣPy�r0�>jKr�^�:���xO�ӄW���@�#�y�m���g�o+��e�	{�_�"sȮ�6��u�WW��6�}� �o�.u[/��F�2/�s-:_w��y����&�a�0���O�}.|P^h	�D</-�0�0`5\�jl�˦�
�m��L]��Gu�;m��X�;r�t�2%����"rM�7���F��A�#)��dX�3����Ɋ#����"�\�� �lq&��a��|�:�Z��w��h�$�hDy��J.��~��K�η^|��O�Wx�8�����.��y�?�´5n���U�j�j^�#�;^��2=�}}=MS��e:8������g\f���mf�U����ǯ�aJ�6���' ��#-�{Rz
� ��9�bt��[�����=�u�F?:�1(E��6tY�ǚ�O��	�8�m���I��e" �. ��+�Iq���3a}l�?��`�V%����d["��l�.�UvB$�'"�h}ۥ7�g�^czI32�]�����G���p�v��H�����������M�����t�N�� R���u���T,I�]����jB�n<��#�n��zD���t�!�=˗n~d����|�>�{J��:9ݦj�3Ht��u��㰒Щr|�@="�i}q���/��� 6���=~�w�����9N�w�.��r�z���#�lc���ON��4���d��~�me�=�zTo�#f�ꈪ�sq��;�>u yV�D��]��-V�k�}�p�h�H��m�Zi��Z�].�s���GR�6������,/
����
ҵ4��������y7��#]ta��Vk(�+P<���An�sx=y� ��~�Z��j��s�.�E0���ߣD�^�3Ϯ'h�5���9�>�u;[i�'��XH�Ŷ�3�w"��!K(W~��m���X�IA��(�΃K���$��S�g�:���[ ;�O���+d^�Y =^lw5�ǑQ���� ,1���	��uG�|�ɉ��)�Dy�;�a�î"ۡ^��p����t�q�Rڭ���qc����ҍ6	���ټ���Q������w5"�ÑC���&����|�k[�Syy3&�V�r��qB�[�U�Q��63=��4�&y��2d��	��ba�7�	�a	J�ԟ}�F7+��i|Ȝ�'�4�&�u�[�$_��yw��>�⤡��H	^Ę��|���3�&����4�e�iC� �fh��u�h��G	�'��A]�~���]�1�<�?�Q�M�B����ѠnE}��D��K���e&�㕶]n;3�i�T
��Nw��𖹍�����B)gn��yxQ���+֋�6�"x�rq��﩮:=�鶬��.cl��#/=��
�ׄ$Z�CE��Hp�(�2���{�9���l��s9sD�H6X�:�C4��AXeV1���<�;C�^V��ç���P��*+��2���9@0[�&��o55R��t��B�Q�2dfC����yT�����K�^S�ʧ���/y�2�?$� ��Wݰ�Ż��[Cn� ���e����𶻞�Tc�Gu&��d�*�!Rٞq�%m�o&��ɒ=�L6��������$��3A�[�����g����qX�*xM�e���̑��B�,p�m�x��4�3A1(�tv�;�7�V��H�bB,���jA�z�x1�EJ�<��,5*���&�5֓����lu�E�OT&g���M�e�;�eCȵ����F�&-dx�2�����&�Vty$ ��q>�� ܁'��O,��J�PW�d̠�+!�9����,�#k���*A_�*�J�b)RԨ[](�hv�u��s�?>�shW�`Z����䴭w��T���Y!��;I�x� F~��9^�Bas3-ev����̖���|"S�_'��wN��3��KnW��0�FAsȊ���d�r�a�
:��ۀ��̀����6bi�5<}WB�{g�TcY
&|�o����k�\rU�38ry�����#�Wp�+$����5��A�Df>�O��s3jc��R�j,������bȂБ�]���`���d��?�V��ʚ��M3�P���bҲ��{Tl0�:[x�l:��-��%~���eԠ�>��ȓ��d3Of�P�,���|"%�A_oqG��*���X��T��cIr��hg�A��a�つ�`�eؠ�5Z�	�T�%�J�=J@U�S�^�ۉ�V�l� bW��It��+�P�j��$ hK8#𓮍�z�^�k�dk?�<����J�W�9�ɧ���
��">�雊�[�����gO1n==�uV mc�N����=�k}O�9j�ԶY#��C����!��懀d�d�ÿ}[�T�4�m�a��,��I�������#�_V�VvE�A��	�l�`-pr�����F� z��g=�\%;�r�E�@���X:6��9<���+9��v�����ڸ��c/�1��;K��X�WI�R^O�r��M�wF3!�v.'G�G�h>�v�)�k���)O�K�@܊/�f}p��o� �
7�h
�{���j��U��rR'���x�M~�y�h%��?���QZv.9͗�]�Zܗ�7��qn���[2����Se��e]^m�b���Ĺ�7�9��_V�`�lu��ުg�=Pg.N���=��L�ݤ��̽��M`�S���� ��SV�`e�ȩ,�̚��� l��͐�L�V�F����{�b�m7��fD�� *�[�#$��J�H����#�~T�*1-
�g�տ<'�t{�Ѯ�)�"�q�]����	-.���0|�㔤�1m�Q��L��BͷCt�wW�_?�w��3L��x3����*'ͦ҅�0��t�bM���
]�]8K?����w��
�Oȣ���mG��ǝ)lLm�"��4���iR�4�i�d����� A��ו+C����b\��D:E�ܻOa���_/�x��*X�*n��.j-�V�LO���;a,�"�B���%2�^���B]�^�yQm��Z���zH��h�<���Ӏo��F���� m{��x	氠�[Ձ[��,�Gыw#�!��s�G9�Z���A��k=�Z���'X�6���e�s�K0���v�����]�N�P#�����	����Ft�� D����CHbu�9u��P�`AT��w_���<����J�
���0D�����x��}��`�Vs�9v~5\	�t� ��EfWl���Ulv��j�U�3�1������k �`�D�qϜ�^�+Ѭ�蛾�m�9���Ӣ���\��V�r@hT0߮Ăӄ�2�G{Bd�b�zG��$����;h�_Lĳ4�u�����t���I��}�"=.�F�ʡ�w�UG��M\�@脐�H1i.�����5у����NE��͊�6�g��`�E-�ƅf�#�v �������Z����^�s�f��8O�q&I@�|���Nӥ��%��<����v��ӥ��8c�7�-Z^��)���MV���9���4U���a_s��l��w�����D����h�+�)S�֪�$	/��ƤZH"�Hg��Ot�O7�na���G���׍A�Y=�QC��~�a�p�Y¸-+�h�kH�c�U�P�xF.��6L	��.Wc���/�����Lh���[�D�ʍV9�$I/?y����o=��u�%�
7��$L�To�KN	�e�ClTA���y�� �d�cx'{+}�#U�fqf�hm�"%�t2+���[�\��d��:�0��m�lW���3=�{��}G���pC���JWi.�}��b�hkSg���\k��a,]�r-4�'s}��`��J{����t�r nN�qN\�,�Z랾v����dE�l��ۻ�y8U��wP3���72����}r�
���2X*!���¶̺&�Ͼ�#(j�颛�:�(�3�B�9�Z��� ������AN:�#dZ�M�d-ʛz�.�K8>R ��he������������ZA���˒���70b7Y��嶑�-�X���,�o�@��.��(婴M{�v�S�#ۃ-I]%	�5�� �ۇ��5
!��g���9�OXJ��p~�Q L]�ýղ�#���Ί�F�(�X	�
J�t�(�������jD���+�ϻu,k�	7e�J}���+��Y�������do�;��7���V2����V$�k_Uy��Sj(H��IYj4?|c7�.l)�"P��W)G ,%��F��/��*F= (��*�Y��3���< �mYwC��L�0�<؏C������������ŗx�>��m�x5K���P.9�bh�8�FՉYK�9Ň��mX9��~d�k*.�@��ʎ:J/<�߂��d�M������-�(k�@iF��b#!Xd��&�[�a�����^�m
�qr$3R��T �Dk����U��������l�(�� .�f�yE�s�l=�~�'BT��؈XH![]
?k7��`�T��n"q'�f3�D�rX��F�\QE���+|��>�,�(I�n��3px�<,���\[�2���@f�|&��Li5�-=#��w�ySQ[aE���V~����(!�EN��7�y{*��L/"b��v����Ɨ#��~�?k�ګZ[���i
��K)���:��t�l��VA3��ZEJX-Z�z�r�_�>�+��*�1;%������4����S~b_c���r�.8"%h�pq>D�ec	�b�g2�B�b6̱���n�I�H�wQ�1�F�0p�?�W���5�qM'���U<� �^nJ�5p;`1��׀@f�x�.������AM��7M�hf�A�W��%����C�����9��s���?��o{�9���.W�sLR��f0�͌RT��ߕ'Dt��Y(�$wM��E�}�<��;��jM<�~=� r��d�&�EnϏ%2IJG�L嚢.&�j9d)��;Y�6q?���,��-�< �rS��u/�sK��>�ID���
����e�Novw�>>���	Lb���1�������2h{��F�h�Y7�r��3e�}a�:�����&a�M>�-Uz�UɦDo��5�f�}_�LNa���8�ݘ��0�?\�j9}:p�M�_�s�X�F�zh(�֩��W�L��<cs_A��� ��l�����U\\�x�Q>��XM�(��|�*�lR�5�>�u�{gT�@H�b�_:�)7�O>�W��:[J�k$�^� NI����7���7�6�*��4����C�j��N�xC4ת�2("�������C�2��x#�B���/��}���߀�z:K(��S���gQ�AJ�5��������D��������$~���%#�%U�@RG���
��+W���4n
�`�Ձ��o(�sc?�����}�©��#b��*���@
0��yl�_n�_󑄘���${)؁a�6e���rZ=����e��w11�*ݩ���KL�\�0lb۝)e��i�.��`@?e`��(u
�BQ�s���]��~3�tNSGͪ�$�7� 1�{Z@�1�|�����g�H+��(^S��h{����ݐ��/�[������k�~�L?���g���t��{�A�!1�"�d������jҰb���b��� ���	Qn��A&����[�,��砟�&�eT�/MLJ nk��c"�}J��cB�����Q�_�E7��[f�_{�p�� �%-eers"m���A����7�c���?��,#�l��r����7U���qNm�_@ �%0*xّ^\�� ��
�U�G�W��=-�[3���{Oq���!�����zp0�@��T�u��ws�YY�F���j�����q���o���%���s�8|�IJ�KOU��@��0!�߂�U��s��׍Gl�%��PPڱ��!���ҏ�~c6� ���R!Aq �y�����&sM�2F�~Y��W�W}ɐs�ڊ� -kdk}��$*fV>�aNM�*,�'�r������z&�~~�0��}Q�}��%Iv�A{��)ȃ�r��I���M@58;6n�s�_�+���;ƾ�Ilv�Sf�"ZQ��=��1�(�<*7;�1K. T#� �sR`L���*�N������g�{����,�#K��ڌ7̥;mt�i[�B,5�غ�y�A���Z�mN����_d�}�P'�ɩ�2���δ`�#�� ���M��a�<1���:C�;���`b�@b�u��}ҭ+��J�v�*a�&�Ɇt����$�}���L��x�Θy�3�ѯ�����7.�ɪ�B"	�&zY���.�\V[.oξ��#K���p��mm3�u�[���sG�c���(���Z���̧O�ϳV0}��'g��	�:`���R+׭Iq0Ϲg d�����f��VRB����۪`7�4��O�i�)؅��˱����?�s��7�V�Uu�p?[׮g�����U�Ō��L�r�r$�m��2��T}�a��QUo���7'qM4�"~�G��+Wc��a�Jv��b7���P�������d���2l)_�̪�8|�󎀐`�'}����
�9/�P�Zx	��ϿB��w���&� ��Xz���вn�R�kt�r��Q<���W��Z�G��`S;�GD�u�p���*L%���_�W�&a�Za��-
E��!#�;�L�.P��std����y{8�?�%�w��� �Pk3���q�}����r(��3��2�?�v�a�)�g�d7�Y ����x��_�����]��)#�<��}�6�y<�O�K
���A�@�G�8c�L��S�R��H��[��.��HTu�U�7@�Th��P
t �2�VT(� �0"�?1���N��O���c���sά���Ы���1�������=���?�O��͔�c�dXNw{!W�/��V:�9�ͱ�խ'0�l��O���h��4�!kQ"��_6��=�2�(�%�>�0�:+z4~�]Ū�j��r^4��x���"�l(�##�ґ��k�Ƙ[G������ ��!I��
��I��/����P�u��0tv���:�7{ZM��4��y��_Ȓ4j`��4��eH6N�i�=Քn�����T� �̐�L��
	h,u���* 6hE2�Gt�S`�F���O�y���"��D@m�������t��QU@��(`�'�HC1��w����-o��2BL&U�>�����ovj�#�/"֩�=��HZ�����\s1a�5�0~�v��]��a�:Ƹ�\���}��Y��,�i��Nuwԓw%#3��+]8��(5~&qݺ�(��O��[���1���q�L�lZ�C7�$��y��]J(�g���YaU�ƿ����
�sO?T_[Dg*l삑�;K	lȀ%x�_��_��/�g��-4�*�|�0W�_���+�%Fn���1�p0���@�;y� wIb�tƒi�C���k�Q��j������^���:Bp�W�A 1W���q�xϿ�Hc
������\m�)��g�1.B���׾�ӝ�,	*5O=IT�U\����w��vo�587r�2+�Dt'��A6.���(��a��q8����#!�r��U��"��'ˮ�\�?���X+������� ���0��s�\�UZ��m���a��Lj�NH�������"�W�9+�)����q�����l�|�z���Md���!q�����Ԟ�B�V�V<;L֝�
�[����OSvC��:9�j#�j����fY�J�C�鹽��x�oP����r�{�i ^��V�4k�C$������_�1-�
�Te��ٓT`����_W��,�:'1Gh�_Z[msx V#4�f�	C�2>��]6n%rM��F�U�ƽ�Ǳ�&�*#a(�û���a}4�7ۏ��X�V�Wk���!��/������W����b�=n:��,��5��Z݅N��G%��,�V��F[Q���s�]��N���J����d����8g�L�!}��q�9�����Yo�k�M����,r��5����K��n�˱����[S�.�-~4G�8����(C�0���!�vɳ	�F��b���u��eӍ`��^d]����Xԣ'����x�G�=2�(��B��z��[i0mעŗ�s>���NU�3��_�Ǿ5�/P��;J�9��+��d�:��N��|�
���(�oZ�a��jI����[�~��az}n��˸�d`�;ǽ��Rbټ����5�"�s�ز"�"=}�HD\��(:G5��l_��:q����5t+��4�7]e�'���L����0�?+��$�߸G�"q*z���'�M �̗9�w0+#Q?9��5������Œ8�{{��jX��f��ie�_1I��~n�*^�t�ɒL��?�bxզ_�v�Q_����b-on G_ˊ}@�D�"�F�~��n�>�D�Ja_xt���~T��>��5Cb��&E�_Ӌ���G�t��h<NK%$� Ɓy�ت0�ە�&����:�X=��?4���S�����d�Y-^H�۶������_�>LʑT0�,�=Ň����P��<n�qV�ͱ��v����x��ó��+*�Pi�P����Y��?ABo�<;���C=4:�R�F����=��sH�'�9b���*jhP����&5
y|��uK�ɫ�N�4q��k��mFƽs1@��%Pd�O{a��|���U��E;��[^a�eg��fN1�a+�e����ܹ?Va)�P*_���N/�Be9� [Zu�O\,/_{�/����ͣ~p��e������^P��A�ϔ&�G(��hFL��F����9T`��Y[���p��j��*.կ�!WIރ�M�굹�h�#�h�U9��d ����D}�uB^/�X"�&T��쏻a��'��
#��xcЍ�"��#�0�!yug�
�g�9��rR��k������ ������Q���VFp,�{��@�d;�?��1�-V�Wla��
T��i(,w�cr�7��a�X$�*NHX5,O���R��|>Z0�-�l��<����؃M� �*Ms��g�����^?�	$��6�}�6S���ht���/cS�3�ٓ��̯>�
<O]`��+��:t��t0�E�/�S��ԥ�vL��,�HK/
��l��`��ԗ���r�ʤ�Q��ZFLC��%v��'���B�ZJ-揻��H�
a`��k.��3(�qEx��ch���%�ב��M~����GG'����WmN{��2�ǂ�g�����:}�(A��vd�΂Y�PQ�WS�_d'��?)�}w�n�)c�Y���.�Z���T���c�D�g��c�q������x�9�uw5��5{��zӄ�웆�|��8�D7��ѭv^T�{>o��dݼo3kM�������w,��_�c�_�"�3L�H-��e<+=�״�&Ӹ�uJvS�KE�x/=b���:Ż�!�?��8�^^�%��e��S4���-�
aX���������{H�+6#S\��Y�s���H��N�t1U�x��@r���#�I�i�-�5�} ��A�����*�d2���>�9,�Nݘ��0i��wx����V�5 K���ݟU{YiM����d���c���:>��HB��/���rO��}��˛�&#�3�,<P�IY�R�;߄)X�-ځ���	4|������$f�p��f�&�Mw3:L��U����F,bO�_�r�L�#�YM*GG\l�B�A�2l�,���+�'�X��(:�$��~�9�����+q�ZO[q���j�)C�k��A��\��je�7�B�\I9�|��c�)�Xw��3�\t����r;��^wL_�/ĵ;�!Rsc�e�^�2	2�Yy�Fjv��=o3V�t�BƘ-�Q	���M׫�W���}/k�#�B�#��[c�I�j*E����*
:����x�� �4ڗ%�[���;I��[#I�˻�mF������K���`ˋ�,��c�tkX�o��-d��4=����+��\c*��
o�0��w�Q�
�@�#��Jl��5KX�ڈ�Z�}ڮ�ł��S���*�}��1@lΛ8w@�H��0�%N����0��#Z�]����R��k�-�1��|YZ��5�5-9��c);�?W�����f�5(�^�sxg���\�5��=5�v��=��LS�_��"ӏ��]A2�1�>�X���ة�zm�+oepR��Jf�3Q�:���N�2���̍���¨��&h���^�c���ڨK↬'@�FCl&�FM�a]�p�����[\s@!�7�ّMI:��qB����&3!�JGd����2��[��+�p[�1�KE��Y�' ���p�Jp�8�P���K��$L5��d��7��|q<ʍ@�;Sܰ���f�H P��.��3��&�s�҄�%��G5Mu�?����� y���C��u�/i�����y�RK/�~�Wq�V�.�!�������{�z�?�]����z��n"#���Q<����w�oݾ�9�尵�6~�/�Y�9 �Nc|c�{������/^�sX�d��A�(/J�8�
�3����7��1O0bx��K<E���\cz� {9���X�c;q�mG�l��1�����S|g�Vn�{�o��NA���*;�K��Ԟ�Yl����HlBU[��{���
>]/���䜨��c�ȉ����z=a�9���5]�b7���� `m�3��Tw(�����Nc�X굝4��:���C�We�2=Zvo\F�?���Z�Jcm���T�A�r�N���A4(�ʾm�w�>4./���dV�б�%�����!�D��٘Ay�Ct��8Y/iY%��Ā8��8�\^��NC�וBdw��{���n�m
߱u��x�;�:&4ϗ�+j/.$���ǕM�����["��MV*� P~�D*|�Zp���1֨/��0�壮�푸���<�}�4�N_����M�br��#y�7|'�� ]���2�;���1�f�����l��Z`.�-"����ĺΩ�h�W��Qf�r7sD�`�D;7����r�T�#��)?�����R�sψ��=�&u���$T�ͽ���?����EQaI÷�S�����7y�s����Z���\�1BD`�{��ڎPd��+B�n�|v46�â�j�o����ߕ	�7m��
v�qt\�ٜ{&Ios&5��~w����.�G[��\ƏR�\�Lt��m��3�\�K>�d�#驙1�Vi��>�������YgT�9EE�/�I%`�@�n�j��
�+�z;P�rhr�{�>���:�.���v����9u����m�_���	�;6m��& Q�Tu�9�A@���
ph��D���X�R�4��C�diP_�uJ����@~G[��\׻ٙ78_�O��6��25Ƽǳ婻�	'����hw��vY�X�n&�2&�8Ev)����`A�ӧjs������v��*��0Y���<�&�\X�o�����%}�����	c���`[� �K����~C�?�����_�7T�-�{}��:Ӫ���_�*#`�V"d/�bbT�{M��dٕY�T�����0�$4����O<ԭ�:6[�#�
 مa��;�
��B�2|�5�p�

Ϩ7��ܙ�kz#�E���5(&�����<W�ȃ�-�:AD���AZ��$d��i�~
��J5�~�k�ʡ9������1�Mq�ɵ�&��aTI۷7������'��nH�=.�22�Ko<(g��o�4��y��֐=�f��#��e�$��Ai��l�d����(���+/$�W��đ�_�MQJ~e��Z���F�Bd�f�T5�oئ�g5! 9K%(��_W�� �H�w�h#��I��ݒ9c}��M�$-C�T7��4�:��R���>�l,��!�I��s�ܟ�x��v*�߰�=9k<�ԩ���PP�g[]<���;�23ln;���N
4~ڔ��s����"1OCL!MH^���5��G_y�U2~3�*3����U/I�.�?�J����O��Wj[�zë�B�os���ΊkcCrj5�T�����fx c��j�bi���(t���L�&1��/����u�T��Q�����2Yt���9�$��p�׋�rV"���"�Z}(ʱ����|���n7�@�đȲ�Jǜ�Z�g]�ݟ�� �«_�Sx�>�Zk|8�Qк������r_�D]�� � =c=6��6����L�& m�wG�_�;v5h��o^�G{�"F�Wd!�����O ����a�v�[���1�1L�`��b�;\t$&�������(~��e[g�j$"s�J�lA �"��F����-[���bE	��6
y�ۂ�I[�Aٵ�5.�3�0T�g�Ҿk�G�6��ꃃ�`��D���[��$��,Q��V*�� 6����8���!�;��u��))�)��Cڭ��zы�T�O��:h;�24/-M@�.���0tF�4Fԋ�'ɩ�X�/�7ݤ���y�����zQ%f3���#�=��}��*y栅��!�F$o�9�r"�dV#��_n.���J���?D�9��*�kt���?��4=	��w�%�|�C�;""s`y&���|9������1������a�gg�?�����Z�5T������;8��d�{����{@+S>P}�N�c�r�Z�+�x�~P��c92J��RK��ɯ��Q�����#�$�a-i�����W�t��ӿal����޽�a�A4����!�
0�b�<��/���>�l�j�H鼩a��Tl�����6�~�`��.b>g8R����v�S��qw��O�X�R�+��=|��7��ҢjR}�w�����,�jb�.8�����B��h3}B�+j������V7ZH�� ϫ���"���9�k�>���C�%F��J	�{q<�ߛOe� �}����8��x|'kQ�.?����fT�nʲ�����9�ǿ��|{k}N�������!CY�CU�t�\�T3 if��6��ŘW��r�Q+�b�@Ȋ����!�%�����9�l���RX9+@,�H,f�Ģ�15����31���:O�VӪ@(8ڐ�K�iQ��_܇��p2����	'�����9��jؿ>��?���몧^v�Ua�ǅDb�Oy+j�����o��p�i�
�2��O��T+	����ir�=�EZZ!,�hl��|�N�C�xHV�k3;Yt,�f���W����ۑ�g���!�C�`=��:}BXz��6�{*�'NZ�`
֑��I�zc�u��e�ܿ�V
�~<��>�Zl�ͮ!Ȗ��zٞ���?��9��+�.0�<H!����W�J;���l�gCm���u�d����S���ܿc�KZ����T�^�Z�@i%��S��(�٫��� " ��V令S��g�7ʭ�f3��p����rwr�2��sT&�,`��g
@��g�a�X�vB �Ў�g��Y��]�Z�Q��ƫ��]�7�!Q��Q��P�:2*��n�.�JwO�C���n�4*|�46@�v�@��\F�B�9��k�i��+D�
vZ�
���6�o��j%H.��ç:�st>�hz����l�T�PlIg)���XG��˄���ux��dt;���%v���avr��F�@��ֺ�>�F	��sn:@��_b�K&?>��
uB��)0�<tX�W�KSҥ�ÿ;2�����Nf�<=lv��9�'�t���\�'�mU����ν�L��-]p���PO����s]ֵ�34��#�g[9�g�ῷ���n)VM�XvsГe������|Ƈ87%�.e'I�d�� Hit��ㅒ�ܪK������p�$O9�,���|"��a���^<� ?-.\�p�5��ְ��=����Jk_���n}��E��_G�a� �2�8�]�pK�Yӫ/�;�P>T�v���M}��p^ܖ���Ɓ`c�YSJM\���������LgQ�i�!�¸/��;�(4������E` �g
��ȉ�SU"Su؋�s�D.��M_�>��� �P����i�	���ȓ�4�j�`~{����a��u��ذY�����=O��B �j�T��{:��ipY���okO6��rU�
�!H뻝f�r��a����#�=4º��z�N�U(e�[q/4B/r4�FQ|Kg��v觭�b�y�%��b+r�%3��|W���Z�M�/�P-��F��S�΍^�y0��-��jn��Dw���?m��Au��Fa��Ps�9rAR(Bͥ�ăj��z���Z 1 |X�q��v��j���r�Dq~�OO��G�m���)���*'��Ȱ���pKDB�suWx�β�Ɨ�+�T.$��K�PMBI��6���nO�䄭�3m�V�	�Rb}+LӅ#X��[Φ {��;]v�z^���j9J�z��j�<���R3�{�f�D� Q=��a�4}Jq����v^?}�
F�����;hwV7\sz6�뾋UTXӮ��? rp��9��jy�m��%��Gq�C�h��¸`���-���`�r;���rΜ�~��M}e���P����U$�q���;�"�9xxz��2�+p��7�������w�ч�֩���k$M�Dv�LV��ke�XS�r�9��M]����|����ՂN9�1�VJ� -~0�>��!f!"�&<Ѝ���&u�̩�@�#��h1< �P�a�	��h���/g�Q�!�-��z�����ՏoYQ﬇���VbLI5\�A�r�rh�A)��^3	�Sf��~W����ժ�aqq��vE��^ܤ�Yp�1��;���J�~���<�W�r\��6���[��G�����$�x�o�W���r��Ő:#��E~�5a��'cb�T��r�V�Х�L�
[�z��Nk����au�؛N�%|���nq��$��֏���*�"_������Ua�՝�
lA��
Ȉ�Җ�'?L�C��]yt��8Ϻ�t�o2�I�K������ud�%Y"f�Zx��� �X���<��I����9i��J�V�s{� wjY%�� �$�Y��Ϯ�[Ajm�,t#~�UV���͔����F�$`��"��|?9�c�Ng�o!�b����fa�tOU}���&�J����seM�fD�7v��_�U�}�E��,����(�}0)��3hsk��X��+s;�9d�L&�E���o�YI S����fj�31��8C���ʂC��R3t�g�`��6�B����;a���%� �G�RER�A�!|k���]�r��f�%v�ID�-����>�g{�) ��_ĺ�W"�8!r/G�3.�7I,~84��)\1@/�}n1!��Tw�8��f����`�	�'��m��_�J�7��HG:���!����=v� �1�*�#:TlҟH�����d��|�F^���	��h�c�Zt9:���X�2�_L��2��Yk�~��S�q��O�j藲�.c��b�\ƻ��5ݳ� �pZ:��
�;�����lz) �ZE5ők!�ڡ���o�84�0�7��2 W\z�붵@,OOS�SQ�=��Р�Ic��߀j�uv������ �/Y�k��H��k���߄{�>Q<�qP�� 2�9I��2�k`��#B����N�˴I�9�īcg��*�7%$�0xY�p0�F:�R���Nv�/<i�oG�\ �K�Rw�=���΋�=�L>=�޷���4�_��������	�2-��P(̖팺�
��s`2�__�՜S"�pUgV�4�*�r���'���4��ȃ�q+�K��;t��Yho��i�{x��qp�&�(h�؈��L��f�&��<�w�����ln*CzPM��Qw���%Gfڥ}�!�GV�A� "�\�O�<��;�v�셲a�*��ƒuv��q(���8L�芭��9�TB.�+Y9$���&�Ǡ3���+|-�X��k��i��Vn���OW���#�1���4�m����hL6�	���R����?����Sg�*��ϒ�����g���Hؾ���ѤA?,u_���VO�t8U��>�i����'��S�(�`H_��,=�4KX�^�u�������M���&$N��tDË����jǛs����Tv�e�H�wU�&�=�%��b71���*���#DŶ��ހg�����+�|J�WL88����~����=��&2�ӕk0��噖�@�5��=�ܓ�uwa��$D I��ͿF�[r��\�x������j��a�q�=V�Z��EV���_DAE���IV��=��2Y�Y�����<��J��ӿ4@�$Ǚ��~��^�DcC �Z�w�����2�~<�A��ƝO���}�+��;[�Y�)<h'�=��F"��&��eP[x{����'���,�����m���s��~lP��l
D�ά�o�u�����d�r]}�j�MP,�ޟj�<�j+@��b"Fv]4&Z�J��A7�$bm��CMz�qy��K�0O��T���+��pE��>�}Je�c�����!�sCƶf���5���Q�0ϯ����?�%,�>����t����	�����_l�ۼ*��	�M`���b�1t{��H1���S��A-� vߦX7�d6ȥ���6�[�\����Z�^�&V�i��v~(s�z�E�u����`=��c@��Fqz��ۉ<�C�b:qD1�����E�.i�~^#)�z�MI��G>D����?9���tU%�v�"�y�}�F�2G4zs	W����{��?h�q�ߡ�1��2͝�����^��
���>��H���0��KI��O�O%Js��?E�8�^1��&mP X�O���-�C���/+��ׅL����9$:�>s/,��>��=$aS*�!�V�`��;�'��Qm������� �b]�:���!:��*H\|�&���H��B:M)t��M^���C�J �f��!�B���|��s4U��9��A�4([����m�ZW>��>������7�S�Iн���$�@�NnIԐ*�g'����z�
��1��4�*L&���Z��Snw�(B��(N�^w:3=xJ7ۀ�oa��#�^�,*�aKݮB�2��`��2v�G�����}���P�BM!���sd��[
(W�*1����`�wh�OF4�����T���f��������bX���m!`�챓�wQ� ����c�	��������ՙ��?چ�n��ϫle�-"��|�f^���R2���E<�O��ъ�4,'-(#�J�d��j6�6����mvbT���?�{(�9���A�Vj\܋y�I�Q�~�Ը����-τ����`*[L�%�V�.Һ�tY����k����#��L/޿6�e�'H��ڇU�nq����>;�l�a�w��ZH��+����l~�����l����'��0��X��Bmn{A+�lc���Z+3�9���z˓a�*<��,��UˊH�u!��	��|̡�%Uͮҩ�B����z��N�:��Wb���"w��5�D8ė�p6(�k*I|��o#<�%?���VGG�+����|ɸnuB$GW�� �� ��d�g��|S���NT��n�.���/Ok}��:u�vjY��Ѭ����!����&�M��^Nl;s� h������ ��j�a��t:"�t(���k!2RV7��80<�_�ն��Q�������M�.=��"x�����F+�*��/y�ӽ��$��f��|���R�����Ar�/{/�U��ak����j;:S5nU�QY9���c]�܅�a���" ��_|�q��,���dW,D~�3Y�̓�e�{7³«R'��\����#�c e�G�R�!��^m�!\�S;��_S�j�&�@�����z�fa�ϼ*sG��*
�!���M̜u�R�r\�(A�L�#�C�\#�	7��q�^��;~��;,q��-M��R��������Q%(����:���r6gSY:���{�҇$?t��̼CY�We����U�����	���>�u�<Cp�||��t���
�(g�J�������x�����O9��8U9J�l�p��@q���e�F��lc/���U��է�$x*8'��q�5�=���](�ƣC�����=�,S��SM��bET�#@� �fxLx�Q-�.�����
���Kh��i�`�@�P��5)�l`X2K�q*z�_���G9
��j�F	���O�rE��p�w*o�ٚ3!pʯ_�`p��xN==�a)�A+����^�pב��3&��U;��\I�� h� [�-?ٝ����qS�;od�F����u�kS6q�� +���!�Dh�o;�
�j
��3�D���ĵg�f����YЄ_�n�Ό�tq(5Q � VF ,B?�Ĝp�>�B���)!����8�y�Ty�i���p��>�Q��c���\����g��Rӓb�#�wG��7y!I~����Jgv��������د����F�+f�������|� ���`ˉy���e{t�]�x�b���I ���N�+�����)�l�ò+c�}�K�q��[��Ckc����	,���~m�V�OQg���&�i��HUp�M�%q�k;?�����Z��%��Rȣ[Zn5u&�ʒEZ��,L�
F�g_��a����N�+e�ۦx���W{�Z얪�w�#��@Q�f<F��'��0�0�H��?��O?`�<�GM[cX�dP�NJ�����ZQa[��-t�q�߅�D�N/��*˷ꎬ�O���� Q�{��o�՛.ͯ0@�u�8�m/[�Zhc�����'}4�U���6�}����7�6͋"cDBhټQ�+>ZD�.Ɓ��ҧ� B��S"��B$�p����/��S#7��x���k��ۀs-�/�>���N����3I�+����d�Q�Z�ὄq��oNA����
UF��ـ/I��b���W��b��ݴ���ʽ�2�Aׁ���{�0ke���Q�j������*-I� ����/��kTX�i�|pY��>���X�Сn�&�3z�}��1�9���i�e�za�����@^�Yۜ<%XYhB�g����&T�"���U�u9�I!A��v�K_~�O�n���*'>$p"�\/mc�u'��֍���?z�@�c�`鮝�;318�� h���D����s�яC甇GB��s�q��{�7H[񬙼\MDcCa�'q�~��.�J�EfE���?I��;�6R�ߒ�*:AL�T�X�;ә�5 +��hY"�3�V�<���;�0�����dS=���w�!�7�<��m�k5�g�;��4�dޕ:�3�TH͝%.Ӏ���@4��M�7 �)�O����q��h��1` z|����j��3��>]��8ͭ��^�����~�h�m�G��t&�4���YQ�)W�ieU�1ҏk��mwH#2g�I�~xz�E��g��m�ɕ��^{�{9�4�ԣ}-vP5mְ�	����嚸3v9�a����L�TY�PB1%ˋ�xG��ac���z��R�nw�u�����3k���g=��dC[� � ̴~}N���I⛺��|\��E#e�/EnO\��"�_m��t�l���@�-\��	��G�r����ڵ���,��?�=�;;��M �^��A�<6�<�٭���m��G���Ù�Xfx�Quu���X0hm��1yP�[=�G�E>���j�U0DU~�S�f9�Ҝ�K|��^zO*��[���V��^���o��/����"5͏Wp:�ZT�c�λu~FB ������͝c�O�ZxM�bA6�cz"�s�`;s�oB�F� �GS �L+k�7���:Ӄ�sT6tJH�Uq��������K� �?P|B�9�rh�"$�I�N��yC�<�]z�o���o ������ۍ�?�6W�?#��iC5�ݿ񱵗��B��\1�X
#�n?�����L�]:Ů�p.�4�t�|]�T#����"gS����bs��S��<h����re��[��4P��銬�F� �ga�k�.NE���3��foL+a3���NJ�D��4�<G	�G1���AǨ��9*�y.�rդH~}��*8�ϏAŞO��7����6҇�K`�l��Ѭ}�����V't��&s�T�!��?��:I05�K�B�ɴ-NTj{��.-�?�L�����)���JR5�>�V����6�(d��|��=��YpH�ڢ�]�|Jc$p{�|_f&�� �(��{���;[ߵ��Rg���
,Y��V�z_,}��k��*��vLQ�Ƈ(\7 X~�S�<��'+L��l��lځ�߲��hǢ8���Y�D�$(���/��������oi]�:�;�E ����R�h(!J�y��d	������^�ON�����\'7n�Pi��-v4����	�4��`�O#,&����C��¥� �b_�lD��B� �AaM��i�w\�Z���Jh"�\=7��9��$wz�����=a��f���!����D�{�!ܿ_܈U�N��q�xm�åJ�b-��^�,î}��o�r�v+�]��2-�ځ�bI>l�F/"��U%��㍆�N�d�P�c�
��!��erlL��PHAx�������~�n��Ic��L�i���*�1�����<=����Jߔ��w5�zTY�2�)�V���W���$�ϟ�z�G��#��������v�(`mVW��|P�w��z��<�y�W��W�H�O8�Gۅ�R4Y��fa�T���)Pj��'��=���jǋ�V�=]�ir�:*m9��`��)�5���d�G~�͉p�5eAt���UZw!�$��v(m�W�,��*�]�E�rv�����x�xF��1�j�C���qY�$��<����?�� �qR��4�����xWtz3�<l�a�B��Qf9-:ǽ��18��fH�er�j
0Q��=�&-^Jx+;�2́����2�>���U5�D��ԋ���-
�j�TO�4;?�4�x�g��(gαe�q5��})��}��[��C�Wyp0����ZJ|��lS��nE�*p��h�}���ˋ�)Cb�����k�8�t�`M^7�_�]��$x�\�b��t����o5�K�?��kR�(�wčՠϻ$+�����z��l�a��_�$�\�G>��'$��
��ȏ �2�*պ�F<�{�q�X����{�9��8}u��ڥ�Pc�G��n蒐�(��h�>���?i�l�.�-�4��c�?5���$U�_K��Q�=O��Q�N�N5ckX跧5��s)��V'������Qyz�ltK��[��q�p&߀åXD?��F(���^��5�w�5,�LM��6_�+����rЍ�@�_����?�c!$�b�d:�z��h^�:D��,M�������z����1Mh�G��^l�4��R�J4���o��z��R�	P.V���p��F�V���Q�ED����u:!�oL@X��~іys;VBCʤ��z	�a��}�E�Q]j|��ѦK�Ҭv��ړ�7�F�қK4��7��ڗR�םG���%Ґ�e���1T�����	2swp�'"���'��dw�z���D"�Z��N�����������fƛ���U���_'a8��8ǋ�d��ڙt��&���(���2\��
��c:D>�FR'��f�W���#�U�Kݏ�тu3�11��޺�,����1�_��_h�����E���&��T��Z�6_��Ȇ���ɍ=; 9�-�7k9bKV����~J�<D�ޤ��M5E�1/���6�53���Pqӣ�`-ub���%�F��(�/��V��9<�
��c-cF���s��G ф���̈́����s��H��P�z:�;�T��v/5.��c�U�d��ɔ�c��{%��.N_�����1�&x��;���]�X��BѪ��W�ӝ@I���OR��iUw�W�ΧɈ�U���"��"�Ē#���S=R��wʞbK�'տ%�K�n�ș���}����r�bW4�Jym���]/����m�:��KF���|�qpb���rE��/�"�7p�<�Zn)n1+E�C�T�ԇ��}��3j�#�J^�8���F]+loOk+�]^v��|�����7ۈ��9��o,���'����oiM��8A���+��;iL���X[��z�!��ՙ�|�c�X�۶�]L�߾���<�~�BL��4��Iʘv��C���>?��~��*W�7Ona�M���-
��hŗ�t�`�%����Û�&�t��v8}~H�G>�����f�!�E��I�w���X�h��S�*�{~/��C����* S?�X8�a,�f�Md:nճG�~�G~��ŰF�(���ܬ����}�����@�g8���vOD�rH�s/�����r�O<�M���Ҩ�5]q�h��~�s��h���rp���R�B"ߘ����9YWO�,5�����]�ާ�����<?�C��.�M��$���o�R��@'�(D��;�lY���bs��Dސ%�����uڝ�A���G|H1j6#�]C�Ec`J&������PxP���p��"z�F�J!h��&��pFv^R�t��V@����`泚��S�+��d�V
��0f[윎���J��=	a��C"ơ���$g7ڗbʻ����i�zz:��>����nl�����HY�����v>�L��B�cU��#�k���\{U�2�1x��wzk�(]|�����q�����9������
�Ns�h1�����*��\����Õԗ��Ԣ����S�2IqS[��i�R��<��:o=��T�ԫ�ئ��~�	L�x�x2�v�׽:�E�cQ��|�i����7�G� c���8=f]��j��@)�A$# �� ���o�g��%o.�����B�<�������KF����Hぴ�]4�%=rKQBb�`�f�������W���"�gh�QQ���RP4�/(v�G��"@6��:�˯� dדNj� �΂#p��R��k�}��K`���:[q�q�'��YVqj��d$�e$����@�I��ʥ�t�myg�tB�u�}��{��wvZ}M��N��5��Mxf=��n HqY�V�̐�����z����g��o��֍�y�d���s�:�e>��N$o�kI`��6w�0���|�$��I/�mw!���P���o9���ȅ��C{�3��ZP*�[��S5:��kh��Eu޾AT`Iz�?c�����5W�&�հ�Ǜ���i�!;�1�Ԏ��4���� �֨'$�n�TA!�Ъ��9��ҙx�"���=�I<�=��3/>�{ �',܎AZ��q�^"�G��xzoy�	U,)���WE.��C�j!�qÌlݒw|�":(;�c�W~5D�ɴOH ��5�|LZ�5��*���\�sv�)FkӨ�vT��4�<�%����+�T�xl6Ud)�^�#��Hu��WA��j�$��	lۯ	ID%9����Q��֘����@ף�;�Z�_������2���8�fG�pTU���׽}�c=���hدP�u�i) EF����Ea˳�j!՟�Ye\�#%S�^o�ً��Kt�o4k�l>���"��ނ'�<\���s&�ܲ�Q9�T��V��>��g���9�5L �q��=�F	�E;�ىI��v��8�s�'��������۱Ѳ+��b���?�\�Ȝ/�K��Ȱ�HӥO�?ߏ�5~dx0�E?�<��0&�k�M`]�I��&K4�%��2�Vn��E��hu���h�ˁ ��63]��5��̶i�(�����<��ߧy�FZ�X!pM���fҼ���Q��l�}4�,���ўǰÊ7�" �j@����9�>UO��p��6�p�k���3+zƍg�i�U��Xu��Fb�
�m Z˰�;	Y�	�uӈ�ӓ��/�pԙ��u�ln�`ȩ`0���bu1�+9	@�a�&�g��6'�����I�_�'`6�-�Mq�f�����>���~��k =
�8pZ1��.���;%a��Ɇ�|=5F�rVsӂ��Qn;r܋�.a����J�i��X!�ކ�-�#YY��e�Cc0w�ξ�$�d�A`Ԥs?�×uF,�i�̫Ӷ�s�ɋ�XI�Џ=m�_$ő>O�Ҹ��J���_�zd\у�U��\�(��w�jP��B��1
|�d��q"��Y$8��1Wp�����8E��6����S�nH�EԦ� ��,����S���=�yR&�����.1��hֱN����# �D����Yx9P���1dq���eF�8��ۯ���hN fn��s�b4�9΃�(;4���|8�o6c��)c�j2�5*�W����Dࣕ���p]�r"�����ZO��mM(8��zY<�<�{2�~�Ұ%mB���������@��9Nc &������#o�HR��Z7�
&+�Y���EL���Q�Ṭ����+3�D�g�7���zS/,�9�����?� G�9VD�B�Fx�̢DM����B����!�ހ�h�E'%N��щ��-{K�"�8��u5r�Y��4�T��VM��^*��fhx��0!�	C�̍IДR�%*7��4�}e��)L��ә�)'as�'���	�7�)�ް�Ǘz^���4}}o�|�7=�A��?rMH¯�"��y;�~�[�9��3�6��F��$�N:��uZ�sYsJEd��I��n��5�w���N�8^�h�=<�$7y]	d��z��i"�_V5%K��ᳺ���)��
�^>�r|�G��b�,��M��v*�\�܊%4�S�s� EN��K'Z�'�Yr����C��&�r�f�
�U*�.9i��V��f����D�������'��P3I=�ud,��Z>��⣪߰��f��B�.�!�Ĉg�NZ�r�p�v�u< gro&-D�H��!�V�p�������LLW��(ks>#r�т�0����N�S{�b7?@2�C,Y.��:���
8� <�`�]�X1���<5�8oE�m�d0��w�b����/���8���0��YYCX���B�)�D��Q�>���,'JY�aJ#�� ��=_Q�E�rd�9t#Q;Q~/7Ww�<�{:RL����d�
��������+o?�1í���A�؍���!�?���e��qXĸ~�3�Z-�B;�X�'6�5��.V�$�uFFk.���)'i_e������Z�T�k��N�bʾ�|�]}>�o(�4�޻|�o��(O�B�fo��ؒBH{�<��-
�nJ;���C|tc\�w��ǷYr3PҏE6`�#�x{lk����`K�>����n��Y4�.	�J��ߪ"��w�ǡO�$h��3�]
�{�$=�D&�������X6#9%?L$њ���A_9O�����P	S��n�����C��S����)���<���T�/��Uܬ�q�r)U���ExB�Y�:������5���*�L@h��������,�6s^��q�;�nɠ:��_ԓI���,C������ar{��������_-xHC�\������f��贅ӝG.6�O�0]�0�"7+D�Q􆥲s��\���0���
�4DOG�^���Ĵ��u�갥>��������腆��c*�5�{�t�,��evFE��L|��?x'����flE�N&A)�op:�Swh�9:�ל���mx�O.��^���E� T���\��q?��A��e/i��V!��O��q��n���O�]9�W�����m��;h�&�� `�瘰S��d�w����Z�Gq*�`ƌI��,�j��JH��u;�W���:A�S�J|^�[uFĐj
�������_O�XU> �D7e���U�mR�:JN�����-g�sn��~��Ty�.������ I딕����A�ґDt,5G(O.����fǊ.�"���PD ��F��t�׶3/�3�pܓ�K]��|�
f��������?[�R��&%cбN��m~�K?z�!QS�!��w�4����8!y����|��-!"�n۱rH���+or�%?~��Ig�F+UH��A1{~�Vդp�^�o��i~2�^RR�VP:��?MQ1w-��_��=�Ƚ�Ƙı(��0ײ�<+�ݗ���`zl+ӂ��mA}!�m(�]�k�I�O4���TJj��̸P�"�F�dN�a��)��R���{���܇пR�.T�R2�K%0����+\�a�(A�S�K����[�e�>	��C�[Z>�8܂��'�)��>�����6�ƿ�h�(�Jϲǵ���!.J��A�3O%��Q�_��*�T�nX��ԙE�iu�ɸ$��OU�����D�\AI�e4���I>=q�� zd�����e�5��w�4'��3����u��7�B���l���DvIܐ�3�T,��J�Q��!i�L�" }(�e�qݖԍ�q'150�檋���!e��t�vk� �0�
�kh�䭬�j� ��$��*�NȘ��R.p�L
8��mM�[���4m4���W����6$~�?�.h�?�Oc��p��WeyAL�����H���g.f�u�b�;D�<yb�� 4��b��������к38����T�fM�|�m�=��j�/�*ұ�����(���?s�R�`�9��*�jM#i���q �>�=����!��[O`o -��g�8���W0qҳ>����aKcP �8@/ob7ekK9� �E���P]R9F�f��(���cN6hZ�4�ҧ�Jw�*	��1�;�C�K��2؝A�9�v3���۹(����ף�o�ہ�=!�>�fY�J���=v�W�ړ�[ge��UB�;}��CF�j��g�5:��?�S��t��ȯ�6�׹a:�()��6 Jܸ;pL7tcUc�1�B5�=�Zoq=�4�_,�4��_�4�w�_/'�=�*�{���+�����M�3!^�|
�/b��qU�LT��:ۮ�'�����t���-㺢:�`t��	*�=y����z�Nf���o�1x���Ra&�,�M�o5��栯iM�vd!��vc�� U���!���*L���0z��g��ٍ���3����߮*��d�xA=�k��ǎ�V'T*�dB�^�������&��P��5��@���z�V�<M0tw����@��W[=��+i������ަ�	����D�Z5�\�9��ʏ}	�ع���3��lH�RO�zV@1R'�Av,�ǴbH}��w)�W������� ��r�_����WF��Qz<5�3�l )��s�]�U6q0���^a����j}�Ȗ�lt�����F����4$/����neEjI�Ceb2��\xj4O���o���h�����-}9��!R5����9CFhw�5бFq��M&�S�3d9���C��n5BN��hs�,o�{�l��Q�X-���`��/����I�].��	w
�d�9@37׽K�<�\Y$�H�U�7�f��Q�{kĎ��#}\��e���b�Ud*�bG?��-��^�V�$h�,����u{�A�n�/�z�Li-^	)y�"�1�a�j��^\���?�(k3!a�$���
�v|��b��Zҷٝ�l�Y ���� Y�q���etC_��ݵXH��1��F�n�}���4�^zIjB�'6�B����^-<^zR�
´�p��"X����yC8j��v�����
k�[�S�#�Z�U,w��<�� =d��Ll�����~��`l@��2^VA�R���xʤ�Z��z��"����+,R˂n%H5i��Q����@kK�w���0"�4�:-p��q>�r�&�݋�~_\r)�������j�+2��Jhġ7������.ś��眂$r�%|�ۍ��-��e�~(�`�kaЖ3\�c�	(�tw�E�A�/u��۸�d0��*5>V	?P:�C�y����E5S�.=��U�j'���=�>��#��tur�VXz-[�ܚ�!�R6����2��.��Ll��{8 �)&�~{�ĭ��x��T�b�B�%GFhC� Rbf���zv�Ҋ�o���eܯ#Y�e����l�L���$�2�\G^�Aۊ<N�2-���|������~P8���r+�� ��F�3�!��9*�2���U.{:w.;���Ɇ��f�03�fQyy!%���U����I]�����0�_�Eox{q�Mqݣ�I���N�>��E}��Ky��V>�$5#�A�!�a�Ɉ�����Kp���Z��CH��K����6K��w�r��qLs"N^�eR�L�f��|(�3���~�#�/!�Ty�$�>s����A��7�Oڠe8��[*)'ĝ��t�I��F�kŕ�a"<�k����5�WD&@�vl*u��H��L���΅��|,2�'�� D���[�
~M���9(�F��CmE@��;���˸�p�\2�4c�I���yPY��I��>I�։Q�Co�i�
1꽤��\l�Bd_�Vq�(3�7�n��Y-]�^���	��6��-Ug��	d}rx�O�)!&��S�AY��t�lOzS3^ǻ3L�vЀV��S��?�̋8�ظ;���3&3�����[y�JbS�,5��x2�^���J|��e/Bz���u����:���P�XTi���w����z��KThܹ��c7��*�C���q8��0U�� ]z����$J�'D�=<����!��}����[l}�M�	�����%�	Ȁ3R*��C�߮����y8�F����&�N���4������&
�#�"��"��-�?�G��2���-��/Lج�2�Ƣ%���8O����c
�r�nYY�G��yD�@w_���^�y���QF�v��]h�c�a�~�:�)�H�L�����B[hy@ `�Iv~�,]/\α^��_N���q�����v<��ĸ�YP�RK�8_�cI��C���-w��J�5V����|��C��Gc�:��,㹗�*���>^ b�k�����ӎ�p7��^n�/��>!���L�Oh�#��Z����E�B���6�����01��,:z��&�:SR��7v���TS,n�vB��sVu��T��|⫠1P�}F# A-z�䕣���|�<T�|ܜJ��F}{2uƁ��y��Z�B��C;;;Ӎ/y�� �Ε��ճ��f�C�~)��s�Y/���{�K��Hl�<�J�i],��s�n��0r����C��<���&�u����|L6�0p�"���S����pM��Ku�9�&j��HE�� c��G>o��j_g���wNMʎ�.��ڈ>>�h��awi�� `9P
r�8���JFu��a<�F�ҫ���8��~�<�������WVH�s���-X�<?��ٺ��&D�D(������+`�,BV�f9��B�������/.{�`��2ų���:C���/���Kyt3�
_���wM�h1��R3&�J4�jwdv[�ȝh�S��,��z "�����n�M���NA�p}�L56�0K��vݷ0�(��5ys&y,�B#�W�V���� ?3��}7�)��im�b��3�;@�A//���=��n.��"�0�*�6�z @�	у�B43�<�fx��U/��7�`y�y�c����l����7�\�9�ޖ|,�� �=��X�J�[l��Ű��9�
|X�I��
�5���ۯ�'�z�5��*:�OJ�5�5`.J��-�b):�?���q����}��>?�i�knnz��T?�����*,�,k�)����w�칤��8 �}{�ȹ\$� Wh�ˑ��pN�J��RlU�y�%(m*�/E���.a�]+����f�n��	
�7E���@���*hk��¢��� ,���i��\�n�s������m�ڂ��n�DdՍ�гRu<=1w����h#~}P�=����u_:$8d�N v:����n���E�34r��;]���1�& ��d+<�(A.�B��b�Ո��𺁗}�L_B�N䰡��[������ժL�Ʈ� �3��K�a(�8��w �;�.���u�_�y��fg"/�YE�0��x��-�y,�l�\P��7*ez{���|�~_��������w�G���ި�dA�J�rn3�R�"����{�F"rϐR>^[���Z�Ɋr6��l�c�<Ok�̂��g:��+M�������̈�;ɫqcD���@���9�\slW�!�V�E�x$�a߮碤N$i��W+����=�{v��Ϋ����UO$Z!ۦ>sʏ$�ϗ�A78_y2�Ӛ9������W��$����!Sɹ.��R@SR/� �?�5T������O :&�I#0wA�[�C�_/�Z�(:��;��1.�}��:ߔ	5��c��Bd|Z2�@ P� S����x����{�]�N�[�$��yٗ��m�dWӀե�5�j��`�>+�dc�r���8�� Jhh�TV+dٰ �Y.��"t�WՓ[���' �&����*��/!���g,���|3a���(*G�"�drކ�����hGnk� ��
_�����7@	�2��*#3�?�x�$�7�	;���G)�>�f�)�҄���#�%	�$��Clo�f�L��� ��
�Cd�'6��>���\6����%�>�����i>�0�<��Gø�H:�x`���Z'���a�HC��<�Rs�I���gc�S��N���\b�y�j`"�_7�?�s�+���FF��Z��<�()F���Ĩ�M���.+�t�*�JLB�n� OEB��(�"�:QG��TV��`7���o����e׷ng�L����L����A8Gh�pZ�ھo+�uv���?��{�o�oC�d_�:4�e"m��ط�;�+!Ԛx7r%�[u�����6Ѻj��|�H{�q��{��}����C�=������O��>���NE��3ʸ�7�ct؝�v���Fa����� �>Tȴ��h��ʢ�^.B��2&1:�M/�[�\
�s��@]�H�#�5���\$����U�$�5!{�}����HS�����絳g���������K|HG'��hˌY��a��O�K7�jf�N��#3Qk��<��BV�
�����>]���o^a.I�R�b�B]��aECp;�'�,�G���Gy[i%N�Sވ��Or2��O�� �9���Y�eZ�h��G����p�� I�?wS��I�*�'��A�6O�Q���HҴ8��8V	aV���z	�Z��"{���bT�ZbV\p�d��5Y�VH�)�c1�zT�(dd��Z}�jќQkc�
�	n|��5��#/�՗�X[\蝻9���Gũ�&�5�U[����ծg=h��Cx0��|z^��T݅�L߄�峄��k����S�F���H�����s+q}8�{��HzBM��=��S��[<�'�n���R9߾�33K+�^��g�̪|��)�b�����-OǢ�Rp�WC��z(K1�l����I7�䩻�;���H%j�D;��2�!����_��iĦ@m�C[ْ�o�m$3�g���0Ύ���n>�_��K>��\�}'���:�7�.PD�V[io�38�('a��-_��N��!��M�,�~��5�d`������čTbPJęƹ�Y�����^i��YgAH7�<p� ��x'Ū���k)���9wA�<�U�B�g�	�S}�=t4��p���
23M�sg���7g��3��+�G���
�e\9���.�=Ab�C�����:��~D��+W�Z4/@@`c�;n�v@8�/�S���:��87���.�>��	2���mx�ͱD)��.OhZ�w(~:[�tٻS)�� )�ń�1#�SH]I���U�d��o�F	�Y�����b~��s.
�Tt��i�J@�ʠ���g('���h���#��T���;�(E��q�aև7n��z(C��}3��J�B�����H�6ך�^m�{Rn��E�����t�^�`�L��{�o�3���oGu��g{Yt���0�Z�V��t��^j���RY!�ڛ2�E�ѹƪmT��G�A���s4���z�k/�%�d�]������Kf2Y$4�؄�â�U�:��f�P�nY �T��e����~��r��}���a)�SKL/FC�B
���%E- �Iίa��_�o���-4��ep��]�����7�����NU��r��G��o�90��!+�ba�����F/ڭ�R�Z q�h-<瑖��4T�eC/�_tQQi� ��t�����b�� �k�a5`��]���y��;q�G�U��(��k�h���+�*R�ӻ��)=��A�#���d\p���Ea�Y�F�Б���'e#�`s�٭hr�a�5o��ew��M?��5��1��I��If)Y�ыI��2�錕<��O!�����l��P���f.,�rK
��+&�iZ��g^P�^�eT9�����Y�}$I̢���	�d���Dz�x�F�f	M�a�3��P�1�fCp5����d0���Lڏ�V��D�\Y%���=���^��0��қ�H�3瀂��~��1��8R�������<����q2�� ��(\���B�T��|���x�IuS�M�ƾ>׬,��G+`�;Lm��	1N�®�V�U�2N�^���!kc.�ڊn>�9z*[�-�%�1n�T�@C�`"F}��������׿����[šk��&��(F�d��V&
�<�7�Z:՚x��1Uʂs��x����`��l�N��kKw:�I̋**�le[�sr�v!��0A�w!rYag�$	B�NY/�P|�����̭��]���0�7`|��rtI��=<Ӓ�k�/�e[��@!����m[�
��7�-E�IЈ�{AeO1�;>�{PYV�m+:�zZ����ǂ�	�f��d�]ᕯ�)b�9Co�OU)Jn��!p[*A���~��T��P�1����-_����c?�^�:�!K�}��j��-2 <D���VƠ�rS�]л�-g�ᄓ)t���|M�J6pafs0$��4��H�ʏ��.Z��)a���1Ld0�`�=�޼�lxξ�m9�Ho������ڗʤ朧�L�o��#@�ij�M������7�˅��D�U�]��	����<�&����{�-۵q�be�6���i���R�  ~�����A����RL�Q9���$��)IY\z�&�5�A��`0/~���_.{/(��*_W��դ�l�����5��=����;x,9�{�&)�+	7�}NT/S�I�����0��JP:R(WN�ԏ��s+\�]�����h��� �`4���pd]��eZ�0�`>�(d�k/��U>s�J�����=r�:{�3&N���]��?e�&���=r4�E��Bsܐ��&�����j�H��W^�/&C!�ŭ$.Ν�I��Qac��R�7���[Sz��S�� &����pn=�"b�x 	G�2���ש�.M���e�������`}�ӫ�Z�>9Չ;�@#w=!d�����X�?q�i�~��{��h�����[�iH^;�ܐ�� �0/f��?C��TE/�S��,�6��.}	��F
mI=�7�%���x��O|�K����q��2��E��e��Φb��,g
��o��|j��?^?ur�@�C���s?��t**����<���p��}̩�h��2Ӆ����Eq3��%ȏ�᎖�1���o��+K�5�}����31>p5��ñ9�kK�� v��ڳ��$��޽6y��?g��Π�-���v&�b�:���9���NS�4%��fz��6O}�!�,y�:v���6���\CJ.ƍZ{��ػ��� ����]�����}����G|eh���})
��!�Y�66�1Ԍ��"Y���
}���}�.���pe�7 �g�[��X,�1s��\��?�NNTy�ק㨹g�G�
J�g&�k��875��M@:4za0���c�h�O�Mp���5q�ȸ
X��f��8����mU�HN8�/#ٹ8s���PvȚ�O�!3A�-liw�q�#�� ��P�����ę�h1*��6�
j���p�W\���'xL���C��M�R�#3�Ʀ�n{���T 
f��y��@��`�>[��$�"�qd|���>B��!aYv[����A�s��5n����:M	�U�r�2��+>��Vc���4�j-c"k��5P�)V�EsT�{��S�a�S>��);�������݇e����V�}C\u�x�ތ�Ϫ���� �g�
��
'sk�kx���2 �3tȓ��D�Wu#��a�x&)�I�d�1�B|6:E�g���Ax�2��$���W$�U������,�h=1��s�v�XSu��-;4�+��è����?d[7L���V`O��+���������[��'	*����oyXσ�͸C^�.�i����u������n�czX<����ɳh� XtB��Vf�7�s='�O(�H�	���>ku�_4|-�ſ��D��r��IUE����(X1x2�Q��ʃ���dXmp��ڰת�Z\��A$G�,��,�z��?���U���ntSF�����H��[E����^�=��oɜ�|��V��iM��DOt�f�:�KA(��b9D�/���>~yޫ�h��5�A�Go+�JE`=-�4��ZSŞ�
M��
�!�C���Jue<�tn0&Lr��퇕�X�ׄ�V;H��7�wO|��h���m"0��[+y�Dp���$@\��	+8�0GucR;"��xR�3'�Q�?N�B3?��k/�fH���p	s;��8��Z�5Q~�M�tƉ�{ڗb��h9T@��L�$Aa9(���	���8-�E����W1r\��J|p-j��-����UI6��
�`���J���wwgZ�D�p)��r��舨.�'1I\���J�4^��S�P_�[i�U�^��he�3���)9���	k��2��hƖ��j� ��[R�ۓ*�e�?�K��=n{�'�{�ǖ�!�m8�?g�{�:|�Ç�Qp��.z��� ��v�%q���r��������|�ĊgT���zeܸil:���(P��q�H��q��yF~���G�	aN^M��ʯ�� ���5 �7O�?Z����!\d�0ʔu��rM�㋾Z����X�fx�>@$?/���}wE��=���hYiͷ�o�{��c̜���O� �����=�I��d�+�`���O	5�y&�cɪ|�)eiKO��#�J�̷ ~�_m�6�:��Ar64M�������������c~'�$J�6%�$���!4��r�!`,�������k�b8&�D�X
����n���#����WSe�p��eKlSd� �_@e�su[�����s��$ژ�o��D7"V:�z3�ac��'�u��)���7�Zh���;)�������e
�3�M�Lk������z�A�`�����*80�,�5��-Æ9�mꛑ�*+��r�W���1~Im"���@��v��ϰA�EL�1�����ao�Gv�p�0��p]E�X��2F��;���?1���z�d�*���X]�0B�mr��DRό�*���|�����Wb��ƹRi�����j�y<��ʩ'-�.z�	�A�?���!n�ؘĒ��9[�j&�U2����Ho��\�,P�{���h��~�
4kg"����}�1��Ű�<�kO]���A�<�B�$�5����DDNѵ01+��ù��������	�vt���E��6��8���/�M^9�{d�Ay��4<Po�g���%�޹�.b!Rb5�uZ��ܲd��O�bP��L�/�9`��gzk|&���J�����:n�,
^�hj�	R�ѐ�xB{��aA��ۦ�J7� K���E�);0��"4�vʬ0�
�	<0�E���,f�jm~}ezJ[E\��VX�䤁bVA���Q�Q�������7�p�����="B�zƧ��W�;X�[L����
�E�ӛ��b�6����7e��D>��X
�����W$~aI���5+W'X[���� 6�VP�]��+v{�����¦8hw�|ڰl�)�O�yA�!@MZ�u�3�a[��P���4�A�nx����g���;�8't�<y4,�W���P�{�J�����D��B^�u�ϔ�;J�ٰ-m�c����O9�����i���/ԩ�5mw������@�Ǚ��3�9V�,���Tٮ��bH��鍖�[{����������NN�*O���e.'�un.�U�9�#Pt��y��4��Ö���6*��>sS٭��A���׺uN�m$��C-1vUa}���k��c`A$�lR����^�j�(�%u}�$ZCÈ��(��d+Q���@�ә�|Vx�S��.�3R���Șc�c:d�o&�����\nnC�٢��b������������c�P��ԔK�{�i�W[����
�;���P�9m;K��~�;�NYH�a��U,�.O��L㈖K��y|YPisS�M�Q��ף��ɤ&Hgڔo]D�����%FQ���tN��z�I�twD:���JҖw�?��[csj��b�U��t����Ъ�����!r������iK˦�x���d��>`�?z���"UG�G}f˵ÊB Dqv���A�ͽT)ސ��+�ηC�xr��x:&��޼���ION|�Yr���3%�FiV�B	V*�3�SXEd')������f����S������]'�\��J5��$C�]�h�(��n�Z*����T=DV��e�<�p.0׊۰U��C��mҨ�a��JM�ܱcy��p|����2���0�x�T���2R��΂92�Q��'�Ee�x�E�ɰQV�	��F�G���b|��Z���OI(@K���>�ieє��~y����+��iaJF�dE����bK�����=�� )���|��+ o�1��+�! C ���ӼS�k	�uTg��)[�sYL���`�`�[Ǖ�
�Fh��\{�}ʣs�+�r�(�Ѐ��M^P����ɩ�RI -�_�󆐱q�7f���K�(h�d7椇p?�1N��L�
Q�u@ٌ<�\�v�;��{��0JX���#.w�.DC��$���PH�9��@�x-���%dÞg��uS=0η�.�)�m�MO��T�Ue��	��g���/���'���%E�df��Gg��-�+�B{�rs���{��5C��<M���$-�
<���;Γ������T��_�}��SP��^��U�ډ��R�p�:���Kf݀p���ņC���N1b��'h��}�L&��:��=����)�o��Q>���g:"��s�BI���.�h<�)t�a-?L���ޝ�z[d���fovT�Ƅ�'{��QgR�߳m�;�i�Yi�Œ4U8�4�|L�2L�MO�F���}E��lt��f�0sҳy��Ӥ]?,Wyj:���@��!�����4��|Q0֘]��0���ny������Z�%�$�,;��e,㳮��L���2O?W^��k=�he�����5f[����9ت_����Zx�b��F�0�F��:�u�EʼQ�0�ׇ\�f0REz�$x�Ӽc���z��v�]�u$.ޓ�� ����%;v�hY=[-?�Gtд�u�>{(���Pp"nc��}���BP�^D.X�`�R���� �1�U~�1(�� ��\v��bBD�#���i�y��9ٛ$+g������������ĉ�>1�#��*݁c������8(m��D�?�BI䥣��-�~�,9��l��\P/��a�Ϲ�V�@D��fb��mN_Tf��'���П6�eY�ދ�����8k|��\�����q�>ll�������%�m|�^�������;��)Õ7�v��[⻽= |�!�������E�>����k�m$5�v�h�lDT����G��|�G�ϑ����,Uc�4�]G���o�f���D"	���h�D���o�r�x�cMIB��t����m:9��{ؿ9�����������0��,D��{�B��Aa���Mf�j����A�?��{17)�G~D��#""�����$����j��Ȃ�-R����C�_M4Cl��{֛�Y��r+�adJl}Ɣ�.?q[�=N��TjrvUԯPA]|�F��/�?��������.���[�A{[����wAA> jN�:�"!З�BO�QN�MB~~�\�=�����9A��}�
o@�t_��('�]�2�����j#9qf�U�i����?�R�9VD�>�͡/GZt���%��@����)z]���'��f��yݱI����Z'B���Ld\C��@�=����d�.�x^oC�1?�+&K�+�"�`P�P�xH���3�Y�];�P��%�A-�lY+۷8��/)z{�`+9��}*�5�y��QL��>VĿel�� ��C�$�@�T�&b�V����I�g�A��5i���v�x?��S@,��O�0��/H�̢�T��:'/	5���4||�.{��<��;�@�%"M�j�}-wiN���nD0�xb^9����Q<G�61�g���6�q�<O���@\��-��g.�A^�y	!��H�zyB8:�{
�r�&)$�5/��ėp�~[	�"#
#6A7��m�f�4��$e AA��q9>!��s���zE)ܱM�DuS���93�8,O��9���!�q�LU�,��I�Wu�F~|7�/ϑ��jtߊ"�I��9fp�*�y{D���YPE/l!�%U��ɲȱ1��̽Q*A���.����\���wKy�VF.��޸�!��-R2�(,{m|���}����1wѭ�C�-n����a�k]p�ߡ�W�����1�x�{�J���?D������iPi�����go�\�n-~�)��"�bI������Eq�H��c�!Z��w�>w0�@�q���cO�������� V��DUT�f*iQ Hn�eA�T}ݲ��~G����j�HC�d�����Ŕ�gu��H��\����ey1�C\>�g���^�Ʈ7��N��7�;d�)�X�{
?��F�CW�,'g=���TCel�CqJc�>)\��(��\�yX��oIO�������Ѻ������Pl�VF�Lz��qW���(�-E2�����jЪ@9A�� 5I��} ����ב��|��Z��4 �R���O�y���`G��K�qb`�T��}"D���C���>ʨ�0�-΅�(|��
o��b��S��nǶa���KS�7�Dc�T��G�
����pE��o�P��Z�:J��,֜:����G53���o�G�C�?��
 Z�x�=�u	�Vk-_��i�&_�6� �y�M���d+#�쪪e�t�D��n����f����N�8���aS��(r�2��h{I�����k��/���(.��UL���>��#����t��5�{am�h3���� �Iup��d��N���9pi�ڀ\�4�ێ2�ܞ�#��#�1ѻ�&��"�a�]7#CD�=�*y_�����GRR��O�S�y��Xd�
h��w���W������WB��_[>*Q���7Gŕ�y��T�Fp�F[�	���&�a�E�l�"t'\eNO^a��m�a=�),AͱG@#�\�a���l���.^���9	�vΪ	����\���d�*���ZDH^1:�"��T��s����,a:[+;��(ў�_\sb�!q�:a�/6�o(�j�k���0�Cl���aS��-��.���]��MS��$�Y�	^�2(/T�	ſ����Z�rV���ޤ2��P𲤎�rj�{s�b�Z�N0Vҋ���~8Lį*2$�r����+�,�GbIs�ką�̏�k�V2 %T�c��ZO�8���ŖsS=�,��Pװ6���\Y�=�ifu(��x��sS���8f�JD5O�Lk�bo��i۬59|[��ukS��C�u��I�Fon-+��i��ߋB��Pg��� "	A%�c���O�&�v�y��r���-rK�|��=���������g�P]qO~�:`��<k��{8=@��@�%�j?����W���bK��Cܓ��/�g���~�����F�rU�n�jb�'��dh
P��f�$ь}fvb��Y��F_�<����e�{��Ū4T�Փ��X�N�[���M2���za��_��Ӣ�t��nAF��x�9ڄ�n�97�_�D���[�j�D��ƵP���R����k�i�>��2���q<B
BQ� ��"9��8j�7v7:t��"�i��p��q���mg;|�ƣ%d)j5�J�zK�7���Zg��_�ӄ���ܐ���`�ȸ� tCѯ��K�-���I���dx�F�_����X��I+3�4yS+�I���u{ݹ��s�	�z�䫣6Ɛaț88ȥʻ��b,��.�]��y�L׷S�_��D��-n�()�gZ��ڻZ������E
7a�f�_t��2o�����K.�x���R��ƁƲ����l-ǖ�B��b���L�����,�
/�z�RO)�m���t X?t�>0$�d�d.L��(mk9r:����,5+Eid��G6�}nٱ<pyJ��;oF���V���{��^ O5g���+��ڭs0f��g�h��g%�������g�ʙ�g������s�.s�w�vi�n�M�:ࡖ-(Ts�W{�I2lU�֗�w�#.,'SRf�5�y#<�2�.�Cg�)˹]�U��?���L�U���m�Md�~�|F~BNa2��
$PD'q��d�7����
N9tU+�,QwQ⭚Ml��F>l�7 � C7n�Qs=?��K��~X�U�-�O�q�3w��I-�B��$ k�G\�U!�0BYw��I�v������0�L�-n��&��)֗�ۨ��}��ʭ�9���HNa��L�]��ѹ�ږ�?��e�@���?��蓷ëv�����쩟GD��x�������T�0�N�+4~[�R��)�x��.���vD�)m�	�\��a��g�ᐚ��G�0��j%ʤ�5S��*��E�2h7���^4[�\oK[�^:0�� �i���,��F��JJߤ�+�e���	�����m~�g��i��(�����s�Q4�l�F�R����.k8�:�2E�&��Ɏ�8)����lPzĳ��ɶ������T�養q\��L������?�8��-���F���B�H>�96�u��l�9	>�����p���{4�b��o*���x���3�i��jG�Q��c���\�����a��g������̿��b���)6�@��oD���^�^�?�
�|Ɉ�Jh���4tS��6�_������{�Dkv;��0�V	�+�ˍ+ǋ&���P>+ü�\�=x���T��� �歁&�Av��wӍ��cИ���^4C𞥪��E{�e�98�\-�����2��ͬ�xU6�f��߉9M	9^N��Ս+]�Ԅ�~�*\���Ҿ[�������E��{b����^�m�4�1-u�D_� w�m�65�̺Pb����Y���R.�"Kƴ�"����ˡ脄���5@	!��"*�H�&. ��s��xpBё7��(6�|��o��m�>�'2��v��D��_Ʃ���n��Y_�j_��y�k㪯�����O[�V�T­K�P�~
�	>�q�ء��Cx�DK����V�П���fU%�e~�X���/�����9��n����U����Y6ɨ�o2�V�Lnf-Cy���2/Q�d�es���Gy�{}�S<ae����G�.�ejy��Ƿz���m&e "�K'������5O��.�캄e�[A�`��^���.P�H,�}㞏%��]5V�=�EPL;���NGnd��B��3�ڪ��E�t�k�#mY����ť�=)1���{�L5i�����R��^� S̉��O=��
����GR�x��;Je��묇etUmG�1����},��3!g�Gc�4u�ײ�eA�P��V�2 RD��"�ͭ25JWE���%��Lb][n�1�x9z4�j9N��*�Ƈ�S�;�x���H^s�B\m�("�-�@^�-��y{A+�>uJ��h��l,͏ɤ��!wW��A��,$��UX�,:l*l�>l��}�{'.p 5��%��/aI#S����rT�Vv�1_���k��*m�TV~H�ї��J�Iݶ��6��?m��O���/�<��U����-�����w�7�\ �߮��NP�B_��'4���f�#H<�Lb�Nv�{3r��p�&=˨��?V6��p8��������_I��+k��>z�����uL�=�c��/
~���p'ڔ��,^��:I���)��p\�:\a������>�K�T�:�BVfl�vxI�����¤�qs�2���Ŕ��9|��y��m�h%G���6A��˚Ī+��J+}�G'�2B�wB.�f̯�v�?��5�現t7<%Mֶ0��o=�����e_EƆ!T��2�4�����m��d�?�2-��7&���#!�A� �(u+�֧���򽢟yD��I=c2�j'��]/�sj`q"���+ y�&DT%.�~�P�#.`���*��N�p������_��s�r�!��=���ً��q!dbȹi��F��(3E}/4w��i�a��S������3��� W�1�<��S�(K��O�]�F��'�h�X��A��VU�X�<L�M4�:ժ�*1��:PH��$�Ш���yP?��\;�<���Ylь��:��b��@:s�E�]���t�Pߛ�÷T3����K쁣zd��#(��j}�+�a"�H�Iu���NMu����:�yyѷ�~�m�S,��C�\[��ތ���G���;�y7I�����e����S�>%!v"2;ל_{�e�Ou7��5(��d�C�@h����,�ȹӤ�c�'�� ��k�=�6r�,'g1����Ќ���U��E�"���������/��K���H\���9 b�YV����C��� |��R'�-YV��os��H�G��`�Ԛ���dIE]���an�μX8^��%�,M��:.�R��a'e�{q�l+n<�$=n-S�#�#M��E�ɞ:�(w��z�Bb��C;��	w��+�=k�o��������?=Eۿn<."a�2�=\��։ ɬ����p+��p١1�*�匛h�?��A���PTw�@dŞؒA��L�?����$�a�;Ãմ���ua�BM5h � ����g'�*���`��{&��J/���E��d����ٲ��$("��@D;:�X����� ���vTVr΋*ܻwb}�����4�Q� �P&s�/�t��w������b� �ć����i��N�#��`u���G�P����^1З�l~s��ݰn뤂4<��rr��t��}	R	ݩ�����J�et��}޻EJ4o�Ġ�FqF]���lܬvE��)���VϮ�d;�&��4�W��p���{�~��̦�7�x��澣 �C��|��Oy�r+
3[�XѤ�T���o��G��x���C�[�	�v�?kc6H�́,�3�Z����l@B�������˝��R�6Jz���gЪ1��y��zw��� ��?�j�h`�k�c�}~�o��6�5�=2Y�/@��� K����;˶'m�Ci O�ՕcL������(��˝���P��}�4=���{����y����M����*~�-�9�S�#셸X��XUC�״���/�)�6�&Q�Z�S!z�(?����@���ʊf��Z!ÜuSI�~6	2�9>ᩒh��O�Z�cj0^�06yǑ�H�hKo�1��������ov �!�ԉ�fma>;�|ܶ:���:Um�׊1�C˶�݋�14ؐ�8쑷�6�MMj x\h�_$��9O,�x۝��D�(�q8�0��K�-��b'���A�|3Q=�Xض�V ՟
�;��[sV:8����Y᥼Io�t}&$6���Jdͧ:��,d�Zñ��2l�5A܌�*�q�C�{;du)j��W.��.yM���O?�j)�'��)��;��w�U �^1$��uTA��J �d���@)�/W�.�Q%
68z�­���t�v?[Szpy۠Ј,��n��o��� )���P��� %N��FF}�-
��r����$|������{���iEƐ��2�7u2���ί�l���ܕEJ��[ ��;_�v���ݦm����|��Pe��f��
���C���po�"��k�\��������J��vձ�t3��T� 42K�J��د�y\]^�7�E�"v�;M8���Ƨ�S�e+Z�?R��4|=k���0*���Fr�7R���[P�z��x����r��^ ��P�d^R\��ԗ{�2O@<��le)� z!x�"��l�-��+�/P�x$�k_�|3�-�����"x����û�v����W�uU��'�7��>T\�h>5c|���߭'a�0��,��0�^��tɻ�V��{f$K����|���p�;�x+:��6ɪ�{�BI�F���`_p�5��F#J׊�PVtm�InS�u���山ި�_LI?�t��,ܲ�4c�Hy=v@DE��,ĨYiH���J&����Z�)$�����{31`��V�w1� hqa�C��,��kOH�s��i�aq�^ݖt��FI�+	�K���9���݈{Z�)C����R����3C��k�ї��.����/qm�h�.��ZQp�! ���rw��W��0#���[�]Bz���k��/��Kz���@s��b;^7Q��9c��t鰁J�$��*\v�'�7Wο���".�+��D-�f ���D 5���L��9�]�WNO���h�>cK%�`��P����6U���M' 5BW�s3��\�ٯ��[�H���J0�I{�����?B���kH	N���{p#�&�Q|�|�`�Y����P'y�LM�!�1i�� u~5�<�v��r�c��vŤ�
�I� ���[Ȓ��N��5&���q_���;a�z�j��/g��H�U�h�nVUgk�U:;aK�~#\t}3�Yc�;�ղ>��zyO$��R0z~JjbW,s��vm��P�$�b��!(���դ�9?��=u܃˭
H�|�bg���lkV��ΚT�b|-^�g����R������`ouF�	?>�g��<$�浌��^�j�$Ϸ���T�q�>2��Y.�@�K��{���OK�E��J�F�`u:_R��/�TiJ�}=�s���ω��T��$�I��RU���[�\ �?�(��]��O�I`Q����3�Z߂� �K��8�E�$P��!$��!k���@��D�kR]2���|�%[1�n���۱ :vh�!�[x�;���<��-�s���t~�	;�[��&������}f�~o�}�0�T�ᐓ����6ʤ��?���$�lS,+�(��niI���$"�����I�s* NY����`,B�8X~0���Q��4��Ϥ�b�0TY�F��YM��Z��̙��/3�0�����cg��9��
ɵT�ES��S������X�|�at� ��n�����"��������y+=w��g�l�39zC���ˡ�Z�Kr$�uA�^�c�mxj����-&��C����6Ų��C����I�V*z�Y'��_,��hW�@�p�I�WG(ycԜU�M���C����"�`��Jr2H7�܅����ﴴ���*��ME�,��jL�����
�o:�b���SXQA�Uf~)6
M�T�d��p�]�QW|�8���/�7�$�\���N�(o��W\�E!�"fi[Lu�p�CN�UITDh��:�.P�[M҄;����a�̢h��X�y�e��q^J�/�g�s�&���o�b�[ؽzY��MJ$ H���˄TM��+O�B�� �v#�B����i�9l��\R��G�J`��g��� �@�ӖY6xN�rt�6d:��0�lRLe�� {u��,�_��]ۤ�bW��x��3��CP� G�`;
0P"��F��'�u�4m*	��M�ɰ�C��]�/���HuM�vcX�c�C�h�`}���"�>������!,I�g���nb�?� Q���1�r�n��Ja���F����,����X�����g�w���VB���ڈ� s�-𒀰ԭm�YH��,�3�,�T��ƭ���3���}�zy�j;��=��\�>7����Ӊ�H ��"��s��AS��rɤ$��~8����k�ӌ���siH��������ׂ��վjE���n�e������Z�]9VH��]4�b�iu,�2����'ð5�c���^�\sb΄�b�nmr�]OQ��l>�޴����cmxj�p��#�6?e���gt��`w/���Yp���[�D�~���L�!X�O��o��Y��纫���¼U �Ɨ��t��V�4A0|zz�j��|�k��&�<�w�ʌ� �8}#?���#� zV]X~C��Kah�g�0�0�Kd���qX����)/�/r��!�Snv�*H���W��BE�K��پ�ڡ��Z���#ze�.��w����!����g��^!��Jӗ�j���!{�pY hZ��;h�b-S#qY|��T�I
�'(B��i�x~���7��v�
�^� �d��L泦Erۢ$�Q����v���E����?�WXv(�*^"r`S	jV���7nsɦ�&@!���bY�4y��n�PU����
QVAh����B��$�����_�Y[q<��N������OH��y��S���'���jQ;2��G�¼3��L.ȝs���Z
Q�̲᱂��t�0aK��JQ`�'�O�J
n�S�5���-�3X�������V�����o���e`'/�]�dkBe�~ֶT��X���
Y�0Ti�ѝ�0�jL�ˡ�( [޲MS�x��oR ��>�~��X�]�,��`p>�A]���?��4�.y�Hf��$/Z�%�x�d�����-'N���CN�Xf�7|B�I�E��f!]s�.����Ld-��zqU����V2�W�����{P0�H;��D͎u�H§瞇~��ԃ���%0���%�q��6�W�.*�!����z��躌&����d���8�#����f�#��*ƚ��"��-��<lؕ�E������~&ǙS���^���,l�&��	<P��h�[����y�AqzD$��%?������J]"|��,g,8Q�o%����"�l�(�@.���}
��W�
��?�|��OԊ �oJ�4�����>'ǿ���D��UcR�`�$_w��
�,�5S%\��\+:���D�� �2�"�4����	�:����oi�wz�B���B���Lcg��nC4�[g�}�o����������k��i�6��dw�|N���7h!��s�ؐ�������u�]pU�[�L�M&��?�ˊ����)'����Ӗz�J^�T�HB�?��zn�K�v�ODY�?��a�#T�+�Ody�:���z��Cg�$'�^�o����ݑ�����_)����^���2ZzA�}�0���.�u�ʊ>Ύ�6�4<�lȥ�
�W���8,WuD��o+r`,���Q'$.Zr��
�Xfޘ����c�������� A;���!�����z'#���/��pE�W<�h�g��d� �)��4��n�P�d���"��sB���gwJ��Ex��H����i�����SzӇ�w����t��_�R4�[��[6�(��V�9χJ�,�Y�� +Sy��/�2�d3��F�i���dMR�/���Q+�v���J<[U2�M/�l4��_�_3pJ�9�}���{Z�L���'�}���N�1=�{��Hy�	d�����t�@�fWx��K-��G	���g��e�$A}|�>���&x8�l�Kz*���]*��.i�<�l?��Oa���I��q�����̤e���Ų^|�����v�l����7u�o����~���"�1���P�K�{ƸJ�/RWNi�XV�Ww�� ��$m.�4՝���Úsa�T_|�n�f�?=�e���J(�����kҦJk5/��d�_�!"�ᣐ��^�Q���ql]7=�an��2�p�6C�����iC� yٷ���6u�1y,�;�W_��7cZ^�?���^��K�h6<��P�^��ևnB»xf�kA]��i�vD�s�+�����˰-}��1V#[���	ˁQ�ߓi}��8{kU
�`HB�.�����ҏ��i��J����������G��$a	�4v����]	�kACX�U_�vE�*e�I\�����x�9~g|�7$@ ��e�;����VQp�[��<Z��#<���4��*��dN�	���w$�,���M'�'$����Gx6tM�M���Bzѫ\�/u�W0��ݠ���Aeqo��(�C�z����Q-hw�r�{$���ނ~�Y�+�_?��
�q�*�yO�*
���Yq+�"H��?E��uZ��ɆV����y��N��+ŷ�ow�/}m�ٗ�����QAbI$�k^�5.���{�ֻQ�pP� 0#M$V���:'s{N]��[��$aڟR��3���D
�k���'�W��S3����K��お `8��}j��7l�6Toid�bdڊ_X!�*�������
�i�H��Lc��/��\o�2����SP�Ǒ��)���t���KL��0g{@=�3���3\S09D���"�hR����u�jDά�{u��gy�~���Ł'�xDJ���F*���~d�'͏ߌ7{��8�+Q�բ��E�c���%IhYW�\v���ȣ�2�$l�g��"�6�2������$��W7���Ǡ��$��,���o�9��Pby���t�������J=�7DX�`N�e��309�������~&��a�����������ä�W�t�`،��ePc(C-�*,�F}�@�t�Dq��S7P�6���a��d���Q�Ӭ����Ac�1��b�6�A��70����OƦ�w��k��V0P[":�sE��ء�Ocf�'���}�lw�*g&��F�Yd5E�����I���u-�����=��χyڧ��(r1���w.�I�+8�2�����R`(JƮ�p�ҡd��u{[F�hA�lv�c&	Rξ���E!)�(O䑖o�G�Ik�x5O�W0�u�Aʭ"l���&�������������R� �Ķ����?�Z=��NM���d�Ҕ�Ej.�,���������*��G��ˤaT�r��%���v=�����0�Gg-���g(��3�&�$�@%�r1����q.��Z�|�kJ5����d�?���{���es�4(diD8�6�0R��	&����
��eER������+djŮMF;��j\�����2D�K!G_�0���L��I�'{���PLM
�	P��@	��}|�3Km@�|k��EܜD�ZC߅���K���s���k��@���Mu[��ǡ:�r��ި��S?!�a*6�H�!�S��Q��b��rvp��J���
������0-22�kכT˕�^�"�e��5��P֯��y�r��A��@�6��X��<�ɏ��=Iy#T� �]�@�A�����i�3��S=�+xq_&YZ�� V�77q��
�����b�Ks��� onH�}͈����~�m�j�،���Lg�c�2�N��6����l������A�#z����kjI�{U$̖��q��*I4p�TGT|+;_��҅~���o�[���=�m$��!�Xp��F�^v����Ot���@m����1��8�~K��i�̠�W	���{-�2[�`���[�7Z�Q���*��0{�[�l��z����q���x`�[	����w�PFX� �퀿�����\͸}
�'�W��M�XT���0���ea�t&0�t@3P��pܖ����].Zk��Yr:ǧ�P��bY�F��Ģ&䏋@��������&_�Q��*��Y%{x����K�����2���H��4]������������o����9�T����K�C��ed �ĥ�Y%iR��/�b����k�C|��h�'��+�TQl�S`hBwF���S_�,�6mG�]��,�ؤ� ����5�%oJ޴����[�� k~3q*,�"l����{qPv�/��D���=���ΗM��P��#^|�����д����*��L�.s�A��EՂj�p�������[�S6��t�I���@V�G�U�94�%��S6��#�b8k�1o���Wl �D�Sꗯ�#�6P�$j44��*��&[��o��@͘3��=-�ٻ��Dӌp���O�%�^�A��4AoĎ��K����D;թ��g�PM>b�9��YO����->h��ʒx�{�o��)�XE�Pk9֨|��~C��U�/��`��K}�'E�hь�	��7Y���e[�̏��2ѻ�u�j�DIK���7V�W�Q���s���2�e�]uQ�`l��kZ����s����[�i��L �ZlsQ�=x%"���X��I_��b��w��0��鳈���S��d	��kT�d3i�9�=P5�T�~߭�RY�9��t��"��ETp-+\��?��`�!d�g_iC���PBa
�0�J�)�!�)�jm@8�k>N8��q�[U �s�=q6���v��S�8���MK��4��8ay�i"�&T��R��O��}-�Q.�e�p>�3��Dl���.��-d�u0^�i>>!���N�`L�`�<v�g�����6���U�����i��j�C����h���dtVц���@m��mJ��{�j�����V;"*r	"�h �ȸL��&�|MȞU�$�M_8[9�aUIG�+��Ħ8��a}Ey�:�P�*�N97 z%,��H1?m�X'��}e���x�Bt���Joʴw���Ҩk�)��Yy	�5���|�s��������]�%����Y�]���gU�KҘue*{抬ZF*�V��(�V����Gq�8U�Xp�����M� ��8�@/��|ĬX���&I=>��J����j���8�-VL�a�����R�A�O	܅q(�P�X�(�&����Sm��.����� �ڋ�
B��S:��%`|UE��mH��7v#Y�v��^��p�(�yǒ����"	$�G>�r��mt<�/A:��sf�l��d���c{P�Jg�vV̆��ν���9FI䌠
F�
IȻG�K�O(����ƞT�1��VŖp����.����5˦*��{����k�ʏ
�
�� l�7��ldQ�F��x�.��?8P*_jIK�Oc�D��	Jp�	<;l3��J�x�UȜu@�z�Qr)�͈� ���?�.%�Z`.�����`�{�8�~5jЂ&\?���9����W%���W*�?p�]�#z\�vZO|���U