// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:28 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LqzgeBguSzNC7NXMO7D85fCpT/eNUnrTGlxy859gj4fuAbHmVqsv4Unm+slXYlCE
pKtxF8ipSKPGFkWWwIk8RQVABexfIwk3t3Wf3OikuBZpBNLXGSvFjuEpXIm8gm9h
Tkx47d9/Fs7q4t0RlHkwTmMZLvsK5xAVdd7Nl7iwUaQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 100720)
Z9pfQqEuuhO/97TE4GvaCyFwdPtkG434MS3dQqxNAWodamnE1Fkoro5q7z3G8Fvh
v52tHtH63gyP4NheDaI/Eog7PkeSg1Krg3cUv4NkZ2Jinc56EaLQNtR7csAbAmYj
PSWCkrov+GM/EkxKIC0+yvjf8YFIfgQ28ItlTXzyBrFFrY1UROmSb/kirHUZCZ5l
E2+4QItWAqL2AtX1a1FY/9H+/4gsJzlSlDM6ZAwc2+Ab6C2CgENeqBCl6OvDBDy7
RWwyE30RiidzxknsRML703Nxlc5es7gX2+qnaOStCtgMc7TCaMjrsWS7U6hUIDs7
uHX0XQ0hdAa2pxUcmBZgqRX3U/zIZcVc6aV34BIZIX7zSaTB7q4NcshO2xw69ZQM
OgiWoXjgHR1gjyZ39h+VPGEJBRw95GakZiFHpdC/7eT8pUFUCpcB75KXrge3F7yb
TtrUu6M4ykATbt7/M4t+94jBtruUym0Iag0ga+C6y2Ownk3LvaMDCs/l22n6jChQ
2bXlJt4EzPpcDHHfbQklikn3fnn78tcyFXCeSF5gMHXRpdfSwQ/t913OOcxRBwqY
JOKOtQ1INiNPHAxBg8154IdBi5L7CEtCK93jVQjGCC627hpxHJEv2NYHB0zT8GB2
7t3BC+a0ci8E2pGAIA6LGnBuSyB6K4h9ZPd/G/0Ofz6affjb4lUoxpPybJ2bmHWL
BdAUqC8+00TDA6y7QrDwT8bs336R6NpKJFJHG9W+XRWBKP6xq4MrTXdYeOMBle1I
tQhzZIrW7VyKr29WiN/x7T1eZLRUQLlD/dMoEs3ivYjpjBe9f05xLGHjW8H/n4JH
tP77Vjy4UvCgQ6ucrT5yXjIae7advN6xclyATu+Li4EeSxOSHL1v0Vmuk/Qpb09w
iWmaeSTbl+0iYxC+GcN8AWXBbwdCoko+jNJkKVVWKKN4Lf+TRCh5H16STF6Oumdy
MkgPi7WYAjrIR26rrDyDMWBZpo5FiwzOiZycpvMokZMKqmDBrUWsMvicKmnlvTEC
dkgFGHAJRTLXjAIk8j93wb1+DQsl6HKciCANhW7pR1InTAiewYBL+kbd38JSX01N
aAgKBMN95v0fBfYYpOIbh2r0EKwCSCXOSXnRPNUZLHMMCfbpv788cFq5B5dfYr1E
VLZ0rtJPMX39cglIBS77I9zoA81wUQQTDO4SeIY7cSn2eMRZqre4MLPveycV9Qop
wnbaez0vxck9xkLRfEYkDS7zkP+OHkvVqCJXOdjQ+8o56SJHF3aJX6qiE3vGcJ+A
P9tCEeY5LtGmp9deCsivGF3RC7/H+9n9ezVCqHL/1axIkH7GbZ5nEXRTY2wmwzup
i1PuwTtKywkI/TS9TYZbxq5n57B54SbU+GKX0r/5s0fsrOsuLoEwDa+RjIPpDKV5
4UlN3rjONH1N3FmqCR1fphgHQh1UWHCgo5biLao7y1JWUfjQI2vfy4yv+HgcyVZE
SnBl5YNGHQW8Iyp4kXIM2OIPaKH2fMi5w8IxfH0qz/bg/GRpKDaavK82bA4asfNl
a+HObOG4pB9R8XqGca2f2J/2aORhptmxZLLseH5fliGWKEvl52/Qk369McS50oZ+
eKtLoeKpvYsMuRpd6fUwwPBltNb3wPqLA8IbnisKwgGfhPsk23B85aokoURZ6GL8
piGxGcxYjpnGrEjA1zBWU6mmQpxEhMRbaIEk7i+7TKLhDtDQjBKF7Y7ROm9Fpvdv
DS6UUNHj2xHQ2QwoRduvgLYlw9HFmx0sDJRZO6W4+VKe5URhVK8NtmEaIe/LPOXX
r1fJ+XD8ucyzB0S+9vGsRvrQBvT+5Pos74RJpOzuT3p+H3d84/jD7NmoHpU3n+LA
wimpKs2Of1K00mim4qQeAuLyrujfWwY93eLLcdwD1kqSlG/TQg0baVHR4m4yRK5/
/qEy7h6pvPxgVQQzwZVffUjWZxdXzrzu1+gZc6etFNDgb0bQPh7AdzdAlUcuqOqy
oQHUeMFH0y11vUzg3qz9A6RLJ+J9wYEuWCcf0T7OavALZnLJEnOmZ9M/30NE1Io2
omWcTk6LWrhMav7QgzRjjMIj44H/dkp8T6+ePVA1Nxc5h9YmpCPq/sOOwPXri2dX
3qk/19JamjTPivERPQd0uRg3djdUszoHg8YW6qiHRAD2Oca9obLLF9P7nS+Y3hmS
coiKVFOBknuhxwmOENqRWvWlkBHc5OnaIHxhgNjhw0y5EpYW7l+QP9RmfkeMav7/
YT/Q/shQVS428Db+4JjUSMzrHMTvX2PEsrFX574WLo7//mNR5PBQ5tps5OLxrA4l
zqXoyvQTNje5W6w+SyqrPTJhOovou8xSV9BpwyUkGLwibSHO0vd06Y2ea9Uqt1DB
k+JS7aNzcxTBhUmRDjLUDlzSgZQd2NIx+93Wlp4HBG2rVeoFF08MdID3FczOZx/e
07o/flSr420+FxD2emEiTsn4PuvVmWN0LfidW4KlpKBbzXEF/qf0PPZATQhd0Cgi
+O/rauPnvsUuT6KhacwHP0jYuy+C5kDCHvGU99tXGcy8q2LW2GTkffCcW1mjpqsU
Hx+JVzZmTx7cdP5OPyTIrELeq0F6Pqq57IRjhmt9+HSH1AY6siCP7HDo3jEUTsYE
wOeN0qcTaTJLrb3KKNQzwucaKgFQSVfinHFbFpaY/zWxarnRhz8OIF/KQ2dnmm5+
DPCNaPWkZYPHsWe752sbwOS+E6pD3E8yZmUYoVw+wdAitCXNUJ74Vw3zeE3e/fz4
1qzdKxoOjvBoxjkfKB1WPxF+ESHLY/j+b1tNi4clje+4OZ1zWDN/m3HFxK6czRCx
GU4Go9gnOka7ebbQ/C4gLCeOOImvjVj+k0OGfe3Zw58xvprw0Lg9wVc4aOBR/a/E
rukegpjVW/h7E8m4yOq/jZiNB7KEgWRHraT3s26a2MdXlj4eeFhP6/eUERZzYSSS
O3V8nyzVH8CtO5ewfHl6FXcoNQrET51sRdjIJ7UiaWQ11HfjVX/bC6i/hdVrm2mm
GRcYPdefgrle8of3z8XPf1jMJAbovrR3dZhTVxHSe6J7rPSNwnaF9qD8GJ7K2WiQ
K/eQe5qLIxZnLFhrwwsbm+avGTngLnPuvY0hxscRkqM7U6QlvbW8bOztQOMYEo+n
bP4FcvNvXyfRbDbm5cLgYzVYn4Lyhexgq0BJExXqR33+Nig32EwTAEbhD1W0XvYY
1WWyfPmDik2Oac0eWbduAOM00EcQMN7pO/A9oEnIILHCPVUMehKGjgHIqpAp0bhZ
VdIkGetvWUq6wlTxgJ6sTMe3SchTRnhYBeTH1YD3gYJ5G6RBuRUTahYbSWZIBO1I
LOjJYUV9WjJVrJGeOZadC7+MUPsTarbcwNvZOOxZqE2RHrg/fS4SzjjP8T5H9e2i
ZWKy8Nwz3H7Xmhsapz8iXeCa8Q0xYljpNBPf6dPCRPOTtgi9RQunXQw4dYsaEsNu
TuB9B82r/O9tTYsTQ2DFCuDg1/qfJaodvDOY0PrMRtWmnk9Dg1Uz9zAiuMib321X
/oPNEO8yeJ9yHhQkCrXj+16EG730DG3lvL7/DQZvc/86xeRpSY62hUt4yUKwZuNS
v2rFR09YtSx2Ji6Z4YBTnK5Ymq5/27TCZMwleexmYMmt1AgBEl+LiQJRQSop4y3v
Qzg/1H5p3seYFF4Itjvcc8dDKo+8MBPMGEI48VolvRslFR8iivQ/AXONpP4ejUJp
NOB5piLiLuntP4MghA2+SbvLwsvsEjSFlC2dH53lcL5wUG8nFlqOQE9Ge8g+EieA
t0+xBixPCl/R2VkVHg1nFSVSlfbjWyb8KGCOb4z0Dld2Otz2LxdgqppZoAaOxbbA
SFDUskY6fxVHt9MEOIfc1zAp//yGQ5rcdxSDvyM2n406HwItQaZyKi7Mf7yaRm+g
W0uCOH+Q7IbkBSaZJ2IFXWjNSxvNf+YVSD+R3BGOQ3Rjh/RNn+jbPIb6oXR7/LUK
yZAcOI9RIzP3is2ft5GIHjItkuUDxA0Cz2mT1t/S/I9RVKeHk7EURmAd23wYoIU5
srHDr+FI3kFBDR3zaanqZs4W1enO8eq1vZhE2aqNWbcsb3c+qTXnPSqdnB8SPGfl
aHwKiarbLjyQHaw8oujQZEc+YTr/C2g7Pr2LSoyXALhH8ro6Lph5/lcmqVW+TVXe
5RdJW7tItDWSfX/uYw+fHYaH8nj+3VxEXadh8LQGfJYBK/qvOJLg3MRl+6q9Lwe0
RQp8nMdLpVV762/Zx3KucwUY8vx5NBF6OdOYLQYyoG+9kuAh+5slSf/r7hvk0D8q
5S1zaQ9npCwEG9cJYa1jCplAo8XoXiZpFgnUV86oPD8kxJzKjaQlfubQH9JYXaev
wUB9O0A/0axpySVnyZ4P8DLL/tiUKgJldal5nEzZJoWFPrdd/hki6VeYFEBdAJGw
x8PSQz5BUV0Mot1hi8jxeRo3BjTiR/ILPvUY+qh99s1s5YbL8M/LU0DGAYVWNhKo
GEFdOTTDN+cQfAMOwlYiySm/XzXO9Ho4v/zR0im96yiVnVoGJ4itgfTsi4bjwOGg
bCPDERON766rHqlcSQYz+y7f2vGi/yVoYHcJxsny/IluWPhPasaRtJOoZHln/kq+
c22OJGG4AUZV5AoRBAEMg8PVKHUoESUAHQW2dEYiyicYL4ZFQvcxQa2k9To+D355
f1DROvHUjVLnF8WAm4P33T+Nqzq2wI6AYPLbtcwBnr354vJKWXs/HeFFvumK4yK7
Y6iQzEmdibyUx+w6BkJWHd3w2XITfAFKa4BjxdJJWnrUtPoJojHLu8O5HSVolzYe
U5x5QhTi0n9cG40uyIps9iecaEiCtzzlsYYzv7rEySpCRL/qe+0jmA23+qtGdYTK
BU+fzH1p44YQkZXH8kHL+4L6o1YLVp7DGqJdaHgWEeSQphHRykM/wtnwFotYoUwk
EEv+WAmSjtVcufUj4agwHMPaQNcCkgKUzJ1KcwAzDRWmUUDZszw5YqvHLajupUtr
brQWjryPmHtDJn3XZHazjB+RjdHWn68E6L0+9diGLTQjwx3EkL3fYms67BV8QaTz
5WOUVVDNkoInh5tBBvro/WPm2puCYzuoaNNeWUCjtaW++8Maz9atBop++yP873KC
ovLH+dUHF2swQ8oVIDUs1NM46eQAlLBfqzi0S5LpclM/K1NkrAEMDyrc13J/ZHUv
m9AzhgVj8lvuUZu3xhmy3mp8Qf73wIfm77nPB8IuqbqPILVlaJL3wpTiGMSjHxNb
9/xN0vqy2djLeHdc9AfSMMrw1F07o8A68mcLF9mI9isAP3mKaAshU5m/InTpewot
bcm334pXHsssgVxAa3aSQ0XC1ww6mLqZd1irGcHipQp2qrM5/3jATuZ1lfl8GdQL
Nnv3wNzo6WlJAuUno4H+YAlD4NHAW4/mzAJDhPV10Iz2sW/Yp0iWFOVd9j7Ilcvu
SXBrZv8BiM/GySVatvD+9h3SOy787ddl5Vu8XsSKpx1+IdB9KUkaD+XwY60483VW
UyYxF5OpgrZwULqf2d1CYGn6t7pTVleX/41Yb80B6jVDd+dWOYXnpbx6wpV5RWvH
ZPAMr/cN83n0jGswVDyeFO6gtdxxIP/aZvI3zvWntC0ZfQjISVB+05yL35V6Klwj
GkHaY4I2NkZcuWf3y1r81qK5hSnCmYhLg5VNteBVImVwBtYxjkj3yaj8VK0KB3Fa
ymNzM8Kikg5nDtLpj8Oc8K+OhKxe1bYyIUGVOSC8OQ+ia4PLzNOnPIs4VTKsuXe2
861WpSkSv43/aSn1V6+8hRSTKPhmF014/hOBTiaKsJjw8ua4zMXm3PbCibN/PVvT
se1kiYmQqAvYca6qmgq/3rbHmTEh1ub1GD4KlKB/hA15tyDRvv9p3V2gLvw6TcxU
SBbnDqWrC/UCcH3vjX141M6johIsRElppTyW9nI9waFacDVtDSpiFlgZnmBwNAOm
Z2tBSWAEmSGZePmPuGc503gwpf9gIolViy7MUeHDRTUZfZXVkfxnI7XdstAmsEIQ
wtHCDRSgVf3xNsF/89cOwJSC1mXHvGVyWwo2x0AKsI2/8+CbtVDx4SPsIK4Uusw5
GhhsgxVH4fNsEln76X9TidHM1jG501hpo1yz6VrivyeoFR6lQeKjUJkHUd9bCBhW
EsYgVBD2/QFGxHLSxBJYzFfiucjIaGuLf3JUkArBXPeyV2YcWkNaDN7u64IZPemp
AsQ4kzi4ZVyq8m8J3ampR31970u5NO9cK19NC3Do39XTbEzSBYkqI9zJCs3CShzT
RUhtsuvY5t5nrenGFSg+2ucD1TR/lxsowr9dn3i/aEEJbN8vj+adTSBsgRkHGahd
cUPXm/YPku++6OAeSlAnl3P66x6zPsoZA7arFgQbM5LHeOGidorg/EBXJXNo9AES
3HSdl1r93GGqGJRCz9LClrp18F2po9yVbiiTwI1WR2OBOAkRmimDXgnB5WVwAi7j
0mT/CzgsJAnmoc3mmeR8f1rFeSXsugzGmFxTtn17rsRWFmnW979kY2zUhYSD5X9S
f5zJmc6sMbE/wLGDjNZL3LK9y5nNlat2okTB8Gq7XtjPCdsiOzmK+lCaOuGl4/hK
LSKrcH3E65GlYoYouisEMgeh5Up26JKVV6jj9M75cKgzKe62aywNqY0YwrljDqrY
l3GfFribfmmj2yKtDZIBjI6vKRqIIbAhhm/7mO9gKztdtn/PJoOiHdCd60kiL68b
ayiSoQbcKo2IvZQAyYnB2HI+BwiIlkktOJbaRDew1inYfCSti9uH5Jz8aZC4JrrR
6cycrzWLftYMXXG+TpmJUir6J/578wmEST90Wm+CKznEn6W/ADa/jnt9ecoMnpEp
U42vklI2Ke6OUfWT7Soa854trYLiEVWCJOvBlJ+9peOGgOGL1a9fXWY35D266qlc
xJwxy/5UMSQDOXeHRvTPQ2NPkjFhbjRXrh8cbSnHwKWkGFS7/7LSaCSaiJ2ZbbYS
WMkhMp/eCgqYLMeiL2/wlKIQo9tGWq4YU5QXX1u6G45kHC7b+G1pigV4h8f0Ym+G
jzNeOR5x9TZ64di/zHtwIWpYvhkOpr6uoE2KINgQx2ogRgg3JCrTI4ibjrFGPLOU
lEY7ixTsInLDRKVoKhPMIEu7pVN82PiHefKwu4ICDCc8iZYrYw39y+yQ/6x8jIw8
Q0s3KID0/4+CjyDiV+G+LsVKW5rdq5KpwkX3tdvtf67O7z1xRJ3FGJcSdNJJuBpz
+Fs7XFuC0ZklnzaN1k4gSZLfhDFdslrv+2GB1zq5XAGhSgXGQe2d+Az2zVFR1z0E
o98m2HYJmNg4PV6I2uGrhZzu2ei28LynkdKDWcSetzMcaAAyIO6DQ0ek3ogvTq5Y
H5yqYu/ceKy5Omy7gQox6gifF/nP31EJ7Ada1oC4cYUQNDEOYVMtolgOwvTUk5uP
bvnf+WaE/nJkHPL3mRmC50J2LyjjO2TWHZYH/i/v2/2Idprqy2cgh/tyjHjUbeQu
eiwjxFNlunERYAh0OFZcQcc517f1mG9YfT+WzoC2aysB4yDxcU9MGKenkIV08Gva
1ajRDvLkZ0GF6hGQuRbLWxQ1nd4m2fF8dF6DxxHc1Lwt0vsld9EBaJtF4rajMBjj
7DF6m+OiYVtAnpr0sI3ig/20pCXiUkWiVylAHD5VsYwgULPKO/wpqPzb4M2J0tAI
Dsi6HwIutZJyMuFgQG4ig9z0XfKDVjsqE+tUEcKYWBWWIVhAcnWvpSETgV73rDja
xv2gAii2Z1pCYco9F0XQo/KiJHTHtZTR2KqhZG2WNHkT0OoaXXbZmJxixXTGfWI7
vRmvq9W+hDox54fB19brqPF5vhafNxPvNEKvAMpJwLBFaW13HAhB/OgC1cZCLY16
XRMp9lgr456aLfnGBpWJa5uoNMJE13KD9lhkvBXsNHQYv5Ya6xrAvp2fAof4/0nM
QwO0PKTA2tihEdrwk84BGGXUWR3j0MehQFXKdee2qcgSN701SmiBxHFAoQOYy6gE
oN5XUp27gHJomu9KRB5Euw7CCVAvMoqCMswGwSnetdU3LY/Wn2PcgCfW8HLIBasx
lr6NPSKQcalzdDwhL9a10U30iUlBY8O5N18akpGBsFn1QOHABym/rv9LbMncioTa
zbGv3AaTahoRJvwznQinU8qa+bKucCmu9t7hpzoX61w4aRfYM/FCg3GSMlt2L62K
OKA9NvWARcKfYoo3PJ0OLKGhj0M5Scx7O29FgqYJRFTP7/AoRUkt9dfQ1kobS/sX
PSwqY9hgng8h3MaHcvY+Lk5aP0vV4hXid79dnyJJ+PEDvnakifnhdQW7lHfg+ney
+rGZWoYZxPhrjnS+ifDfn9bUol2p42ZBkZULjWM/c+oz9dikzPr+by9GJ0FIo3xf
9Y8XiNsDib/YlZP2EydWCNVi5jDA55UShFMGxmGhcwHiG0BjqS6MCfhr06QhMuBS
F4FFQUzs9wIM4SIgtIGad1e6yhRZiGvpvivmGI78GlOIM/Uj8M2PduWxuglaIwXD
W85SdUNBUBOLDth5YlUuEtmnqK10X6ZTlH+o6P5sYj4W0XOZ5SxE4TmFpgMX2btl
S0RSBoSGKUh4ASp/2cjRV0gsUWSCtIWsYs0hXt83at23WjsSWKzJVI9dJsd70i6a
U6DFVJQ3J/XPnZY93VpKvqbwNWtmq54+n8TUs/0IOIRN3kcGuv+6n4V2BVoGcQGZ
JGNA2q2useYd4VZiI2RuuIp8m+v9tlYeJDVJ5DBUJKkGJQyPEQ0Gqq+4VhIOHsE8
qrvrsP5d3HqT25Tu0GLtnYGCOVdwklAKsA9JHl2VVRFNWt85HFjL3XX2p0gt7IDA
jGLaZK5BZ15cYiWsM7xpoymPzVLfG5zW/42NNLDBZPE31LMPq8T7eeiv+TXPa2AN
AE9d0yqfsmzkJzrPQl9IRS1Etg5OSd302GpFgJQVK3NMt6UW5HTK3XH/2ntyXYGw
kjkm6pzpTOlxjXtioxvYd9qiABOA1aZ5FtiN4TRs4YDY8Du0gXRTSuOjB3j7uEPv
KPf1mDukpEV6XyM0NrQOSj+49SzVog33e/YB23e+OnNHb7YGJJpEfa6PHMbMZd0N
jzGS47fRipUdVUl2TZrbrSv3lOeQx5mxSYjQEL1Jrz7A8DypJjLwJpnVRUmFNpM8
vRk7ZBnHFXfbElL81IIJ5cKhQsLC2KwnG9dD+xVEw8ykjWzQGYHta/JIbl7CJle3
PCCbZS1ow1fL0DEbzgiUQfrsNGzx4h2Xta0ePVdym8o+O+IUsOQ5Qmcy42Gmt0K+
O8Vs4OvZRsBdGHJgZUgvsDIZ1rVlaYy+mTW8ikDyQ+GWs09Zt9IUx/RNBCuKMIQ4
X1T401EzSHaHPeGQmPe8ZzVtaihnX76AqBCFbKzAAMGqc1hdhbDRjwn1EwFbZEHA
0RbTFjkR+DmylLRglMdrASjwmDqJelmrIjMH4HSWiDYUImIeFhbsKYDnIYJ7As+c
l6ROCiwVSXyCjniOnjL30OTjkMXDrYGqdODgddBx+rBGtoj0Vsxv4BrI/2w0JZo4
GPEW8vt503Eb+d1E9iY2aBIX1CWdgtTNATj5WKbhgfxkriMGv72BjNkYRe/i+0xx
nxpoiF1mW1sIIqzpZOrKP9uU0z7jH6uCxiPSOyRobG7LXC+jFmo9XGozQdh8Ypvp
6uBkr/A4WSExbkPe5hu2Rv4HwUXdvWM3+0NKAHg9CW04guUST2TbgSOUIiqnnUkL
JhQaeVmUzRZIemVQcbOIPNq8fz/s/3gDHBbUY65GjL8oUPgibc9dplyoZ6cg/A68
oiw8hJLOPWI4ua/5hp0rNL//rpjUjTLsEGu2xqpbPqm7BS4LB6AqUzP5tynxkEoj
MV9snT26LSHNGMnWXMvacugr/L+/WQPPRbrcAAnoulIpL76r32j/q5AcNkDe8V6i
TmrYFZ1P2iXufDyHqaWukzX9xDLX1ZZwBYyQiKpQ+o6SD5pSE4EtPlaJ5hHXV4ip
TalnW0YoQsZjCjuA/zdF5iJ4AzJw/Kb6eXcnYlxTSBVDHauIbfND5Pm0aKiPp9Sn
BoF7UDkkxmNE+WGVCVnGboRy9m1GjH+UM+5CI6lxi30DHvO1pElOKz617Dgv+xu1
DbB2cWm1eSsM5+ubgMizXlf3+fVXsJrFaBc2U3NG+w+1VwDBCg+qiZEnfElIu9eB
u4EOYWeyPrMUPo6Q6+WuSpZMCOja8cLLPDMaKs+J/3b64oCcMznDE25pciwj+XNN
Hid0bk2yq/JJ6VfSKCQndovOyiJoceuB7eHFEORXN3qdlJIqyj+2e0NwjN4DjId2
KIJR8eEoKHyEvR32+tR6xVPUuZvDdHQwe2BL8TrSSYqBSF9jevgMvfjlTc75lKla
rsohGQ7hatqJJCi0f61Jsk9fGjvPhI8pOrdwXKD39xb2ccw6d/E+4bnWkhGFK1Yl
4wPtRY24WV8yaGE36bIH9bUGygWJRCsdE7Pa+tSfWjTdNJxf1T3xtJh/uUVyeqp/
phyDgdVMS3QvefeI1iMnJ9Hrplcuy8sHorOOgq6UZao87gpbzGQlhPDdIBTUnbX3
iVxjyoowUt5RsIol/0c7nDg7LV2IdVFGCNNuoIjR9t1DflKoT3D+qlPXgJR6FSxW
wHSqC009BGahplEpJ3qoOtzSAmjek7Mw18pG4ZdRXJMMWysTn45W0upILjn72E1e
BSAduxOzftobpOlGyXi/IbUU8Nid9vPDBVaOVn2ae2f3Pre8NRqiQnxSgK1AVWvM
IElW4eB1Zy0YKy/VJW/QzNuc4lEW0YMAIOiAZkMTlWdyy4ND+3q2+cSPENkQnJLz
E2brmFtP+PWanv1WMckauaT/tTZmKY4Crg9aJyxOpe+mbyEjP/2SHSGajCroreEr
rLCkJOVXXZo05jIUNEjcbe/sVyTWVGm6woBjXubWjlF5qaEjajOfPzjfbcDz/c4J
VX17hr0s+SLNXLuDin3grPbSImp0NiVjB7Tcs/vRMoACAyHZBdXCo+IN2Zf1DBT2
OUleiJ8aHjtkpzIlsRN/BSeGUGATEAE+XJ1Nv/H4BIRTIqbClSsVjbtEEDuR5CJe
pHyQHdCBi8uASrcCThmFxeORsB2NpDpcyB4pRz4NM7DZFJIgIfpS5LnI3suLnToe
jaiZ1uSy2Zec+U/eWoRmjY3hrdFbHY/dMrDfR275Lh7ApJ5jZgPWUVmi3FnZfPXs
6kdN2bQPxbNh7ShA7OSGafZ8UzUMLNGVW7UXhBmpvUwGLxhjtIVXhawsNkIOFL5v
bkxS3/B0YVyNuq5TLDw7X7Fw3bpqvZoEOvs3GFUwuwfVWlomn8eAvIIR8aDH6ykH
LDeWK4dRJ7H3SZNjNJlVBXFqFSYbsHpVf/RY6oL/H0vM128yrP7I9vEAxFwfCx64
/Y3qlCqNCWRk+QdhqvPYkaRMDP+WoNG955mcPQ+SJcNhcemm6MHXhhBZV/Z80JB4
7s7s1MKrjzRJVdlOLnPpCYgmt/Ufmu2Bra+kvYBL3D6OlacaPpWpgYLZjaMn9Ya7
f/J7ZtyF2RpyZRaGapCzEuDrrFWvKtvR36l083WvMK614uboAE3P70tIzXyR7pu6
58zLleRDS/iOvrbt4W6nf4KyudW8mbICePRqBloXcxSUp6st3nXJmEupZioEW4DB
nDgUBvQeOJsEeBvI+oDcE7spgVcEAIBWALfJDkMZtw2zWUJ/1UvX5R5hS4mbSrMx
eWzBDwws62gVRNj6I/vECwymRF0vAj+cnqk8rC2mE7W71yJBewjTNI4fMTiOrYZ8
bUc0exHHQGOYPDvioCq11EOGTrzrcMXF9IewhO1Ueq9dSgJTVgN9+3eTZGb1rUED
hR8I6n3mryA4nEwSE9eNauQlZXvxfLtgaZEBl5y7CbzpqNfpiQZv/Xc8vuhI4MbR
zJ3+MOm+yAmbrIXlc1K80eOPvEIMWkFSH119igAenurNcj+xp6ct0bGJwwD0S1gS
p59+WSLSHgriQzpAclCWbhieqfYmNuMxckOaczxgUt0NdR2xFDm152vzkOAexB8w
9cvweP/lVDI87DXEOTewAjtNBXl0wJEy3Q/M9ruFo4m4wqfbjhMbKVNBC1olUT3p
sNMa6wHQ7iJgTq2t2r5hC3yuMjKk4Agu+W6mF8fWUpWFR8FXHh3cYSzwYqMlOpbL
hxgPF/dxcsA04fOyBeNc1lnRe9QnKvc25QE2lxkaUaSABQ18CJCSIMxZqo+V4Udv
i3EmvNqDZry3GmTkXPXuDBHUAvPZpdnpzUVeKMQa9HUsadfDDqkbMizpQq0c6Pyo
1Dt5M/7mvETu28zrvdnmQcoSB7hdpRxlZU1M1fXuTfNQjw/nc/toIzPBUX7jUZgy
dlW7456Tq90Dc8ZqRAACEbBh1QcF3WMDNzJPI/0uZiQJgykR8dyP6xxbzTjAT9ki
jVGpseloEtf6uGjJ2MxALxdNvNW32cZqVmYjJMIzSaKe52YJLdUABxu/fsmztkQp
i95wFC16cGtx75rfKb4macwgfWT8Wg/5YbtMHruU/B1ZnWw6/K3pFuP7ocwFOeqT
fdR4L14JdiM6ryDYEoLOlMj5ZNVpxpbFQVC3htU9yjwPa4xqeERtZSkAvXFJml5t
hqLO3gp08z7qwaI/y0X7qDFr9Axmw6MAiGk6mkJpvsnQZllyT7CkCP6MxYFp0qrG
Rtdk60Ouk7FQsudQA2lirve76UIFLT/zN6mvNVlIqKKAP7/zar2Tr7LrQw/JI6kc
4WsxH4n42lAOm4nflkVCcuSDlXoqu00/NEoK3D1WH83tg3Licm//xAUQjWAzcSNE
e+RQ/wvrfj8CrG/Qs5czSZNuDUKh/vtNbMttcTUkQUCpbOaLAybWl25WygpH0gYj
Rjt9scRAp3E2dX96/KmNwOoygjHTiDxW6eonDez9DKCqzfw2mMAA1qtPTKrX0tY0
KiaTbhG+4AL+ASPQDqaPtmAtWtHc0ZO2/Dwzeeh9/8EQfsCk83Bf+qBjS6rX/3K9
bp7TzDKaclKe/WTdm9G4Sj7fyVbh6K65UPNwlj+zLE5iMq9HkVgzN1RwxgKfncib
A3wME2pDUp0/AXNLwxwZIh55zbnPiNqovgeQnpuRTocMX8TNf6SoiRkzrprTEUIL
mgX0+hqsVSe3qAVkXW2sgY7hQ6pEE/bzdIk0buXyIGa6zFqi1Z3NMM4bO4IGhIPl
CQnZWyW9+MK7OuyNltnGehdgZMVUyOapP64G5ucV3I+Ur5cgFbEpBuWMQNh+AZy6
E10yQbmmcoGPoSGKITmH18raeQZIynaTNInVt18m/4QMMDFqpCCxrPq9tSxIMMkg
lIGr908P1vpefnuoQgYNo21jm/dWVR4UBJ4ZgFUTh53xRe2Tv6Sg7qWeT5qAIi50
1fZBsr8Ms1zMKLkePOC4Vt4xFrY6nvn46GsOWI21KnCv28bCN3A8VN//BZFBax4t
Ue1/w4EiFPmgSCuKLs+/sAtx2xGpHI/GLWRU3VYQXKLug5T4/b3dsR8vBvf2nB7v
anZPOc/0rxnq9Q3/XyhVCQ0AnqmVNY7qZWzVhURNznV9hhNOckJGioXTwJmK2SM5
cVRVxe47WgVFrP4EM6UibZklbxJ9eGr7M7ezi5etHqdGAt+V5dYsfge9eqf2Uwkp
g7tBcCFll/CEv3tR6DSei8oQffCkv+V2HHrWDW7QjsL/sYVeAAuMG+oM8+pEmyvr
B3qKLwO8Gmike74+KjB3tB1i5wIRmoKWzUpfvvtYvBif8eVFgvbl60FEjrnIE1L+
VlW1gaO13A1NbQOmbzlhLEvpDu5PISPmZvQM4YIHiT68jj4NWIotsDfvYLo2pjCJ
jVVmZ+X4/oNurLO0Jqp9sUUyE9z22Yeg0JDLdgW69fryRgobE8PSIxN1TkYfACBb
LiJco0aSdGvy532rhr0cThyrPGRD8n6Osem0GTENwgKgRV5xJjYZpfk9jQUxMOJ8
Ea4IHEKGwG9/iGStO4crkavj2uDY6yacaaE9Ajmh1IJIGG24j/xO6pGTRfrrWWA1
taov6Jd8UUqnkn+CxT56/7jYJUbkQHPVgeM7dykpB+KXZscYVgiu/53zf9/pucXO
UDC2T72HhDh7og5oCZTJLRc0Zz4DlBBODqSqrjqfuceyq8BacRx3QjBx+IgWGPwB
LEdiL9jIvif9WZYkboDLvjohClrU9emwRKF5IabpIxu0c+jndzrhXFASDsDMolSu
TUDgGYRUhZNaXU+NnTCqAJ+7CNNl2pz4H6JbTYZIYTnf7oNPL912POh+Uar70FZD
OGsTYtJ9q5536vvKXtJvpyR201LYpwUaAnqx7QtFLrsEWru5aV6CaSi8eIK/3Mpu
HyJBEubO9RLnLiBoD4GuNw5P3WECdGHAbDTw9LTb5/GtllDTOjDLa/6KOrdhogtk
Lursijqt2Kn47TtfHuQJbVGL5IlG40Y3FQqgoBQoqFcrJQ8yOs46maFKjeagSYeM
qJJEAG4VZogMrkZ9x4+wrUwZZNQrx7GcH8khKePlcdTaZcec9B8musx4EQyfTvqu
F1SsVXeufAQJXesrcdaXs84AA3YYQNEPpWrTbsZrtlfEHgnwFCkbwr3fYgRg6JkW
ogXQh+hvMpqurge9HQ25ry7nRPKrUkEPg3z8aaByGyfBdEma7i0L6dM7GUSqxyU+
+ynPzK+oe9Clb/luJ7IMDxxvhSmNE+Jb/cPIWPj8StP1NKcyTvtxuH3tJYTw8Ac5
MrliVdDb+AByJIHaFG+zG0L/R+cg8XJjPCADF/7Bvdx0Kf6pg2r4kREdq3AcBXNk
j1EXW+ZIg06JuxXd6ZF/V7aghM3V/CsnmPIh1uR4GZzKrcsSJfRREsNpEci/cllR
M6qsi/YrQMmWRvfGKjlDb0ArskqyBeo2VwLEgtZ6p3uaHYnso992zi0KjFuwbZjH
44/HXNpFV4KEIyBuuqzYJaE6xbFDtQnGMi+FSBGjBuY9QDYFuo7G6qXDshxdJOnd
Lc/t+XjOEgr23TJmHfXsaPs/gtCmBGcZ6dPPn5yAvBxIrx3Wb4NEV2S4kJNmZ0Lv
w0w7QEG60tGCw9j4ZOCWqpRQVtoDaeORD1Uhvf2m+I25DCpx+ZSEK85c7sVyHep+
vzkM5gyv/XyXmgC97BuvWW3CwQmnP9+bLZwbi9F7bbucb6Dn06HbRBruk7nQ8+sn
uHq0fGUNwJr3gnrCamYmR+LDZtFz/81a2UTBqh1emhBFEk4xIn2RY5lQwLlP9TnR
Edf/b8gB9cmDonzDxwtRQMTJEFm2mMesv9W9d3JgUuiCWHz40JR1FQn5N9PB4Hqg
yKms/illEVwZMgK2bCgdEbaY188BNoSdUV0ADWBjEfghi/WjxELfG3BI6RMsU9ji
mLDCQsXHiBgZAJw+3CxY2GMJaZf5CEmrc9iBLY7wmZrUFCujFcMoyNmuh9oEhVAv
4p90x4tYPOJv1jPGDh4m4QdbIvHoxJWpz7CF+wsKsTUBZQy+xNdvB2aKC63jPaad
T2FSsr/Gr9QCicmNSxXgpd5M32uebkAWoLv1vh2G83JvFqRKkDPbRm8L/03p+8/B
JRKS+AWpYBP9kNA9Zk7LWeg373zT97VZzMixa0O/zR4RsuWC6gea67pWMIqwoUBB
XqCNCpSepYprdpFTDdMpfaUNj9aDscxeB6vRU3M1bfLDvDymoZRPH8PRQWHwc5ZI
+FAlUy+bUh43lW4RbEzM+6rQsbnq+AodpYvC9xlt/El28E55ADlNp+29oOq4wGYZ
uTVCnUIfwkGCZltuLjGPbIbXokjgNz3EigbzPgJgTY/Ds5TotelZn7cYZYHG3viq
gH+U2GtRLxBFSvHNUpQL0j6+8YRh5XhbMuXk+QRDgieepMH24TCFEm47hyu/gUY5
dXEzxMleUvvzyNPiR6czmN7VGUsgI6kPrIoOtlNIt/lwPrbuyMR2wDLdcgwdepxk
QVqyon8wwKKYZSwrPvra9sAzsX9bjjHTVTOsW5FYvRFnPwG1eLCj4lyUGU2Kdpn6
KQewosB9DzaREpxJRjujNu0XUWylu1smlR2keDv7g0qx22r90hYDqWl1Jmo6V2qr
LE20W5E+4rU5b2aGcm75Jv3fjdcQgRkqw9ibKqYrR7rmeAyU9Q1nXOpoSjKn4ULu
rGKDalaI91TskGIQhBCoMpCPe3tRlkWXgPL0eYPxGdJRQLWMW7x5o7/zPE/hXbw+
f3aoMIzbNDOg98uFYvhrA4YEHndHyMQ+1dfZFaTudqyJoaq3yKc6vkntt4m9tVja
bqxIDDelIuXFRBi9UDH456AoJr1hvtPVmDttfKuNT7cwXKGeqoPVavZVLn58h6FZ
TKx/SHCoz713JJg+k5XKGmCpM8AaZ4DtaRgwzgyeRmZOBml4iRp+oTUCcNdcCz05
ipOdVZbziA/tGfwz48JybnK0W0Gbc/eiOBlKZ2jwrzI1VZhSAUx82VD4njXpIuEb
g4Qvm+qixvnfZll50zgKrsy9+rPfYZM4ZK7desWLHYKo1wLH3FVLYK5zbMZjjhd5
AEa0G5UFMDizlDXCS/ZelORBDTUNgcXpLVxOIWQSu0Vsg03qVLjMlC96a5V838fm
mDR77ivqlpfROBg4vRuVC2jcmD4DiFJBp7AWV4nkxBJMNXaDHmrL/qLmclivZtRZ
79GHnV2SaLGNJV8bpvH6c/6Q4nOAxbAej1PK1rlXJT5CxPCgIGGwbcWPp9K8bED5
gY94oVyAfmTBjVtzDy4Z7HHIHEMOhXeEbYYkLDoR9ZkM0wdhMTKCvEkhIUr2i2ct
BWwOoU/X1pPHxn7J24B7W9lFpRLXTI9Lpd44UbCBOxHruvmuJuKlUM/qHEZU9NTz
1F76/ToMhDVdlyf3cP0WYjz26kL29ewE8/OJt8xuYrK+nM0xkmN1scQ6SPhfhzZ8
MqHoREy50W+I5yoxwoFRhpl+XpTopfZw7S5T4eMKemgcBljzor4MVd8RiHEQLpZe
bsGYvlcK21MqQCUJmvzS2aslcl73F5ViBv4aA5RsODj+BJrtdjHPZBaijgYFWLhK
XLjaqXtqzA/6dNxe5KIU7htb8tnqrkrMxEGhZQHbnZUCxQ0ivMNq6T2On4UnF4Pf
G9BNSQFM8scOyw56TzlZK5LFBUbD7RcKRzaf/SSmE+OZvwjqspwxKmiQh48QAYGB
qKglDzq4b0nqYefUNkEAxwOOlLdaszIvUqctT0wXNEwf4vhxnvaep+ALRzpmQQ1K
S0sgNeL4F1ZAFrOdmStaR9D75uaVm8kQN+YRDAeMRTNLy17X922Tycm3zcfDZnV5
tZWh+Dhik/SGZssjSOMGuIDAQSqlqm2MC1Lx2a77OZvAkT18DqoS17uoiVVAQQio
vrZP3VOuqvvYpSe6OhEoCmRTo3KT6jwSFkpLfKn6Dy3DXDL1GApPnCoVmOdyJQFq
EO4BnkZe8uPs6iches9+QNCmQngHXUlA9TqHBixQv/rcOEn9Rx32z6fAFxKxm0/B
OUJr6jLL82/IPD6v1G+VXJbbEsvfJnDFRkqO+oWW+MRILMKLDA/lOKvqJJ3CFCcI
1v25VDmp0C0IbRSpidO/4agBr5X/vL9MUW+IAzJdTOrawagCuBymX5bpQH6KhK6Y
lZFRoVYdI7CEzdtys3kQGDJFpgPGhWTP154EXn055CzjFa0K2FOJdsj1jT2pll98
tjorzUwiNEq6H/jdB656TzzpOgCnn3pTgyjGXnoxuKB94SxVptdWHzJgB7Jr2mUK
tbwyBSG6pAi+SA7BfhUmuIU5BgTY9fAoqO47+XR3wVh1qKixowkdbafzt789v5//
ReFW8Wp+dNcsCcUOtUAeP91xiX1kKv0U0Hz1sp2Pr/lafwgMld7VoDnDDMU6bBI7
fOH0EITNuKW+7KXASqXzIcWSwhkIQzX2wYUY6JO+xNdBpEp7V/9T0qW6mRDa+L7/
4syV+ibwr5pOoEcSTP/Qf4eCTLCjtT52G8EcAIRR/Xu4WUttJdAzVkRF5QCfLNp3
t69QvCNX5n/iKZKIfHn+CU8lX1yXQ9jNF9u36tcfrVDP4nhOw/gdU6LF0Wh6kTv2
1jJTOVEmQ6LXvspLwadA1BgCN35WAIoh5ncBkEluClctFXd7uQ401R7Z5qFuVlCO
aOqfOszusmhNprg4Ll8x8uvDPII7OynvRhF+AwMeRmjkODck+L5iaKfKeUt1mOo1
UBQIaO8M0k9Yh4X2Q53WbKhvgL6r4H25zm0SnEtQzN6ZAjjoYC2qgEJIGde0IkM7
pY32F2g0YoYCzV+tgBl+bjoM1DbQlZu3sd3Of3NabfQWio60bKblp+fHT3d7ITzc
KP+ezari2e+BfXKv8ApEdFW/Vv6+6TQ0HL+J3hkN6ImPIX6sLQbyTQnUHbVkZqtP
SDMCiDwRUFqualBEo+63fYcPR/sEoRxyv0oTFnjiy5/xYxSO5J510dMlxx/wGHGf
rye5aCJlEkCr5QuobBCAmNmYMhYU01fcAdRf7yQj2gDlfID4Ig7fBLMzlujf+uRC
Gzf4tw3yz3xCDjpWJVAsPMtHF+tjaVq2WA9LQ3YVIkCQ21J6lPYdjFMgGCxxmUXI
OsBK3y28jhvxjH6qnyhztevi9aq6/lkwAa8ZA2kem3RbEQLViUgse7f2pqBOmcLk
PtXJnN2tq7ABa/xeJFtMj6J/gfRnq6mFJgsHLeWpTypLTiz4fN37scj48U/mg6nZ
a9I1cGYeX7j18TZKxZza4JajSrXh5incGexIdCCowjnwbwPG72mKxoj6gN17/cBP
VX3HmKUWbYoyDaWbQUGsl/bcSRMx99IWP+kObg3Ljt22UWWwYHoPh9SUaZ0YofKD
KlYCqsTCnGEh92TqDThu9G9c6FYwpwKgfsANEXuiswjb2kVrR2MO5Rpliu2pVJTI
qnu/2iAQcjhqxXAfc4qpRsct+Jl76plPfzVuZ6gQA+EJsWv+HravmkSOXhboF3EZ
Muu5wlOETpRlGTAGm1wc1AeUZf6BozsqJaGnT5geaFbak0MQ+2onISlMhIWZU+Ua
z8Dh7bGBTyTAjcNIC2hSyVlzttSWHRSEQcqQkgLAHFh9QwDhf78GXohQYTZzPMEI
XhMUgHxT/M0IhBxFusRLfi0XbDhJzf8dt41iNSqkQzFuudN94GcX5xDnusX9IkRq
kZCno+YSDu1tobTyEcJv7NHb29zQCDNyanx255JDWqxG6W2cA4Ea/F063N/i3vcD
KuZVMU4Pt9/USX991xrOCXMVPnOO5M0A0Z7Eg9piXaElPURlY1KaU9Z4yC0jdLaX
j3bJ6PLZPUo5gMujITWK55o5vBjp4S3C186Z/7GVxHky+wOJ6w5Y8RYB3oxW21D5
mxZboDsK4Qe60bPEA9hWkNOD6LhOAicZsOmeqLlC5t0THfOZFg6YwwTthFpUflg7
/fbfx9StX7QS4K7DvTpPHv4SI3+UH5qxbJXNLugI9CMAfKoYtp0DGAc1mLm236zv
cuJlTbNEOHqglYzOCeCst+CtFOtl+HsyvyO2Q4KmlaEQEbjtxKGpHS1xxfBfPwuw
c8LYqyjlSmMI+66ETRxQKwuJbBok0OPUlimQGVvzRY+73sejR7uNjIxPwBwXbTT4
TbZ4/btCmSUwamWC/XxrdxmMsXJw9LenIEwU+8GyPemJXs4SupBiOQLVY9/ky/3A
kpm5RwtYPFoqm8K8corgnBH9fp6RPhWmxns/pT/AtsQIxqG8pBhtNFZkIxdIbzPu
dE0ph8AyfyB6Dh50l3IiiJ3LK4+JsAhogfqiECq+HnsWYvEhCFyU60eetpGnWPY1
D74HQ6ZlHrQi0DVHxPgJgS+ALXLjxOUuQLnG+V/HxDHYQzp0MgJ9xd+P9AzjJnai
v/t6UK9mv78zjQ346/vrdxZJywLgEU9F8WDtKZTaznN34D7ef/IMFMBvmKYO5F9Q
8AFoma/bs61pLLw4lD57XWivftY48KLUG4obrp/Ofm+C65oqB7HoqULSrtlyZlAb
q/c8RIEKs8hrH2V6vA+Z+st+W+xRDTg6tVNoU6pJqz0VX4kkMSXgrSQG3EfmVC2H
kjXf5Xj6pwR0SDokWXz7H6cd8EREypQUQP7NTqv9pQa28pxeOli8gaHM7vOxt7pb
VW8IZ/IV6YkU1zmiQfXLptK33njnZQYtCEXtvh2WA8Adl/UufKJhZv2zHQneuI30
DZcBdw6vtO+alr1P2gkQkGVJ5Pnobpp391bCLcAhWUJOmcKLAi11u3x3fHVAJk7h
4djZKEOxdWUftEaGHlnaC2QDNUDR86QX6Wm1kQdKbWhGHDBAccn8sVc76/B4VL9O
XbO0vgFhRX3kr9w58+IShi5f1UuCAVYCwkppNSqbok+5hxn4iXhFbvFBJtVUGe8H
Nua/4SllPYyCLI10AO081qX0hVtwGborH1QJ4VZbc903JnPBsqudAPNq3Xf5jqAH
Nd4piv+W8qkkwO1SsGhDuE22sqAisCg59OGoY4tlpIrpG2s5q4cSdP36GX7u7EXI
IF643MJOM3vGrClx5Vk4hAzfvsaAiXVZa64y0F0gHQ0jFJ5n+chCweaUNzQgAu5G
vMyrb9IbxdrPSI02WrWWJwI9hAe9j4Xo6JIi1HAs6nkv78X6TvsO2dCsFgH3VZfn
lvT4T37axNaELOCrKwrhCHtRJm62KfbV7LRi9Vq1b2MQrZTZEWIzm+BHDSXq0Qnh
FtiDuliomhqKwU1nAdH8cijAHyIddRN7R3FxK6z+vnzlFTZXwxJwKfj3yS7XR6c/
JNjBgJGA/JlBFfih+0cJr2SHy4hRNH/Zoadej/3JWXHJG4peav+CxOH0aydrg2tP
zR1oJTNqWkiN6LvYrXG3I+Kj2GlqaSUVU+EeOC9yyXh0+2QrytC953FDUVyW+3YF
jGjC71TzDh0rk2VvA86Gd3VsGUc2wk/nqL6ceXOYwoXPi8P7/OJ60s6mCux0Ga8W
K+6FWep30pWk4uzdipPpyYfcbKdcZ2Z4vsQGtCJyG9vxbEAtXaZmhO+RlSEduGpt
2/narS7BXjigeraOZ3446VZRAXLmbm3KsagtgYZHtYu1szAwUYXlyoAxMGE0ftoi
RfHgt8J2MS8uVe2zhVdoS68kgXjp3qG1fzGXATIMtaR3IuqsTIaSGbRI0zgepIij
7unVrWME8/owhnfvN95/s15/Fyp7rRROou0bhwl3rPdFDIkZGz444knCGmgnf+/z
cfE51HCUfTG3OK5eKm3c2I0SWOd7KGKz6ig4BEiGXYaRUcIs3NXIJM2AMuKfSmA4
9abQxb9n+ch5X3arEIoilF6ZuShi0o8Y4ihTOKKZDSXA78W8a4ZQ07Fq4uN5q8A9
iqPl7zvpPuHMqwlGCjIZX9P7145ZzYBHHUUjbdqF7Qm1FdwBgOmu8U5kYZUVJlvk
xOghWgf5pB/swvsrt8fmNQ29xPXnLD7P2MQPPJrHNjURxPs1hMKp1/8Tn3OYQl80
ew7UF55uDWhI/SjrB8lszn4rFwNgCt8hv5i2HYCgCQoYgkunMqdm+slaDXMb/Iu0
SsMZCoqAAn0EVV0NQ3o2gITndEMCh3D2A4tRtqF9+tk87U56StpvkqUapJnlq3CR
PgJ93RidD2kbeM8MQo8eon4Rr+tyRpa9+mHSRGkbtpzz+CfPLxDHm2/PldYm72Bf
9DJLBqWxzrRA/MHKgObRSc5YigWwa6F+9DSffxz9gRd+MkWzpwgfezbVzhSM7iRI
67sXUhmecN6ACjp657XR/edBS8ft8qUI3ewOgTZZhe8SMqQAIfDo7K+L1FGRTUFb
vJwGBnehdyjEOETzGyJBv1zd+JJLH23MrOhfTUzyqwG2ALqaifP/o2kwHo1n3/+2
sCVjCmMJdAfA7EnmP+Z5uNjP9xe9jgQYMGGSsYBuUQuk4/Ylkxl1F5XKy0CjjS0R
SesI/jxMbD6HdOkNrD/N7UbUk5H0pIyYAQy4ApyI/anLVzeNCmHBZAmjqS4wP21l
Bh9LmzncgmSUdtUJ0uqs0bVi2/G+ETAU2WBQrO9qH8H2nFyy2NOXsLpTjxJeKS5b
u717lqnlt9zQHwuqb92IeEh6ZdFF+3X73Xtq7F0zX7WwShT0tX1R8I7Co95c4kJX
IgfkiRZW+RxXnF/rpFrRse4OBEHNJT5g4vuQq03+Nl02RrVCsxy04SQq0VKroo9c
SnL2TFn4F0V+E/4akPokZshSDBdhXaI++L/hCFzPd3RjiLNugJgFZYOTRCbPdRQI
U7qX3eUdyADOeEzAq0XCuJ2+NwQmXUIuRfLN3CgjW5z+REm8Lk3OJFAkIHs/a12o
Huy8hVQ1eMsxbccJuXNVkrWXEHDuYXKhA1bEJVSsmfUWUVYC0AYbWcJf7jegAeuv
eaq5gkGMCpbeCb4Kz+Z47yLhYLBDLpMlOaWwf9b3r4Mfs+g7K0QjP8TciRCWn4Vs
SMGmPz1DwdFFVKjRtjjlMpyUqWpBW8FFt+RWTMBWFslBxY20wKU1YezEEQxoim9c
dqxuhgROo6FWw9QuK2yDmahYw/nZmL9V2ZZQzxujA+lyCWFib6AZtd2vaZs+GEtU
MsW+DVO4T7JuQzGWOXCC/SypV8FSDxavt8kuBVl4qFpln31fSfU4wJodY+bcHNoD
ZGSdKrIjrDNzdsBFZE67xx7YdjVfLFFCU58/XMYtGSpRhkCykLxCFAXl5sqB9x6e
BYWteVrYb+CSh2Of7y93IXkVVi3eqy2f4e9KN3Dqly1Aip3iacnGmepBF5R0kZWW
3K4m6cAGL83x2HHxUk2lZ3hIeYccg18aY1dYCf21Q7ydrlFpwpklHzOQd3NDvgrJ
+uWDWKkkIYQ//HNZC0V4dpDgmcvU09ybwccFIiMqQXhbIjVdhur8PyfDwt/KF4W5
UnVQ/fNy0J+xk+4OQagA2iqSVY7gyEFZntKHf6uTbiKh7+vOSCopbZDnEQGqwiXU
WPzdJ+FHNFjslLP8LgX5AV+5X3M4+YLphE0s/Xq4Ygzd22DMSdycCGD+YL6dHPcm
3I0wS+TAlEr6pamsiYRJAlVIK3pBnbZexwWd53RzCUjwIbZUmaW55c7MYIRa4vK3
v0vDUs68BDfKlut3MCy7lwIZiX+ZLV+QIHsLZGZGBxjk+nkewHb+oC0Ns1Ph5M0t
XCIVzwFBshFa3DC0b3TNI2fUDI03vyiQKRfva8iHWBwy78jQGrtnE0FAsJR0cmb9
d/fqXclS7gxHlDi34+rFAKiBICCiHYKh+A2fj9Xou5ICrVZboUqQWFpQc6fIZ2ki
PCuuazdHEZeYUEnTIBUUGgHTJiMsYGRrUy8ZCSXJM+TanuYbTMcINs1ftNpEFeUs
nm/OPHvZyrqATjpcgkxPLlIceQT4pFJQpjtdg3jaGg6ez4W5GxJgyzQA/mMweXbM
/TtVJYkBLfpabrlA1FxiHYQ4/EUdZfWoFu4mz6EaxfcivhVxrRKsJve6fsk1N+ui
UANLcp96trW/LGCiqlxPicjNGh9UORYQSVB+HYx50wbXq+YtywlTdp/Pb99wMeI6
oeE2YBuvZns/9zHyXEU+8z+kpo6eT7CWVwg9EPH4xVQs2mcuZAmZ8o3hHNedar4J
TRVhg7zTqZsZYObdwVn6/Ka/SpPLe2YD6DNPZl3JX0v1vLiPLUBRvIVYAq/ZpVD5
v5pItP7IgqZWw9mq5kzrG1lYP9CJAu4OiGniULOJectnSuZ2MAVJPQMWBI17lc7K
324smdfoulypDDBwqKRjQ7EP6ZP2NoT5LuY4FxNt5/GRwxger8fEs8/6rek6OEqX
8Lfx66ltAyAI9e7mb7CU/LUSpvuAcXYnQGjQoKQmnLvqfKLANN87jKeJ5FJ/Nv+7
n6RmP0FDKXRWzAJoDZaWWz3RFuv5EakPvQgmIZVPfXrowxMIVfQdP1/RVRAd30Lf
2vdhVCHmMm2m4rm/SM7wX3e5KMB3lygmImNPblN/Rak0N1YPnolRiPvrBuUOBFzr
6d4MWnolo4CaNX3Z+MfalXrMQmlhvBSSGdM4nLylWYtlyIykXzJcMJYjtgvgYekj
/+0NtBW6xDKMp6Fi7/QLon1bCfvncGeR5ahkEIXr4c+YAw79JADQ/L1i/wZ41y4W
RKqf+P28TbVfmFfGDvBOXjrSebjf1Y82XwS4ev8ju8dIdT6ZWS4z8WcypowgviET
UwlaOADF3nyH3tRxc1aLdAf1XUlzvPfksDVYJC9LyUUK6RIMKjHQGe6rmMPW0igZ
b/qKpXm2UsQGSOChvuEoNtGZPD5nG8/l097GLwgLsosqzCivNBDeJH1VoCoh9CgG
K0v+54FEgThlFO4OJhvDfAEgD7GRr/G5BpoFhV79ipQ6ITNnFiPTOwX8CrOuDnnO
cmRVEi49J68mwUcVc9oFz/DouzajhMc7GR01aoih3l2KwHzN7SFBGOg/nSFwC7P1
2ASoaR84xPEttWTIq48IUmwxjUlz6GTK1rHGAkoA2EegLZJ7YzXH80jnGPwL2AeO
ag7jErss1wtlv+cgos3H73bC3/9H6/AqlU5fnKMEV1F5LTxsW6HDlZor8mgLThtl
v8NnPPKV5jqLV13i7hxpabMQkKFULsOii7Z23PPNjSDFMCH93KV8/caxhH+Tv7Ae
t0C8iVS9MsCgAU9iONMfuBsTVabnSk6o6386vV3ZH96p6ttxIfvq9JZtX4nWuKoc
RhB1FEVBv4LIbfP1OrG5842a4XziJ11pPPmBA5PRXA/lfVYFJyORDDV8qOk/GflX
qYy4zSK5DcULUFXtVi+ZJuU3Wb6NYUCdVZpX99mIMHiF5a6qIFR1M4y+OJnM+NY6
8Pc/RrL7ZxQ6rJCv50kCAS2FV4G7qv+k7pvXpck+98XlxZ9PpLLoZGlGQQ9cDi7G
cXNpZ1N/ur72kwTkaQFzeQaXatIwtQbdcTaapYMNjvopnLQPTP7aWs9Oo1bWbE4N
uUcrwx6ZMKNgJqAqOLl8nhqFT/TEOP4ityyuvAjmS0hjBUcQI4RqjRf8AL5fK58q
vDqE2h3CY2qoqDBK5INxskbZW3togMgAizUROXtCnGuhV8Gg1t1rcf11b9XFOLmF
Ej5DATU5IP+yivvoyCn65MLd5FzQGrqo7LkbIPJLKI+HWjOdMiMcB3LVPcd9A8Bq
DPRZ5bYDdW357T8aPgc+ypsDoQwt1mE33EUqS59ihTyIVx1t+10v9nLmAmdZb943
LhRHGK1zsJwQWhad/KPUB9tw/vuUtOq8xixZtQb4GlZ7avoFMjYD9HGRr3uGaipi
M0uU4K1pSKUkHsXx00+iqaCA79oQboB6K01zk6eTMuoE//PyI4djs3UM+jkTUEuJ
5zHgMAJAywNUTXgjqhT+DLMHYI00g3pOJapzM5CMyehRpaYkRH1spwzgB0lTRpEG
JwT7MF7gckLvTA27AG3U8fHB1/0QqcKhmH7v/AF2fl8o274MjVBBUSfXnlYadOuU
27cWlLNtUda6YXsA4GdxCsRdSfgcBTXtYMULYdryKudc836pEvlZo0ww8qsYWGEy
W6zmfoA4yzd01gpvDW8ve45+Vu7f2Z5kUmf8hOvxDU8wYM7JxNPOBWDJlOuIND7Y
i0lqKbJGYzuncjzsrkHYt8tK3fIbEIGxzxtG/Fn3iZv5jZr8DtTZZ0npKTp/rK22
eyr/DPpuLI5Uz5x5GsyA4G0BUjo4wajmQliBXt1FtXKivQnu/EpFYWMe4qwR1Jt9
J0G2gcqv2uirXpteW6keJQfoNA3W6zxlwCpQzSH42DIKSKPtSHMAdZD/U6Z5WMsM
IqRdlT6OujSg+pQQX9WLaqqwy7pUECHyyrIGCt4bPv9/5H5cZxqsec5qQOO4Teqi
CpO+JbIXa4ndjUSx9kFVyR9CuV50VdIFH32kSNNFKuKXTZLtL8nbofEzBQCDfLFq
qcUKuhsCL6gWTkcudajBsVEv2Ppwhpgphbcbkhj2JSUJcmR7SXUZeZGk5mbvwQG/
hx5A4ffpU78ZWMeotWhgIDqtXZz7fVoJS7OY6jrE6ICP41yyG+qWtsGQkbJHV7Ax
CodhaUBmLIf71yMPtItBhDn9/VdDsxhaiggc/+IV43j0Ue9/V+Ejc7Oh7ucJ4mXh
EcAzaKQjggNJ2nNsK7P1QZezEmDSyOyM/n8fPm4ih3scmv7dvSeG6QCqjjoHdVUB
krPK+W6ZtJtShN8qNWB2Jm2n9MPQfU6J1ucmFaqRZfSZ5G1uADtxZlAOkZ2erpIm
FEUF0FE7Qa9AyoO8MR1mPer9OdEdE5FkbLiliaXOdS9G9RuEOntV/fYe/2l+72bw
HCssWixNG45hdAjvPWnmK6TqyoigKiQi1I6ND54a+2A8FF7qozUCshFA7RU8eeQV
e7mQld7Kd6bY8qXlJHxvV2/5/f4RA1TPXWYWoarc6NA+fFKQOwkgPNLJb1+H4L0M
ao1gqES7QfdwxACTxEcAV11M9rt3yD/O/ofDG6i5k4kV87mKXrZcyR1dcj3L3h+u
ugnm7XwBNbbf57rXSr7oBJsrsT4Amcr7Z44elEa+a61cuRhW5zjhmhas1uTPWXNm
K25AwR2Y5NhLYgmQA4UnCNEejH5yuMnrJOFkVAOtYwQVD98X6/3CxOkeQmojRirC
dOp8esstFKi9k5y1mr2PtoP7CS0/dZQQQAhIHhU7x07y35rqFn8uvKFZECoa0Hdn
/nFjwxTnrwUgarAkRz1XZBGB+ipK0uoU16GCiHb/UGQd4x2J1j5dKrCJX/X44vgU
mlfkjuxGz4+8by0xhDN8SeAAEfD3ak8L1eaajWSE6FESDXo9wcNwawAhlTkaCN7s
tj+Z46XHNC041DP/bmBwqdff/OT3hwdKP/w5j33AfzOf7hdhNreFo9UxxQi8aLkC
uBEXzCBFbBXNZK0tE/hKTKgOs0hWtdQQwvLnjTEHIpsIo0CD4vbExmSOtd4Tdh5e
+QK6HMdTEwtCe8BsptYtn+vtOO3Uxw4uvmDWq7GKS0M3+pvsbM52uF9RlYg3hsrZ
G93sOkzeL20km3huSmFUdTMoKj8DJ9Wr8wv/NB5rQY2ubHyDT7PnsjqHhdMYQWFR
Ja36F4ruwDfGXpwayLN6ilZd9hXuy8Mzs28eSSupIJRP9EGbDpjiAQOMBkahYYfB
iB6M5CcB6e2tA8xqFTaa6v2AzHjdPl/D5Qgs5HF45ND4L7eae4MJBRiSmwAEtNVP
AdDavMo94iz3KFlnl3LK72MZb5BzgEGwOSpjf0BDktimOlCor+mb04G95+8UGFO6
Il4x6UNr7JsJ/C5gKd/deFvIid0X/hyAsR6zRgc7oP9fLrEmi+Kzmn8Jxftz+fwV
fkiIq/NuJkk4dTsDtKeutVq/p7JZjDvfKaQYELiJlYl8wIWLvhJvv+RcYRiUHC49
7L11RW56d7XxqIgKaArdSO+SlsaWo8ii+KWb14tUHm2HWqKCXT8ORVYJxbD5deaw
1Q7wFjoPeIXZUmHPdQWNwgUcZsAvgO1frXJXncBEEir87k0ZCM8dibIb0dzfGo4/
v/4GX+jcK060ymHmmgDVq5nbmZ/oRAZFRfMbPqexYHCv1GfLZk0n1QLkVyfJJgFF
jT9JjwSn6ab1XgpuQUjG8redh93dIiDGWnqEwJ07uA9nTmfT8fp/2GTCxkkOY4fO
x9Q6clb5Wu8lKmLXH+klUaP4rICPz7QT+jlJVFq3srRTt6zAFDFYrXOpM8VFqGBP
2hhCTtOyKCCLjTdbIO51z+ooXQjNeCmbmujis4Fra0Wi0XMOWTVCi78d20D9UWOv
Oxqj+Vx+pN+4abGBV+qB77bBxZ5dKSKFwmFBxcx20SZlYDg3oOsjmRriS8yD2q8Y
IQKkLm//fOzybU9LwG3xXZQvybBKOzWvND21RDucL9DcsLykvvlRw0H59PxYNyN8
psjwbccrC0X/G6Do/llLiPU7qp7wbIvBqgwaVvZY/Pmfa/Vi2Jy/Ort9eXWfgrvH
0VuNB2NjTylogBwqFZOYsovSQ2U1KKLSocvrK1nkYqndytpsvrNNO5gQpwCxu63r
T0LrNOQatfESbGcVqPj63S7/fBno8uRnMXmsrVFXu/X20VrsILIMB/829e9LDwwq
L7wvgCMzE2G5FnuRrxGLBfTQPRITGTR/fDq97qD5o2j8IYiWmHpRVEbQs5IzfrBb
L2f2RGC+YdQGNmOHzZxoTzE/iAzeQfYeFScuqdHvIFrlTLKv4vh2+xPmcVdMEFXf
0i4AK7RWUZK+XMSPRyLKK2bV1ljkpoD7/YAZGTqAvjnutFQsCRL+AFXBvNr3xHHU
Ey+XwzFyycD6ILu4S7wWsdRuL+WKoFQWgSwOuZY+kZ592u9AdQXt7qcLujFZtZz4
iwpDuBmb0IRACV3adY2q9fQyGcsrgY8R4lxmklQpT2X6x7rNjWOe55r/DUiSSve1
RIBx+yUOb4ibiuN8mdy7ekmpMNiHHSsCoD6Ng1p5qTdW3EuQf+yZj6MEKZkqplVW
WD73Cx6Jkiw2wtva7SdZvP6WUF9iYs5xlVVw0kja4SvoYG6BWakOHwsALsyOErC/
4jJYbmX9rL/rKEgdwGdP34Flk9O1mLks5Vb3F5p8g78P3z/Di8Fx+QJP4ov5JVc+
xph/GrxQLQa0mNNNllCw+G/Nf9W3UuU9uD6jZAQuBEEgYzycqZqqNGCFJBaTLDOV
vMwE+7AEr3iRLvBWyh/jVE/A9U52Yj4VGEZd5pS6J7VNmWddLr9P7jap4R9nXy28
IFGiRpEKdeWSe259yKkhu4dY3Y8K98NnJtqcA8DLA5BX7B86U/JMzzT8pfJ59h0N
ZXU8Sabl05ZHBabhMDBW0FNUeOEl7Pw6imky4fFBhpHOuGP+RDFU5+tuzS+N2RH3
lpjJo3wY6lzNZy94SGhH9ysWrnqbY5i/qQZmHjF/F+ZwoVkcs8t84RSXJyAtDza7
rnCzhhj9KOaovqq2ZkxqLP15w2rJasDwX6xihlzJf0jz+6WlloYIe8DIiJnpkW+G
RxfukO338xlLiWlNhB5+8AObyRx50alZ58vaLVmRAkxWlPyB03seeGSlz+EtN/ae
1EaeP77qTkFRPolXDf3gdnniAz8YbuPt/hr7zPI6l12XNdY1DzXvGecgY5haENwe
dCrNIQ8KutKFlrfyJdzNygT5E6zlOUIRk0j2RQZ3/Tlsb9qw5J/NFFgdWKKVF1mU
wDj0eFrYsHiwgZYr2cDdmr4d4tWVAPhwGDnjOftNjyeKUc6lenOrqnA9Mn/oWHkK
szIbEkjaPeWFHxX+X3koTbJh6QNY9B0cZ3978tGH7s/R5Lm8tLBdUTPfJ9NmfHX0
lNehFuC05KmS1oeOR8eKqcUMBLLpwxhBtifznfisW3uEZSi5snqi5bqrTnEQpbBV
0bvt13BlHK816X2NkQzLiXD2SWIo038spgHFEzw774iMhyhe4UM3e9U+nTzw9sBt
e2hYAi0JWpMAD/mewds/I2pjgoEBTanXTZId9bIaIwN9DMKeNpGEwhDWMcVuwriG
zHsKhofjh9hPsRvEG6iUBoEGtZR8KCLzmHIk8sNB3imuTNMR+MfgB/wLCrF0sBgU
JVuPeN7RxKdVMdYJcw46uSinciIwH+AhKaFx5xuPTICbQLPe6hYvQofhGcZ51OEp
EPwcEsjhi0+HMt38oEylz0ohLEJ7mHbNwF7lXDKPZaTDKi9tu+lnSweYdVmna/n2
5LG6r9lzUn5wdt9pu4+KpY4O+NcLA7IwLZE6YOWdsToe2UK2mnDUU/edvoAZucl+
WnAf4MyDQ2VDFfs8SVQQ9kqcmFZZiz96X6uY+FeLxXWEzD8lSfaLbVapfmcFrfqj
+UL11SRnMXdoc9pPgmIULbaoyw5r4Q4ADyUE3q2XfxaDX9uKKDg5xzQrQikzcw1H
1WqzexvdQt41WBl/05kuJpeQniVTjtjYR+qu1K1YyZ3ccedDnvI5qBQJXGUqEeEr
4nTlUE6vcjLLzOaGInv7Mm3q0CczGKotSCEarh0SsHac5/18gRpzzNakXg4RtZ29
VHMKrk1QVDwT75Q/0DMRH0IR/HSfEUl7F89jJvJvbamXfKM6kJ65qZs2jUAG5bqP
Q8LGlR7l+dgRBEU5hfoCFCcRSEvqjYR69C650WTN2CkHmUrt+JZ8nRbOtU0JiOUQ
BqAsYUuxF8oNxbwE2bJWQwnRiCfAsAp2byVXXHE7iPc/izddRUBGZ81uDXkSAfJi
F2sylsZuefLMSpJOd3w3PvwJsPted6bR9bGRftoSx7y74s+X1K7OIUrXSr38p93B
Jj3t/wUNBKuefBhTAO2jZGTPKavlJW2ZMIcIAXIdgZ07fUUp5Oi+vnN36HCIuVIf
vjHENUXVV4GroswqjYfgK90ly64/Sj8VwdDF4/p7gbCyhWzbnetGuecl3d1K2FDI
5KrBNf8/ScbUyD5RkFywrCyN02uCRwfH4Vh47mD5btOmIQRs8azsPaNafK0ed10A
zswJVH6Cs3wQdW39Q/68zRSzv7HxAMeXygbLa4tyRI7H1TDGDHlOugsBqiJgr1OV
wzZUodJlakj6TvMN6/aYdTLSS3j+MQiY9jAulipYNDf3udbFl3i9OdtP/LJMCFPt
S5ERhWqC2QVqL70ACt2YpYMP37OI4KwqJ92hvsx+h+cxYNzNgExkyT//7LZJ2DSN
wb6PF6ILI2YE+8QybXr0+YZUsezCCfs0BsLQCDGFsZo6VC8OlU6A8JVqJx/Fsb4r
ZTaGvHH1NuvMexyrKS5xuJDqqBYN37+fd+1ig7vunt/zg2jieH43+7QHsKye6xIP
x7YxM63Pt/0RzWolIKeqXU/pkV3YiLne0L64QdJn0LMC9PKr7AFbeoTYOyx3PJ+8
FEKF+siU8xB5ZjHsjUkgywhnbJbmCgPFXqcwJZFxfNG1mY7bkqSi0NlD/AUbXBWn
CMCq5ddEvo6tltn2dGHbijarkm8dvJvPX4bDsYto99/uFYPUNpeucHpARsRd8kbl
IqgA9wAabai/jkP7A7rxQ9eZnLG1VvTHB/ipNVhDPBf/Eu0jEzTKsbL6vI3ZOTXq
D77dHt8kxx1SIJsznDex/lSM0JY3oH84dqQOlIu3MwOWxRMtyIOxsLHcYZCKJWDj
fbIidJNG8/DkacleEnjowZfzm41M/Lc++sbUCR5jVeGdkjM77QIRnSgZ2lugx8vs
J1p+Mbx4j8KeE21UI+TtNvnyWxDH83MMkJHaQK2Z04V09NyKsCDS9/a4OAw7/4XV
ADTxBUCFGGyCbc5amLA877fg1fTT2hEeEZe7qq93gnTbpPWYJjucMhf8sEhktVDT
db5LHdJJUG3ovNFAKP1aXmnYUUnN0TNdgr/xMFCjJa7kJ611WXXZFmhAH06DUBqt
8J7/z9oKMTn2qTqjeJfbd2q4HgCU4hz0VGFyGz34RGjwtMFAaA5tcY15xtC968Kt
sHrbQroJIPLcJSv76oA/qIDd4HfuSt6EyBHRI4Z70KwtxfvtjRm7YJFTUcl7GMnq
y8JgywJPoPNmBoFKCy9BITRE/BoIOaazFD7/ub8MvU1f/2qL+gcBSe8NFyu2DBGJ
nYV8ED6nYG1GXmsg0bTsvYrf2P8Gk8KDGnOxpLjkcX92POntz81S3eYRWL3cz4/r
qLi0pVF/nvJI2jjOihmYgf7b5qtN/dIk7ogsdUR1xEXJLAaov4P6b1IzQXEhywjC
0yLkrgoo1OCz3Lo79+v9e7BPbbEfvp2kN2ew4Gu0OSqwe+sr8LeDegjsXigxXZ4Z
ZO/MrUGO2XUAt0B1uVCyzmh2VLOpiNWZLa5/jmvZ9/nbPiZ91g8mdT5FAV/kiL75
lVJdgvlbRdvDx3sQvooYlj7mRnkds1XiB9dL+Z1NdQ9ZwS4tZJOhh/3wGNd8WWAm
Y7u6Ai1Scujpc17FmRYxbnp2dPTEMQcy3E0vK0a7fUvDb/2NXd7yBHEytoQ6MBRV
Rw5Mt5kOq3U2r7NDxERI5ahCGga77xVFilKVDlw2y6RGMSXMRTCMlQbv/vlK4sPV
sjVzYZVe95mSsk9QwUrdLeZ6sIwW5jxkZ11bXsw7KqAQxxe+QNRPSz0mQndXwZ1x
X9mm9pHG6STIGagYwbv4dwa7Ogr1lOzuu//NiLOG9cUxoB4/GWStDrRKqGs3NEOF
K+7lw5fPnDsFfei3s1Q5WRJQlluKqJPAdXHLEF+ForCuPLfwV4kzg39ayOeUwftZ
wkEY+UhjZyRQV6uvHbZzdIKYoVr/UlJ9CkrJhdLMRe7TkwngtOW3WAGruWzJPHPL
vjQLfCS+kUpEPb1ZhFYIUCfAdJ9W8wJ3tgQrJitoyMT7fC5bk9tdSY1QSncP8y6y
VqYGmVoCiooY5NW0s+E3oI7UJes0ivFH6vaBRmQ7dQ5FGRsIYhZqNT2ZtTm4rbnX
D0u+08WH+Vp10NtzvmFDsv741YN+sGMZ+typ5ISQbi2qZ+EmxKxJWAP+LJFlPC0z
9JH59L4pyxrTQRfiXSogDAyh83ixVyI1XPiTR6SGdRHTxA23XrUkejwkWH12P5hF
4nJgWQDoXkUL/sGQGQT4vWSTK89FD6TNa8NscSagIYRdz3O8b9SOgSBn2oqMFom+
uhwyC22Xffz58dlnN3CyNO2FnR6S96uA1v7ra6KM2OAxIbdeI6Rg1c3QRgu7qY+N
CCHe2IcFzuT2QQ2enLazW2hS8bCUn9v+PsWNTXFz8H/OsCnCGgXnXBVNOD2htYVV
iMHk+9srmYWAlvUwozcnErbfmLQVG9iOqDVHtL7/EEqkFTEcdTF88iiqyITbSe6n
2BXkw4oiHsYr42fmoH1OGaS4Kfux5ZpuQjU0FNMAI+emEGW37GMM3uJo7mAQQCtp
tRxlmJgy2Xd/VLZiYzLzLgrOne9p8xerltBKvTmlreRZAhgmqncErljbBIJ+OUC6
sl47yHfAYm1285vFJYBtMA/a0SmyrYAAkCYlXXlcvg3px3lW1kxGuQjQU10wDJp1
lUArtAkC+46Y/Ab6pVodflhz8DqNRfu7BGZKkIPJyud2Wu2ptgp8KpxacfxQyn5w
wnglHvtHmEJLHDoAabkcwOdgYeSCTIHpViZkEUev9wKrkfCMSayKvI+idGYEYZom
UNAniixD+HXq2g1IyM4yRPojW2lnyrIitL+R2nXyY2hkliHRkd4ybNJQXs7+ldXh
6uJBhrfjA1bBvs0++EFcKfzkvE1dCYfWpI6udyrqH1iqcWvd0hXmYnPgdhtY+F/6
V+/z0vmbxalH1r3p2FyiBeAdU0va3lldLkM/75BypDk2LaoRQ8ZxOSUE7vfbd4/n
qi3eTUyNOKxRcmKNor6dKT62135lXlIpPTIl83qQP7LW89T4NhLGGz9o0UcJCGe/
Wg99eSfQtHFzhg5oWLjRVQVchgD7r26VNHvhoa9oyuK9tDOfVfR2CRkQX2oTdizY
jqiSjDWeQz9WigyKDzkwkIp7XNrLajAKri+SQ+SUPTKxiEyHrUIXXz2P74nNOn2T
FvMnAk+182Xrpm0UPmC8sO0pwJvcU72ri5nIb/YYgyK/74J9Yjw5SdPog3q9pzuW
UvNpOGlsdC2zOx3hla/q4v6Fn3cPzHkn/EVAJvkhVPVOVwJhidftGoHkvvKNCjkf
0R8uP5UUKaNZzjh0fZmW0jxKR4thsvCuQXFVhGlAPG5rStHl//idEhcCBfFUAKys
y1EA52qtdP66V1QoS+XOTfgBg0nh6heKc7FJay7qwcSABR1cDu+DhqfBtaskFGr1
1UTT91ThdWvenKlxxUVt0LDSxJAtCkuhBgY7o6L7cxgk0tnbgGHwnYfkGiIopvQA
hVxIjq/1Q9AEtVz3USdrzK8ooz5LcryKlzLHI9J1OgMPbyMqpF+RFT4HOrAwOsia
5Ceiwc1ndhrC/NcX0oq7nlmQoqfdOOHXHOMlDDvtTcS7f1xngVhjlhx12KhK+FNV
Vfo5wNw1DQXmpdWTNg+VRrO6F14RZir3khA6WvuUbxZ1XrUzb7jSZzbXv0f6pffx
qPPGfh2EOBsl2EDzB1TVSMgAKOPUlrN3RulpDByp9Z0a3g3slvgXRqE599R+sFl+
AU//S4Eu67w6leOgVtEp6mkxmVUhKTJ2F+VlWdkQkgtx2PoEa3VVHMjJ86Ud2Xt+
Voy0nqyHwjCzfCUHd/GpH+s0XIMWTmoKRQG5rezZsKq7gh2UMzNXSARVEaJamUS3
qzP13GciVyge7SQzgjNjj1kA0z9Yo9B1UeGF5v1i+DqKWIeuIR0xy1oMMy5xg1w0
9784Ium2CcQqVkgekSFX7+Go8iL5dMZ3/RBh+/TNzk/Z01jmGUKKkIiYOvjCpaZR
Dps6u1jq/2HumHpVO+OwGxnDlsQbgHPNz5vHUeMx0C+J/lTDNnu45r/jrt2jz5jC
i7+KFhsbvxkB2KyiY3kO6Y8i+VMCnVvUCsCLLd+kjr7qj+SfybWuA7hJLKdNt4rl
eZBMIerc2x8BDz6bgB2C08xwG5vOR4voIW2dIwXlicwDL17KMGRbSVc2vK2AIF5l
phCaXIG8J88fS4CjHcws95XtsuI/uqOenxH2sj3A1MlvsGVZOo/nddHGQWpj711X
e7oS96pEsqCTBkNtgH0a+/pKJVAr9hASZD+LGiqqA4hN/hYm00FTutx+AZ7cqsG5
j3gDyiH5PLYTOqpWUXqe+tTxwPxzP805QWh1CINIYgQ4+Vd/WyRiZFElTMPaTnTI
sdQWFJ+UnHwrKXaFSI+2u+G+PdKUpyf/1894Zk277vjdPRx+XQ3qPG0Ws9njXBj1
GQSqjIjhoaTb2lji0C7gF4A3jb6GTHeTUpBLEj8JPqwFkv/SnMC43PHBSXcoMFkq
AKIDVx3lNDqrX648yUCuLmBdneWZaYM2ucRW+ieJFEsrCl3LTqAMBV6ft0H0cj7t
WY7ED2Zg2V4kScKH0G6i6+RzjyiX0clZIa08TVL8UT2aN/SiEh8QsSD1pXswUv0W
GdKAAJTSQ+xTZUtNTyD6YA/Hh5kHqGIqTyoPTk+evA9NUYrM58ljc4+iHWaPmVQ4
Ia7fNKjRtkvxvZcKc+b+PxIAV9rDc+3pM9D0CibF2coGfw/FvhM+bpLhPmnVwHNn
d+HHO501SRQbxJ5/445wWH3OIWNgTfxAUCR1zY35p6jzsi4AvXSxHAeq6fhfVZwe
u30mNrNocR+tEezoTeBXNA+1ChPzC16ZFwlSMwqlLOsexrHCpxNtt5b2jEkinmKq
z9y+6DRl7vmItt1gZLgPBC6M2bzYUQi4cea6VO0DqIT39l9/B+Su4vWV59junrMq
5dtCo2nyAAqdScXNxPBUOmup37VCzsz8QMJedKfnzQh5IlwgktotUkrbq6noEgxZ
fC2B82YZB8GKadKP4C/2TszpO75ciVw0Y2XeZcYClc9LGezf/frkZxXameFTTsab
pAGlD14QxRxkrOgGmxilMp5m38FezCaifwY00hzaYKo9iJYcSKEaEHugy3hg/MnF
8zFFDO/qFg4fuQjsPX+2xi4txpYBovQc4ERqqCC3cCHXlqQteXCXwMIWdA7NqKMl
HagNf7Iw7Sv/txksWetUSIoom+9002xaAHiBw+rpE8bQHH40qoRQND8WEVafdB3d
QXILZGyhMo6W/AtbZ9jZxhSMrX/8wioMtXpW4BYcuVNVLYLmeVzG9glxTFusi9Ou
QQQXvFVgNRxi6khBL3x7XYtpnrPnX5ERnT5Myo3MIqEBwK5yOyj3vcVngGOWTNUR
xFHX5UEQBC+mERBy5XceDDWyyGFgnkbIUrhG6XL0uCEaUTcwKszJlu3i8O69cSNg
H0XMxCPnOV7mmwkBZsJBqr4G2FHVzpyNnkyv7jEyTnYTlFVykB/dsM68mKfxsNHF
8H/K2UGFTJ0ZiKX9wIfEyU5jxkU/btUL+qYloHzM63lkAUgFPZGQlz32OKspIxYE
lfVRTv2uxuhUnT6GSMtZBK9kUCVMXReb90OREwJsSD0ZOIfbVRBKGgHu3ZnFqVM/
hAdlJkK/2wDKdKz+hILxGGiaI3OVoe3WqG7qCjoTBdX90O1trCL7nT73+aEhZswV
sYotBB1NYNEp+ifdYi+iiXzGFJSn+so+3N49aYzfu5opSFzlejiTgrDGiXb4x/St
jn8j7ZpNRKh5Cu0+A6RK5ftcrcLD/NL2/GiIvE4I0z3wrn6Z7SOgkMd8Ts4VmCn+
yl16KdSQHgXsYP47mBbyzXu6Z5K4X1GjJf9lC2+i41TF3fJ4gNRzKKqjFlOKKW3V
OVKA0hGyGIm9Eh1nt3lNhBGDG6Cf4xfNS2vmw8xHQz8nYx+8rkyxCFrqcxLb9fl0
dBbjBfiodwK5mG2e9AIe6SM69V5isVv6/JmENBwhgR6drQAc5UFn7bWYju8PaW2c
HcUuL2MX54+sprlwTiyteLbufAYkKVq7ioH/6kdkFZ3oMIZQ3gqKOlgVwIQ1fWq3
DN8iizHgwyScQXRBe614EdLNlClhNDugZRA8fIIwItQqd5biRbV1c+99wB7u0hUM
ZUGqhezt8bXgAgtFqaNq8khp//cNHRiAJgW5hiGTivDBflWmTZB+JRA3FaDBNBvO
MO1CFZ0eTzpjX8qfAcRYRbK9vATqn4XbHhqXhBVDzVw6WoUJ7gEXlDSjuO5ENMCr
IUvk0cvsTjfCbp0OAwcNjmtRPVyyWF9Pwd358casVHbcBK+YPbKQlHHd3VE2Salz
DLwKBaffAbDsdOTxxLq7vV2PARkQSmXxwYzboLnzlUdasFj3P8RQWBk748md/0iO
bVvGqJMWl1BYcZi1HvLTn5yS3UMEFDFUSZQeS0/J9v3O7irwuAAf/wBL9EU1IQed
JQzRjiV1L0ksl17KX4ZMfml511JrORgdVqU4FkzyL4+a5u4e7z+igofwh/5rxxIq
zDhTXYGBOwRCd5m1ca0iGETjDLCRvJTJ202NxyGvqJEi+wZE7cpluZii+CNkZQnF
TjuVQRLGSzb0r35oJPoK+GMLRYzNQn9JqDBvNPU6yPKOMGGKMITuuppX7PIiT9/j
envCk9ivDmIWuxE1gPe54haOwDRiWpOnQRKKJrvV9h3NTG3d8tLz39JvNz1LjIvx
Zn3S1/s1TI2oTZB7qKHptFTrgzmxrvx2OTL+4MGmGj0QccOfWJjvFPmMxwMXD5RS
XVsAS4jrm7UOBaB7QYnatsCE0S5H2MDuaVHVR3ARQfzQix1ORfGClh3MBVWaIW83
p7uHrOxDTb38vLSqHaZh67zj9kJ7QTSbBFPqN1szzux+Iq+dwDoxx45bgl07gV9o
DTHV2GtEofgSCj9/dRYNBLZUttUssDqHdK5v89kZUGPQKI0gYQou3b9UDc2PFRft
AL5tVfVlkaoB9xgbiX3sh6mHekBNpW2feGV6QP2nrIJ61ZE7AN/YFpCrOFeba4jf
FA1HFtsujjKy//K/opRA6qQAC52dAMujEt8MkfpfaiHolK3vBT+QBfeiVPDp+6fC
lPzA9TVTvY90LTXiuwe4Ug2aAO5MS8/SZ5DAyYtDSesVLdcMwCrlauexd0nFbDD8
CteaDZw3F8ycoFPtiLnHnrW/wlpdesSBqbyhN0bq0LN/hbAywxKJpGAv+dVLOjlJ
2MB8cpO31C0XU/Wiq8RdeY4ql091oHwkKlgmExft3rXEw/Q1lWz88WkCpfcNMc/1
sa2HSTCtcDh+cnSxUm91OjCa/00aT5bb7vTEjXGhTQCAoR810kuoLbPlarLefafY
G4plbr+5Or76b2MKsr6oktfRZdpG1cm7Um3bnD1hewg8zHDM49rdINccEdkPNX83
8QvN5iaBgRcEduPlOObnDGhR01TFjeMZVvJa2nTrsGvK3TTAjyDYK6FlxzShAIOB
ZQ5GCR96HCULI//0u0dd6Z2NyMnCOcTaIiwn9zBQrm56uZMJjQAaGz6PZ0eTxZbj
k2rjResjU+TwIsk6JxBZtfKYVl5tFqGJ4D0mpWd/u72QJUnntSXncPGf0o/CHTRI
Z+Se/L8dnG9DD7rO3oIR2JGrSGLajaNde38hS5iORcDDY2mE+BEA5j0wIWd2sz80
nXPt/2KkRcGfk7VDQg5Q77MjOyuL6Aw1+bbMvs9zcrp7LldPJCIWuzxEhwCzAGga
9Jk0Xo7AyYMo8pPzcZygUH3t8CFKsqjXpvFTXDuRb8YEk5cy+eZb4GdYryvdM651
PsybGRTeETW+1nAN4wDcY/B3MBSthCWO8Ns1MJhsPbCJsWR5JUPi12GL6roXzu1U
oX6N/0Ws2kM25FkoH1Aew4j5nly/k8R2zTrQhZJXvuvUJt19nXb3K6uNB/Gs011O
hGI+JR4qvaG4FCyDKNRAeaKERc7/NXH/Dk4SQG99XCeWgZySLlgbbHKF1Y8IB7hs
G/bRyB9s5g322Z5jyih18SRa1YDB8p5wnVEGLgpQc+ysGGZ73auq8k5/fVmkN5ev
Nqy1QXhXVic/JNjoI/iJphOVzjLss09C5Yt6n+DT3kev+3ZOC1VdzGCHyswgXW38
L0mKEDMmGMesvPakTVfBs6kT+BN/SReXLnoui93Gr/NJpKXH8whmGG1zj6ytXn5C
EVwH6tZ7OiMdwtEQMfgl7mUKPY15zIuh/nhR/bY0MxmsoRvKPfJahkZBETaY1iu2
gXirifnb1gRvGrQjrhEWhfvrLzk0mkzdbBzq6NAr5jeMLEQH48oDHdaD6NEzEQt3
LpJIwWGjJ5Ka0tpaN8eWd9PAzOQ/5/paZM1Cw2o42Y399sTpGw6HpRjfTQWNI/dQ
fIsDtzZFGJFo5x7r7WUmjdfLjcrtWCJYjQ0ZowPtJB8AxK0PsZX2avG3NWAYFRjs
5kWS0+M/v9hv/lBX0bdICNLQOtIsPlhPClHgELu85S/KrPzt/4RuVHM4v1AFlYFJ
+/f7oGF5S7bIFji4MLUWxReB8+mNx7tTnEPQnZtnoxi0UOB69qX7kMBB0vv7k98l
J2/cZPaUgtqkgPIJ7Ig7DhKCPDcJqfvPjLyg2QqZERmmeFCCnz3ni8632m4NqhwD
yChe6mRNefGtpFJ4hiwfPTmhgGgEXoSknjNtmA4ZuHZgC9U4l/80ZnoZu9nzS6iy
iIJ4tgpBu6MaC+/4rhY9fjJWR535cuJkFnoV4F1p9vHg3I0IeBnu/j2reXtDbmWz
1NNCaPb5fEZPLoKEQZibc/1ZrhWRXB70o4zRJSDTo4yEQl8i3T5eTCVf/cwK5m+G
dwfjyh6LjhOoTXt2DaBTDdgWckUGzTexsr9hCzz2GzcCWHDriQ6XCmbiluI4bHP5
MqCtDMvj3qrHCgTEyvrBm39Lhd4QTVpQUymrWmVpOPQmd7IPrh46uv3T0DtVzzfX
5N/DlPMBYmILZ0GPy2AT2Y1ArlLw2Q/s6Nvp0OxGl8inwzILUzxryodAzu7JBXfM
AieVFUWoWS5v932CshCfBHvhulXDmcXs0v+7vt6ugmWMKCaUV7rOHnM6FWPwM9DD
W2jdJ7KcgG0mPxwOr91ARh8LPlH9jjRVxGknpXDVzgdxRd21fGzHEnadK9PpQt9E
GdIwjO+zsQTeF3H6RHwWCOM2/ckpGwtzgUAxf3NVyQ7A1JoNLwTohviExciRKbxf
ITERezTG+XRfQ/mvEAhmugupVaWBNhRUnAdZPKgFKo7gqCeS9xok1OOU5xfAtcWm
jhhATkoLlrXoYaZhClWc4dcOB9kMBWHWMhywXqY+3GnDBuR4ZWx+IWayuIG53f6L
qp7PmIlGgH9dRfe1MrSFQ91C/WciF7bmG48PfTXNofhi1OAVhtqfwXqqiOxfLD+V
7cn75NI3rCQxE09VNai6EK1SgtzB6Ki9vW0MZ2B7B/9CCwxWAH4nMKAyXSCAt+sU
kvK/MAbziW1GeBG0M2qLwQUE4eL6vbHcb959A2u86Q3xILMp3iOaQ9vqBlTR2N6C
ULoYtY/00Un4RyaK8eqIW6C6q9bfVco9JFX4p+QDXI+QmmfQAQJ6wQTZIesPGRTM
PoMQW7hD6fywFmX42rzrDLX1Ez0VIQ98+XwjyGRam0qcPF4eoNHy+JG2K9jA83mP
Y+U1Fi0QtAy8kMn0k5b/ufODLj3/xzGmC82YQi5I2h5jcBnqK/moimnIpenyYw/M
wcBsyG0o7/QYTYrW4otwT6sgZDX3bKa6gnrFiBAgkF3Cb4CuAjEWgE7Pryse/f94
Cvuvth3vJFk7lV2fySADxpenuub5YFBMSj3nmUt7kCSMsaOrSYgzKv/Y+0qA9M2f
ckCwJhPXIBDUsKZ0DmI1jvXdMSCZAjU99w0ChqIN4pUKcTalA2yrV6dUCM0tyjcU
F6g9im5saxzeFUNtL9EzoNCSzh9yqrxOAzxi652PBS+G1VO3JSO711ZXO7q4C5ns
RCBSt42OqJPYzJbWEqFGQRjhjeNeUS0N+GY3oU2I2X/A+K/bPq86LLzpzF9jz4Xw
62HqZ5Sy+q+4L1BYEz8plu75dMmdyA2t1zj1MRdSE9Plj7ncReBpL0dNPHugpYea
u9pCgQdWP5GKd5t5sNRi+OC4tF+skQRsFjJqr2Sy427O9ZrPfTF9qa8bBqxPdmBh
ImT8cFWMzNrtXrP9lOz3dEC2uPZsaI8dWo41lss31keikC6Y48ippNpmnowdf5xE
m7PhAwBkxrZ1VCaGAYGh7AMK2/hIdXGALQeYTAbsvxxHHP3VZpO1/w2qfl62AKs7
qGWE3p2q3FrNpqRo4QSJXFD9jPnL6dV0/H9ZaZbI4+m9g5svwegHKwNc/md/qAHv
qK85I0VYrDM4gX8lJBDLiyvRp+lo1onE9jmhCjh3vn5tBd7rFtFa3fj4npcOu0ob
9tuEr5Kvlh8a7zV24LBqAiLU9bm83VH9tbL1Mbk8p+iG98inogjuH2j9IPfxizt4
MuqvFVrYuw9uXaANlr1xTKqLZn7wnphRRNIc7C0vFMlHHUUbercTl6CdLK5pxUL1
ou5VfvjQWowEHWmrtI39CyYWXIegAx8+L1c42N3q9mzc0jWopCtMjBXJCkLA12X7
rnPXZnvQymJ0jqSvRSemjBMEPFRQ18E4DrsAN8qEv6nH5dHtVA8glCHteUVs6cbY
iyUtPzS0L6f4ycr0o7yxHQb4RKEZjKbhxG2NCQoI3i+2WY8j0SkRf1rqZBqKdALi
3tOaYfo4RyFxEOVufZ4Y2JDGdJuG+yrtdTaNGKx3RGdA3U9GmdGvP1kHhIgTyKJl
I+KlqGWreKosANt0AUd3D5isa8m7Jqpdo+xeRy35qHLbmKLKsGc+/VOq8hl0nNZL
PQyxB37eYK3sa43az908dJ/V+/zeSx64xDCAHjY3DYpj114LeKKFbWJVpJc2t/nK
jW5Stn6dlaNKXEtjru8Z02bnbJE/kIEpsS8cnkaaDnHUv+X5H7U6ewIoRdGKP+b1
2K5sKW+GU49pyMNgb2jnX7vEFRvWizgl01R5o71YAcx4+P3QcnMEVEG3FbEPL7eg
Dh6CrRTYNnunVTiEmolYPZg+rInM2lXHTlWmLMGKhidcJXv4IIrJ8f8OdVWUy09v
7Zc76oNzijb/kLaKKeqmFb+8Dy5Zvq9AQhSnyr8wyc5faGMnTi0tQCzX05xa30er
uYGB0r9PqgjQxSP6xIzvWTFEjye7OTJA14yR/0oLAGHM48KJSh0b0YVSv927nYVg
s1gATZwQfmXcF93mFIwehWptFcy+0rl5UQqDjxJxGdAL8WOUE3ylONy+Xjk9yhyg
Yu1wCuTkVUeeKi7UMlY7PRcn8hG9xJcOH3qfon7ZLTJyR0TdZXu0t/Qi0g+415u6
by/8EaLaPzv+qrliMQmMiZNQyPfzOkG/+QDmvYmItqlPV7/kpHwMHwL04DY0UFif
lLy2nkD3aDe70talrynIKlubxv+HmScDbJWaFPDofGhrLWPtUvRqnfWEE3hYRvRI
ACj2v/HQj85JqN9iJ+P7Coj3F68uK2Xj7vi5yWR0vQ5l8HXNyPniCIrMps5klT4Q
rwGrAnWxg38WKiVVdTf7gRX4Ja1SYcfrDjq0y0F0CSJ3BetLvNO66GfnoQ8gOa9t
7ID7EyMgLeDa1nwX2CpKOIQA95klMPrlTrxJiRdXG4EmFEs8eE9PYPPkmaSkkU7n
rwklOyBjb0q4br3+12MUK4jqYCTsd2julY9uQgnpFab4ucGzJR+JxsflcDTQGp2f
qdobaQAxqLl0unHkdGLNgcVEDMTCOt5tCATaiBA94+eRqGs7IuKrISv3OSfoe6kz
wYgwa1EOGDi9IOpsfy9MQQyooSEbgG6vRKYc9DDpKgguCTWIV6WnSac1UvQniZ9F
DTaQzjiSy2DS+BMULEWVMX8D/ov7QtJaqPC0FD0ft8CkPkyikX8qPNxFrGf45a0k
tDnljntumGtC3A9yPeu88SIvwKFnKVSFrF1gvHR5FfYBz1C8siI1C537oZhg7sXm
/kkTn4BNPg2RhC+AIBAAWyNB9yeTpnnYRuYUCJTm+Xw9UiP/I6gwvBCJCM+L29fQ
Mdr6wFhI7aDXuhQX8yARCq8C3AmkzlTk/6YLzSt6Lw56+YIjjoJc9GkF5DNAg6Jt
ehThLARriBoa0F5JnJfNVckgi9q1PrbzBTXmZ6CoKI/+4awZde8ScyMDw0FtZSJF
bfKfbpVKYMZSkuQ9SZGMqw0/yc+xQurIpVa1yxerR+FkQ0ygdxhTd+7mlVUUSpiw
ZKWoC9Vrp3IzayqEfIbmCZmzbH1nFdNT/i0fTAoGIIugnmjDXPSoAWGmPD6kU97N
nNiG6gG/3t8pfP1FAKyRptEX6M9O6tSBZy/PuvWDCqxTTPKAee9gDdF+Yzvqpls7
E42upxhvA1LClEmgPy36YRE10UkViGbQjOTgEpkKfBe41fQZOtNRcVxq5L0ZTemW
3L9mfhLxuy8tyh3v+I1tgEed3JjCdsTnSlWrNXPVVqOq0u2gMmlTLsavGqOnAHw8
sAyqsl/JHCCcjliEl6YOkn166xbElCMubAkgTnOc59qYe+s2FKrbTnvFp6D0YYSF
Gq1tR6venqUtJ/854H4uFhwixIkaiHv57WlMta3WBSFppN18tyjggIPhjF1gAJge
SsNdQ61blTz57Rthuqe3m2HaLLMoMB1creR1gD/vS7gfUl2l0bOu3I3dyfufXTZr
3NdNFwZ9V3NANNLmbg6NijOwhxrkmDqUig4kUBBVFlf6JE2JzjEFfDl/1BXEoXE+
VonJRyGd8885GUKF4jxQdTtBi1wCwwGuYvnurD7u5n4D3AcB0xjbkF0rImmgGP5/
Z64KTPMhQvBNAYF3ov+VzLJ1WqN2NFgoRPNnQqd7isj6H/y9pkB33LjX3ULPBkI1
CbCQ06YgF6FN/yiZ3MyVbzuWa8xIwjzC401A2c7IgI29yu288eWq4o6xQBM9qm9W
l4MrTd2Bl9SoxKjEtSoRbofrXIhVoCw9joJRZcHcOeq/PO+MWYqQo2Otq7maWfov
WAUvBCpHsxpWEwa1gkTebEn/GSGr7AfjLie2/kZwdlOavU5j088gaGG+a+LObtYk
GfxkuMw8e6Bn03ANB3AHNtD1HUNJnAUVvRoHfnxjm3tJXMjalyuNd61SoN6jxF13
neCkUqu7BIrLV2GecBv8lKL2dIZ1olbs9Nm3+au86xKAcEXZlElI5XUG0Nsaezkf
UjWJV1SWwyGPoZ5eWtJDhDP93Xw2y2DO8E679+F3p0jUPU4LwSMbt2pnKvXYfkNb
u7Ls7smWU/Zt5jhmRM7r+O+EOYrDDN8N924Om26QbsGMWFfjiUGzF7kF3ytyTvJ2
DH40Viwf8t8H2HURiLuGkH9L0hVqsMGnzFTnP/s+d1Ofh4DsDkO7NrFnXNNaLe4U
p9PMPGrmjhwQHSlYNRXjnO9WRBip5BljZBKwUopgBS7RH6PpeHt0bqaO+IGxg5mo
yhFfpjHNKTUnf4gvjCKDBJ9g9tln0eFglU805sjIf1FWi20eG7gIQEU6EujAyGeH
hyt4aaQ+PXnsfGsTDyOJBMtrNXSO4b5KDPc16vkiGwfS5whWHz4/SucVWGt6xTYK
uGWudgRBfg2aIz65U+tw5gUnDjnateL/JfrAVlHUEnua7n8L12gNZyTjdgPk6TiT
TE3mSFM3A868QKeQbcPJXQ0Y7hqFjm9Rqw1lwaaW7NUmEg+IACXoaHNpTuFpj0Jz
bD2gUa/oZ12hGMV2iL29rKEU9NePIghydNFPsgbChKveVhddQFOqy9S/eOSSc9mr
TCY6Iu4opL+dzfTPJp/rqJgR5t0ZfkDst5yWAhTNn6IDbPPjciKMb1tpS3rnljpQ
kJESk3TIOmwEEL+F/5mdvsp9Gll+7K8xAhZf6Ucjss40z2b0NFnvgJrM290imdd2
joq54LyImMZPuyIQiXAvjh4XlCYpv5P9rLor+ATphYfuEq+11MDnMzeJQL0vTIc0
NJU6/i+9eqUCkvJgJyEvnztYqI74Jh2lvt+ACzgs85esr2a4+tJiVBludc6ud/cu
VW3/c+WKGEVSBdaO6P7/zg/PHQkQdpeVemR0TS88BHen0px4sMdDXxADQzWvWaTu
Jh4ooyxhahzUZkjDtH6NWFL+zS0nmo3DLCo9JfFwduZQZwSKFut3P8JOIqsti7YE
8WnOw8pAV0FoRPcgdDkonMqPT1v2LWevphCcY+JgLUBImQpRznueBHqYEgYb82Bm
g/IQeOcRtmKoXUSzr3MMPbRyFs8mfredKJN+XnHPdYk18g8YhVlOTQWkB/ye+PzB
589l1vswwsL0caAFM2029UsvzyKNla89A4QQ/FASUHeab5vYO/YZ/CXrCpTpRpYy
CDGgBs8+YKMN1HUVeU3NmdwrscqhDbfiFdXpQwFdaIXwUlYdnjE0TAlCG2ajh6dw
gAQpCVNt19u3BAgYOeGN92hmSpbGKbJhdq2J+eNOGm8IDIdhm3UCsOewjG7KPDmN
oYhWD5TNCebdYUYLc5ZhaQGEQLn6v8ISt/bvg8XZ7sKneB9fiTVDa21AyJnHzyHz
u2V3godWYGO5wSJYPHxlIx7pS6Uo7km250ySSidFR6CIZWbtKL+w3qWRVdTJesHr
wHl/eDbKUNUl/3LCH8FDmCIvDSr+hnGk9BZxZSC4+JRJoGpnKRNzkPCM6QoCPDOE
k7d2yq5wtt+rqqfMkrXp0lyZ0fkL6WYkCvO5jUNiYxJYbrA+pGGggdLnongu1DlE
QwQFuM7gxqnF7O7uAiTJW857rett+2HbojKBAVG4ZVOKeusT1Z2kdFmQQGqZYHc3
ASLlN1Ltpb7EKOVg/ioo7V/8WOyFZ/q8Qg4rutKoyMh7+AY72ZCdNJUO9NznOwwn
sYckiddaBl1WMVUb1fVF3c6KEH2y+qCRbTgljoAO/Z3DyfITwO7tLnXeDy6gnVax
6P82XdA69uS7III6LdvJJoE1QZUU25DW6K0oZc2O453AhOwAmfolUA/wJBg/yV6I
R6hl8rk8DtppzaSJx8I8UllbBjnHT2zgTzZ00dkm3tby9la0BRKb9/oEhllzOVp9
sfGNYVJIxSnPctwclPvIICUwX3PY8OXVqWetxfes7i1tVShZ/Tb/diwR1HzRSrf+
MWqUreuuODJlXUyFbDT1KYUamKWGQsqc/OStmk2WpkqxfLfWfHfkYal7KkahZKHo
ihm9H9LMAi5TZdeSp1zf6E/l+gyZ1jK7RnO7vdY7iRfB+1Kr1mcEom018cg0yywO
jLE0FVGbhsWS2u3UZfQWFzcfPNTg52Vnv0WZG94EU9bDQAzcRJY5XTbNC/baVphr
YMT957LIly1aySyICggUiwyH2hnNzsqy8O/8mtyPmbf3AwV0TjkEMlt0kiUutAJP
cNsFyI7qQC26kcrjAE2g0C+CFa40QwHzm3ik4AMDqHuzslBQSmSi/S5pkZVrP95H
kzGcSKuIoRMPphvnOuQWeWfQS+TFn7TvO3MEzVkaOgZsRw7GyVgc6B14u/uVlyFT
v/xqYKFb64Y/Ga5g84z61Ahwb1UC1bUXoFJTBhz+o8367KCAyVia1jPD7WAO38Mw
XektebDyhW4/P3tVwtVygXFL9DiUKM9M+pahjcVQTubu5452BpyAP5dWNfAAloiN
8NfbQ5a37nCzMVFi09r5B6u0KYiKJiHFpIZRxP/xkRbjvTOL6TQl9V1Ecm/COOzX
J3HVYcTxuwwUcS/Pp1e++ykeByuYZeVMhjdHwhwwUTjgkWdBmzvHwQNQX84IY25V
MoGvC4tEFHuo2Y+z0ziJkCiQkjz/IDOpQulpJMvdLv10JtURFrjSog4Q17pOFcel
EBDS1cwAyoGabg/K+OxgIOhqTQDJxvwAajgVWHu779Xo4QjCoLXS3U/7HgFAMUK/
KpAZP53BuEyj93a+ykcKgPuaNTCJIa8lKmevS7N5+Iy+g6JdgMbwLN5PUB/rYCoD
Agal3+1GsDzfnyFmVL9Y29vK+tI2hhTjY15bP/Mw821/HFdnR1Aa89PEcfiAwe+G
e5YPX9R6KXiCsO0MCuO0+mCaKIry17fXFV4g5W7g5mtuSw9odLNZE6yFN/w3QEPb
RjAHsmuo2yQ75+kak3FfwPlu4p3m7E+H0er53y7Xb9is/bEm4sytGAZ7mywfFB/z
+92NX/JcdeMSdl/sq15hFeMOk57eeRA+O0cMOfO31jTep9nnp67GXCtO5crPu1NN
rUxpEIUPbDBukCcUo00FR2H9tMu0c957NhFqGqqj7Z6VHCYA0AVlIqNY2ZbBuyLp
Mbz/Ag3EKZwOL5pdaSguQX7VwQbemPrUl0wGEE93+FsGeox0TxDkJFO04sgU3jTg
igRG3uGzF32YRnWqJxG5aZL7LJWvWzPDtwHvZkxCrycnu3PlLbUVVGYoR10LllAM
5qEuTOZX04aBx3xSLGiq3AZrMd+2nkWKpM+5klN07tBMB0I26/znGEhtzx+lJVgS
pUx/NcYvgHWxcqWGrZ5/xcX8oQnEsVtxbx5KkE0Pg+lTrwG5k4FDrsors5Q2bdSV
aFSgGAUx81QNvfJoWcaSPyH6391jclj+MCO97BbCQgn0prpOqFDdgNpe1/+/zkXc
Jy2XyGX+8H3Fs8/y23Fb7UacEBs1r0Kmur7xc17axtSvnAXeGWFY7lUKJdFSzRRQ
/SKhHEmYo3RY2ZPS4GgvjxYfqY4sbQjfsXP/bkg/tZ5SfPVwD0q4IxDEZ+AmM5et
DgOjxeaG2hofQW2EymRvF0JidyQWuibpQ1PiJJ/6w/ipuT5kNKdqloNguvOQ7AHA
RRNanGiNHweDOKbPARa67KqSKBkUkzBsvRI6QOcmCH16AYDVuXpQgShj7SkUQd0e
uILYgSBqfipXI52srdSKVeIZi+TI1dTeojEPKoH5nQwdL4Wm+OgULberbHJYaxIX
eNCIDUpSRd4oyiZpz+2ovNxv0xmJueQusZHRUEgHaWgMwfcJOvm7ymvP6tBt1MPr
8iBXl+FQxEmCIib5vsxwetcUN3WVEnqxQqdXYkMAiTnV2mchKQ88zmPnH21aO9Wp
M2nd8YjTAgOgrP63MIG1t5fOq5O3pwTia1ej+bXTNy8YRwnYYyKMOFza8LaCXdHs
lF/J5hXWD7VU9V367J53hxEuFQdf+mAUFmCr0O/QvzCNnA5hiK+lZKkWJRlnWY+Q
I/mxbwN+AeMMQqEo5B2T7HJAh0I0l1cyp/UvsPPSv4g8LbNbIsrxwZl8Xe3/ymdR
g6ObgP5YSpuHEwpAgkqxtHj/keKvkMIFrygQnVIvuyxoweYrM+dOSbsK+O6qlTnb
vieoV2ZPvFnoZIQn0UB6GrJtGVqNaLgk0KqBMBcpsW7k/NIi+Udum0GjvX1Mf9FE
bVvcaK7jJh4Q2VEmvDqM5X8N7L42jl/z6LMRJKKmyzH8lIb/hqNrfCUgggmvSweC
5gay1ebkeBytoBsq6SpJRD4s/Fq3rw0G+zuq6WP6kz9zDUWZPEZS4ytjr+7LWmos
EhNcZYyznYL7taysD86WwY+VPWqdasSodsJXJeOiQh22Ucl/1SAiAKYG/SabXAPu
USyaxPvagxu0r9EwZj5g4tPmNUvUeeXvIjthV+txAC4lhVNkt/9bUjUZVwmdGlAc
+SlH/rtM5z6bdt3kqRsyjdVXVmgydpsV68dtNPc2U8O/gPldkm+MYlr8YA00rnv2
heqal86BzySjTfgNB/zXTvrYFevTvZbouMQg8b+LiEdLxWCnnix+Hq2367gpwZKi
xEx6IJdNxvCSPv7S/PJHST4Hl5ezRJ7FLK5Li0Woh9JPnojzE/zwsbIzZdpOYmvi
2i9oKfI2NBV5tcLPprAwBIC8A96Cr5CZWMniOc3mR5ssbuhg+xH1abGehoWWjH/9
bFZUoFYlrxkvp06b+uxO3yiPq+Z4IHoRyvXUSJe9XZ0bcnNIFZzlKQMEv9jfk4SD
G9SqDNkrLsYvo4YXEgDpIgcDu0maOBipa0LT/TXndl9dx6+NTOyk69zUBWLZxniy
UuVLZKUpfo32fOttut5gI5TLiIsDHmZlKmxOps73zXJfWQfQWrxU7tBr7iShnqvM
QhTYaYLapG/1oCnl5hQxWUlNy1Yp7DTwMVTgHLTosaBtNDsXEHckup7VrhmPPL/G
Zf+uAz5pdPhV85vZzMrL2L6z0jzMUG0m4WaJ6lZ+suDoodxgE38/Ank+kQOqzBeo
ukoHdN1yskMlFPuHe6+axPZcgW8dG6YtPkGFhWfnvZLKMMVV59GTXRuZH1fa1dct
0UOiWDDkqYG8Z0plKFqP6J9fZajKCng5XcSZtUcx7gJ4C1jSBELzaLIPMk+ucSbq
Dj4ooWDtPrQlHPVvGHfq6/WdW5y43pDdZlk5vX/VN5f70iPprqPnuNL4OTt4ceZ9
Uc0V88cyRJc++Z8wLUsuIPV6vd1CLDSobpwhUPsbYBMdpzbnoyVextv14XIpqqc4
qjDZSLZZzfTRJNRPq7PFdknS+gy3zlEGBTSJfPg7d40fvwy/BXrahsvHmcltW6lK
/kjNFvC0yQw5K5ndSRAnLNYbht8Hn3F7PASwCycnibfzH/sAVg8/UGX1Om0YGTAW
JygQ6p7NP/2t6+P+UNlZK5ZS7Cfqb0CozyCGHqV67vHb/46j4e6EJLeGDDbTZw89
J2bn+5F33p8JKLOSHY5BlFEyBxip1V6Dsb36OACNzlYEoVsBOwV8Zlp3jHyObrH/
r827/2Em9a8MXaBFM9kYwIC4i6IbWjw6Q3DiR6/cXP5h8O9Jf1OojhSkQ7d77u4b
2XC0aPukFApS+RQ95rK/IM9CAmFoFwbjEEK2wV3TBxxwoZz6mnV5Wo0LtkZwHr3l
BIclg8VlT2iKJk18dvoc8EcSrhw6nvcuY+wGD5o95rVpPt6uvmTpo0KKRhKMVjTM
iSXQmwGsvKFW/jTH5eFF+iqaO2cgQQfdpMZ3EuxhqiBzeSQnrZPdXgmqvnqndS1+
rEPY+8dmRVtoLhBGVCd0mRCVWqxIeUzQOOiVpbHAZag8UTPaSR78POFLmvXVdoAY
cxo31LwhnZwiNOrIXWmI5vsFfaRvAseMiLkbuGt//P2eD3KLbZ1q29wftZjy+0vY
7CldnjlF7GoKiURL3H2njnRnNaNNPHRZM8DLJjRnY59DuVYZqJn2IHfzdfno6Ffg
Wq2OGYiBCCr3fHmj6xa198KqERRZXb8SppFgCFrk2dkQO9GvSuwz3jIAVPySOeG8
HB1WK4/o4QZssaOf/wCBChx8PokgsDv415oepa5rdXE2eRg73KlwAiS8qGwx+I1j
njQSx917HhAF2DhoaueV1kL9gwNBDf0Il1zRKg90+2FJA5oO64PuoxSL7X2HWDGy
511P4yHFSJBqT/HWAPsf4GVbXH6NNP0kmIj6lqV0PKCWgREAFU3Ssy/pzJbPYKbM
J9ft8FnQ6WU77ev6PCa5hGqNX/GdSHqsicCWv72UQ4AxchDJzQktk4q/hOFImy83
tUHIpSJ265Xssnh3UEg3a9JwBDv6hmmzVI0z124EYCGg4msz1Jgwslfu1hOWTh/A
1o5nEUQPcfyySSIk3my3ClPnl0tOgQAcozkC6jV3GLz8KGEu9t5HECOC+bH+iBGg
RZio3bEOnJxflc3R8Kfi29MyJO1o3tOG+G0Hu4F8YGGDwq+TNpFiyMRCQh99Ii22
LTCghhBVO8L17dIlkXJuzmyZ9hC7arb+BiPj+NQFmbIv1xHEsrZYXvyF1e5wIlUG
7i3f+jegjz1KeDdpd5LyqA6PTuy4e/jrpzSfn47FEsUlwUnyM7O3AMRogGQf7JAI
1S0nEIhvEkoM7zkZFEBmB9uC/s7PnFqv86Di/w5mi9FxNbhHXt9I3IlKn7HlLib2
ZJItaWiIiNo/rDCcxdIO8xmbEi+lka1I2putDLC3VSCLRhkZjC7pk1Fl5v4zvagu
OgkQkS7hN21R0VwXBJXPCE20ECm4O7FFwPEgC8/T1idHSpD5iLcjySzMyGooB624
yyDBud0s++rC2dygBtRhghQi64WpjxSiVyfaEcxcd4EKjVo8ubWDTa6CXoW1LgdP
GXUtlsDBiOwy0FT2fJDxReDXYNJI6pA8EqBv8UcvynbQuTGMa1yvRHTtm3trxpeM
7b2/6zWlzEZwzbbuoHdOlm6LoOSibxC5JKSs7ddXrq1lPL8+IjZkHPOGqOCaLUtH
seED5pmPwnlD4SDqW9En+dTibvN5Eh6p9U2oXUW/JJTxX77I87DqWuFPUyVO1WTy
W6xc5+n5s+Jt7iKY9ebtrEKdVJz9SiDpfOyIjBmXF7mKhexIBqRwcAAO1+NIb04y
d7noXZ4BUpIHjKavfBlqDKIAVSOm1XAEyJWTsnTFbV+bT83TCgDYqfIYC2M9Rsq3
jJqqXa20Xex2Ld3HXhHWL0A/ND4dtRsG2RkDpaRdUeFZOgl1l/jz32e8HVvZ6Gc3
9yQ/IKq4nEpV8sQsPROc5PaQ+qTiyzpdFN7F4fdjEwnB9HsKrl3sZrra4Eia7Xke
QPmS2KDvj2z9NkRWY7ARMpzeLQhUQdEKQ+q6df7yVQBOtMvoRDT70vgry0j87mJD
xrTwS+RFEvV1FnkKbv53XKFDNGzWJhKqyKUhC/jvQ/3NLWw+w9e5TA/ovN1Gja7U
0NwGRPzs/tlQRIRCyZddpuxJ40hp+7QYQ1acdJIe8NBiopdFLeVnpnhY7v4n5HXR
vztG8hKOteKywKCyS9cFWRMS3DfhrsbUa5DE85AMSvmEKpIL9pNe6yDU9R69i2ju
+teBb7awP59So+Bppi8FYOiB1vPiX08PamIUknikKoAd311oIdTfIHo7e0pB4bhQ
xqwOKucMqwLzDI2yzscow0/1upMBxCufCCHgXY8bDEv1RmKDjWeYVoCOlo9FhsHG
Q6VA7ibzedF+zxm+6Zz4vhMdsvKjfJihFqyPhEWTNZfiAWINmAnc03StxhVj3g8Y
2rhce0IhfF5vV3wlfv+rYS2r1rdiDTrT6K8+maiUStfSHbAVMaLlhtt4RXHkEQCD
7hLRNeqYRF5cLM5+CVUqk2STyR4CaiEeBPTKj5ZiDGDfg4bZlKEaxCAMoUMuzby+
wAbwcSCGLmyuueFlc/vGSJCvWQc50qxpTVX4HFIH6rahLrYe/0T+gpaSA83oy3o6
QA2yUG4O04B6yb+tg0v8w7rzqBxGRDZTFbY50PNi+CsJt4vpAhsoRaq6jySiLmtd
YWSitMy5xrVLgP2H3CxDlkWyPiqazRGCw1pchz4uRwEoyc/qHlCfg+KZJcYZL8y3
GXEeCkdjE/JOsFxhG+xPChVljcz32pPbIb03MKnwNrlfvoMZRzvUct59MaXNJJL+
p1VLiBo1QMLkdedJWAEtAbFImbGgR9HOApWAieIlfLizZgT0DHHjtWgNL+jZDlWM
RR6PiQWIEwAzfW5H/FMCTNvZYatjNCkQCbfSoe/AuLIjsQ946g6I6XuPFqRvnhj7
UWqw9A9MbQcXwwW2eNwKLK7Gm2o7gmTkr7EinhZ9Kmg5TnfBeqE/ULvLYEkfWdwq
IKkXDv3Hlnys0xQOm1/YAKzw8EdGz7dEYviLj7Qjv75oPECq7xxZVcP0PKSv3y1W
tuh3zaK8Y6aNhbrkgFop6y8SUhtPbdFEcByegvoVSiQumH5q/FOayv7mCXwug0w1
1yhW/jcwEH/tp1kDprGwXTOVWIJ+MT81TriiT/QmG4716eJa74VY7V9gHClt6ipm
MNSD+wkjaZlQS6s4RwLg47LDQUSdkqHqyh9B8BAZCk3kysKJvGugNww2qiy01rX2
E5RFnnAwMDx7q4acISZf7kJBiokqqQ1SMqWeLljpFbFbk+G4Bzww0oE4uzHI/LTy
Q4jBbm8bCNS/07hI53nu5C0v7NbV25w0217QmdCJQHpp4wQSK+K3tIMOtZo0Bixb
uE22PY4ckOnyyLcUdOjqB7MhlzZ4ukpkDFnaLCcSb9lmXJ1bPVueUnsgaQqIGLlf
75dK8Qot5A9+ov/Zq+TpMFLP74/7akR37d96Dwb/gBodPHfMXp8IEOl3u0+M7Y7e
X0q7Ab9GFOsfzrHaRXHQbRLgTxn8P5GaZAOfsCKWTZ5a9WMjnx7yvQZxed42VuhT
TuEyYeLWrCZUu04KHETqv245O5qJuii1zPtzR+1LAKLboMB1iX0ZzVa5yR8MgGIX
rKpzkRPTjiwXVGGbZCK2+Hhc/rL10i0DdLknydUn96Ymg/5a6pu+DOwiPDVjqGOr
1D5RlmOFzJJNaeqdPFQXGmpwVoxGU7n0qA4cEmSEpDsMj5waUqGMj2MR5O/xpEoa
K/7XC0bEcOdQ7hNi7oxOJvCtRPxqswSh5arObwZcE4yJ8hgtB6+5IMdGNVI54+X6
gJI0YV7NuWlP94ZiVApiu+pYX2YGd6yGcNltaZ+B7ZuOSgECfXselHfnMDLGrapa
X86+T+U/NkS+BnCjCUDg0EZq0B5LOofsWIhY5zEJmbY35M6r9Jt7awKELd//nAwI
mInIUNt/nn6tqu45g0Kfko1f3sQrSLr1N5AP2xI3TePXix/MuIrhIKiPMliwZM3o
AbGiMMvymT8RQ252bnSB8sTNejBTvRzFQFBi9n5ZoMzaRiS1MPHCOBuFm6qDX2cJ
qhArH3mFXOtYi42vixnbcZfJ0fA2VhC6cqcuxsQbknN1fwsd6YCfWmxysFMuIOAj
JVKdJL2bJFR9t8YoQuVzJy4jF4EujEoLhHZF131emCdhxzuiBb1zZbrDEOu+R9Zd
cc4LV9cqspkzdvxbGzdvXZeFnz5/bjnQCrJevqewNFmdYHm7E3GPbW00hZx4hCz/
uaQbgp8EV45Rq8+fpCj4F1H1efCnj6yGycw0TzWwgVqkCKwTVFnz8oeXYBKD19xX
SuKYGKNIP1+FZ2KnvD1LPOXxKhDSsXolfLYzMgcHDCN8HGq068boh64usd37cc/z
mfF4+i4XTK2x7yvvftVKdjuIw1FjJY+s65Z1ahXVcK9msbdQC+AkPqrgLaMo1d0R
Ey16JQjykTNb8Iry/RAtgv44DQOuepA0TFU2xNBFfg0hTSSIrMz6s9kgV02mZgXr
03iYkuQfo0OAATotAQ7G3FI22Poy6RT/fHK5mm/0nNRMWcPAK7hvffPXhgGdeh4W
0ZQk+vXIzNPmV5vZibBrqymY0TSVKTYUyEMJxYNV0aHIuTWJc01RTBJXEWzvOXV/
s4E/EIf2adJD8TP2VbS1YHoedBR6COQF56e9EOiW/j+lg2vrztWqlNlrZ+ICeRJD
Cg/u/kwP6f0j1fSy8R5EJ0Z9ILgsBQPXKrNHJx9sesgFuPTGUeR/w5hi015OvO7R
Qp3MiqIdJrGT03YQaYxJAKdAaV71JV41TYYKpf0nRkgNq5IIdCpkLdp/f1V/XOSW
38mtICtbkgDoHRsevwyjCMKeWZ4MwXSUu/GLNLuclujwCQBa1gVb+YaAqpaBekEK
KTeAl74wyFxPE0fDWt36E4OIFiqANEVeV1a8xYxEfPfbuZSwcS65AciqJCSauk/E
zsw05WwlZJgT9uhyuiOpATZPpyF0dORCZID9LSb9wZz5FTsDkhiMpWfPxLOM7geI
RhTdPgJ4PwqdmRF3YcrNCoB+TGIG+vGqd+1H8ymMsJH+jw1e9lUYWD6BL0OD0rQr
7eBKDklRb68PGhxBLuxLJTFf9XN3JUiDDwgu8/BUQJaRilrAmx70sToybEuDHTu0
yrjIcQ7nEOSTs0GEq+8meiRYEuXA8xSv9LLnNDxZaIB2+aX9fay/9aRKQ3mjs8Gp
+IqS7VTM80mHvN7o2jgfCBOGEgsof/KrZ8e7qiipN49yGxHWtaB0A1yYMOIKoiBU
6Kwfo7SkvDrSQWywe314wYUeE4O0hP+Z90IpGeEmiKTictWsVcHUJWnOAasaZWGQ
QVs2ZWBrrMlvxPn3azGSHodCwSbLSipheW6hlWRA699itECATkzcbNx2Ar3i3c4d
fF4Ptdl0K6Rk3c9pgTa38QluKIp3LgY2fnNYkO1E1jJbeu+8uS3+kGumNmzQhcr2
8UUhC8YDvHccV3xc6Ht+DdRK8RhjMU/slH8fsvaEMtIOUNNhW1yjUGWF2T7S/wvf
4KOl0SJAlChQat3nENPpk4glIczukxziewO2SxsGh9ZXCOlMoFcxZkGGiqbSh2dY
GLL7xl4B1OOZHhqv4/Qc5VJkYt9AGrBOy9HA6UP3ga3u8QKu4wz1f3WX64spkXSE
lfxMsSmXULWZeUYBc2yu6rEXwGcZ6VvRCSidbvtXeJb6v/Dpvxjv4f2LfOfzm8cP
xAvaBZ/mL76NW7VU/7iPEX7EdTZ35CHAUita8sj5sxqQ7TzpTEkqEi6+4jyq1a+o
FAaLuyz1drGgDU1/WXTrC12keBdp9kkj3lNr5lFh5mAFh7JGwT2lubqW5BS1Z1F7
sxPfSB/XRQc+c9icehnZIfNJEg4ki9AvKraa9lzGZ57bVK6BYeUvjJ3Y4ABOEEca
zV3YJbRzc4tZWHl7esXeuYuwLhMTSM6Fp59BApyAzw1YPrOwIb4pD/7bA4waJuvC
UVfBg6KtUoXhTPNPfTxGOOgIr1N46nWPTtcNuSwqSDzRQsM0rmsB6pd2dYvgygWk
gr0My16T/e3KkCS59LQVlUZxnV5Z5XHpnEM/ILEp4gLyXWV0KgAO7UlpwTxUUyW4
EhBv//e36GUx9eRJmJ4lMeExiiu+cjqrqQext0dj40DF/UM/IlBpI89tRHCx5J9K
RTK7FUxiitJVsU3SYTin1gRvQaOgcpOZBWwVG7uqJlOuklJ7AG5Mk8i0uT5zDNyw
MI5MKq7QoKfvGiGk6ZQHrPK+HcTYJCDWoSFrIIrtHdiBDzkXfjoGvcoMj9T+FLEt
cj2Q4xYh83x0rIzbL4vMzu8Jr8Sm8iWrMA/nTl1L9IXdj9Cr6xMIs3DVfso7txxo
8YnwqxwEKtKD9NBqiQOedIY8Y5nDdHE4lgRJ7SMxMPSS+dsw7ap5KrfJRI/lA8Dz
h8x0zo1L+TtWJ9+bxK0Vk7B1x/7QESyRvonjCI9QY5jf73frwNJNIBibmSFSHdm0
qp3Ij6+1chUjNMnsMIvZFxyR8LYn+/sC7dHKw3rWeCWRXVuL0622kq+mG5DEggRn
x3g/ocd/xdmmbBIOGP3hFVzGrZQrDojUKs/pQbTM//bxOp96T3Qp3LJZBC0Hy1Yh
ZxoqdTVPHxZgfk6L84I8dEwfBz4wFXc82lFYwXQibngx/DKkBm5nGMZihP4IGZk9
1ytDzKHOI0njkvr6w54THPaExJ4czeYf6GYruI9qWIiCROgchVlVwstGwz0ewejO
vcMbMDa6mhftOq3BpYhrsAOYaow7VKwR+dZXRcpvF1fAGILLeVgoxB7d88b9QmKw
h9SyEQ6DCTbmxaGXMwMobsdNQq6GRIh2IWI7GCmy06iOgTUcLniFpkX9MtW0rA8P
gunBt6PIG+QukCnjd7QbXeM/9ZqTkz4qxZ3A6Fo0gGvK4xRUePhxwTEJBTUTY2pB
PYes9wbVthAU0Ve7LJQKbPt/sDISKBbeelJo0B0YhQi2AxXsv/snyWeCTEbv5Obl
T10aPTRoEWSIAMaelrQG7K8boswpmQZQUaVJMY9HahpFw0lQ6aaBorSy285j9fNF
5pb2KMHNxhCaMz6Di5fjuIg+fFcMAZEI7sEgCAxS6MzFQKWsivk0sVuMeNJuFh+p
9kjsaKCkuTpIh5HDcsmAcooEeh/AzZmOduoTgQ+krnVBZCIv0o0sQAMi/GzemOtt
CazdHmKZvSO9jeO/PvBGyXMruvNTWtvo84c8MKLKLFs4XgT5zc+n1JE83CQ+BByD
xtTefHihPXX/GoTo8Oi6wgTimuZgopvrY6gubYQUPrusn+cys6wX1Qa+ZThFTY93
q0uMjBIXL6axi9Ih2t8838JiOLnQmH9hUKF4Y8v1vlQUpkEuK0C+Jq22qPfzOuvr
wkvDQJKf6MR78/CC+DjflGTp6A+rA0CGnY//imoLtbZm7RzoqHoLvmGABrP9wLFJ
6/c32TDtD0dm3ViUQRuhzWD/KGcj8B9zdM74IAa5I+rJbaEMCwS1MkXRU6YUsmPO
DiInm1HYXJJNHaJayYQ97H9hTtQe/7+WAYrOgKthxE68y+pSxXIe6BZBOaYcKLvv
z+ixjEhgYKfrQjbAnI5R/thcOmln4XZRn9CR1rNt913XYocAHmWXeGOpKvW1wR6n
kek/EHmONUGW/g76iUjpC1Nz2oev7Ek6qPvFFG2LeSb9gxbQ2R+svF8z/TMIc34k
rnzwZBmAtSCITwTVhEP2wV7R4hEAwkmxi/kGOs5GndBumWG6rIog90tVOtAMvNX+
r+z/BD5i1mK2P1kkGgQpbG2pKmwUB3WOVf1KqRFkArb3QUD9+vR4Y7q+3f4ecgT1
5lcRGB57/SBTA09LoRRzjnZVeWd1S/8BALnm8+PRUpanaJ5YeySyKFJaxer0WnYC
dgsEtDr5rH+AqMeK0Iyv1HwnKo6ekxzkOaK05uJJXDStb3ovF4Ea5LTU3FU1hf1V
FPg8vwILswxgG+OsiiPP2p5oJO5IXYJSE7RFNfZ9vNGV+8wzrjmxxQ2SvTid0rYb
ZH3dpkMFHrhonRNz03s5XqgOZwXL/eNi/sy6bcKtooutAcNTMTR7QhBLiX8B2LFs
adhRD3IhHbU+EgX775cBq4OYfZZSW9U+pNLCZ5n2iSAmqOW1wgahEhqvX8lRUXB4
Hnhsf1gHXRxYtaMQtlEbjvfXARvRBmOeHNVRts1GctB5nDRhA6X5+B9UWajmfsVU
OlboDH/Yb4fbyeF6Iki65LeL4xqYIZ2dnHXcsPAT+15js++EUAp4lo9eJ9ww5TGj
TI2OZxgnOQaoKO57wnooYd+ZjLFDfFOMJ87gg43CARzwVnAusw52qayOrZppa3TN
eQoL1ezPMLKp+okQmZVYjNZM4CawOjkij7jO1+8DTxmrCTcM+2TPGNEvPgIVfXna
eci0fmKBwoLyh2Kz1R7fhlRjlQ52Wl2sqFIBoWRPScG2YsOgaGUreJrrWzMjKI3L
uIVY0rThfZ3boldLAvwkTRdGdeDRVjSlqWPAMQo2rvEJq3rCVTGNLvrBfGieBwiN
t35vknluPjqQWith8Q77yclmDhm8q0qpDLKziUxkBXwAaBYqfBVelhsm0X8+IcVR
fgYmc3GNHqcFqme7hzHh6R8r6X40XPMHyME2eJOThYDaWNZ3bFzwa4A5QtQSunmj
L9Gff6OTHlMcHSwz13cKfXZW7RbMeVEpeAEYjXhdI/67O4YEmiR40XytllhLFUhd
D9s8cRVEhK65gpcUOv9+VAFj9eWJ6jRyIjL2Gn6jiLs8dr2bipxCxJBW68dnxvBO
VOEDK+pKdmjziM3bsl23fYtxTOPVpJrq3CQdJomL5je2DwCR2kD28GJ+q8sH7Oly
tFCnygHDBBo4GazS/typ2GdXz646xxdzVuzPSRiSCPGX6PQL5W54MDLTXCPFp8aa
/FP6IBaa7+G9maCNDyouhQmg4HLSLzqCSSfxNSXGcWkvfd6BjDhAo42js+R/mQ/z
9W+2rrtCKJJcRr2j/WET7BkQOy4xVE5P112Z01Mc+vMFGx1/7EFgDQfpxSMTpoth
YJ1l77ZD4MDS07tOgEnqXkJiwJX+1lWet8qD6dr/KVCBK9vXDLIYCxGLLXdTeSqz
cAR+P5SOMtUfIRS+jzP2ljcrYMahmBoACUhJ18aLX+qMiFKoyQPn9vo36ns++ncM
6HZW2iVNZOvzs0tm69OV9OPK0IYVaFTQMVGdEjMR2Wntj53RPXN0Y4pP9lItRofK
WAEu0t+BB9V4VWKOegsQzkfRE+YgUoGB/IbESZDAzviQWMHuUlY9930W5aJ2ENBl
4lg8rG4wGJh8ABvTLTdhKktp6d5U5nktGFJSG/CN91DZCYyxn0xlxO1a6//QOR2A
IODQv/v1FvrV/HQVlFsvWOpNpv1x9n3tIAA3S02BcTN16OqRCu8jA4iHsf1hjpf2
OU8aX+k69XXYicdF3ar+CFlnPyZf+ZpbwJr6MrL0CjPWuRtuSKUvyXWe8X/0HbWj
FLmEdG3wrs5yDrmV7YeAuswfWwRWltr1YVXPIrJLnQOHtmxf362o50aZw4ozEONQ
d8P10amQtJTq/BNM0pZS3rkACtbMSqcGiEXTsBBU0eYQWzf3gJ36OMePClbeq+KM
GNqApKoaJXAZIVlXpSmTGVrcq8dJLtCk2nq8TlSzWwucD7D6Rm87P8FwdH0a9Ddf
T+OKQ5bWmmZeOUMWPQ1i2Ff+GNaAc72zFO+CEw7xYMc/EKPQtNgj6LELxTV3SIKn
Olipc6Hodg6m0riz3mzPl14S1g6zLgjoxip+bnhuJTPAYs3IXE4lii7pWc4QGHQ1
TnWKIyUWd6fxMWP9g3LG+SdWcvr0M2P/WNVXjAbmwXcsz17S2PljC2zLZjDT++QS
8IzjHBZdcSSEGhB2t5os72lzzP+4+GVVTGeSmb6AxmGTPUsZEe53cf1QqJRaT4WV
BaNtXCrnK5gsDjhUh8rmjbUNf5OS4OSrhn9iRWYusaOF4Gvrzq6a6qlgHQljkqL0
ScYKCUNSiNdsyfwEII6a2W4NfUIjAKOvxAy916H1PRih76NLu6+mlvST5rCE8PUs
qPhBJJaqHThi4t98S67FaG3qfSmBDlkhn7ya+W7B1GDLalV6A6VXD+M5810Cnr3I
82iuxVnFP8q4UIreq13Dq8VglNTR/4RDsH4HALKlwzVAcQjGrzTRL50wbfuT3Ra8
V5e0sSRyyz0McH7DURhVhy9Go4z5P+GPfhizPxgKR067jgXCqiWlRy7PozknRir2
cYBVsEaF6TmMcB5+VrxWtvUGl5zi0gGHDtYr2fFIKXM64xZXp+MDua2Frbn4tBXW
gjgBBRlfpc8J2Cs4cdHap6hqAoSMzaDpS0UfQBzkbQjDJOTZfsg9i3IFY4/1eSW8
CXode7FoFiwpKeRUiIQVqAA30QMiAWHpYzOLKOSDJMjjES4HN59wjLUBDC7oUFAQ
DEW4n33a9U5+eD5Taq32Mza8G6U5YtMCvbnWiQZM/Fbha9Nc+zGmAElEMhnlEXfk
+6RI3L2CoKIQ1aL1obVYTEIog0R/Zlb/ACC8+L8oe46E9VM930nGFZU9mwswKRXR
e8KDfdyhtrq7OxAw1duW8n6M0/BykMsSJa4pyovp+oYaz/EdcSQSDjn1rCEjBaR3
Xk26y92KlYv9yQ6Pr1QimHSu7II4POBUg0ng7zktkAz7JMHp+bVl6Nu4viv/5YUf
vEKnUnVv/QqnE1sS3kKeQdW7UjdfqYvHlxvfQ1T33DXvNcXmrClSQysXLXv+W7G+
F3Nz6lac658V5+EofGVVxA+9Sz1Wg0xe3mcn4RThNFnPgoLu4dd/nPSzfNWKtiQt
4OPtp+A50qSFWo7k48aRfimwGhGQRG6dWiV2M7fqTxR0P4NG97SnkLfrS+FLhHXS
UQ5h738QSfH4duLOaXTjqOqRdg/zPuXVy/6krq4fPYNYWnswPdniRrrE2FE7PrJz
RjpKOUfqwA4pumhKCqbDRFsvsHf9+ML+GjVTyuK6A6YrrW9Qi3A9OEl4Rqq+AbLD
OEdWavZbfQeUlbtdoR/fodzudihSTMDJeiasLlPR1JjM7JBa73oQbZBdYdPmF2VH
9F9Vj8GKadOXTnbrZH4k8z0PvKSXOl7z7YKbDafYrDluNp1YqaqADRzAcj8PNNNc
SnYtU4e/dZvivQdQQndh5vMLrE2nXjJEobaZe41yQvpQ/I1UyIfaUKJ1IqY4PzyN
Mi0G91fh43Hbqq39ppbcTeiYUyDk1G/U/frFSQMZRDaIVE1VDiRRspzFHqz2FzH9
4QDlw0SZ7xfTab9BGP6gMozmDSA8U63hdEcb+3XKBQOE4mYqJooCKfX/0etMHKnw
fTDMcG4YBgKzh0gnvL1lrShy0O1iVGSUhnGEkxF+G/sFUCZcNUCtQ7oFW8YzjcTR
T0PxNoe0FYRtkALiWdQtuo+4QnvQLGvhmUbuWtJZi9I77km7/zAKOTNOAZMIhk2G
ngeQ5Ay+kIn7gKuzyL8ZdT+CbyRKD//IfQpz2u3oJZzbb+CblU+QlT9sDteLCnyB
16hfgkXfce4Ujkl3F9Mt4SipVv303Bgo7ipf21uk27bUt8uoYmqo9EIdQlyXtNn8
EzYD76VIk/6/ruN6xRxaoWSEmzwkg+Ve+gpvhMym9U5Fm8QlI8hKQxjKRjxE8/fK
WodbsBvgxjiP041H6rZGZ5aAjVPkoHnPaS6R5+0ZSoP5BvPuRRkTqQYlAdE4SLbR
I7mT9j8E8yzRJldNfuzxoiJBsbgRFm22UG11sKatLNh88ch8aMdosN2oJWGKmMJw
GPrXRjhJqwIXHdQ4Q1yKaqjlSZyi5XQYVWjAjhR9xrKv8L7D65PoQeN5pGtncmKl
m7Z/lI8ABlxvTGWpoADFOSEU0kcVy3crG7+TPyjh/FbfKOVLb7VSPvBRXGRtrDsL
4oZnqOrSiwjA4tOyH2YVj/fCYfDofm5mIpdTwerb18Xkd8BBT8XxlsI9tGWeg7er
HfHwwfu2TlBOupJ/DDoKCp6HaaO5F/Sonj3TPZzoiDJq86O6mU8p/uLRIDrtBWoq
zHmY52phZdk1USQErD4dSQUs72N1oolbT/scKSiwOzQwqXbl4HcATIq0qWh/t8T2
b6NgjUcY2/W+K+LTvjqZvAbTfncNPb0l1+q8jZc1mxvY1WNRlAQi3G3CRIet4O2I
JeAouzRDW46dtpln11ZdR0uovxRKBjUaVtonL6XxFbbEyIc0i1Q3BIqToNkHgORY
TUbNYW46ulLnl7gq+fl5DCk/VErTbhiLSDYPUKsKg7DK0zf7Shs2Uxe7rk0NOghS
id+Za8hhqXF7DiZgWTGCCQUL77shvwvPjxMyR4diSrdus5mUTQ2cEH4JyPBUQ9cv
aM6O+DTzbAqB69artd52/x0jkxNMkkzjPwVrtNPTmORs5fckxBoljSk7c+OTVsrb
0/qEPOJGbp8ExN4eJa4eQE9DRoLBM/lwK0pSIlLsimHpIMtmplyVQtK3X599hAsk
6r5VVCFf2t5/3/GlrWn2vFiggnMup3NFX97m2UHDHt0vmncRlmSr2XgBqb+/NlTc
FzCKh8Ly8BkcrlCYvlBV6P9UFvQD4eugvUpLV0/BIdzkSvWlLKbUFL6RcT6kPfVF
PsQ+HUxTuvGfiSr7FMKGqTshbpzinc5m8Ne+FNp42ncY/nKVAsCZ9oihp2Z9poqr
NtoYpSRgXvG43FY1tPyg7z4tP7V7HlWSggzi0wFneqX8oXVcLNCZ5OBQ9Z2O0DNs
0qFw8aCnGs6UvSMrSv2lIxi1aYgWSu8H+BOXQWvMr7pYqZyZfBCWgtQugMmHoJe9
rOsQMCVupEc+nHclYK9akHz7+mCAFgAFWKbkzTvtlR9h4SPado8dqUNO1zBnONbr
t6p7h3BdHNNIUCQPYC095Hyb5lH6otCk+1A4euWXAr38OiKmpsPlxTsko77HJgVg
fOqblBlZsZjh6FqqZnFpJHVVerj9wVmsclg2nKUiTJrMHBA4EtVSu264oHi5Y4QU
9ip4i4543bYVhLfT48iKSpQ2+kiWYTxBqJdOl3Jh7IbBhaCZHi/mM9r8BdMn6gB9
sXU9IeLTr5s6aqz3I1v40QhNn3usqosCFSHRez54Q+3ycF2iRExqRWdkIbcslJEi
VlKjMVPpgh0YpTmwB0XIA5Qk7YzxuFC5Nojgqw3DwSmUkTK4Gc9PFXtBKeY00UsS
+PZTuscqzAlCr31yYbT3v/PchiXQdDlwrnkLulVMHiJHrE+aCi8lIlFU3exgjjiK
40hrWM3xYq/KOPVINfbog7FsFqLQlIclbcG8E+Ue5vd3vHiNMQ2NxJK43PS0nWlW
hTkI2f8TmGgCxCNoCOXEDlnX/3PtE2853s3iZ0FcvyPLF0TemSwG4DxqZkC61GC5
tkxDV40Jo+llvOgKoCnE1J/X1kplNPJrPXQ+282S4dh1Aqqfd4S8rIL4tRJTnF57
c8KG01sp8NW/ctM0haGz9Yq5vcEuC1lc9LWfSjQ6DojI5HAyWwO30mtz5ug1LI18
vZEVt68V8tKojxb4tqltm2JhWkyN/ObYXyDBmNuIqgps0aeakH8jhn/n6o/qmiSE
sicD4PiMqYJ/vbt9tZ1gkDhTCEEeA86hZuMxesG2on8KdS3HTL4DPqtVOL1F30Rh
KKwq7RUK8ujX5vwzawKap6518VS2b+/sXMbyzOD4/SPDcoSkguERMoxuInUmOrKZ
C+QCDxqJ67i1Ka0zI/Nn+K7/2+9ejxFP8+ePSA+l6+ZNS3rS+fH4wETnjHCBGowu
HrTQm6PdjSc4xhf5VQWOmqPfkoi+WAHWD3e3MbRsJDK4jDxDTEiYj7CX3omfcMHZ
KDQjuiFDQohjllfCbuuMNu6Q2IcJnNoEQH79weW+lRcHObDCtlMCM46G6TQmB3T3
dXsEpVcOxVMI2nHAXFqPuppWW65msQaKLzfRMHnx7ywPKX+ZRpAqyPDBJ6spUqeN
Spoh+dJllrgaIdiftliSeZ1Hzxsihm5eN+h8jTDjRZYzOzq5uFBVxRSrkz3/p/XI
cO+9JpYAQnuq5GH7b+HswXJcJKMbNYb/qw70xdJDKl0mFYDWGF+5C+So+cHu/DH/
TzTT81fSBnPTTP2or8VmDuIyWSQNItZJQovrscNlamOaueSKTqP6mWrTnDD7Qw3s
iZNj0H6kJPV+Q04bzyPWTTTAmi3Mdn/5tIxh7fz9c/XWATsfEdEz/iLGlZM0FeUN
cwNa5LAg4IYraRdSnPYJm8y9fGgc0USmOKNyN/eiGPenUyWp/uajVdIr4r4UxXJf
f2y7oLA+k8DuAplHf69q7rbKFakz+Z87sa6k0uyu0yZjaon+XdRaoZxfYcgQtj0V
MXoKmn2cqOKTHDNBDN+5n6RNf3RqoGbvN7djmJ7oJuvxL/YLyQ1fHgsRT8DoY3eP
lU0hph+lqHlHuPYt38I1CtVgMw74MABWqiCG5AoBnEC2d+vwJQTnBdnz6Oa4k57c
ioBKr6HpHqys1PznhutjxaRWrkRN//wB+28ysCxh85AW6wDAaV0KRBdSEIkSqFKH
Oa3pBkXOc7HxVVnLK+A/o/ypt0x6/a/4rSLQNSRPwyAovUZtaYxDXhsjrxkP2Iip
4aRvT4+MIBg4XHqEyGYRJ/9Awx6qpIQnitMdbTkyZKRFSwoH+9EUlsQ9HQx/32Pi
uUJqCzH304fyKdtQgOsJ/zvXpHYWVm1mFur7kZD4oF7h/l6LWvaZ8UYqOeLON/jN
qly1OdNJ6BBL07bEIvuIaBqqfT9hiV1x9U0to2Cj29Gr5bXCpV/XX26+cTdQ3BBw
jxk1qWoLZPeYoX67PUDTSryf/yDLg38xXlyu+f1pHWyEoY9NRmQfr3KAD3ABp6KQ
jpXyQW08rM2heDbkWVSFQfM7mbQQEnku8534+f9ToNbs72Rjvp/PLoz3VANIeDqX
CVMs6JP2tTuGylJCG2yW46uU4Blh2w7jRh2azGofE5qY11FkykDNlWGvMes+xcsu
mVGm8iStugz8vY0ivgWeIdntafCgl6mmfv8VnxKkCh/m4M20ZSb/54MTNDSHzck5
tt1ueNweuqIFfqmt5PP4zU8ZcEJmzO65ZNY/MyrHfIKaPrNGGilzznq88OfeEiYZ
dKbbNcz2MqX+fHSjs+QfoDzuky9tXbrGvm2u3OCdzE9LF4HfytlIsJGlgZYMY04y
uCqUBV3rQvxwfc+PipLqd9/ylXdXTm0t3k6woqSKMtrdVwj0uL2RG681CWIf/2jD
ZpwB+XYBTaG7cTeiNjNZGsVAzLGWbVKuIrxbMmBlFbmHd+ye50CDeQfCkLdChhJ8
TLnSw6TloELm344gtsVcy+tEIjKH1F7nW/Pg1ci6gWTSq13yMzgIgua1BBhNjmsU
FRvMNHcu24pe1Y4nrcZxUZmpMbuxoBijekGu3pt38NcjFptLvP8bD1AGPeV7xQy0
uEfp8LP6k+bc5BfekAOXq32yQmvSCu69PMkIqworRvJjnyzYXx733TTQ3tA53RnX
NHBVT7L5k35RwIXxg44R1p2R3ISbDgciz85CxUQGiYUNq0nEvf3yri/LiD0cq+xG
d24qQZvtudLKIgPxF9J6SqzhoLJX3skDhAMxrcps9GMlQ6csR6F1OxjoXjjLhBVy
d1Lr98weNDetATzYDGIxrHevoTRlx9hF0dHlXabWHuC+j122XjrpoAgo7ZukV4jk
pinnSx/3omYlAewovGCiu75dfsLXBI18N8T6KmPPSJAVANANkj8mKo3iA01LB2W7
z7wNHW1OnrQd3OIPJ8C41SFW/uIxIDN0Lgg70C261rQnq/tpynZ7xEfesC1bU4RY
YSZmzKAnvWSBXUDubw1ZEjolkIQSc5T6/nK7uMT0hfJINBwGiCGMUiwIpezcuoBi
r+nffsQpnXOf9fde0zXDIcQ0b+0o49suew4RwYZ4YmsUOfe44tH8frUzi/5HmwmL
bSarDmhHZRqqDHx83BPq12NF9094gmcz9gwo56y8ANplciEi4t+LpdcdGdX6OIFu
fOicTQ+GbpU8pQEjbtBajw9c1V0wxrZRTPp0/+zF33ssbskaPmMdeyE5TvSZoS3U
Vp3zfT5NvdT1Rn+lqxERPXhce6xlPsIF4wqnn+tAUReTRtF9xkcKXz2xf2REzBQs
29juKxlCl9AYHLPw6ZYk+LMnn8bNMRNtipRHg11ZgZta1nz4Zdk2SZMcV4ns+xCD
G1ZK7zXloTontvrvnPGlrG9WUVmH9yMVhCwuOUQ2orvWtQHR3TTA0RLcsZ9sRVly
o4vMRRGjOQ3hmnu5QGVXZJdKi2tUCYZedrW/71FoksaqA/AvXkho4cbvD+o43r9d
ZkNWax0eRRWoo7Kzqj24dTq4bhnj+kFeQomTy0pOC+uFBIu7vosz6LwwTuxBiDZl
jjRHtNhlgUjRtzyLaKbr5FrwIRushqVBLexO9JiYDU04VMjz6T3CkTewqLEH8TGt
PWl51pcchbnKp9oG1k0S8VZJ83Df0lmBS8Ooh/iz0zio1uBkiwGk4fgBLr1foX14
ibcocHmV5VrriGRic4SX5uVRd9uwb+dVjnFj4CQLuv9xSrXoqg3Ziw6oPPjVht61
4GolF5hudh0/HBHghyEaSzbmuIOhJWxs2OM2gc25hpVxhKGdwlYlyhwN2NhzqMc2
4/8UZk0wb0995vm9wsJS/J5AVEML+Iy5hbJTNxmwMeFuj5k47PJEjfCZIg/y/M4y
1qCw8oMo5xhpczuXGdXy3a2vMnA1xzuqIN0gaA2/PWtgSTys5QERiRMMLKj42URv
JCEWd2bOeAKKMnUIcu8HZamuxPpaHih8r1L1NXjQggVA20F8CQUO5NVBQ7c6pLWa
MjdgXW7NMSBuyRZ4TqXse4J0DcvThzSLmWqjCzo+8qF2c+gKxdqVuCl/CfyHog+W
ciqAMSWzswhYSXSOtFv+zVmiNnhA1wrAL7zWQN0xp2LyC+iJV1z6u1vHmqBLrfZ7
3VwW7koYNsL9/ytvDpxROz4bG286LMdTfzZmL6xtfCzDQ3PiBoBLFBcgw4kK0Owt
eVFHGd43r0v1VdQxuD9yWoWF+gOcIVrwj0TzPVZMydzjxoASmAXt/jZ1/kqxc4m4
zMgK58yaceAQD967f4jdHsLFcXcacOmHdS4HsLmaa9CQO0Nmq4hvcsMDL7rrwfOW
NV95DzHzNbo3q5Qz9hF/+yicZiUbsondq/nG+9bcgFjcgRGLqdDiBnyFLTJzpn0j
D8I6HOrZgykshkeURcLDv9THtkXbMmgnqdSvopj8qMRH/EVI9ntJwDggFTl8tWzt
L60V0ltb2ndWBhZy9ESlsIfWzqBIUc/f45ALpPbwHJXeaHlUgoZoCHNtzL8/SJgb
pfO15yWEPaz72zz+MtXoH6jK0rKEScMYCUWNNDZGtR+G8fnNSYeijKNJj4lsQq5J
B0dKO97y7diTGBnF5Ezgj6UlTKF9mY8TR5VVPC2jckveAljHLa4d5BN27vF4AauG
IkFX62PSYBOQThD7N02aP/wtmIUtrHx3/hssWUc63kLQ2Q1p7S7z3Mg28Jqph2xb
UyYjXr9cFWulorCVY006togk8qOH+4fVW0DLvlRzWBTxFyEDPjduXjLsz01hI//p
pw+QY+Z+J7cHfx7tCQk4SyS5PAg3VN4adD/cJQF8IvC8tvlB6AcuDCxAWAFxVeOL
d8bCQEPmgufHrDxJQChu63TkUiywihzpbgNMmctbuwQp3Dxhhhki9ATwfjdYuSMD
ciqK3hxPghYpmQ7+DpouZPdF7PbfU9jAqOqef0QVp6QQ49CkV0pk4F5kdsOSdC4H
Q+jia59DYx1ORrMlPwvQJ+xwPzbMifMO9JswNikVB3lxN0Ybm6lRg41UlllCmwbe
jB3ndJvjeA3YaFPb7ck1EL3m0b3N0VqUJ1b3WkuPDKKwns1W1SPKH3O0U5fmWTRO
b9aVSqFM4MqfcvNnEGAtgQ77vkIpXsWWZI33zSoIeArt4pNZVeiHWNYBpGMSKpVu
Sh3s5i2T/LbqiamWb9PyFi8iwntUQk2REkNMiVzLldnwjjXnvcSyQ5McCe/Kx+wD
2QSv34UC9Al77c+185gB2eS6cpIrMwJy3Sosip5PPgTG+QGVaWLIZ6fqd1wMfpEf
dAEqJCRduw9y6AXPFM/Mos2lt4hwUaAXdBFCJyIoRrtN4+7Cr96dsydGkLuFZTX7
xMoKDUSpZFSqGuQD92+a5JRc57wVgRIcX+RMcI5bkDeaMD9kDNVbcl5eDlNCgISM
yNMqR0Sm317m5tepgckYQDqinIxkI06zU0Zd87xlsMt/OVefT3HwL5lqRzbzU8y/
ykduei1Fwh/iEKJDwFPnbYIVHmPwNIFRyGnqzsZyIiUQG+BogbLv0S/v9h3tanVJ
CrVJgiiLZ6+h492WrM6N2M6sgdh4VBKlQBS1X/g8Uy1G0HsgWOzxSjNx5LOJ9WNc
yDKsrFvngaIR9USLr8+ia/JG8oTINj9pM8ln8jNHmybIrlyB+dxyzUEX37/IMsa9
TMNKlQ8QmflrtOXl1gxOjogHI+w/T9SLR2xuupRmXeU//MTbAw1lhfLgBR2SFz7v
jEdg4joopvM8t9BtwyvFAH/HReeYyR4XJSjb09GPByin2sspYYYrn3UQWcJB/1JL
MZO9lZ/Hl7lCUal9OrWqOstwjTKuw6fXtb8dhuIGocoWVMkPg17M30/w6XhjNfqF
eeSmqXzSKY0LZwoOISUG92+RbSg4T+PTf87sBYpQMAGlPQUaQ4BNrMkKGRgumuv6
GanhYRGhXyyECcvlHMH0U3u2wp8xisuFWbMS0Vt0okYgY/O/rINvm2YktjnZ7UvB
Yn4RNJHoIQiL7J4YgdXAF5WsxDG4KRpHlCeTPtJVOfFAMxoFtUSsnx1UPmSIDNE2
MKnDuv8sStvOYDBgZwxHidLO8dijK+EI1Ntx+fzb6tdfNDn95APAp0PhEbJ8HqzH
xSp9fq90vdeqWrmLSq3eDb6Fxe2gM9KHMFqkN7mdxW33PH7qZbdQJPANwMRfxriP
a2EBHlffCkxtjAwqOthDHUQhtZxX1YXKDNNW+VEiDAq6YHy/M2Ji1nmBMEj2F3dn
HHLsx43dQU4mETqexJojHaDQIG40LsrcjZ8egFSUy8y999ia0Js4kA5yx/IQxIvd
DeslrijAVo/yRLaKddleryRprz5HFiagCBfJ9+qwDB6ZsleFxGM1yamvoBGORiR9
c3gwOnqe8ZNiMKXbrPs3WvieQOspLJRV+eda8e4nuPAdxFZCveajaQjhMpdGK9l3
cbLLgcCjnLaqocpSH2MzIhoA0DdArhtcH19S7JtlJNQMXecF1eTt0u+2ZV3yReZL
jEHBxTJYGXtKiRTm5yYRSYl7o+X9pnnikBlL6px5S7W0wMjCJzp0r0qTlh2TPWgH
ygBUeju+txcfDGH13DQ4r3i/dvK2uJna1xijFvSfgb7d924ISKIgoJPLXkJ8pub3
FnmbL8jDv3KeUqiwCHL+vb4ZDLBj8BsammWvsqW+ecx9kMOvI11srgXbSKS7Z5+V
VRewPL8M1/BeSsJzhg/cbvTrO7PQGc39kG8u90d6NqG6sTrN7gZRyu7EqejXgpaH
0aYXRVJXyAt//RO7UZ1hGcV3xnwlmCfQpszsZqDt76CwNhnyANtQl/Jua1anR+gx
k/LfQqjyTF9mNvEyVGmhqK9ZrAqGUZTgBy6bZJQ6KCh0bc+USFQAULlQe2pdk9do
NcfVHDXTt+CzUIEvphyAc78IWeaY2kThzEop5ZjuHnzYAxLAkYXVhu1wpspiGgGM
7UWuNwOIPk3LhZVvwKx347Fh8sXHZWP/15VfJmGtaG9iNUFeDTqoNeIlv6GrCZMJ
QxkRS1KA7M+sqDOcdMjTNxyXHopaVH8JO8kBM33RAXqCNnoqmY0LZUyUYATrjdSi
AUWu4QTU1Ch0UaIXIfaqwjhcM26lNTSgVz9jWIR0m7yfaa6XWxxYQSqti0zeeaPn
pqmm0VShmLO0xM6yZ8fh+QMqZU9xojxhBeCDIuCI9qK3JN7rg3hpQ/7OiSxziZNM
yaLGrJJT6Non5d71ZCqE2ND9iJM3QbJ9pH+G/ODqFFuj31Zwjmr2YVPeXHvxC9Aw
TuONiARHWBzFst6GqdGTpNztKhY00JeEsiIbmunZnHakHsIvEgnG1ezdRJQgj3PJ
k++nOzw2mI1hpmPgSqK9BORg748Bo3eesiqQtv7uD9YT1flBb1iGhzMC03F0TOn6
Yv4XLfSnLbIuaZl2GQlx3dRg+UDnvoUDDd5hoQxNPtsxH6/z8INVxKc7JcJPUrj8
FJ/Kp4Ixz27veISuE2F61GYbRcN/NowaEykXZ4if5bHIbV01xHcgWvfxXaD8A0s/
Rog5t+bua9vupC0bs5uFj4wItXyakXPYHztWGXT8jKaMn/YOi32eRmEWD4a35V6A
ZXf1QCe8ckB0kuYLiRUdPu0aLB0UrDXeGGvUDH2JtUKOMTylkhb2sepNLnJkM42q
DZiYUHIMa2Fp9GvS8M//2bRnjJa8lW3SqIbCPE7EvEWGTrGF5S/BXRZL0w276ttD
66Kaw9l61YgESc/aDN+eUg3RUam4BSpkfDrabDD2Sbo4Bg8yjkhzfR58E+SIlk/3
3VssWNQbos6vnDvvFipVWumdCMwfrpP2skl25p5+HfpzOe0ikNnkNPwcMsgSqoXs
GniyNrK0dsBoV52bFkfJ8VNEvFOTwRZj0Ep+Zy29aUl5pC73CtWib/TFSTaLNUjk
VuJymuAsS9C53ze7dD010adbkYNgBXssZsqiHCRFPcg541AODrNw6K2QkhS7O9Y7
2MAkUSnP2RKU9XynLsomX1aE9jpGYcR9VnHQYnqdPX39W6GWMq1P5A0Tvd+WUIxB
C2Y4Z6/CfxQPdXcKgeCxGBO/RxMEfLYcy/TImMm0h0GLIUk1DRUvSpm4N46o7qwU
CD4XPlGrscSzRfED/VkIKzN9jHrFNdQjHq/Oap4BKrPmyXl4ZLh8b1zQOsaLdZeD
eVe6EzlBBHA0bNJl36IXRpBZPKqj/jY9nM8/bHi57z23NywLBas99DmC/C536gjz
kiumBYsZrdj9tEo7VhWBuIPcKeK9w7bIq0V7/vzwIH2uCPBMLXdBwXy5p3P34gvJ
XJDM7QZLw6V1PWlLxfYeenuHR8VVbYuUKeqidxjJ4zyZLsIhOY0RMavCVCypAzzv
sLrOdNeQjdotthAptZ7rQu7SLgsQ0ex4MToixa8YH5lzSKxT+A3E8q30nlEmMgRo
AaDbs8yekbyd2jy1kQrWfkCWdBDdAgOyr4uW4CqWNvEoklCWb65k7x/WxpzyqA/l
TQVh8xbpnuBKp4YK9VR2NJQPDncfiX6Tuv2yZTMuaMoffQpU0NehEojFIZPFpYIl
kNeu2BpXhVbG2iOpd5TYxi5Bgrr7+6JAuh8FwNVqNEifgodIUpg3pkua4ZamiYVj
1+58k7V2V5TdZxHAbCxZ/x1c6QpEVyFdsNW16fHk1iLS7lMhB3qaXztww02QNsws
wt1hrkKYSY3diYG9kreNQNwSpyjVqbcDzViqnPLFqBIQEAZHGhF7Y68uYS8g1Xal
nAj4UwrWnKHMu+zAHhWxqY4GYR4IWcekfSffHhuJbepBM0CWC8WD/RwzzBc3uRiT
GXDgohceP6q2YBwunYmE7KHGn+FdxtsCteq1JwuMAXtBx2SVRAeTP+MxrfM+uxU9
4w0NsNehoHu1KhxYTgmL8degtWD1fkK5BubBoxDXYqmFYbtXt43SHe+vkytR9QFd
WEEDKNi6P8BTcNCi8W3d5zlK9rYIx06gGwQnhRxR0GyFiFL3uLnd60HaWF6pdgZB
qv6g/wehT/KG+FsizlW5XJg3PrrEReXrd2BPXSNT6A+m9igIZwC0qLjdB8xmxGl/
PbeAJUFZunFwMH3ibMIniEuzS4ktwvz9wLt+QxPXoJkURr7TXwc5LQUgW1kpJr5B
j3255DaeFl998U1HlbfgT3zeNcarpdd9TgfdW084068O28kxS8rfACCb4+GSGCsl
vRJMXJK0oRzCDWjl6Lck5FaUW0OPAwhHlYMlRJrIkA9DQv+QPCGoma9jI9RMNcCg
AjeTDLnjmiaR9c8B+WE33stdIGrGsL59694fnk7L/SMhlsHbcINlk/Z+v17v8UQT
NrdgXNhNiwvKJZJX9abrHZGKVfchOD227Az9HxxqVtfpDrWUhQTTTsdAmz8suqUz
JcbXgpGB+w8SVHkchsL+DB59Aya1qgVmx2ZrwR8t9qpuJnloD5avanSXc2xeFqbt
6NoXQi3Xobk/6QfZQdF/j7MMzCUMmx/675MG7Ayiz78cmdhY4ne56fMIwThTGBF1
l/E1mICjFY1wrckjk5xRFakUBKZwd5P3qSFbkSEnGZfVlI15mLuh6XZ4Lh2Dnv+e
Rc6uyWCZ7LoVLp/8yAz7w313Q6aW5iz06FDloGZNP0jcHDG0KYtXoN2ORFoRtEtX
JSTUGk/xrkbIFaamlDdKiQvWMGFvT3dm3oPiPyPcD6IIIspH46nQGZiXgjJIt6kW
d8qlxkEx5lbP2FFpkAJtavSLdISeMZOPOhxjv8l3YT/s6Wd5fmanpve7G5IWR6ES
AIq8+SoemUxeoQTKywvhacJZ8V2c8dQbpZsEsTktNf1Pa9EoJb8ywJjPQXAkmTif
JvUJC0pG+HU+nPuGNmKBTAIY0PWVme5EJtuNFLHVm8OqEs3WPuVgf4sNI9+hSJNb
bs8R9JkBm/o0oVFOHXuBWAFa+TPQB76DEzLKOPCVrzxTagJkFi5MnMf3raMzgaCy
TqCA9LHWYvhJaBe415jOeJhvJ3aZJCwq7a1iS/UY7IYK0KUJkuCkrL2zZOl8aQui
YgV3ICmsm25SQL+JqHRjGlAiGuSY2KKelMpHyDCW11Ms/DVmLQAnrDCWHix9eQr6
WAyFh1Y21WOqzxkV/H7SvJ7au+hIdagJA19aLBcNggwxrBQ/ZNzBsPsyPrJet38h
4AijnpKQJrmgvuGJvyCkM4xUt0jSk81e/iGGaHF8au5ZvScEWCS9z4KXKn62qQx3
o5D9siyXBH43tJUyhGc7W+XzcWqyS1kQY6KuOBY4A1A4q7MsnlY2xAR7fBEk8QFP
/iMc98z28Uc1aufTihIx/26WonRN5JqOWbFMDmXQXyRhIJBWav4cmHQ2UK3+qNZW
5K9yZkqrhrRdDD5G30ICc5xqTJoNH8RhnaQzvI9e7fyYbCrE/IBcnVoANjocIH6P
oHiAYhsSB/YxZ67mFPXP66Gpp3ZDWX5k5NWGVQvoZbuP917iBKjcff1Dpt2wuMFg
1bZ2sIXeg0uIliwHCA6dwdhhuWpdXWZhWb7RJZPZK2heow/PzvvHgjFpduH08wCB
i37wPjin7tXuFsDPmPzTcmwMGAgCJWvvtVgzwDH2XZWMoky4comqNkj/3oGiWskI
+QAro5gFVU9K3bmyPd3wHZMR+dM/wp24meBs3PQ5zsTT3el7B/x/4Q91h+GLCEHu
48WGo/oXUfB9hdyYeXvMVksUU+zt7tpWE1Bi3+lFLYSAiPRKZ6eZ61t3mFHPQ3A8
I75GdBwtlVueKzft5TYb/ILWeZkt3dc4XvXLNmtgsFA404H59PtB2Xb73ga9SZk/
JCcZkv4y24kn86jJoSl9/gljSEGYQfhHuG+mZ+JhaShKuqs7LsO/2qt7d9dfWiHJ
oGAslp9QvyOc2a/XxiVplyUqbbwZ7vA9FWxaXX23qgij0ghIm3J9EZRrxD6t/YIt
vQ/+ojci7iysiN5MjcY3u98R+nozcZk1JOHtPYDmw63mwKchHMpPbeNnLFA02OVO
oXdHpuVoY/dbjZ0679qE9mGP8r/8lNa6oiQpKHw8LGfrJ/byFffEdtJeIaDKx6oP
W22MU9OoTM1/03qsUDJOeuLyOI9o4qQH/pDnrxiIW/Uw2Dqnp2wBD37nJ1OJYBBp
r40opkyClYQX4ei8ePkh2mNEKnad7mLFcPSf3exPIfeY+VVybNeE12/cP25n4zOz
5ImnY2DzskTV23AHKUH3UV4L0hW8OomSkTGAZbZJKuCEQjELbLALmNHNxsC3Gdv8
HCeSm0mJnQUsxyAVy0bmm1pH9/xCM6C+PqSIuqN4c4ipBzsBLbAkwWAbZpuvrzwW
FlMRG2lUCtS8LRg8csC3XTRkonDba0qIE2pZlW2XOCPOP2lIm6g9h6S6LogT564S
1tseRjUWWU8byl4uWWr69MD1eeX0ayEjkQBKV/eZ1lcvjxSxRdNtPW1JNFSAPIH2
KNjtRNJKeNDk7Lf1/YskiTJaDymYFO2FBrEt+FhyLh71NvgCXUARUdakNQnfIGVv
P8Pn0SRnlfQVo0MrfOPRDm4sxivlBNNNtU9Q3kWtlL5w3v7p8HSGCqv4Q0S+rMKv
kVYY1/F2cZmHtaBb1SOfoc9/m1vVBIRDViBc56hFe2q+skqf5EfM28Sk/0opKtnp
q4YqK/gS2MHaDv9uGSOk2jKsLv+sWHTpHkLwQeq4vnFoyOIo/fXSiMLUpgst8TYt
Jftri5da5pXIRvWsW07PeQqHf881570sWa2L1l0/CClBW+9FzX44Kn1UztvQ5vaj
7rIZyCnNzAdSXipekDIS8ts+2rqZ32cZoEUiL3cbI2VgXV1oiWfm4dO79Ol4uN18
4vODvliyF917QuEV6m239DSWebWDHuRrcfihGS9gJUXee5iyEOAK/ltrQVFkVUo4
Jb79fFMj1HQxo2019prjM8ssMn0Njw55RA+YjQjAYEY4Njh7PhraXA0t18Q+iN/+
2zQGDTPss48hDWQ/YXfDvOlUWRu4Y6M0TRyRjCMNVYOupNqcCguOkjAzXKjiRFs8
Bpaag2A9wOcpOcQXbjVuLpvSWbje56kcWt4yEiaaoNo38HW0bVK0n7HVVCicRhpx
KNcO0GFSDmhqDc5HM3fEBNKyqiGfnbmdpDN6SW9FjY0+eMRHl+pIgvGuhCM+02oE
Lv2qmgMXfCZClO78CHevNFzxie8F+71IwJ5fdHrF44zGYzVnilK4hPzwNkAPn76P
Zh+YQ+VKFnb80iQHglGl8kEOGLoOwKH+EqMvET6aWL5bZu4pcLx9msQ5Vh9B5kYb
4gwrVf5/Bhjxj+/b2yove73N20Aw+/mgja3rOHsOq9ia8w5sdzWPEgJWA5hl7Ysi
650YpjZpdsd/VXIdwq8NQYpwPK/ryj6scwiNbTW/LCshk3oBcGJuXDDBe0PIF6QQ
T6RYNI/VcQ23BGJSjGs+oJL1IvBdW0kmvPdaOqHPNjwwZXpWt8Ac/0MKgpeN3SEp
6ZcpVbk2ak2U3/0BkB8CwgLx2awsJWXl4mYEaEPbsQrDXDfpYSianYMGd82/uAnF
PMeNDm2OI//IrdrT1jp85gnt1C1uYchxfrtbTckWUMu+RhK/KZyj2GWKdrN5jNlR
NRN+8M+47iZU/MvY8nIQMCnqlHwdDtUlQCcrLsxE9mKd2LBBGNtfFFHU4TRt3pY5
L/5X8/lGA7S3ejgTGj4vfWkcnrR3AvMfB2c6IPSYT0rkOTElkjymfAgsmkYMHqSS
eewZml4igtQ1IluZ03q0CGpFW9Vg58fBRqbFPNubi0+m8QI9wRIx/u+HDiakcvJ8
q7oRAQEUjlvTDeyiFsL9RCC5HOcwPVRMJHg6zvKztvwNXSmIgkBmDOl8JdgA/5pk
dhqlGPKwrr1qvMNRJHT9LuHgFm67k703RqMsPJsk5l3xA2NyWaC7cj0/gYbYKFsM
d+8jgrorwyZAJLVYOIp1BNlJ8rEZ/I7voeBI+Fc1Ll9HvL3s2jrl5to7PkgNOpsQ
/3+fu7zswc58ywy2mJ+p7/2f1Y8zeUjavAMdujDiQkmb7BiN9TSNneXoEfkOkA2T
F8xXOFg3QnSw7PbRTaG7nuztUKNw+gTlKvt1Q5KFBgsC9GJ3FcnUS99/Lezcn4bP
c2Z98MCihNpCc9X7ahI1Pzxaoqi2vIuD3y/PAijL8DibwXyhbfGhZKIajR6pqPvV
kJWkXAzLjgoEe+EGK3+dMheQnH1rJCYLqoHPW85aYPc77RA1KmKZGUtoSKpBOA6R
thVl6voWf5H1M7mDafatoE6Sb33Q8zh6TXiTJNh/iM5+s2MMVGlSagN8A3KX0USA
7xQZ3a3pQmV6mUnj6MRn1ipbFMTM21sFbPrBCJsj99ObF1kQIsAjELLixFR/vKnT
itFO13sRCWdtgqPrkQgarPIZEQgpkmo0jRUMkrOCMtK4Kq163ibG4mEN+pNLMUyz
o2xH6vaXAlIcxm2SpvtGSHy5VLRUa+gqUveZ7tFoInlYqIWYj8eoHuTeM/LJyG4n
bCA3r7Cv/1SUF4b9emHQ2w8BcLmmMvXG+NE3qu9txcmat0NpKaRUi2Jp5WVMcU36
vDOMY9TEWUmzx4a0tfWEY+9rZNYg+9Z4xXyGkqIYUZSROuIpPQrX90+Ux+sF8krA
Izx2hAfCb8GuD7puHTvwPXA7U/yPLmETmDy0hB+f4joO8VM1i6P2o8YkUKvHzywx
5hX+Fk7MG/6U/qG+D19gMgKDmRBMMOjpxG+PXqTXdshjfCqWltp0d6quno4+Hinp
PDjktoSEf2ZZA+7a0hzK5G0Rh69Qqpfmk3TjOSvKb8rSqEfuzs7BBtyeFPrGHO7N
FTsYcAA9uee2oxuNtPVBzpBPbmYYUJpfCEYKgT8rwMq0TgW7P+Wn250RhOK6mHhZ
jVPtV4t3iYb6hAmnorAoiN0CrLL7G3OXeNgX7ZXk8eJX1ZtyyTGqlZKQJ175cXx3
YrBS/jlpqfk5s2IFLwTtG0FZrwmfRM3N90gotHwIabdBpAQHx7ePg1BCOzYo3yDK
XpfnjxT6Pnglh4DV5tXePQGWb4F18bsNppuYsQxLdeB0ojaLSI1oxsm0N73e2+bf
mibztoKuvTUqKjbQh6d5X20cMDwvHguWo4DpTx2/+oNyrmeALPxmqX1qNUmwrwJk
RX70/At2yWLyUVmBzx1gMQdgcc269zdVIkIVuI/lg4HsjoKS1KGTwKBWZs7ssyKX
E/O73ex0t2TmOfrAzrZqs5o1J6Xh0akeKKsGIQ4+sicsnDxutsG12GoQgfQojK92
PgBi5eW4rUjApmdkj1HEpwGN5qGg68x9nMHNJJzMDPgvK5lNiyN1WkUAf0Otyq+p
jHZ7LjDWb7zMVd4etvnnIC9tHISvXGmtwr99ve/58P77fjpyx+2BPQIqNzekWb53
h89DRxTnBwaYKx6VV7BqRmXiUfwZ22XneBE3n9p4+a7MQpBxb7Tta/q1J20tsHej
gOIg++5jyBHzTIcoKtpYcSnSwcaU3rkFDefx+E2OYS0B7DzRtfg/iYxeI3xvy160
MpbnT+vM4uBCwDUOvHXWiNDr61piYPn4nhqldD5ot7uBfRo8fQukbn43Vm2nSD4u
r+EJLqkeQoO3n3mvLy6J4MUqS9HpiUbS/TUFU8rbsVzMBQgOlVR5bHn2KzeHTDp0
TN9aMxOQzU4F+iui4cPpY2e0xIj4EeqA/9d6HwwfODuZH2ST8O+KkLnJEML2XUnt
GjXKPU3ZlcOKA9M3ehjGhtYGIf69rMdO+x+Pos428c5Lo6gYECEplYEeCqM7FXme
ojthzDYVcWARPXSzNm2k/DSBKaECWL/h0YXSTmAh8iLdZbO7PJErHcZwANCTZDwb
V5KNsFq9aNLiNWJUAqIO5St6N0Hf89x244Qrox03EIhjsp9L6lYeHpCvSR7eUfRZ
XScuCSO8Jhg2vRMLPbAv0+WFjP8hohjWrUA3QBqP7dC667ik2iw4B9znBNrLx8+z
W777psp9YnsMypjhCE7Hex4B/D8V/Lw/1ZhB1RelQkGbjik6NLWHY/T1wDfss+ws
BtJGmbD+SF4m2kl/AOsdQtSNYBWmoKKMF1Q77+LLBtMsH+BnvFs6hYRmr8m6onK6
133RvY6auzlWTFQqbqQaJQyF8steIxPC2YH6Ahzck/j1HNfMij0IuU4yqSt1yEuQ
+6QSIsxjiN47kha3WpG6vCaKKXlpCnOen0ef2oNr54Yg62LSlxTfywu5ADdv6uxe
n06JQhw0rebA2VlS89UEeLxqSVOhmcH1OXTlEhWrEnuGwdvxROtkB3sn83H+taQZ
F73Ax02u8Xoz28UwG0hjMkX0+1YApLk8Y6B71BeFxmsfT3p3zHPd01Y9kZC2a2zd
QEzOx6j7YI783q1r4IXycRqkdBVgwZwUykGScdf3v1ORDz61rZAVdzGcv4Pn/Gyg
D5rQ9KqpP6IOLub0aThGqtzj6CwgnK2Y4IEjoNS7hwnG6JJVqfshEblMQUsFUuy5
5j/ErZAWfFUNrWyLWMHjDqjCpQZl0H2tcfyfMkOHMo5AqihkNbcuyz6s5jdIOmVd
/hOB5VnMMGnpBIKj8gTHcbYnqZ1uGbQqMrgDs0MBA2nCTkpEsnJMKQx6DOdRsCVO
WHgPn6mmQ48sYjBYPNu3FxqjJyf5XmxfsxfArrrhBeEc7PE2f+ufGbdX/ZCsIbLp
YE7023fZiveHVHSe9/2CP7U9uxJaMQsLTfCjoeTqX1vgjhksrnYKbWSLPzuM4zHq
sHhvBGinrm45yqecEw7nHANxKGL5sLOgBHmnwwxnhaMBj0EgB9vdIwAQnSZp9UC/
8tMVSEzUe9brko0i3pDXHQZowzYv53BqgqwMcKB4FZgEPdO5bogXY4ARJqQq4dUT
NLc3k0Xv6+yQCqatcQkVvUlKGq9pYznLRNSp1VhWmCtzqFfMpgfNuZklU4q1TXAf
4UemVWV0/pep36ests8UF6xrAdM776htDM614NgDhYVnKWnWkH5d7V6TvKEmrgNZ
1DbHXSX+srT3mPkHJ0BGgRxabd+A+3zw6Tg3i+9xZkS87G8esZIHNZpcEyRdb+cy
fGBMe9E/73wofhM3XiPtEG/s3ToRrW7sMb3o+cgE8L0cH5YXvdJxAa+F8Q0JkOQh
htG37LktyhrJEU/uCzBFeZC9EOmQTnxxwapxDC4WoXcsNmLdlX7z3onkDzjNOuWa
iBJCuVWmrxVAoD4JbQcOnPHGEVfZcHvbDc/eouUpvrSN9R3d+YvsbDaDglhBNyq1
X94P1v1O1gCMehEIY715w8YHEDMNBCQPMtrNaEB3UiPg17xRIBXDOUp8M00DbC3Z
3uGOeedAmM+X8DmD8IpBVlDhb5RewRpaeGnw5FukUYoTAZBeOchhyotHq5bww9u7
pUx5KtLBMHmzWQqmjOadqDDnVkgFKhcmAB/vmX1EvmqHj/k4rKGM1IzriQlMbcjf
KLgXdueUL4cxyaGBuqTfuJ2kwfyQVtFc3MhZ+vPiRGWplO78RCMCdsIuftt4z+Bn
8DP8EpP6/ernDfgKtoxcl1VvtPdbeBpLkpv5ERt+1PzKBI0HmJjSpHbBOmgM9jGz
pUv8kVDICuGsxHuLKZeGezjZRc6EYHwjayErB12W0SXd3rNUIoDqqzI7q28Yu+2W
4Ilw0rkab96IM02g0tBNZbItaqH8ebXrEYPmljub/HW0lh4mCKaHFGRZyC+EdglT
/P2kIhK6FS96qaO/HqJF0dQ+gGEUJhtcdTgDtsHQcmKCFVB+IUkvWvDX2w10YYtW
fexUAsquvxzTKGo6KLmJR4RQcmaUNy+w8sc8dl6HcfKfQZ21u6j3qnBOUZSHiqNN
s1cynTqaQw3jbwgpqLJJLdkoTJHt52fZl0ia+VeW8XBreLZpsl/sOn7jIoMx/Htr
j4SP3RBwgpe5zACxTgAxu3mUiz+LnZh7V8yUXX6hRsaL4eXbApJwlPdUsaqpAzSI
6SamrnmXZVyK4VMyLyOYk7IAFEN99AhLvnI6MbKsO2lDnv4L8hMMqu/MezZ894wa
Kkr3P15L43dPdebTLx7HAWkUmg2UUOv5UeDcJecpVvHz3cHbH24QWQDPnkhQ3M7/
P5gkPdRdePn75koLM1FDaAZRAdAKh23vTY24Ax44tj8Y9XXMovnQg50EK4BnzsE4
KdULPJOLeCdTdkNu5cQvpSB9V9sEYMbQQnEX24N9dOD2sPBNVzmQ1PsBH2g5FghB
nPOWkEK3/9Vx3rRlq7YPBI8etQW/LeDCjSJODsTIntfGL8x4i7GIJeRGHBdmbmhv
rG4Xg8QruM4AgBoZuMqYOUXBIYhBPA0IEYlyB//1+uJ+I7wwH3bKAtYCKsqYCCZM
vzD8Lt0iglX1L2xYCK0d807VUvq3cRoE3+bUIy4vTVHp6jmtvU6aqmoYZ8/iH6gd
X/Wd1BBXaIdYIt7xuwzMrGOLWc6Xnh20A0EnVIiEFkDvDZkBIId/gGr3bmUWjTWs
g1OMK5QrB05G84/fsGy+p5SEnV8+MuZOjG8BKTqsva3p02/efa65uUiEo47uIItE
rHYobwMpfNbUc/vB/zuHhQ4g1mzWzdIPqxhUDuUEOWaFwL4hLXgbq05fIXNIMZzC
D+FG4RJeiuKtQJspETym5Kr1jXXkt/iF6cZNvZ0Y2MNYUT0g4ij5r60CVxvh5MT0
pA7P/XGi1MIGdbyLugBhYbMFMGfMa6Q3VcckpMt16CFE+UofBvcefclyiOLFSrO+
28D3ztiEqxD1jxEnPoRnrUMRXDJ8uq8VSB2zZhYSIM7zGrbhgsOR6byv8D3Rhnar
arU3uHYx1H0y5hcvMKNd40f4oA86/A/0mJXcsUxPKNNewYOcTq9G4Y/DHIDe5Q+2
nyJO+fJt3iPlgA2w+OS3RTHC+jlCln7ky7W2f7jthIt62HtEMzmicFa0+qQIXS9v
FemLHGteM07NrbpREIlISAv6rLo+FIdoWh9IwTmN8eX8VeC9hOoqI+4gXOcPubQA
N8y8sMoobJCO7mJT1dFq+RejDqU5wyfRNsRhz/oxc1ZvkNVWwZTZvhKKvkrgRSuY
O39NbPcJv77BXNAuHLjcBFc+1meActJXWhy0E2oqVXIp14ZckI3luSgANeGRMyT9
Cl3RtAypreid4jusWO1mV4Ps9PqIQeabGTJFTjFJglPBmbhrjOBVOO3sOK9cLVGn
vaIzDE5YVhzU1a+kS5CPh878aH3Pgugwzh0fPXkG1MBvbvq3SWOlJMQrfblpWxug
ghg+KGFN4jLRUcqBsJwnRutGaHwXVyCw0kDH6qLXXrlYeahfkkKExc/2slUppKKh
58pfduCd/J62SHNmatp2xN89JbciHAPBByFn0/j7fCh3edy90iWhxsp72qw8NmbX
IL+LWaMhscn2yyS8IkMrbrH42SEwhQir96k/wg1jTD9wub1AoQV2fV70CHLRh7i2
BebTXh7XAD/y5dihd/WiPpMIMfAfxsz5LeE9Fod3b3GQD2r5Gg2g8n3i7NMPLF7K
0/2tddX4rAPKS0IwwM2Wx3ANcdhKyGO1XWlf+ViQFrvwcwvlUfBj2qXV6gyU43P6
k48IV2gEAKVBMKtASND3XjOxFIZTcBw8qg4m8e0qf14sDvmgTbMI0R3tI64jAI9p
zPY6UCvNBlUVBpGkJHd+43ebW1+DMPOJgyEA4gpc//YC8ED1k0IPbvnPqPpcbTMe
b2nLGM1/TYNkmsPhCIEjwkGIVE0JYBX+mwPBbwzxh6CHWWJyJ8ZcKIXclYjZl7l3
gQgvO87VveEIx8XexqyQj+45HRK03eQLB35SIHHrVv4HDJ6glJ/kGxNJ3F7S2xvH
e+YPoN9edbLJQydu4jAk6PgbL3Qnt77ueI9XNZMC0TzbcfLL6ECREA5G8oEpLXZh
K32sxQ8MxnvFYQwLlQIW/wfXlkZke+faisn3N5LrxWP22WyCI6Sc9ve3UeyrVISd
GsI4ndJL82Lg7ytf14ojqtZ2Rtlu/sp2HUpjEzCD3ziDlg6GjnZjYM6JU/qy3rT1
rTNDtvTANgcXJ2DcGugo9NjiUl6mhMgTpYi4Q3+6ppFelJED0y9hk1ekWKqmHuMk
I8OUE8lG6uCyXVwgSTsCOF19t7r43JRpp0cpAZ6IRhKZOyhlb0kSY1OA8x3CbJ7y
cy/ablggc4seTgBPSNlOB/bb9wDRvq74NzN26Wfv+7tSgecV6Y7tOVc8eiulyVU1
D0q76wezshcNa29q+6mapZfpF3rGspdnDy34IMZrh9Z54hFah2aq4HQkSbNBdDwf
2bToGZk+d8u8p6WxYpnQR6vSbCAqmMass3phPQgeT7WmAiz3ezIUPsrVP62t3eU3
uu3Mk+xHwrNhj1ks+GRDBnxbH1ZwBkVo+4ZkQ/0I5P8xBU+bLnIPARfD+3CgVNlE
Wyv1CYFz7YEMsfFacb76CY8qFrAG8V2ZHrRlL7XOEbntPImnwWvi7+XMzp0VKyLd
duyvs4XPP71J46Ru0GoRN1Fz294HUXW8b1K5YNO6DYq9fm2gLmpP4V46G5/sncyw
Z2MfRvW6BKIAxUZAOhPje/KxJ43QrltzGHrWc1/fPqtjABPcIZuiuR3XntU44Qn4
mL+RlPxG72cJxCKR/TlnYBfYGrJZiJPoJ66Z46ba5IVTvn7JDq3L/UUHCn47Ly5G
96y+e/kttxu05TFnZKj5HByBaOYY2TLvExe+crV3KtsRFeOpxXXfZPCOKjhHu184
qH5nwkUkkDe/q/aEWxQ9bbjwA/h4VmxYxXDNwWSEjVgfsRgh+uwL+tOCOiRJ2uNL
fj6wlU364kTl/FE+O0YBmE7fF8zKXhyj15wmABSziKqc0VbwkcHUf0ZgXH2BqaOV
CIouuzo40lXMy0/V75EVyA0vWkA46wFjR4fKulw9WPIyiDrl0rv8DH8WlrfnGeGk
VgeuIrfKGe6fuZwo4ic+hn72GMhK1NJAbMzXik49RibmZ11Pjm64EL/R/uRqusJb
1ET6dc1+CTPE15NhFFGhNYrxKqh4ZiRmA6pdoCIvdx+3DHp63CSkBR4QvELZUPih
pXG0exVqUqcZm2FyFW+F5judBexB8gLcwpU0U7zurlm8tYGjhMLBJAChytkzB2B1
9AboQbbSNKlXhOOJwB5knVllU05lQKKA/M3HYkH9uyN0g0KQatKU4Ay+iru7EDk6
LjmMXXyzmWZpHl4rFFZxX+Y8XRxp6VJozpDYro8ke20EN8IUkVbNFg8OKEp+pltZ
cnVS7KwRSkoqC/cm1Ou+ww+6Oed2vLs580A0xT3j+sMTK5BCZX+nTdsy/ItYmcKl
KUJqjnl+C3AypbOhpLZR4SaI4Sqc4NF00O1KidSc1Tvw3Vw0F3eS6695uesxUv6K
T3ycceNK15b9vmjBEBDcPBzqDw7DvAYt1yp0GmUrCyNQI0oKX6A4XB5FIs4tutcv
+SpZ0d+jV4ymasXkCuJTVqvRaV4tItkOxry9KyPjJUhtyrpEhiwjQxDiTSz740Gx
f+kH5KkndvNHs7GUfCuIxYWkj6B1PBzwwnAHYy6RjQLzh1P0vwh75+YzwfTsEtN2
QuDYkzo+YfnA9gTyswWHhSCAIWjOQ5/eF2NnSJMDZTAqoUUvUXDFjszoZVgsjzOj
lszJyCsyJLB3bbX28H1kewoAEPb4DKFtPq3i/FLg+QyFQA6qboNjUN7IOs3h16G0
ACsp66BsQ4T+sN3lI43ipNf5YlXtlwzCS6AQ37TPZG88rXmo3kKCebGM8TDLmCpw
oRJs7Wpo5RatY9wT03Tljm0EYoC0QFpe+osGspHKwI6tagPMK5AcI+QxQNIxwfU+
yNerTmuAjcmLS8xdy6ZBddOWPruQIH1cfofhR60ORCQJjr90tIS0M6V3oVScYiP2
n+qgM1dXTvahAy9k8jyHLbw9JGQZmqKlUg/StaD7zr7HRS04a7p0YfOdEbx7LvzN
/CiSTWTxuN+u3rg8zLJNXd4ktdFBn0WxIrsxmM7zWDn/Tt8nK9MC8Pn1NWNk9x0z
yeCP6xVp5MSCMbr7zrJYJJMDU3s6Dy7zA5GFE4BTnNchPg+ULcLBGEubEbKBTvc6
2qNqr+d316P1h6WambJKbd0ZZ5mg0BzTr0vDEFDDu6CLJ81PPzyDRlTCNvo63cuD
zbW7uD/V+ICS4Z2V7IojHunaom9xiTnbFh+tnPGo8f5I5dR47mzTtRE3UFkdSVVs
vuIwPswWfDMaUwKPEbrmUrkO5d+Qg7jul5oCvASUxcehOWtRKmmsPfH5JnlNi9ip
F+/YWWG0iN4CxMQDPSkJ2s5EZo9P95nWwGdDEgHJ9vRlUUeBryk7ULdgtECyGu77
/4u9zfqo79Ccfuxv6dVhih7fOhV9gexUbPqwJp0FRcIVRiFyLamhgHWvB0m/2yku
m+xdQCvPTL5JIpvkmGhoWoZLSFMJtxW6HDU7T7gSXou4ZXT4NkgCnh1Wl8S349kJ
eBg/ZuNdqpj/wjUQNqkdGqaXoQphX0WdojdY9oEuMzY7eJvU5SrPJMXoQ25buNVY
H7ninvkSOFEKJkfyhbfa38nSZwOWiiqa0OLuv/KAapLQHO8ytMEV2oUoKuMBGHUh
FZRqB9AtmKocwJF2Dw3VmvEzruUhgl99LSKfCopPPUHbFOnmN6Q3aSyB/yqw1h9z
tCb/xhqcyXouYXr73CnNtcV3w5t3izGjf60D1l756loEptPpie+cYUj2Rsg/FR42
dCtfNmZByzcPgA1XGACz2HC+XBDgjldP9jLE2+6LP/pj0w4sZDLUW3fg/09KZjgN
t50w8a3/U6puGKEaZXGn3YhNtJZAY/AAT32ZSa5B8lrxecgCF0Qe9pxlMM05+wUp
edlQ5DVyM4zgBGopM7Q0X/WA/3VuGsrKnDVQ3o1eRtSmaawtZba0Y8BPG4WBD6yN
BZWZZis+CZ0FhLXftEB8JOq35px3pI0Gp52OxJKkvoKET0pm3bohdPgvhwA0pkge
hvnkAwGSbrTOVre47AGKEWnkkcSKIFopfRe/G/VYmmGPdvHIewWuBS7itIDTfncX
KYm+1z0A/uDoXTJlRoMEuWP0NPQ1fbDkCQ4yPM1Pc92r+OdGskXtnNB9d065lYop
cbRxQD1gtgtqyOOSzLHn5D4rALbCgjkTiQRWhb3TB4ZoT/FEScMUbUucMIX9zjS6
EUIXE+J4UbZs/NLRquK4JTFf4vnD/3T/09eAAXC5AJnx/ld07pG523KgD8zJJ4EA
mvKa203LCBKsaQ/wtM5Q2xS3bVCw+a6k7G66Wx8//XaAAkS3H5Q1WN1s2caHknbs
eGFJCKQlsUFLr//oYvVfwBACumdWFvQTWoMfWKqD0DhiWKc7tGAGsDoN8nlqXm7K
DiPxYtllngdoU4RXch6jvxePydes987TdHQ35GAbKQogLcumMsymXGcseToAwnxg
eEwLckM10F9WivOvXnckUR+oDDOKkybhYElfzXOwfwrO/dpX5vJw34Tp6gPm93zs
SJpza7UOVd89E+akU3LIgKSCTH1GcH3jnkT2nk0ANSGctN09Ax35lENrH84bEdKJ
7R4UUhNbWGkY76gzqSCr2qP2xFasEehMjoRbCtmY27pGxPJhhX1iJUEFOLpriq5U
BOnPDyLAR/DVjE1/DBKpQeTWXye3G5wjBr7Liv4QWkZKwJ6pORefTaSIen0dwqib
vQWeBKEHN9sUIrXTUQvsaZzVrrQtaPP/HJsPMk2PLNL2hyizBdFFqolGlLAQ8NNN
SYTD0Kb1WDP1PO9KYNp8iKvILgQsGoJnjwgqWnnROiR6pxlrCc2EYKUpjxmzLhXU
LDQwxSltX9vQuObo6ueeFTsx4sA4lZOpM8lxInuUZcpcNAv7ggA7DyzLsUfgwYQf
ytW7Sp9Ei/tYuOZ6PaN7sK3Av6n595+4TWxMOXttQHS3/OrbHz+IKwyFYb5BZZzf
M4xf0gO4ooa4lDknMAaCpYGCk0s9HsFsfIXO4InsQUVIlTN4xMNt99/93/QeHZaJ
rstZ7/8s76sAIXZPxWc1b72Y/nSmATT5Ue/2um8dUyU/ZkKG7+MpihvDN2uFRBSq
dFBN1zp7gAP564q1AK+1THpm0G8BPRfztpGhgJyObjMlWf1RiDFcdnolSCvy0VzI
XAtQ1wWq3UJfIcOnBTokAylfx4HiuPyr59GgP1UuMA2Z0eKDjbmIpIIH+/wDxv/8
RFVvCiKWEcydLIINPAKAAqI035jB6yFh7WVrhh3LEuzKH0HkH2xrkaAjccc+Z7lq
BbySEHxeMr1W//lnZd7YtGc2Rii5Qpo6FlwBETjMAfYTqVqBDXe3XL7a5v5DR5OE
NFQAgSnlnoKuZYfWlLnwfo16+XiaqSqGmYeDIIacmRVZZMnKcw7LaNYOMaF6jKmt
wpsYIOtKQW2TpPMzJNb2atx/4HFnWlG9RLDFZSBRygnPam36LkZ5a+7otjjFiiL5
7YoAopJzyoW0fNPxoFsJGeRpYNoYVm4rFMXWJ5a8+w+fouz5CNzxWZY7DDsh5JD+
1ZcFQZT4rMYhFHyqpTtr11YDXr3BI8Q6B7Sm0nbPj4vui3/REOvppF/B97CMfz2n
Y+vljx08wNR6pTFPxelOAWszpJTgtH/e5kEZf64KDqkG/vDlbW7y3WnCv3Z10DUE
XtrZlNsUbBxrV90q4arSn8002KXHXnta71gEpo2FGZpVBxnvFgEtdTNT/0UlfXPB
zrNaH82H0KrthEX+8madZMQRT/zfyZSTA6kP4MuxPxlkpQ0nzHtz9yHsWyEqBgPg
zfqfiIRLtPvl1HExxtTw36Q6h3A/mkRE4c2XB1Tqqb1aKWHVt31n844unaVD6/sM
DxadU0DbdUPlTnzr08b6jrLf5Zm4Jl10aBg1u2U3cWzQ2YTTp+2WEcCGjTU68/Lt
IRwIZBJV6eOUlVytEO8M00y88r9AICVKE2OI6nDNxhvMzWzTZjvunuBaKZKx8zKT
JhE+pefiRB852BJzkyKJWaTz5lSMiqbKgreRmR90C13czsb4N4ivud71rIZDfzmV
YMB8dw9fQdoLBgPTa7Jz2dzGBIz5qR4CISJLmZah9O1pddXP2OjlHpufeke2stTD
dL8UZDY3GrzLSCaJNc+nARaEILgXZCPOq5knN03aMFwGLFus7gxZ3aT7G7wUI5cs
OHpMoBZrtBTLL3hCPXLGnPkpILUhEfzsyYyOrzBQKzziXHGH8i2Gb3hQPBbjE5Am
A1ZmhA9AHIaFTS0aPA1ylaTeindFm2EJKdnd1Bf8yU1XkZxSDI0272xl/0HM4SW6
HvW/+s6rzZXkDxakzwMvHLO3YzRE+W+culP0s0DdqchUsUgFZLp2PvVq6ouW0HAP
nRhws7ZlgJVZW2J3p8Ac2r85AjQ5br06ISm/E1UK2o+UdxqqtYHKqfc4He+DEXNt
LRPGA1JI1TzhnrmLlMkaS593bI8al5ME15vOsfoH4C9adMFbL140YUD7tizzD2eW
xMhYrZK/Nr9gNhZfkB1uK9Q4BArWk/SOENb6NgzdUkw5PUAfkz/nRC0fb4dFAT2G
QbQ0jJcyjgIKXBuEQgVrUewB/Dp7BLD2wOFKsVwGQTNFQfIj/kffjDZNtoO4XyOM
K/sFjR40XSGwKp7uUgjFgP5BESsh7/JnK0GNHnqEX3JXXBheFd/p+aBj8T1XLTOY
7ATS74BqXUABshdNjxRxjJs/DYgh7DFure+Qr0z3LzbRjOw9ANmirxbrLDe5VFA/
UfACMUvnwzVK5qrkiG8sMbNwloLCv0EHSe1GDp0U6OWbY7CSC2daa9qc1IWYvm9h
9973JLHrIPYVOIeDLilvANN6unjQKt07wnV2iU1YnDXWgLMPRtn2CUuqnbJdTtSR
tnbUyoFR5+IkVMD3wVVDZe+L4biUaNMpBnmQB652SVIfE0D8oqZvHSTaUGzb8Gh6
vDbKcbHlxUL5OBbt7MH3C8hVgGJDYhRdjJQ+n2dGrpxU1FoqtaLak+8tz6/FCZMH
qwZeLTLhIEtB/+Y7ktu13xVgrhL8IWbftiFuKbaWIVg9kofQwgqpnSkxWTIrf7s5
5gFCbmNPBhgm0Ljm/uH2lKwmDYOLcAhHgRR/Q3ALR1OaF0BwQSto3BRE593LTkYO
mOkbmWNnVtgfBMJacGugOjhQ8Nr11ugTRFopnvvjnHry/50nvnwJitUUAgKJ9Oac
kVCR475We1sZhgC1rci8X/fyX/clyaG8mQi+pStdVwoipnw1c6wQYfKuJABh29ee
dmhTxlUQ7EecW3ls2m/e2Al/SaySN1VB/zgpFvcJI/u7Pn2e5tRGTf7T7W8x1CCh
JbxnQH08JF29xwEeyMv5aL+IOHUUQiOO1i0Q9+2D54SlFIGh1vKCKfodtrj9uftO
7zbhr73O1CQlzW+L3S10UaBT0EK5O4V4FS1jeaKYLsehT2bwWi7c0C6MImw7n6RN
Oozp63HGPpCdxd1gqvz3WYU2XN4Y8sDW0UcU0FjxYrq+9ezv++oYQejMuMcc0G9E
DYS9L+NmcJVsZrS4KZu/I4Qbk4wpHPs2mb0otFZPmKoRlmaBB++U1l/k82sXn1UI
qQtIkJG4ybIjoDCfhh3zokP3MY2kwDvaP0OAEb0pUjFnS/dangbZ4G0Xi65R2mSK
OyXgGS5hfGuuHs1lnvn0iJNr0zwmdisBOol/h4Di8vF2NPNvu8e4LFsdcIcTGq5T
YlcYZB/x1CkqkT63lbCsd0mJu2s7tUXCfPIUH9fI83Jy9LuIqhBqWD1MxBu6+acC
GBToCg6zK64cBqBQG8j82Np8/u3d4RPRfIVON/1Yr2R++2gp7p4bsHBv1kr3GU76
LdJyHDKsAMrE288DXJ8EKY6yEJxu/JtlzWo1Ln9wBUuVY9pIFS11B4KZSbEvh90A
sR9D2aWd+z7+y13w2un3Ir2ZD8MpSGZsp79VekfTjqTsB63ouG6DvE9p3SeakW67
WYMv+DHrijkf4k10bJXKyEwmZ6GQaSMKJO3rdQOP7rZN/78faxjQExlOAqF0rVh8
JENboNdU/kkGNmwa1FlfD31lEtWcgCoi1Ddn4U+dj8C1d7/j0Bw4XcZeDeIMzDrl
ypO5rqpO5yyJTJMidjbbeyTWJJfhsKyV4lZevNY0aMiKSh24IlYRtSdUPMgBkFmH
kc2ow4p1Cyo4UTaivGhiic77x1ONHMbepsk1SAuxQvbm1vaU70buYWdQc5Ub6Cx9
m+elnr77i6l7I6QqyXWslKsr4G+F7Lsg1S6pBMH8JWAmD3u9rhcAZOylGGslrHAe
5+gGCqaa9sdv3qFHkzjE8vcGNZlZLnjcwXPFtL+49l4o6rCVdXZmjfJfL3acYtxe
q5Nmd0SVdJg+ekbit17BKk5QXayjsAZDTyIQNQ3luHMSJiLWoGdgaou2jDdFtkSv
z3Lw1795Rh8dFVzeou84CpzesgE1T9i9/ybJEJWoyypL/WwWObx2XNY0z+rz0iO7
dQ8zChk3JsIu3mMalpwyAffrR/MyViwElryrdwfzr25lIu+FO3f8Bdho+/oYIuHX
vLaGLegVy3uOJncvZS5N+/Ze7J6AtSil8lUG/nGVsP8ee005VkX64EJ1me2lKmHt
wm2XOJszWL4c765jTLj3gl4vutwA6IsPJvZtEQDyKfw7QlGdmII877ZzHRP7r7X7
ZdYoYBmdRRCs+F4M58YHXNBV41BfLKoJjVZcLH2qPvS2P36OFUY3CgYl1FQWaQrF
XH4V7Isft0HwtLwRy+9AwzfigEPWgdwVGh60bswezFb307MHQPDxw3fWaLT0g29E
M6XNG8U0eTCF0dmvc3BMezE+7ICw3bV9Jn/NUlyxkQMxcwWH8h+iKgRtD3BnfIBI
kCEZI556H0YLN1DtDQ4ihrfZFOuCUVG4rYmzLU/DTTi+Dj38lUhjZ8hMwcw2l5p+
cOyBvBPGm57eMa0PviOkhj8CMDCmPzRcabj//fRw5oLY+SEL9iWh4LQeM4HAt3fI
FtdmoPEsxKZRvBqiBhDoNkHeAwb7s1w7zk0TkjGMKJI5T5BNvPT5ULeUKqOyFMbG
4n7ke1K6KWB8A/AEhi6B/EYdhM8doWxagYryXlAXfkID1smWmCdxcCJPZJCTfZnP
WYidOIZpOFaNpPCDts7sWFnQfnIMOoee2/buFLZdkWz3/3Ygico0aaXAHXzmYc2V
AeTXLcPQ+3ihQUcKjZAiol7SNHt3fQsV6hifUZuqEEPAZYIEdt7t6weiJJes7+IG
abYv7BpG64w0R/XLw3W8rVQQzWFVX/LKMRGUWqJVF2BpRBlTy23SbQRpYLoYDVN2
LCV+0lyQIN626p/EOiSXyNyjsLNW9dst0nCDORSx4r8pHN5unZijoPfWfX7w8V6N
ONDjmdioXMt23pIkGDklRKyXtS1S6wkNmbw1zh9ePquH6FfTFP6Bz/FZx6M//B9j
zdvq+1YfgdTlhS0RuHuY/7CkAM3QuWcMI5FgHsgH3j4KvnPQez3Vzof1027Y2VC0
kpN6w/9iF7eKC4P5dxB+299uLy8h45NyuiKYtqhWsOZ8PG4vjDDQ7ym2DeVZTYS1
VkqZDTad0QD7d3zYLz2IRKdWxkwcsxKvySldRv/BcWN/6FMKjpCw3dhRxW5mSIr6
3wIXD7xfKD3dsVDiJ7B4Vv/18tL92jtpfKOX95dfFOHJk5gT6y731eW8Z6WSI3F3
2+XTArzrCuf4OZd1t0LocW06hExP6uuhRkt3A4sxAeycs/JA2uyKy2ucMqTEEcmK
aADnGwZyDt8mDsAaAcaKfJyfP85zPo8XcIskgUoYE/GbS74T19RY0MerOagaVm/u
eykBYGI0UAwyigIsUhMGaEAosP3Ly0H2c+hWYJLFTyqGHHt9dF4Ub2rhogej6dre
JbNWENUKH8MZxZh1JlwkSqL0853yCu8+ELBh0yQ0b3p3LGi7x4CJHK5oDSJAV0Hh
V6GMIhNhuMMmY0etkb2rMdQEUOtdqutAwpOso8bsZgf4qc5nt203eWlzdPqBiRtm
qaf0MvcFM1oUCc0eba33e/0huOJet/tq55KiKQA0OLQWJ952kXjfSJsXNnh6+Aen
HgFKz4Z7RadFs8rE9yj2eWvtb0wV+0YKugaHZdI3Pbx58rUikrN9MP7DlaiF23Hk
v7Hpqvb6CsgOQQl7q0nuXzYAZz9zuYFHLxthf7YReslzgNe+QTBLy0zF0ov1w68m
hlbZizPGM2TmHSt6MjVxeisvGMq8miLGSDYQTU18OTSWYjbf/aFyAmG/wbew6bGo
tOHGk2iuVO86QK9So1TAY/ctWypTAlNULNe1dLsHWSpTqOyG1lJJUKpeVmxQH8F7
hKSl9kc8xU2hQsGO79lLiUoWBoFRAPANuUrQqW4ATZQDksRMRfBcVzY5KpNI6NTW
TXshz7UyJWt+yqlEgmGvEBYWut2v1K1H6i2KfB3/7tTpVYdqEqw3/M9dvKzkYSCo
Jgy7ZmeFqY8EOqEIGabOA9vuksaieJr3ZiVzDfF5rg3SbrSBISAwgi7kxSJh7PSe
g3dby/dXqWc6DDOnJgFxVYKQnU+rEAhpegfqnWAxKVhGBPFjL6JmHA4CMIUe0X/P
PuNqlq+xmo/3JqwdWgWbI12OLLz5M6qu0Kr8Gt32goUGQka4qYQP6TTaO5dXexyS
+tSfkOpIbSxax8CFfde6xMutRUu5ccOm6VlzZm629huLkf1p5ZGCVA+2TSODhrA6
sHGxLKjmMtFkJj2MoeVWXRcZ1+NBH+8dv0/HPqCw6cPSfoF9QAUF4+Nu+t2RUiax
OU8z+4tcPSFmR7fE8wEdhzUB3GZ5oqqKN43+/WNx0aKI7aaFeLZnCTxa9bLD54ip
rorQxhQpfb5OGf8YlG78cUjDGed791rHQSYcu2rXw/8qOmpsy8j89qlwU358lnM/
IJRWCyCQljTDzBADnEvfQqi3CCGzvTM42wHQrxYNkjAdRDSf6nvDwP2ct4xNWnd2
zm/MezQqyMR6+GetCihZXVCONtPhtQDhR6eQUvLTHzaFZFPNtoF2amdxGa0e6k0l
u1J2KK2jSrUAGYzJxya9MVtaaW9vOhHTvVk6ZTMUPKC6dcIp7j144Q2DWd/JWqMA
yMm0fZQY4hMypy2cu1DHvXN/NZE78lHS9EOMLYhlCAwWq1HnyL98hk2AXlKR0G7y
8exAKYomfJ0cPBuNLOi9kA9b2AzeuXcCSXajQg8SogLKJGYSWBu4eB9QTV6PJsMw
z7hkx+Zyf0UV8GUaSKD4af0WV9FwGzBJPx3avEkLsLzR95QWb1TFVv4Zo3B83rWK
3sSUURqAP/TETaQNDWbu9+Fj7zB/cqExYuvkVQ3Iz4VVE69trDelgndSwKImgMEZ
opb5Mwkzyy1YtTjWaHCELomz4KIPuVXM8nI9MKaAbhPU4/u+Gg3NVg72vNPiZp8k
9AIdtzAs7Io3dsvoJ/kYAqeLWZYC7I+Vj7+w03LSUEanOFvkTOfqu8oJ9bUwSH3W
/O/poo9fShjXpqM4/W/P5vn+IQ3k1iCcUq44/FiZrrba26HYUNYuBHinlYRfQGbz
rOfeM5Sn3vB8I/WsdpoJNzC/SK7FJfe3qX0f8Tyuzh4y5S9te1sGE7L9ZQXltr7B
Oii0gDILVD+FRbT2cUqt2KQm319wmzmIBxDL87DzUjJMqT7Q/cYX35bASz9pv+/S
18Nr5BrALaJOz0NkswmxlKl60/ZnePZq6MvxboOOR3cQp7NusRV3jHM8S5Xk+9aN
KKvl4k76FUbHEPxasJp/rqpDGrIKwUwnCNADzTCrIwPSthaWVyYLlBQlFOaR5m8z
bggkVafL0t+PA9F3k/L0JXB9jx2+TfCWlxvnSKkjWnwXfigDAolwaFydmMs8JQ6V
I0xHO1dq0A7+g41fXCN98oQUjoJxKaTeIu0yZh17i4c4bcwqnklVbBA9ZZzlmvdg
D7rIEgghH3tJgn5UmG8901I5nggRXSiNEfCEFRTsDgmOsVmHH3mRE5IrpkDMoLcs
4KVE3Ac6ihEr6ySrOYkDPh9xUaPJZbB0b4dzEnTl3QbpSmAiavM5K/AQAvynMqO+
ilbyJ7cvh9NHiqiH4zsy7uyJJmz+mAI2CyzLmYgGKJPFE9fLz5YmsWypKZlghAqM
4JSv9pvMfJaQ5m+Mrt0h4qbBytE/jfLw9lypMb3HTCAA3ZE8w8A2+sNjV30O9Lbi
FMI08mE/w8OjiDv/hga91qVh9ceaVJcfSSI9xJr0rQw3Zmf2cVXyD52IidWsumS6
3e/YrQYCW4h+IzSHFpusT187nvw52GmsH9vOK+8samslPa7bKNPl5xCnSHgwQ7UJ
S80mJurUYhh/v7phlTGKdenfRP//xhTzGhR5D282HcMPspmMkQDODdiLY+yQIeoq
ZVjKO5/q6ULuiZ7bYrgfmWBxlGfNLCvHPmnCSKVcL3muFX+4NSW+Fo5RtUPtMD+Q
KGpsHDjyx/JbJRfJgfPhRztv0lJpgpFA0csfHPTIF0bykR88G10DCniriehsICbd
UT6mKqIwYzT8w3SPvTaUP0ZrmRNgFYX4CEtki+t2NtnaRsPP5CusDVWRjufAdVYJ
gfgOKX/NWYxEwwumQo20Zss2h7lXFrJCJd32UP7jL3FXWxKpjLb0MG6QbmEhpgSb
yjtMjaEV3ZfaxHls0yi8X//AIZ5+JzbOJnUmIORzN7qDCkQrE8t3fIuk2WK5BTmR
dIN+mXnvnMRNGM1r8VRKUbnb1cC1foWFpQUS0H6D/oXJwVMhcy8977D1RIL5ACub
/sXm8R8ltspk3vhDSEoLZ7Vv0RS48YrDR5VLJMtalmfXzx7qQKGen2rKakLv3sIl
b5wLkLcdJsIZ6+UOgvsEzskCf48u0kuwRr58TLB0dZw+tWK9nL/WxOMRK/DFTBV1
FUQvp6hSTla1mZy/cj9OqZ4TgnPLv6nFQKQU0plCPhEJQyCjT/Uz2IP5KCiixKs8
6o7NsJs3CW4PXsn2/QOxNr8CDw01VPNBYPM31HerUWY1m+uvDQ6FqvedEuB+1/Ng
0wS+sT+JNPIqoi15LJYoZviinX/auooLpz1cuIve/v0aZVg5qrdPnzmnxek05PoH
oZJIVOW49MbQwx00Y4mSOf0YLtf+mpSU8DZAzxeDjYn9ZZesv9qMvL2ZKZdweWmf
T7whLbX8pVWnjZSiJscKgaOR8FeL1p1C9IBN8pKODhle1IPF/DgAl/evEuUDM3nK
yS1i80OkdriF3h44V1illYH064oQsPrYVnKhd9+J50b0eEhG2JkbDbSaFdKgcwxk
BhbLulFqYijdp4BUkrwRGZZVuUKNtOEOqSG+8zvQDxgJ0+tUVz31E+NCtx74OCJO
X8A3wBw4nzidMSb2L9pSdXwZNEMRasBG0eZulA8HkG89CRLBGKm1HQ6/0Pnr/seP
Yn0peM52zepHu1/cShutH94geIiP7c49qygiq5XTgw63jBAEHZdDjiimXoLHI/bh
ZOcEiGXY85HDrHfyxMPvohrjmR6JLmPuSoDHWev2MEHMDjWLvLbAK5nzE5Nzj7+z
4cO8xauaYWIK+rKC1soUyR+9+DuEYqzWW5F4lSEnwfcywQeR3JXb7ho0ci5ZRZ9+
TlBWWDDPcSpiMNg3rC+T+u/Ua3t0it8KPX5EWtSMH2rBKpWdifSIvXl3LbBQfyLJ
vtuEqC914HNkgsJxYsF3BhqAI76oGvDT3bF5ERadEm8rq4mYIj2FDCpWjZlO/J6F
/yOQObhifbZuGcOtTDwF1mGYzGfPul0jxJzR109oLZ0a6Qelpu72rChUjI3tY7Tr
vCzqSSmSbYgrkI7V8wu9XsV/z8E1W0SbDWUzz0C/ulAbLGTiwbogUsMGfEHo7ave
nY0A2lMvsYUntn18XdiGx6OLEEQ5OvvTqR20etwMQVEVLTnCMBQUztyf87LnQQMM
Zz7sryDbiv33LZWIPJOOtb37hjvliFq5oqxnJGQeFE6giVOKVcuPeXLNhvuX6eHh
4MrZMhmJ2tChuTcpW9o+Q5r2jEHGeMhFenmOru1SxdH26oNhs3PmO+PXwxh8cU5m
0GOxlHslJkGgPOkT1ZffnkukU0rmssAAsUkVMVr47td9tXQB3FO7RzeVfxF4CYqq
7/ZE0TIDFJS81rpApdKbLNr6+BXcoLaw506J6mFvf7TemtXpQsaQ7UQDjxwHM9+C
qnf5TM2j+ktwBnE7ucKfqCcmqh8EUlJJtGTqhc8QhYB7VOIRAb1dWVZxW+FlTNGn
hpvuj7K6ZHAOkhwHr8d9GYRXg9k2W7wir0VcC8fMPQeQixqT9M2tRQuGftvbTnxP
NPOBj39Q78ZQBsIzqZ0jiIThkVPc/5aQcxiDUe/Y/SQ7GOXicV6GRAjqw6PgIwrh
8jYvGEoUhbusz3QNf2ILfDnIHoyc1OIE70auNuAvf977E+HKzi4iFtlXunTCrK1W
Ur7o6JzgZd75LvNw3i+fqNN3cw1AEUZXXiNDcH1avdksXdkLf0w6w1oPWAbRApH1
cd2VKDMXtLqR74ysPN3nyGDVTd9PFgOdAF5dgnzAU0dPJ+C2APWDxgiMidkBZd7Q
KdyL2Uqb37H6ooG3Nvlt6eItQxcU+dRle1NtLNhvwauawW4vjibknVYIGn/KMXa8
NEyLBlfL+eB9+sYR/PJrIR76SPdA5pwtSe7LyRFkn52vGEkInhi+6nFHyizXl+tu
flWLGzWxn2rv1flb/jnhGLWutqc7L1IdPyQufCVAj/5ocjb+i22TjC702pejdhwh
LyyYJk8y/f2mrhSbbkf6QRPzW0IDWqnIVMzgPH+tnkNhGVlpkzwwLZsezT7a9BOl
QSCjZibPGmt5mZOsr7WN2EdpJFqB3mxENi0mcxyXJBems1Eh0jTF9zpYxKWDaXmz
OVL2h753DZSeu6vJ6KeSzPUwPQxvUpOsguekKEXiHnU+aLeqbel+674FFXy+OPls
QD2LxNEZSHcKLSdYC6DeFlDFjH4XTF9d2TPkIqjL5kGAPCwyZ0uC+ZmkV9TBgrt/
CSP8PVVeSeFNaZs14txBlYuskvvUnWeBBASI2cX6G0sVuFV/GtUS+7LpOveVQ8nd
sWczOtuj8o4zocYHIDBg0NZF/YVpyqZNLQsuQRefN/0lsykanUYtCKwxNTXDcoV8
7TQtwMOZfCWvZf55toEAwRp4zOAj8LOds/Cc0Xw8upETj+LKVSOkMAYOu6luaLLT
IuLHtWmwFFreYFzn1EenAOxNMYpopqeGLAZviR8n5VaUX9FGCqwmO6agWLQ1YL+Z
8osH5eQKf1lmpKY+8D/9NkGyltVqEIMoga0dWkyultaUipkxuJqGUbutlYzjhnxf
qf4JT7Ehmw8Oc5dpRNqzTChoDdMTNi85z6IGrVLU63032NDtfmKET1CH42ajs1NO
l4KY5cVYD8qtArkessB6WAIWQ8Pu/FXwGhCrQtyDR2lmDrQkE/XwPfVUosKQSkIH
vtjhAE/82B7C1h1S/Jib/cIpOQFrhbyU5SFwjE28DjC16XyP2GVVNuoek3aSARhH
9dbvH52llryALnPelXgBaaR7q6wNrp2FNsHSnXVCQrtQbR7zWbWrtUlO1Zm6U7g3
EWN8cd18tf3X4wACtWvPKwH1/68YtxFSxRhFQ/ahgLu6BT2hsO4W+zvBmgxEURGo
8LvJHGnbucwfsoXGxNTZyMLd95Pr2xaBe0cFA/tSx7EgpdEOvwBuS5MuE0L6EW0D
ZrQXON5yeSYMVta/B+1QfYNoNfAsrwvD3WxgZ46jmGgq38Z1O/elPsEbVOlPYRUi
3HkIXpcYw+PR/I3KL4ydPjJzq1p9tDvrUzSpPb7G/3pt4zzV+qR6VrG/HjC723Zl
nfTKlZNt4hXqAZQscwXfjCkfX5TIdnRQjsrMKLLkOYtY9dK1eTeDKSd1sFRAa19/
YP5eSKc/6T3uxOHVxXNpic88MrJDW87dKkwq8F9gwHJX02D7o/2rhnhp2WayY12i
N3RvkLPuqBlqpOzrjztmeRmmi+VXXNGyOVrLK9Y/igHXScom0WmNmE1y2jxbchug
uxnqH9H6dYojEt7RQyri4vh6K2tpZTIJYNztRWBty1zU8PizWXmCazYr5vSNkKdq
UvAlB4EKDBsS2eaHFAoT+cT7jzJIonIh6XFLA4anhdCmoZhRkhPezX7srK7N/5oU
KPgm34MB5C/wxljodd/wWF8NHeENsU68GU3TGpTJM6e6qEuePIEBgk0mpRURvT19
S1uvyPr0SXcaRv8/q3qAoSwojRWZINyunCRtbaC9f2VATs8BYROJSaAPNDoKBuUP
IGqq5wguEvzOGUihlbICc3G/xJxC4NuyB5kfEnwlQ1U2iwr3G0Jf9b6Yrcid9F2/
yx5Bdt6YHqwPN3RmXAsmWZuz0R1FoCy8FcOxgn/gaaFiU8vCBwOhkPbOzbeWh425
MqmiTf1VrKqaoGWsO8LfeFJ8RaA3OwmPX84CQItNajaMXE7bD6v+Sqx8LOzD43kz
t1t5xwsHT50Inip9zt3JWsbirvdE8McKS8xSoI0hZXi9rNoCQUxEcnyNGWMetl53
MQZx5lLilSwLd6JkBdxn+wp5QtxCIU/bLBTpyUrpx1g/pYt86dWI9KQQD+IYRhMt
LI/biKAPRKtjLLsCA13+nxd+EYCNRt48zpmloVEUozNM0qtWlDZSwOFiSYRTnyu4
ijLx9uBjzNeUZ995EU70fT447Kgyx3PDIVhFYBgBeSeLxMbaat/2hdMX6/vEWbak
b9rX6NlYGleIx/fsFiJWOtift5XkjtpqirQ/xwzC7cnckHrp8skz724+862YGvwe
NK7XEf5jW7j8E1wsutAIp22E8V/ukn4Ow82m2/RDwYORBSz8lZr6ZtDvb+rxL7Xu
y0J5Qes0poQ3uLQwUWFlfDHRG7v33d7R7IsU6Lb2KahWg5CHTINf9xMReYGlul4T
LJixmMhGnQYvZ8zaxR3tMjbSNrKSfU1d+dtfeTR9i+PigjAQYVUzTA006UHt0qJO
mTT0Jc+EYCQ/3LNe95xevu+Ak4NcuBBWG0glyajthmBGABadk7KKi8tqK4k9C+ag
IKBNuak6c/FFkAjvmSIYyfXePoc97uSRSsPkwujuVG/hD9KtXjpERkkpD2VaHAf8
EYYMnmx2ak3mMPhFCHxC9l5ZjhCGOVIGiksoLWOQC7Ih4JWlXyF3Ol8utREjIF/W
HtZVo8wEYUDf+r1BCP6wHoznC8eJRa6UG43LsxrKBlU3aH9PVIFW3CyNhIBYuqp9
7tAsM9ZRuFuQfaHMMmiUr/gRQVQjQeyyOpBYcMST2g3yRCsW1Bv24N9Xeot5XA8J
B1E7A9KrgTZRLiA/gHsFzhIX9FWmf8XEjbUoKzBpEbM1102kCGrwHX1o5R1Txn7a
kkQO361fYbsFHyHkV6EUPZCwCnzkY7Z2XUqCELB9FYgWd69WSVlErf2W4L5axqNH
vAiHHMHKQqNhtvwrfp1z6Q+DHIHcbizXgjo1p596mHFNuzDiAXCQHlKsbeD9HKTH
cKLTqiAqNmMjOHqz45dgWTqkh7XPV/K4CWDEi4Z0zQvwITofnlaR6VWo1V+1jC3a
dd5hoP4U6wGnRxJr0A4ejActGtk9NcGBNJ4yQqTuPdjDYFLHxVIdnToYERAau+Oh
JEmpRaGtbf5ltAI6cU12eHnRHfvVvXJJ4rJLnDf2uTNblKfZpYw5DfmS7oXUUCqm
P1+cT7sWLnSk+bT28pXW2AB10W0Pzsay7hJkN7wOJN022bkkUt0kRxv4Dv/97hmP
6cCmMsKVFk1fWn/k8KIZ4ORoSzsvFmTkardCMtE8ausr5Oq8nT+0yGN4GSOT90CC
rmPObIJMMm3zLFf3fd8ZyCTj9rkygkvrl6wLDXJmg5lrw0TgwZaB3CV8BvsuqCrr
67pcm0pW6q+BU2cGRXUXtkZEvAGeEWN8Yx6PrNSRD79YAo6DFbaDh87hmwl+5wy5
6DWcgMRqxI4ZzMwFbtS8GHukvLXpZOnKa/NtvKlKVIzMyhQcqgboqjhOzmxWX7ME
so75pn9QTI83+YKg+UUeVM+v1r0hOZD584CVaJBolBFnmblPGaAzxnnFSNSabMPD
CWY1eLEVwFvurB9dIo02CKR5NQFP0mh2aqk27mn+H4Jp+7NO6+dcT3QBt+XvRWx8
T82Hc8FcBicgkWKkTHBMw9Ejwv6umZpDjFuEi4ihURiGuvKZo22fxZObUzqBtaSD
yGtCufDGp1Iu5NeexY7if/xag/s9EJE+yfeKe4KV6qc0x0RInqAaz8g42qhIfLfV
EKAQz0qpo0h5qrUHKGWaWDJLhcNzATXTkpI0U+QF8/7TALQNFUJx56r/qxMnrmV+
0RDVLazJ73zrzHjAHY2Im0A/4iOQGjW7RB8P/BEbtGy/3iOyZGRuG9ErQkdIvQjc
eOTHYE0pLwCZb0SSk9+r3OtALNex597ReebyK9pjFVKbdhMzw4diHn1M65bc8aTI
piUKoQ+B08WiraFj6vKh4lWBFgDVkMsi97c95Axh41I4wZQxYNnvuomjU3nwiZ9N
XLAP8mgY7OTYhbiJO/PkH98VphhXhNtVZQl7G8yZONtBsYQdxZDGGDeddYJEy7Is
YsbkYIQ0XgrMXKELXk545KfAjrM0bs5t/Wq50HkhluQtuFjoMTELzRr5C5RYdQlP
rHb/aXQzlBEfXw3EkmgFTgXSxZ89E5uPAuehn+4n4y5g74aVLAmrIaCODbfS8o0r
PwARvxeyaNDIxBLOTK5BCl4YDutw8dGr1jLq3EdjS9DUkuUHvXfA/GEujFAFPtGo
c5S4ozKCcaK6ybtdd6k4INrKgqbuCy8uhtqpDXLh9tk2aNBAqza60tHmQGKjZgwD
8dc1Ff+RvSQEQA6EB1ODElL1qRZxQQPIF2Ud+jqC9VX36TlWkoh8wNaibA/Wla8m
RxepIRNEJlRi/3Id2Q09VHq2rBm8Buroy+GRZNiZaDAxN80hGyh9SfAA8Kp5gRks
T4sYooSLnqJuCVw6kevUPTsAP+LDFxMbKIptw8Qw97FGdWVzLLTx1QO6v6zEoNoG
PrV0WZ3ESCj4WVL8HmSvKwpt658KBUd09jYFQKLFkJp7/fg4khT9LN8tq9WNUn/K
MeQx8ACUNLBMvY6m0ILsWxK+189FLoRlRuByajNsMe/VjwEothuWvGhH+l/JTGMB
e6L5yVCZvgT6zBURt7waBCZe+z3qlmWo5Kh12Jd9f1O0UtAxUfOKTX40mASpJ9Ly
w2BvyHxt9l2qRJxQqtEpw9xKY69H9STMfiDfUZYIefm8EOmdyPj2M33Z3MoPKObu
J1SZGX56jNeHk6IIoJFH8QKuADXWdsxIgf3A1GKl2EMSuLhB5T3jVEUOw5cyuyWU
1qhBO49wWCD62Fw78i7O4U30F4dbgBVYNll/8G6FRUwggAz+NAVAY2rO/UADtfB8
4S+nTiLpNX4hXyuswk0P+vOFvDtq5FZJUQSAgaHumWsu4iMs+bKwArivLywNttaA
qpqGmOnqmj6wruBxhlEMyRecp6bg0u5v/cVCB9M83xv06MW+ss1zuWd/X4325H70
pH+NdyoaSdCz9wPHR22wjJtzrgXJhGRpGo/MZYNyolBDjR2GRMJWICA498E+tUhN
5/arCBBSK/qEMZ53x9V4uMxF3Mi08rn7K9T1yFMHhIuZ6IipmSRanjP8ar9Utb+N
sjEQs7vjQ8XjY/mO4fNIzS8JeS4pnGYWON3qEaAZV/Tgev3J8b3AZASae+cmt20V
5Z3qYSRgyMw0Ba6QIFv9L1vI/PoQPwv+DAJVt4hUtY5QlE20BNibJ0L/dJhsqvH3
MzQeJFRuhDNbaHu0vcjuj8LeLvAg1CaxiErdWLtQQh2kQFIf/WdNZmORj2TjdFiJ
+gpoSrLJCC8LypjcMxiTSK+Wnn9TTNxIovKalSS49tiUZhxmwHNNEaMCiyVO4DD4
9ojXy6M5dLbGsbMoVJg4YBXk3Jn76QDM+IqTJVy7gQxsfusrDxk9e6z427k3Sjj5
+QyxyeI5Kjdka7idyYBRu1/nIZ4aDZ3ml9FE37f3b0gxgHKK8+oSYXOSAYwML/d7
oJNYEPjQcNxk4ucdOxRVLMzGFIe7Rofse586EZuusQRem1pPMmLrO+HLRgPgPCY4
ajVyHsM8PiglwS2hGRicQht8rPwrUPyZ+PbU5/mOCFm3A7/a15nTMCIOpz99FCCR
J2sQrIW5gHtnrYY70uBaGdosDUXoNsAEO6kgjsGCKhfMUZ5iD7jnbAPo22iGIpJk
uOhnKooB+rhrN8eetCLCTKk/7VKn5PJQC7t860NHWb8bYW8H55j/DTVyyZDEeOzR
KdR+6gY9s6ZwpW9yK5hynY4hoN/qiZGSA3uW93Kon+yXNhjp+WMnKlcCsfPMOLI3
7Dmdv6SHcUzM2dKhyymvC3BogdlXIKPUQfHHBY7tfGuh4sqKaXgirFIw8Wg42WLW
ZS2AjxoFXQAzLJqTaPn0Zm0SkH9r8R5xDYVxwWprmVMsKgC8Or5e12C2hJBgXMdd
gSnAVjAETR791du3HnuQ9PY3FQtdKsRXS/b571MCJtbFJHDlntO5pzmnT6vlGbu4
46SYHRDgr4uDG6Hs3Z6FcR+4AS5jKn/HRPPdxqabQdhHXLSSBUVBY1OtV0L3QHMj
vEZHAOQR2r9JgaMcVG71vhhOj2GVkWXvNrny5tSZCAswC9jxyAg8xyQDXYNpFl/S
V4rREhJL7eT0L+kaDTaQw8slFNZohG8xv3gJO72OI78m0Ta+fruRqqM4tXzMePHo
k0ZcU2plKoXMz0kvKMaZIy+KTGDOsuGBhgO9oH9DbqhSVGX4oq+DdCX4QD/v9jCZ
31r2acJVD6MmjoKjLdxpX1sBuyJYoiba8kWnJ8eDktdM8fM0TgKsSb2g+tUiDaCb
K9jQ/mD01gltcUlybikpsrwzoVizItGUt5ALhzM79mtVaj7+P/n/raZPsHqIg6O3
xjlVkKsOEh0lvrr0p8tMtRGWEDSCUBJdD9x3INbKtb7lykeVwSEqEaF2t8qmkunh
clH7oNfCqQdbjRwsNYtCivkCzqBGp+gUocJKf3w9Ka2AQ1JO2+l4ju4qS5/5R06h
uh6NWce7YJRA5Zqz1zS8ECaBqh8W1d/zBEhsrigK6H/8lzu/qTU8rC5ybfuaydyW
HBgMIUcjREjndPfOSQxEarYTQgzEtYesw3w9O2jfQxhk2ZhZYo2tw0YnOvkmMxAx
6B33jjkqMJzB4uRwWOoZNiSpqx3n6XTluMZOZEGfJ/JMWCWmExxEkRWWxDbOw8E2
nILvYGBA8bsUZkKubAkKTuYZjKVrOp87pRqa+igJhmmJeJAUqNFH7soRBPA67a3V
GioM5bu8eQXhxywGHNdJvzZBklmPRwxYCbxqlBuNQWo1SmDCc1BzQrJ/2+sW/syn
qPbTI2OERsBu/8R3EMU2PQLmZCPSBUgEUoULo/BwGcJ+dHz4cqKzkyvP9/vGIBfs
aKGNJjfI0MGXFcxWfZENz6HHMBElHvA30mwJKax/Hh5FlVvsfNssl4JPpHUWOXbu
R6aEackm3NRCd9rh2RzHUquave6Ztt7OC2630Eht8U3RcOApl2uqy27pcM6Dy9/a
bWwEKPfVcfTG6vGgOEL8tdFcMetXQMbux6rQXWzAOz4Jn9vssKTUyzeeYsv3jjpc
g7ec72kAh/YpcoaO5VQ6N0qO89sAa/4BBaPIAHRCILuoh2IDaa5fd2ftCFe73F9h
6mhZSlDrJPwNxDOOh4WueC/6F5bCep4B5xAhF+gAZa4xFkbExKnLs09u/6ILcxt7
iHf4WLQk880hvAxM97+TuB9s9TdQKJ8UoUWPHnxGqsGYbfMKb+1O625lC6mT0t+s
w+c/Fa8xnTSvMdIvlcuWdSf3RTohA36cqi2mUCnean9HrIa9hVtvZKVeKFmq8BQm
ebPEBZuhMWfX5GlND7lbh8301Nf7aTRul1fUWHzG20Daek2XXDzpwfO/XF6K93UD
NgSMV5+7hxO8/5WvUF+HeWugE6uf5e2Mfp4hH0CgTEtBvkhuqErmHS1Qj3bSb2yb
tQ/p3evbSpRyV93aGvOwcruvGA7k4c/PiKtkgzFyuiWXcU0hZvYnyX9IH2l4ejAZ
Ju9ugWTh9qyl/Aoe9gwwfoVFLjxBmY3YKAPiVQ+T/u+B53YxwGB8lTwo8lAhULcb
D1uv7pXoYlzbB2iXqDCJQisiBdGiqAu/UIciypO7hg8x1gytqD/q1RwiRvGjnJiZ
pa9zJ0t0nnp2YCNVz1Rj+zwBABOC5sA9Bq0A60Mt/uAdQY2Gb5drG7hQLxWx3b6r
XEdVzuiRp1wqslkcg7jSy94zF/xps/XRMhDVuf9ZMEOJN9d84TWdVlyVRhTpGNn3
t6HU7iyTtdaNAdvsDwiBamRp5mOuQkmuPM7niyN+whwBrUp6AZZeU2DsExfXenbn
Pi2pHl/ol+euCwPfvwQDBNmMPNw+L2NVp1K6ac6qTQpavjMfWTWU/Q0GGdOSLRy2
noSHZXIFjfppCMxEgXe4sdNO4fED1qBIiN/XWxXdqYyp6BCiBhtzllpTPFqDoCEd
ffmlEOqdTh6r0sQLrcSoJ3iOmKn31ExPytejNmJxViFZrUuOKsokQntw28Wgafk3
jaxXc0IpH5lAGYrusmXQIVbTvP7B7Oji01RsU4A7YDDfmt23ACEtDQasIVFXUdp3
x65YXj38OBZQPOdbbuV5EIHromkV1X443f/73ql16trIGSJ+k81cYzVOI7NF6yhf
BXCeLrkfXobRM3ysbdxmVaucPCloUK0tiazKJJBMyurD18fHf4hpj67RegPX2PRt
sbuwCtG11ty/TiQT0pHbZ2uyO4hBMRws4YiT84D622bgEhdo8ndlXX52VCDVmYqA
HiNpdwqfcr3NodMruqkbGt9bWnHpIkCF7zCMVYgUPnLn//B4G8Nwlo8GBGtxpiNW
2tvBlKRAiBSFVCse8eSiVvqaVUAuA7ZjmjXVU3JFl34gi73yPx0eWpzUnP3JBjyu
o1cfh+z2VjeC4+G7y7rXjW/CjPVKHw3aWYBfG63Vpwa7q2oS3ss4dFIrGg1iPfUK
h1kfuW3itqB3Qa5Zb/b2Vv8+5sXStrbFi1obFlMwnrffVr4cpjf8byAILyCUezQp
9mqCt0ALaELXZaIMspLopGTDaHslVANDo4Lve65kMgMJC5NBO18/RximB4VF/hjT
el/p3tt6bK223YDNcd0ZB1IWky/Dpc3Btgmm1s4VSa2TgB/lDYQ61STIRldSijZe
UYm08cIDszDQxA3HMf5QsajqZENAuDWSxHP2SeU8qYZYMOoHkenXWKxmSR7XjdRt
3on0UjZ3lca47Fq8bxg84dhKuXgcPz2B9YqAxtg6cPRvV5R1uS0aoRMkQxND9Wx+
jt7L3pwkyeF5eERJyCOjOAzD4GWo6sBED+cJKtHRddE9UiHuBr3EF39j4J/2rRYQ
Rf+cxLxrB3JewUHIqU+mwRJbxqeskrYX+YrMAwfCG4F2faGgVZP4ESMZbGllmAG6
OeFJIqGIWnZxu7tGXHKrGl+WrROmMJ6pNHO6xntrsPEu3UTS9o27ev8SBhjVFuB7
Q+qTIlm3ERrOM9s82lkVcx4HZyE6Leh0K8P7gfCFsUxeuAhmaJDZYzqw6nMgaNn8
Rutdl0P/IEw3u0aWh5JkSTInHmpMXaEAXFpCkym9M2wm+ikSIt2KXTjBaZYVqKGe
IWTCQVOIp/GVY7K4lCLDUdovsqqy5BfxRezGuoKo9QY3la5PlYH3ng61EDuqf+Vz
AI9BZJfZF0cPXC7YX2DujxuonIEbWVzwlqZ/1wZ9vLqWohxG70QQoM0ueruzbErx
usTOMQVtCL/CDgVIm4P4uqtIXjqFrvoxBSX+yOJG5HdrPwObXtPEGmwo3iAIBuF0
lTOLpCg1JRhND1uqOi5//hXbu5BC0O0xbfu949uL58Vn/eXPZ8zACtGMYtEyUoDI
xTi3oGFr+Qne016W4ebPybv2SuCv6r9mnL5pPvhBULIy7uNgAzOBGqMjyB/y1W29
oIw6RywtJj/1UcIWlTf9nItr9bmaa/ySX9bjXoy4iHNA1GMUi+G5hc/KnEVvovWJ
dlWCaW9Eqpu97ZmQINiYvEbqxrLgtuUg5E6nc5KKX/6cYysIdjFHIHIRVKM70X1f
Hoh/FV5fOZt8mWzccXQ6MkjNIN8KQ3LSBz4Q3hrQer6MLoOyll2FSx2ejc2kZJvv
ncGsnXvlNHratLr3EEt0pMtaIgMk1ZXr17KY45RF+lxjy+lVoG/gnieircd8CbnM
YKdgkkcDwc4JVIKyxD6rapY6LCUZfayKs5NW0yY1Hz+4pbMo6a7dvWLkFJ7JrWya
uEc/aY3owE15JWJ+ZnQq0x2HkJNcKPsmwLB2XbvoiG+NgKNCmp+s3xOecHKgGTYy
t4xdt5UiemWfEavY7BNK2lHYAsMjbnBXdqMDDSFeo2qV2nShrXq4CMI8kcMa77vb
xM6C1D0Aq7pB8HYRiaRPVWkq3iIIqxdbJP8kHayDp8qK0bWfLD3dR4xFdw523H/y
xCDqMoFa8VZFshSe0q2Rp/nTd+Q5HXXD7mXSECzs5kXaaUup7Y7riykZFIKkm7yt
WJ6OV+XP8zyCeVNIh7TDRNBUWOjOvz65IyoZ357cg99NuyMpSC09SM1ZzGTzP+Gl
dXpAaoUD/CZZyJpiz4fXZtBejoynixj+3GRl3KMw3IU4puP6+Nw3IzH1rRkyTio1
l7VYqFRVWrOXamJllmEjRR4FQlkqyBP7BbA68rq9PtXClIrNqPctXWwuV3FpAK8t
iLzhy/Bi/i54jDmMVP+DfiJrp98rh1EsvnMqd7flxPXHjRU7rX2OLr1qqokzZbXD
hYnVk+kBPHTIrK9gyK6hXvovYabxP+28Q3fVVN1EO3PChElYeIGv6jDzVD2FTYCI
82njlDSCpLlx89yvJn6+fgjpUUPTKjbv+3jtaWfY7FMU5ZuzOax3h7XyAZkWXsI/
T86Yptl2AxpYKjIYVRgdgvBJR4WllE6YTiokaiFgVRU39smhxZ9VU1fsuRaoOMwM
zfHJvRfEGqRlkjZ9BT5fi9QdjTqnp2YsLohgwWrGjFulJ4C1+2BenyoMQtAG+I2M
uSFm27gm9ooQuysXoDw7mlQCw56sicre/T7KTNxhEdhjAg0XaMH+we//Xmo1XpDs
4tKh/6p/KHibjVxKk5cyQaykP3Wj1PBfIjeckdBmArynEpshnfmUzIo1w2j3MgpR
b1gr4LlVyWW/4O4UPNX4CtAYTe2dIQEyl5nka3SHun/xn6iLODFcwD2/1Y6vPvDs
kLoHoFkX1hw2Tz9HbEtgwL0fxmiWLUxXDdK5eaJK7cQr0W/6J5p66V2QH4Ez/NQu
oGYL4uXoBTTJ71UDAn2CSa0UDhKF3LGSV7PRfOYhg0cbiFgRRI8vuWOCx7Ka4erM
PXuA5/aWeF0jflxJUWxDVAg5qLV1uWI1qy7RRgN86IkrtkgfpVNbmVQgwaMdQQ2E
IUBC9GxZmF3VNqHNJPl4X19gHPuKLCWeTnIvK1MLctorS88A9Jre1tPJY1sALlVY
/H6nBGWOHVq0ExY1XJ/XM59/QzX/vt34iMzieXQr7Md+ZRm0haAHeFdQ7YZ+vdv6
QAIE9l7vhia2cX3xDpU7wNsiZdZu3RVLhnFLLeA84OganSTmr9kfMj+bn5vosKCX
LvlQDNUWxUfetatF+avjeOEkRN7E3q0gE8OSwAypMRZBEeK2FtRVXdbjdnTbEOnZ
FXP0gsuX15VOjlt5F/mEJdOVLZmyzoKdoZSV14asEKDAoHxhsO2n4mEZFNWH8SIm
3qnX3oweTvy4EARMng85zFOM4+KI/NJn9VOLPxtpBxHHi1im/l8Tmp123TnrJith
NfVCA+oO0SDq4XkBM9MG7l1POLEKIA856e9luB/Rgnc4N8Xx+HL8X2dDuRwSNuHO
X20tS6FWQxGPYfLXUVnzixuM3c2jSaQHLB3rVLU7wYBdoWgfVybncrNaRJnjcwGH
N+KKD14tkPGcQG0EZ1xsEw/lc4+0/FlojwlrU1SkLHfqSVcuXdEt7YPXJXQRdSwI
JIzcmuX+klFZdyGnbuEJDy8JFZbS50Ho8S8n5qW2DyEeQ7SpHszPQiLmfGQoswBX
QAbiwP6ZpapLoCNra+RATnr0XeFk6j0HUxAVTc2SG2DFTWHRFsdrnb8TwtXxoqVv
7VCZIfSQKD4fUb2kf+X7CP/4jAC3EPlWq6rb0QVQ9+ZhIy8+fdDhNBhwX+BcFwBd
MirAKT2o3nS7Dm+CKMVW/uidd8M6PTvxZauKWrYl6QI718ms7zzJQAwj5U0kba2i
8ScQan0K2vii7twvwCfJzJG8wFrksS0eIyE+L78OnXhBO16F86176HdZ5aOXk//N
jzl7hfss6FYJUtsPiC1DOQIeJA4CtU3Yxl+MgAojFNq8bDo0wbYqm8vqYzyl+6xQ
7CrizqtPmTC5Biy1K4MnouIc9z9S27a10QqapWwRHbAHdDIbfgPujpKpdpOiTB4q
/ll/3JSDM3wCtr3CxUGXjChfz9LO+ZkGGWXQocnKeOafvsuO3QetRCygEfSOL0/t
VrgcsjM9a/kJJpF+Bd1KYgzGF+Syg7DC/ay0O2VJ08no8tC30vpML9iizSCc1x/K
KmkE/5VmBq14tdzxpW7aEbDm1iUB3jRE2EVi2o/CB1Bbq6Kv0TpkY9iAJqos2FJs
l8z621a2GY/DvSBLijd86wRwULvpYQB0e9MbeNZRTOqhrfc4X3yqF9pTP9JFTB+w
zBU76mrd2fgjIoUDCkyA9x+FGtalnzUF2Uq1gE43wkdKeJ8FY5pooUzI97t2JFMZ
20ZzSzRNmwc45x7Qw3rRbGxBMZWCrwPex7Rhl05FVxbuSojAlSkI6S9Oxj6zmMhm
vXJ9281KZxIjLTYy4IgWVne0KXzjrwHTIqW39MykqtA1LYilrcEz9dU92peQvmkt
mb/JE6NZS+tF7K/Hl9t3SHh+M1K2FTih6/jfPBUwXXyFmprBna+y9vRuBCKTVOeX
86yh/V7XsOJ/JLxcJMUvqpfrJio7+is5sCDH1tGLaW8FrUFyB6MAJePtnXMEn9gQ
v4tyj9XZ+5/DWygU2iXIyQcb+/jbVnqP//Khws6FMqC/UGpj1gDtdYXgHkpLnAwV
5uj13Ky40jCTbpEm8Drkw0zZXIJ3vInWJBuplRTxIWQVjlZj575X1+H88xrHZqwp
e01rud00td9ew+tcgMilVcztqscVpcFCxgbURrD2+Rg9a1ZqxxQIC2xh6K6+Ywpj
KBNRwIVAuBpoLbGwJpUcnnoab6pXXNiqGfaeiJIt87ry3Ctph/gOZ9KYmhkbourL
fY5X1DDgzugyNzcdFZEml/hP6kVNZ/2M/MrXs2qxmMDFXaHy29ltpVv3228YU3Gr
xuSsHGwgRfaMmSkFsKsVTSJ67nVFGCEuMarSu8hQGCeMS+8INorOZQP7LxvHvK2B
r9yVZqz7y2tI+eQXbt7aS1kpHYBAZrla4SSelMJMa41QaTUOx7QXlQUsViy+kIJa
+nln4FXYloXsA3p9PUB0p1ceXEUREam67V14wFzzxRqKs/GkKuNfDGW/ouFf9rwc
ZBfJXVoiHm2Glv1hcHxEACNs3GEivqEP+tC58q/HXxGihg5hLM15wuTUhQAqV8re
ioFCfrlmX0jXKiOztYPD42i06HEMTH3VFo8+Gt5Z3vK46avBiAPWMm7IDg17TJm3
LCnYTHXEeFGWAIq+/Qh8eptpWR8cRLPbLG5cVzYhHGslYrKYl8lGb2QBZ5R+giQm
dtM1ws8jxfjUiSuLsJ7zMAEW7KnF62nt2cX7nSF1CAmBkSOaP/DrPyPDNW/327Wr
HHH2/6lsz5DLevy04IW+rTRKX+bHfX6Bzy3/yjMumFUFYf6xeCisdhkpC/RGUVPE
xutIh4mJign7xFA4QLkchNE1hIJ0jciX9wLBG4QhVDNnQPA8b1+sbe5NYEktrnY0
By67LdxGR+wEl2hsucvOcLXJM2E3ysX5Tu0PHqN9L8rFZxj0kGHfujTRkRySe0sW
6WMw5oc/2se+SQiQipA1w4JAEuFzdSzzzQzgyKUEA1vkzyg5a+WY6tpeHljyBlHb
mers7bWE8o+9P3HGvOzUY7WNc6ybrYIF6hrC6J2zFOfC73NY3Cu4EhC+eJb+yIaK
UsL0Yi2x3XZDX5HOO2I3mSO0p414PzgaQXFLQ86NU26i9oVZ6pNRi29cSMSeBavJ
CRv0yBJswNiPvd1eXdPHa8gdSuRdkcK9XInDDQKregr8j21Ncvkfx+aD6qkOAjxa
IcRjAm2LJJpI643yFnu+NxlAHEjFgBKiZXo0WT5dtx2xuFnvm1gTI09J7TtknywL
lrrWf8w8iBtrcEgUsujx2+r8713XuA7GkOnvkDVxUbCofeDpbLRku3rlamk26/E3
o6kvvjMCKEhSL2YGlj7OeGwLdCZylvoNmViPBJ2M9B+Iw+KJ45o0uFlV9wnb2Q6P
kQd4cCmDcvvleVT9G+IwtnwRDHGVBRHRZKhuq+fPTq2MmeS2B8UH08guV7sllGN7
CYl9W1httnGiVW/o1HtSTT79ch/Cz+QqaGZoOowOMY2mcF1VG3s++N3/fTsVB7UB
pZIGFHiJ4v3g26tkfpMQZTIFLY46tNADyBuTUx0/vOWhRAs24Ctypm8DhaTR2PRm
azBG4uJMdg1F3yqyCkanS87u9jplr/4akWBvTR8xhmkIH9iTHAlENqhrg3+hhk3H
gRjT+wy5+6raimPZ2klhdt7eGmX4vf9bToXVtU56mdZWNmj++70IrafUC8hhgWfW
j7Az9r48uyrIM4ulkNJCbRZUeHky+tFPSusfM03W22b9BJc5ynwpP9XeCQ83nXJs
0tAUWzdaa5CR9M/fZojGemqqTCcASqM8g2XSMF1bS/nkDQh9vxUgGloNB0Tt8M4h
8MY1CtIzMMmoeutbdrgYa7yK3nhZ2NOkk3dEjBX6XDAJj7Yo9adYIJG9DbrfHP+o
hfPGNAQGII2yYJ6V7BzWHMr3mLZK2L/FvhCcaXvX+xyaGSISCkB3dNiG8iM3Ni+r
owAKOvfFuKKFU5G33/JDespGDtdvHDHPKn/n6q0hOuxkZSaWNrv2wFs1RsgH3rLs
O/aJlqGnbB5dejaff20ISdiv0K2V5qwGWHhvyI/kTDQ323KZPnoP7Sjcj+bSJwV1
04hiprt4SCGieVQSgG7Yf2TdBBYR0Eg3QUM1lC9FYNsq1NNfG296Mx5VsN0Qv+78
oTwNP9+BwgnQTgLM8fK2qFlSU+0Vi5sNwfcakV4/2tNZD/2FXls9UQrlsJB2skls
Y8aJDzUrHYgg+B984MXYRc07IE3Q7cSGXtjGXrfKS+bTAJ/Pn54hDUqq0FqZEUKz
vFdLoHVzi0BQqr/mIZu/AMpg9YUXHc1G8qasCM2f68nBjYZSo5WGL+LsOy48Jp3R
21+qcgQ6w9DRX2zQb381YbuGileddo9NBbXjbUSG++AvKIc7mY6ikQpbmuqkFz3G
7r+UWvYg9mF30+1NWYMao+3tvhBO9CkVgWc3vbhD4mcFle7ar1cgSu9+1LKL9foi
/43MwAmoM7+dxzIqcgUYGTYGwbQzdBzy5cdBYeKQeihg4T6k8M3DccGaXSk0bf2R
piI3Rys2mwFZCYfhDrT0Wpa+x2wBVV7opKFxFwOvQdSh6sbgehUBC22dFzlGEbcG
xMWKo3/3T46gkwQEueFCBsG/MuKmC1AQvaYKt9mT33pPWBLmqCUQXQ8xs86E1BK4
/vnkSea/B9PBxDoE/2MnVB4RsOiddMhSE7krdNJ/3QETG2raoSsdrsPlUkpU7qx1
ttne7nu+AHnbB8jOtCf2hIJCY1z3PRIyrsZlahdy9K5q950CIsFeWAVCpktRotr1
9B0Vng+i0PinNdb8Fx//qkEe1m7Q7RZKRFzpUinwL8fWrfhCEuk3jaIqk57hPxrD
1kSoCBbeBlZSOsg7i5pJTCqL+rzAOT0wMxwcOiByjwK/ADpvMkSXgqw93o2kCzp/
+VPU5LL5lD5gGD0tKhZes5a5LhYfkENfuXEwJnwjZGwKFXvyG0PV44pRD79/csss
sAc2mQrBhbFZv+g4q45NvSc/pk50uO874dc01zmsWlsXnzFYTgCaU+UxSkXT3Bok
I15gJV/Cl+nRswhp55EfxPR4a/REmkgd0yKHf3wZ0dWVQ+wMxbSD9Zrs1cB6fAH1
ojh/7TiF1NxQb1Opr8TpZTOKGuBqB3O1Ph01lMfbt5frnK7xMhi22rczKzQLlkig
NVUARx2NjFaIYcn8341yosATQ2aMCyBS7x/AUkA2PVRrTFF7BeV6b8WiW1Z1xqJO
7sGBRb5eqNNnb5LG8irk7PZmrtIeGCVkwYuuIVSvrwldqj+TeZldfOykbSwaTACw
JNMekRzujLaO3DqAn4mxZcCOjfjhmB6UJGwXPD+13mzIQiGOTNQCRwIf1BpBR8Nv
pY9xgZsJLycK+KtGrOuvmDtz1IdSnf8QItezSJKPlE9VPuKhfWvncMoMde8B0YeZ
zbEQEgx+QWmmEh7+Frti1Y7MXxfYKpml2fFCI9iUFB7EentGGc6QFauqHeXTH6Ik
K4igF1ofDgewxMDe7Hy67o+OQlcIXJO6AjvF32XeaNOBsrWxUIUookkHoU757U5v
somUBEIRINFJacMT00jeQcGqEz0WN0/zmD+iQy5HZIr1XEKfQZ7LBqDiA/ETxPgX
pKnVWozAYISXtT5AlpNCa2tiQLrz9ZrLD996ds0qDLipILbJZIgeaDut1XAjptNU
w6aqNSJkmECixoORtqKgem2sXWAt0D2JSh3XRzLWQHg5kLHhNd12AfB9Tbt+aFB+
+uMGCgZH036Ie9yRgNtvVEBniVUpK8Tqms3hisE7RqNd1UfjfDz8X6+YCxMDGNX2
d4sVSIbj91ylzgWJKN9Dpqvv6CKjuG3nC9WbhDf8zmy5wUkLdlNrffeU6Kne3XdV
jTfDSmW1IRbFg9ZqvO0ZE4H3WzmhljEUuvS5vt+xRHjR92o0Rv/HK65Xf909amUU
zWWFSm5vMpZZWXJHuUPtyrnZcOg1XoQK/MWacbvcYk3rJpkSFRlsuIs025gjnqWm
hdcgRHF9YB8Ia1X06UScY9hJXxklBVFYmdUZLdGZ/+MUNwN6O2pyf/kNptSc1s8U
2IC0hY2m8hccHqAoEdQZkvQeieDBKxjw/iE+DJVonFUyTB55IpuJvon6yKqe6bJT
tdTuasTtbkhNKk896hAEeOvuACGER7M3LeAjGqBnsq+yJJnie65iMMkN9sSbwOs7
Mp6QWkU+I6sCBAqf5W7A+3JUucrKS1i4p+7m62vbAWvXZfSRnWIogdD1RZ2LelwW
20wmXM5Xt8GjLV+ZkAtjgKiiO+lP5jju8MY5aKypWVcXVgFSdg9nsue0WO+TT36B
pEqH1d3SjzFEEnK94e3DeUhIa1tYl7ViAVO4hHqJ4YT2pj2nsy/YUm+T53rxJ80u
CWFUJgU52S4+IL2sF+pssN95VvfXWQuL9U6ZfkJCA0pNWqu988aVRSXLifV8LaZY
zDq363sTH4RcWIpPKuvpxOvH8zdFVAjyBNgw/i3PRqygIa65Xc1bL6RGmxmSHZCh
Ol28o46ZpziFpU8LOlGImJe2wmZ1KiLaLWGtRsthFOobTh56TOrk84O99YlOAzhM
XowiNvuZL594gvkXK5tMVSIW112qvSRltTCjlmibOjZPMf26JGidrbaf0WtQaRHw
KCUpHHLom+RnOyb3lRCNIIRtTjn4MRO7kztdNcImgautdfktDdz0GtXgV0kmV4YI
DURWVY50eCUANW4edlYjub0ZB9HESd84yaTOuCW5rFOzlIVLvE50d580bpVFZzbZ
NzIcdFC3dExqvr9w9JVnJvQVueTs4TH6o59kqfkfrc0/qAPG1/yIfGrvnNNvGQbz
r16diuHg50gFBSXyU/vEQY9dq+NuGXZPNRaOX80ev6v77Vz8FgP7giWI6ZcIKyEV
b2+9Y7l8lY9Y6SK+Z98FtMuSm43eDEGnVzaoY6pneGEVhbwfBsgzbxUumkte5V9l
P1kSXAN9s79YOqiCcS0A3J/Mh1B/Kx2GlK7/kcTIEjjj4YQOgirMA1AtU6K+vFlF
7G7lEi4N4F690FA5CJ2X4ZukEflBg3nSZ53cC4hVgZsQkTD2f2BHI5xzP6Gkk9wy
Z2E3XwdzTLRW6LlHiV+bHEjj2dRe1liZxjgJhVf5id6TpO8wTFETGmTjAXpTUscE
p4un/jf5eSnSI/LyeZklGjgYpH11WhgebRqD+udVKACXgPSAY2lbUv5zPQA1p/nX
9gBFdcw4VfoQINVurPrbKiQQvr8cbHW6pWBdwYfiM+oYvBkJtKLNt/dItaFNUKUF
N+zFvqxUt2GGST4IaleTWS2YvAh1Cb6NOqp7foq2fRJ05L8RK+gbBhg7GAsgzGDe
QJYzjWnjjeQoQdC7yOooaE0VamPR6rzzU47qnkqWDL2Np4TS4lOSSzeKGcxfBNL2
ticoav+U/kds1oJ8wxn9cl03n3Rvlru3OI2arxtQ7Gig27huKTBDKgefPQ0c8M0E
VLKX3M2/AV0xp2Ibg5JosXvho5PkpXgZXbS6KO1lM6585L+65Int6DadVUZPqcYW
KY8v6xLAfBDp9q5Jy1eoY93+Jeb3lGthidTTqc/C9xNkNWibK1rl+5ja+0Y/EMGm
s0pHuS0ZLyTG5+4MgJMV6NNM93kPh09O3N1bqNpJHgbWo8KRRKNRa5CIRZVWZSQL
PjV0lXEybyGWEz/z+eMCB+wLRrjm4/U+dv+xKKATUuy+CzfDiLVhVvmUHR2QqOBi
LHi4i6Q2YhbICm7xmIhqn/UDFJ4pR0g9hI9dCaCCiFN3yickPTkPbpTry2P5+3tF
Aay0Stig2VlN5+Fd52pUUnomHVGWuEwa1rtNIDpfLX6OPGfZ+jVYkFpY6+vpqCKL
YMGjfTo493n1axT6kBVb8d5dLooW8fHaZE7HEcnd4070sak/0D1IkBhs04RzhyJ+
s0o/Fld5D4XHGyjNPw3oVM5gCAUZP6jg8H0FPP5dRVr9fvFCWUNJVAjH/rG4hKKE
rj1qbcWiDecsTqZIE1QNb1G9Zh+dObfctkA3aOhLKMZlStlN2CFdgn15dp5+RqUo
8BCxsxVcYQjB6T0HswfkIhJc88hluUlp6IIKti9HbH28kNLPdQxlhQ5aEGQhQtX9
/GqJrW8zbGSTS86raDI5Hk4ZIESoLLKJYYfETz+cepIhs1ozVjRXN42UD/wscPQE
DZe4moq9eQmSAYMyA3zH3acttsRt8QpK3JWGtEIFMyuJ+wIkg7+vAz8bKGzV+0b8
mzsnGP3aLTsj64FDQvToVACJ8j9ubsSh5f9gPHT6fzAbIf6uAUUbiIMuM0Akejxu
1C9y9yRz9eJSjFbemS744Uu4YI5R3tZDcgA3PhBYOVjOe2YJ7D+Y50cYblXWcZXp
fgrUfOq/uUjIl7V2wdSVAUgnJQeZXgVu6NpbnBQnbSbwTrI90+jMHh7FxwL+8pEH
TzFmMsGRQ4wWlo1zsF96Y2VSuxI5YyzdhtsQO6VyHXC+UhJk+IGjB9q+wg9zLOJX
Ga4n6+0FB3LQTZ0sVqBQ26p4Ehs9GKmLbO+3SVy24CVKd67ZBXok1JdBiiv/vzMh
22ghpuocyzJg61IuiwebYktxhnx5hz+Uv5mmypqbXfOgX5EmbncJm8lP4QzXvwmI
tuAttsuCBRPkckSESaUGTSMtvu4pZIudULPXxDBSXUpz3atQ/em6V4H58ZQwnBR3
yICOmkBZ02PMICjH8Nr8r6Nv4oJuFDNqIiR8meCjFgBRuSeS4BA08m3Jkshj8oEP
8O6bIHVtm4nuAbsbqEBN+WT8K5Ib/xSq5o5SpuM5ocoOIUZCwYXNmNOjjMVyBlNb
m3Ri7OfjA2B9Rre7x1y7TrVDPsR7nemNM9TP9Dm6vhMNBFg6URbZp+SipY4rquWL
0FKEFBcYAqC0XhLcnS/EUlY8nAxo01zEc5Ae10FkE7EbqvBSu7WVAEAJ5ZdsONYI
Bf54X9fbvYQvAagSfy8Tp2Ffg1KZM9igkrh462Ty4uiG8SD2LqvFa/4nrycPUAih
CUwdv2bL2hz+HllNHt0bRm6nbrOLs3ggzznlN51r4AAsBvbZ4N3HmT8dfnya3CiX
AIn8i3RFrRK2oGBnN/WfqhU4nu9Cxtr+3jeMjJeXuA7JT9URkLUFdHFeGkmtLhZa
SueQEfEswZy63V6uybQDxknJzGVc03SPRi3qliG+dAJk1wAAARd1y2Rxt/VtXARz
u3jqxLgiI23+EPp5F+bvLQYByhOFUJxESEAVHCbLU9JamZ9BJjJKHjUo0iAjZr3i
LVSTIwh2JdVSdMD/9J0g/Yc3rPcFSAgB07ZQUBLHQttToYwv6MsFhEFi/yhN1XII
NqYsGCWWccUUs0H+WejlO9og6RyGiL8z5HX+lvqFUaxPe/gfKP92fAuFfwmhm6ti
M6qB4k7HcDVMOB/79/NSnFjIIpCUV+AQMjtR/79zNp1QeVgq0qyS8KvYvGpgKv2u
KW84FYcQ7mv8hBTZQalCn+mltxV7OrKSel31O2wSkRUAiC5eavg4tnfCTwhTpKCA
JlIsSdUsXoRIPqGqmndkCb5QqcmkjpRXurd0hbaQdCueAQq/P3tarnJuP6hphHHW
SR6yBg6R+90Y2Ye1PgaQ3lgUsYCzqZ7YM5IcpI+DC0L5vAktGwzfjlk5ZU6qqvNy
VNn90CIxbKfQaej+UaFLiKcdZzdPCO3WFFdDC9gZG04gXI3byKheg2QUQTJIYVz4
uHMtQwvxdRhVwLczkfU3EqP1bFr2rZlP5dAq+5HtDjEH3zCji12MRmOCi8hZfXv8
/D8McQ3fTiuktL+bJTPoNLDSfSUa716iyaRFgyCD8Z9NIXtr6Ht5hPdkq17crGvc
+S0l+Kth4BvwOMLPys31saQ7KZomMHfnA+O8PTuCDwFSrq5FIMHL2LGlsQlW2dnb
BNlPgTWpAs3eyCglp0HloAamAEq1tQQT7xmGqV+XNujfAsW/SOY450FpViWKbqZz
Rr8Vq+Oo8iz8s/c3MI6UOuJmqlec8u+DW2BuxCm5RUHRNggmV6uEdEupxRT1rFdU
ueHTY3mH1xut1LktTsGqPzLgZK/b8LEDzQlu33llVb8zM01pH6EEyrD9YoYusRd5
AHZPvAFt9gajzC8r38ozQ9E2Z5yhLxFn2SQrDVY6hPnEbedU2WC1rChw8v49qc36
VZ9g0m5m3AqgZr0bj8MiQnl08GW1SMBWXOHPrCb0eanj8wXXqQFO4iz/ejd/cmeZ
pjiV+JxVozFLKlbsnAhz9eGpg/nZCBSx2evXf7IppJLrGzr1SAM9uYexr28HwBa9
WRf2Zs3yeuc+b+L9EOEC7rT29X4BfvM2FgYAqwUUQ8a7urQfaHydqV5AotheQjpJ
xXCgBVvUwTjHFSVHUQFTyhsgKiLGi9OgsT/K7Jllnmo4ZIYk/1BcttHKKA7Ulpxe
XgR/jmF/xtVBsJoirxYrqc65RUnQy3aArgc760UazlhhCij+ycws0jvUbVVZ/ScS
fvoIl3VuzUiPOk6BrqEbiKdtqtEckq90yAqlfKmx/ExTWs6TBRsqZDtyPpo9Epee
ZGYOqcDcazseRrxqQa1TNQo7ya3VBYcUY4eK9X+ZULpHs8cd8EtTKqD1CjY16wAm
j8KDSEdzerat33Dm1x9pniwkVOev/hF7vCpjh2YMzO7lsGUChFBWdnQkBA90Wn1n
BWKAw9BbwSioJ972ZNWPZS9ux4CeKB49wyXShOKI2hJsYYov9r73nZOORn40s7TF
6IciGj/2mKzpESqow0qetw6bZ8Bhi0AU4h4UZIeacK0RI1jcVBhshpE8vJaH3120
I4Z9bOuozcZCXxm8O4zkEtWdT9sIJTm9yJJZsByPCj68RZZEwdYH8dacKhGV/gUl
r4yTFCysuDi2aeTMiptZdcXIjVcQDnNKb37tXIMfMq+O9BKejNMEI/7D4GCjTJlT
SdFGQzlRnt9Y4rtdzyYNaHOLjqMj7QNOkFnDRB/7NHJfjhqI9JX2q9VzBPXDb7NC
AKXpE7BMBuiQ7L3I4v1jAQXee83bHGA/nGUEwyqRosy4GjvZDn0TIakjMAg1j9ri
IKTwQhiv5RxbA1rFL0DQJT5npG29ZSwwdm0dklwvbN3j19kuYMiudL5it6Sk5yYw
uQdAhfh5eH4XIoLMOfT5TftncU0mFQAUJxGGd2ESOiliTl/obYRjPOd6oQy0Zq0j
uPM5NGR45ccE/hekmsxOaIMbP7gG5oqglkbOY7wmPMN4ZsXQmP+O5bPO1PpJJ9ch
ebz+DMo/hLXxbiS4fcHJBSIvbMVZ9H0z8BrIT9BfvWwXzg8plpMMA1p0MWeGmzJN
D2yl2fXsr4YuuNnQHzPOeVyYUIBPREAMdo0gSseOqCyLJik/9bsPmYlUPGEn6eTW
UyRlAAOwibTCSCLG5X+wYaxg+ecoAlB7P4iOVsWIJjE0RWIHKbdKbO3X82dIPV3T
/PZeIvJxcKVQt4OBqy+v4G+PIhnffHMH/4fsbi8kuqfKE+RqmODLV2GZxpJzVtHd
IafI5O5fW+gH9Q1ZX0j4KQ1LTLYm8JdP9khTMCv5ryljDo7luILvHpGQGUqYWqmm
1EhrNZPP0bhRWz4ZM+2tP25sP6OSOpl686H+/ekNNtpHNN7LCAGYz5QApUEUb3ph
EpjjQatquOz70VFu9Oeo/x+TTa+nbfqMMwTVuof8eFWTFkNmU0RVy7U445qW/IRl
Y2FHY2aR0PjIakZTGyu/Kz/RpagNcNDnNXIFgrylfqLtZxNTbD/u0MbIykIFCupw
xKM+q1QpJ3n854B0fUpQq9WeldfJOD+0GHrT8x9Sa+B8O8e/Efds64aRWeVm9aST
newtgaJVtAO0gAqNAvzlCW0tMMLZERKL3zxpPyzQjB37WakNe5/V86zbE03bxc4R
neuwI3Pbs3WJg/EgMfQaa8+JeE7hzh2IHgaOcHoEoj4kxSZbwbT3BU8hF75FYcVu
Sw6oAP74Wo/nP7C9ARoBvMvdo8qWaKzQLWwA2DrPFmfHjbBbiQFkP34ACxuAwF2U
ezhXGo3fr9vbjnlBzX6J0gkCoFGFwm8/rSnFJlhFG0SpOLycL4clRK42+Puuudp+
rhbQ23ORc6Tu9QZtKrVzSKq9pcdveBMDzmXR+GPILcvMBtpWEqMGXVgKnuC+MgG+
e7Etype9WoExzi1jlYVv+MOGcsiEu/ioEXSR6CLO7GhH2EKlJGfRuRDZMQVNEgCH
0kD4A8Oj7SCq+/4X5TEofEKEHApIJ+ekI9y+7R3YVj8yKavY27ExtZsDCWH7nVaK
11fEnjcwazbm1VIqLkCJmPpUk3C3vgv/mMZ5UORz90v0NMI6cLJVwj9ZRefE4MqC
7Z4SYpU3QjpVZ6Xx/1gBvvTDxTzS9gN8NReyE6Y7lH/v8JtrGx+AiSdMAPc+mE38
fr6gezVP5ZhhZyXncm6jqpVGygxhpjCpoTtkcWQuO9uZgj8pGPaHXgMeW0se2Mnv
UrElE3/5XSbCle82wkaY9jbp594rkSfbUA8RsFjVVLSkHm/zEA5buw5UmqC4/UAp
4wXUwuO+TEYBPd96huJSFu9itaGWED97gUVoLUqEkNngWSGMKCJEHGJADclzr9OA
Q8v0LbX8nh6P4UaQz7dpGc4Qmef5XXClhluJbdOL+VO5GH7AYdf1n+9kgf3Z/6Nm
0N5FNKH0CPOM/+m2uwch6jBYWRSzJcgAdfH+kREFaJxWGdP0/uDgkVGtCAitjyby
G67LR2mWABaAh7yTIjoYB0J6XJPFNjz142Tnd7KLpqHvLElCbJCcjy2mukEmXPtT
/nyvxkjgoVKhR3p92qRwCWndgfmpXC0+RC+4/n9G76avge0nbl4TYv+G7t65RDU2
WG9VoUBscs5o7s6olLU8KuLNrfXJatw8GxQP+JG0DFxM4dlvSsJGHq+JwWO6e2rM
G/j+lF5QSKNRJ6XJhbb80Vnh4+cA0bz37l1/BOTnryv5T666pqZSf/6ptCgyO8SG
pWIttnz9TTMLgLoB/qMrF+qmVr34vSDU6WgnipNiMxK2RKQA5prGltUKyLRMuBlF
4fraOTcRRGzk75LNaBPqsnNDApPoj3sMVdLc47XYZoBVUSI8Qskm2P3rnJ5QzsbC
u43Yn4wwmL/lEfYHzCZNvnRb0m9781Do7tp7CXUbgXl6RKmmZnElZqB57VpW7oV7
dT6N3PMRn0+syONwWzwr0LbBE3kjSVxPRdO1KbczZuGx9GAc4bOrWaWajmOxRnX9
K1joJ+Wwlup2b8O8FB51TxCvRJyVE/8tJsU86Fv1DFD15rEMrV6faUepWRBEv0VR
ab1j/n1QKVWWmkwnLcSmYaB6igCi6NJdFC4OgXifc+2sNUEmtXd0zsMMmN8U19Ul
W3pNr7B/OIhQMP0vV4Lqy/zim/dMBXoJjy4Vi2iFv+aUlC/Op3PLY+F7mOQ3tZWj
y/USzrHPJn61o6mj4IA2BUPviC3Z3OsXg7XoTHjJ1cEKRlTKDXcevRZ8F55Kreu/
8ZQbpicPqTDko+5RcwTicgiHca2Ek9Rnx1+73YqhBrcBWpM1r3yVPOrXbNJ8kbM1
C2L5jqDeVW/ZQimdh++lxoCU3HnwDRz9Qxwpu8RDP5U9aQZIInqWs6E+21vFrvIn
2yH6KR6yAdaLQHFo7UekFen5X7WPhQZg1VoTjdEgNI4Y1KD7QFELnHzr1JyrutWr
Hn660MfwqbkCYBsuwRV1TfDQZJcHxdbmZzhnjzE79N/QL8o+cUXJpTCXdleFN4sb
LnCDMhk0OS+wiShEEt7zxhj+njFsxw0B6XCAwhZPr/4SQT+4xrOeO0V7jVW7XN97
H7ZkY2T/vheLn0zX5xtX4oCeJlt/QsmDRiqHU83KFsLlDy4McR+UmheQTSIxeynw
/yJXK2WDTX8mDIRPUCsl9VtKQa/yH2ux+NHs2fm8IbgUukz7d0gdVy58yQVEm3QY
H5LMJ9WofCtsLsVxrH8JA+5IHkr4bGpwUDPxDWuvCj1Ognf8WwuR95kn3PH+aW53
HaITQ3cYJhEiFkxOdQxTLKLkn+ZtH2V7VzQ1Z5+I8/I11uuaVon0fHVyR7WjqQFQ
um3YIdq95wH5kXX3JE4U5nSTjKF0CXNYEo5+OkQl98KOI2mK6bZQ8lLesgW40w2F
JiafXI31rH+21qwyZYtwONXhERxFRjJZyNMK7BhFKj9eZUw4tMh4lVI2kATP2uVh
ZJC2SUu/ghHTFopEQKU7A3TYB2aWQHJvFEa1pJIu4TEUOAqB4D3mlSUeUbG+uyEV
azLb/kEirofG/Hfcm1vVUpUoJ0Sw/chvjHlD96WHkRYZF7cBL2/7Sh+ozXVGTYJw
6RzX7iZasOE1inQzDseGAIG0KwF8ohVhVKNpSwTSqWQGdsTc7XlEomD/kuVepqZQ
qQMcapPFWys/uNwUADMT8/hcJ2jAV+kPwOqIqQ+IROgiesCm9Fr4+psHP8xGAg97
XRZ4CFCvfKbk84dSj7mno+Wx6uzZ2ifObw7XHO3e8fWgsjPXe7jDxzMa4BSM3W+5
Q6JPBC//vcobNlKIYQNb7ugBS1VTY5LFuFm8R5NlyISGJTqScv8LsrV+7xIrpAPU
O9Iiio9s8x4y9Ws/xnHby/nf4orK42U8zwQHoGq7zwCCTr+tOZzFrxZuPk0xs0pM
JZ+Kl46wdxJygT0+GcmkkaEc+3BLmXIFJgiKRfzEeENVxMkOqpGQ/6YVy9WvHEot
tIPrMHCqi1ATByVKU/ddSsuVxpfcf+cti/m4q22C+9jj5Q2JQ8sFVYoVmGUtQzo6
VLfdsxFx1U5gM4DvLbmg3vb2mJgVp5wK1xGspiSHTxv7SRVgN9R+t5CyjXvV9ydD
Oh0s/1Vo3f1fVHyuVu1PMPCkTtJkkDtpwdWVS842QlBFhmwpE/xAM87cmMmrHLEg
8Lt7k412VjeXeDmvD1sIuhT/NbMY6xPxxXu7jVvqoaYsoSydMk3Kbn0HmeNdkOGl
Ftv1q/whnGXC7MLIiY6c5kjrkUfpVmfPuJe5vJhPs8IKrwkNgqYJBGSWrAeuIXO5
DOEelxpSK7Lg3IYPjKrQ0/g/HzPKaBB/cSiciwI/K0r7UUNahaacOAAAvk/pzLCa
ayZ/m0aBCiyLEex0x7gj42lkha4BhULogEMm8WNTY4Fmei80QWvPQXHnUlXFT3Qz
9q94T+PKiim0zTrv/Ped0L2vj1s1DCen0AzCNiKuA2/fY1hobsXiEB72pnUm44eR
4bDW+/E0oHMiTJCzH2lvXh9kgqS2g9Q5KVKvO7nYAu/19zdcishoq38VEIwrGiRD
SlUSln9Hy54ueHyRVHu6XuNDwOXomjmo/Ld8B7r9VBO5SSYJU5UZp581UWAJ1hHZ
WIXE+5TA34u1r7KjkSqw+OXLgK7/a60OBkMOWK9RJUf0r9Uz4XUi7XK/EysYMxOE
3CGPu6hxtgiqSeHZakSekP5z3O20CXU6eNkkulfpXdqvfv6KAHQcOw2I3OJwCRb1
lCbaTsgbDTdGqBt9V4CjTPppVda6W8y0hOso1U39LcYH8IDvgVH6++k7jRIFhZWo
LdBW1YFCgpPotoDfGoXtxCqYcBobER47b9UOMEh6e+f+XZec98Q4HFE6xq6AWAtH
4vwziirGRJZfZ8Dly5Dhq6jYmdvKErKA58oe3SM0Q5rD9ni7X3MmIZAIWmElmL6V
WDzTUI9I796Qf92gga4/mVrLJOhkJqkBZOUl1MOHrYfLNJQIdCDwUqaNqRdzCcqJ
3CzQV5X+P4UtqhrnzL91yG2kxDk4viRI0BqV9WjFdRMSdQBD3Ufc7kPwizX8393R
CUGN5OaNHqh2fy98K6q0HIqGl3ie7vEfFFtKZ85yTdo9tRh2Zvj5TY8efJPPcDs3
Ge7ZPbJYZZcwqIM/f231qYjx2MAIFFDV6+7BE1VALTt0qUUBkzyi7nh3Z/vPwH34
9695OVp5RGdfs8J+eSFDFh4PP6nALggKZzMn7zETRkBOis+VlDarlyi3BRPnj0NU
GCs2zKTcn6jRqp1Xm+ZRxOUxAkI90UMnAJlxLz6t5QY7zeozHGuxi7M+H35QDAqG
2cQAy3fyummsfE30xADaoqdqjU/zF/ekWq4mzKKTZ38epSPq2lTr6QLAan4OA7q+
W1WJbYYzvVb+riICpXQKMddaG+t1UwYmf1HYK1vcl3mXyAyLShTtrOJhqxPlSmQw
iCO2KqrjySh9Ij9Tv5VL+jCOS3s5ntEXnYiyCaCrM3tFtxv0SPc6ci2AqYnqjVHM
TYs6uUYpxR80MMyWcxM05s5cHEK/kSu3Ti2emPmDhPSphmd0pHj/dQDElMNE4l+y
tXPvCgzZpytgzxcM2lWAdug5nKunAw56QecOsNtZWBHOOMMX3P/1rz5E+AT9Y4At
HHSiTIPEFipNLMgq45W3QP5aE39yFso9aJECU1f7N7v3X7U/P+9T4XAuGSSoDExe
8VC5LyjjRhW0gflIm87/MQe9bGRDy/dXez1+hkeaObTcZ16wawudMn/H4fNMclx1
GCGkWsiDKcs5zEMN8U7ArAQMlVyBDz202uXQ3GftN59gWv6yXFmo9dddE1Uvj7Ls
n//OcFn2BmRxrLC11ec7tYcP0A2l4nkQF28SIjoROWGooPBIhWoPJQ9ZTvCUsz+s
G/zhpxWtZf/yjCKeiX3c1T1XOcaZxEgGhm/A7VlYVPFp0qLVKViI6SbjEerIDPSX
XfDHmPV7UVtTnqityn3DrzA8ok0bBf0HH7r0Yz0sXRcc497Osym48YTlmSZCmS+B
FCw4S/SNGA5jP5ZocAW8DlAc0/8q+8Y6v83aMbVsREgsr1s1vlmd1JH6jWy1pZL1
P/ybr2viGaMHVm0fXb0o+BpuZhl5IPIOOAhPwDxawa5jqlMoulzmeGXZOcYq2o1l
vKTleZeEKhqO05wmLqxwm0tA1J66Bx8ZlB9H1T+4NzCmWQuCf29nIni6rDOnCdOY
H81QDeCt93XNaOILcor5fdSIX9+qFvyrghyB6jZMhWlOJ5MMSH5s/ulvtVjrbfNQ
8UWdXFx7KDcK+iyNzecgh8BMbbd5XfAKPEDWQOONhhYwiw88vUUtVNxLwyVtC5Qv
5M+bPCfraJnDdDKB2MgT+Ki6Q7OiVnLq0P28BqDhgfQX7TysT0m2475Cr1F/cYfg
xMfZk+PONFpUMs5gFVeBXePEc3fkuLzp9pfkzW+sI1HrX5CUYMhqnU76mztqPfnV
Ubk1FjkGdKhqkk4469kyFt3FyA1AjnhR+8xzwr3CzqX/i1VSzAsOpeJMcdHlFsVh
PD+nt0UkES6S5YmYnXxmsy07L3AFIc4NVlrkzA5Lfm8s/X09avGgni+HC0ZxiAXK
+tv1Tv49DLY/q0Rw3wR0QgMRgLtE3OrH0QixdpHmHytRaFqbDS66C9iBphYSJGDL
cA3vW3Y49rZAcGg/k/fPnZWqghecLtEfGuL9HMNhFfoXkIuf//+sKBh6AMHOthHE
62P//HftXmOuOVgBFzTfanpkGhy3lb9Jf0QyRV7MZ0xI4jmg1U6gmYHmqburrpLB
xn9oTNoRg/cxNNA2cGDxfyZJft47Ap3AQmGo+92sdCceCVF0UgzvC+b0tzLCb+GZ
qb60KMBNd+mZuaalMxxveeCqqU6aOjp9MttCJxhBFIcGK1uImdarBEaNfRMozMdb
GFrOxwEUPFKBbAIFlTytUc32ItDD7q6R5TaOa+BsPLFKQJrAAOL9usOX0mP2roio
I8ne04y4zRxMXyTAeeL3jr8CKrzG7mISkAQxcCr53S9etaTY9H5VeIZGy5L89amB
htyBrOYjsmC1yGGen2xv/5tjoU/82EfGyNoU7KU5ltV4IVCL1jCqCn6WYIyaDWne
8Wq23ILUSXM7GczfCRC8NOkwtefnCyOiTbaNiqZKpdT5oNadVer/ER9TOsB0Xp3Q
eqFu83YVUl/QdFS6gUMn2eBUy0UgtlU9PSN/IbVU8E/k8Kl0SRRpU3r30OpqSh8K
8I+Kjgt/toV5i8k/keE/5cpPjkPIIqgJjGrpr2RC0PkZQT5TO94d9jiRKQQVWP95
UBnNj8tr8AkdiMa+WvsKJ/LRfoBX6RWSp8fm/JQjiYBRXhtndUqJqjLCTr4FgY28
qbJ2Vh8+e2k/29OtCOm0uzKaRAdxhyz5cggpcV2BXt5WicRcRhLVzkNEpVzruYVd
xOAxs4uRF38mARgGW+jGaHnACvthuZvabyMOFVkK7DGfBU4phrA/Ohg41r0PSOUc
bV56Tc+/8WaJImeQIPzO/OiYFOyW6NCgSVmmuR9XgWlNgE5dJwZEu4/CG32Zgjuq
UyOnOE1l9N5SHynBAGWQCSrwOkX+Hf2ny0RwAxK4oQ49kcAjGyuaKeo5yHctoycm
Fiti99hz8B4w2Wdu1PkbETqZ3n4ZHv25K5YHV6QOpqRzuHNJaoKR/7fnC6X3eHo4
0lrpRlwCVkE0PMBW17MYCAifz3PHcVqHWpqQRLx2uwS0v4Kw4I3oAI11tj0W+6Q9
jCLC/GlVgF1Rv6c3L9z49+8EZelTaj0UyEwgVYuzHlmDUgirrIxiWh0A0NYW7Rpa
riGGMxvLAr/14NWPafRUNCZ0nxf5UgOVJI8bIHELW8YrL6FAKvjUZIlHLvFRgs1f
KMEqUB5MmiN7EUMseUhwDAN8OWh4JJSBOEOD37rQPvbmdusIB+D2koOTIKvz0aos
UEo/+aWAK3Bu+XRLP9JBiKpJGHUiwa965Z+yF91b28n74JiQKbO/7i42am8iMeHt
D8dJDKbMqut2p90RLoKUnE3jNxKrHuRGyV3Q/AwTDzDCwjbVDgLBQUWd3mCi2RMa
KXoPPXLjS4sfuVVgAZwd4v68Ee5N3UCP73VI0Ppc3PZql2HiIWRn27tLLYZ2SUcH
gwctSywSUeHtSBseL/jc9KOGUCNDQA6CTko1bvkdui9QKyIsxsv4VsQH+IsUMPzL
/HMRN/3FaPZW8roBIGysmSrv+GNBIxM9CyaORuMqR6AngoRSkFddanBXouejDmWI
T/1YOWZ6RSSwY2sKPpw1HwnfhpfveckWK3zOSAzkuAN4cIny0QEn22OtgXdC9Gif
mJ0M4SK3qt6qqpOnVPbT5RFQ2yzPvhsiWTuFQi7jQTxzQQKhwo5Pb8ofRsvxUZ+I
rvkzJAqZmQxrm/6JHpw/N85Hf111Ecrz6V82q4/hm69Mr3W08bmmHbEK/9KrgKqO
v5SM2pJvJlEfkM/7ZQMaGLsAmDeyQLMxIzsI2B+VOgSbtOaFYi1QPVGerX3/Z3fb
IbVkMEE9pKsSiI101UXsIYN7pQXUdyU+6+N2XWDmWWZP+UhB/wNfCY/qxHrqwA7F
pual5zLvilHaPyUA/B0nxXlTZonmncjluS3YNScx1ZK8/cK0PSsJzFvLNMQLre7U
Y0asPuazuqyBs+urw4aNld3TuDWQE/RX8q5cINx7DVbAzh8an7at5ChNLtcqXfjZ
xf/fE8VscYqhamrLD45qX3b/20fHD+GoDOYsF5OMYkpCcwA/keqvVE9KzUv2qUiR
O5GBm6jF7vUTcw+cKdj+GLfiobyb5ILmb1tm9MoWwKT+sn8YfaKca5SdEXMb/VEo
sRV3CeFVh/BbNHKCtycYA3z72848k35HMp89mVfXKxIaCDuNmTfUpgTdS7IYsFSB
Vl2rybygbRYyhtWSSVD2nYyNzOslPyFwF7ll7M0nVkcaw0IAsDP4aJpgAfPm3Kj6
4A0DWTVLh1IvXnA6I7Gb1H5f6UUtB/ITWsxyyOEisy3jTchfszPn1wHLDtJyv3Ww
jbfBlFFmudN8/gzzEZpmmzkuUYIOdWMnyhsv0+lY0k8mfjo2wWpAC8g2Fyjrew8C
GFtjGuYeLXciJ3/CWsXojgzr+reZnFxtdL8NB5d3lQvMUuibmB5O8Rb3dJCGCHJ/
Qhq2K5V/2UfzGfM9sUGuWnxV27Vyln95BIuekfZGf2Miuc6GIx5XDe1wNyBBf+Mv
W2OZkBkvOeWcyHIWi+zSzsulsovugJWCSKg+Dn+j6ApKm8Q0OnrOECfI2M+gkIgD
oiBmZf1Kf69+WBE+6DUch2zdP+1kEFi9ZrpxcDVTYlQOe8IwnTXtlWkqHSQcOrym
kxhBN0yAF9LVEvzKxCnM9FSHqmt8cVnKtpBTMD7DeAdqhpLMgPzIKEtCccj048nP
CmVxVqncTENf43mX8nUeebcto1NANY2leZLQC83ps7hk9xSyiSxxhxKlTubxQYOh
Xt/UFkC7SHF/YYyY5tiS76PqHrE6th2Yug2n4pumti22Z3U0YlnQ4t3wR012YArF
IhKh+O4ASzOiKAXlz03nFN6sbPLmWKO3qYGH5kcC0ZtIAwpg8zHusdul2Vew5s5q
EysH7fXYLuqw1fxwhQ05/im95kZm6bBHQ4ZkAusSbd+oGbLcfsS0o82TS3pIV9rb
k7bzFAwFqgYpI9sA4TQK3xCacizoBF5Sgqkq+GVXakpUjG4XZxUlLg76uRkx3Uyc
jH0Q+3918oA+jzCpPCkkkYENyHQjVc2IDx2sMCobLaXGTZscLYoSQEoLJO2OOlu6
6UqLEOkW5jgY565TEfy41ibTta2PCbZt5TC4adSNgpejdrvkCLZu+Fth/MfhEye6
J/+LybohwMN/85pNCwMTLP8RiJJj0Pi7FzIqqFuA0mSh7hIO8ORV6uPj3Yf/A03G
iLpUoWqz6TQtW40udqgszrgaAtmUXBKJA9WyyDGmtdfd2ZPcP+GVe+iwEkQh4yxZ
4/cUDvlcN+sIBxnoEcY9QJgc9+uyQeH/bpCz8SPPpGWMqz2qFbDlWKLE8lGQ/NMp
HOTe8LdjJb1W3sr+ykaIFGaiOTvbk14V5lkBeCpSCheh6/109oxRW9FxYkZjuZCT
PWDwT+uAuMVf9huf9GM8gnUCgcPizHv6DMw5p9U9weTTUnip4HPQF0oZ5SZtllAx
b8qfO5746+G5FOe2b+F8sF6fGKmRHXaDPQI2PxZQLG7DpiqW0hl77qI7qdt3gkYO
rpgny+q/fr2ggNwOzSOuWCAeycyLcnH9gSA5zONParaB+fN9gLLRcfSSjhZxNqz/
hSRMtxqg/d0U4jGcHQeYFVpR76eTr/sNis8rTdS20ERIOVLJ3z/Taa40HQ/Is89p
RPoh49TcsbGV7iueepRlC0xnjwliEwlrwr0+16T5uIW7BUw954yf9OZAsxZ5pjxe
8jXqxuyISnnOu8oqNUg0vMKIyPYHnvm4XO8JelUv79ENg04WCQ2w46xzc0mZRTar
onbU8H4wC3PaDeBCLZlXqkUjFsnY76lpULNx9Hgl+YI/T8pufwcRCmOC83Z5EU/Z
tSxp0eByfwpCDIPKcCgfIf///e3g6RIWxf9AdK+rXalOf7GZWL5fBnKaH34brpQL
zx/8RCbTIPySdsgWCRGFHaDlGh0I0dhkEBdBhu10qY8mii/saDFWfnAGm4xsXyFe
m61xWphaUah8uVQS+6ElIXz0LHzQfXgw3uk0JTk3li36+6qRCfgKdpmNEOjAvgjQ
xTcYddLvxua8IfKj+5fbt8EjJGuKeuXHfurG27fFU4hQrrItZZkHMBeeZ4vBO7Ht
M4JCNSRIFJPrOLY6gQmZi/SrtFetcsPJx825TVfuecUN9BGty9EA8s1RCx3ckyeM
SdQdBpsrszU5w3n+vy1SGrNmo9EjLgIdHClBNBESBgGQxnpW1/Upcl8CGmlj54ao
npqL1XYxflto6+sV5llAQduOqhr2+8sZ6MYEhr2UA0RWIGqwQdbk2muWFU2TIHWk
gmr2EnIry7CP1X5Hhp+ULxbCbq840HKzI3dQycKf50+lo7j6MpC+J8ntGMcODHfA
hTzzOgjclmQecYNMidyDtle5xdbBfg8lSZ+LLnc8Mi43t1dyKP9gLVoa1NSWHOFn
56vUjW4ZyAcAWgbUzKPgl4YLhaO83Mj+y+em6nhAilEB2AoInEJA2RMHsB0Ubk6i
gS9xdxEeO8yIXB7akC25k76sFvtfsR4BlxvKrrxklpsGy5o8zI0BNXmSTIhrqxwF
1wVkKDgeeurIOl2gkDJeVzevDEn3u7rJLVGKS5NSa4wo3Lcpi0bIagKWxG7zHjKD
H77pOnt6biRYvAZEnZ8l3u9GhQVzrysI8HM8ZkTDAr7d6f9soWJRXMgL1pt7Qggb
5D2fL02aRiYLa4lTLHfO/aznhksO7jofChONUyE2giXZsrSxqzT4SexWp6NZAm+O
T2Fvc/ovp69qs+uWOBWEPITwtENkWOBS/WnfMYpCpBmpdKzLouv/uPsNi4DJS6Za
tX4COEjGOc91bKPBwDiNmarYm/msUc0+uD5FAthCsXuAb1EjQ13T6wB+1IQo8OyJ
yYeOt37swBAAjH5ah/DjITfVzcewtpsWSTgEorAquz0C75ybrovwbhqASMtyKfvq
fqXGMdJbZu9Z+Yhg5V3zkO1Ts9nSSXewHAcj0WaeX+A9xX/3tm8m0OtHh6Id+1E+
lwiUN6tN6uVWr+ElWMHjU/4IMUx19woKd1wXxSW+xGVFER+nxVugcVPZcI4c1rkL
a948TQg9olLKzra7ZcyiAMqKy0AFqjeqP9EJ3uDhe2I1mCwXqjddhL3jdAhLjUE3
9+73g/hNE9nrGCUoUp8jlRSgS1vuR1QYnQ50mlGQt3k/6O3S11XsydYJIiOcBcPZ
Kd8SUmk6m+QkXyoHsZXTyUIJsM0A04VsTOiNfw65Jx/6ojPJa8HyXHTE9jW++CXU
Uir+IDHf5wbYGY9eu/CSHg5yjmAflGh76woQNBQEMv80WkaPOw5isEMataLadlvG
JtlD2EJIPV9lTjG0aTJ6y7I8dHM95NAQo3R6kkVNCwo5QNbtBuvhTFZVzDuqaIp8
6DbgJmYNWkLpGFLUJZrv1sTaM6wsARPom8dGFL0+tB8r57ZwatXWuk3aPpjpJrCx
/Qb0Zz15E34oTFJIIgb+OnvrVeBnmNxXOZGZzKHF1ohARRXy7VimlLc69YZaAfov
mmwAyPG+45pXqcg/T7t2hM18xdL3F/2hl6kRvQpd/wvnvwc9r1nOZSI4czcg6qhF
pHtRA/xd9mZQ0kF/v4X678S01/byiyq+pRUzwLoI0iXVeSsfdiErxM8DUyqX5XU8
DAyZK3gJ+6fnIzKWU3Bs0dljz0xAOdcmvw/Nn5ZhyF5M4g7Yf3uwCYMzD9kQitGt
TN0qm7/PLia4tFSr8qDMI14kcX+ROVxNhpfa0/o/zfw3fbHfJPG5SbThkDRjyPFJ
fOWUmtgHvQLcnaYYMEwyG+QDELPnZ1PccFNNoRN4a895ve0tAhjkuBl3wn2OC+nd
uy6m7GFN74IIsOTbCYdEu84ywO7ng5ho7Q+Tyyw920dXqLdasmgr1J9xB+EFHFmL
wlPiw0Mub4EdoQW9Ttkp0dTkMaAZXs/VRbFf2yk0vxBRrUZAaLgMCKogqy/ggbNF
nlbIcj4G6XxIBapM8+zWDiIpc4ZtA62SE1sPp1wC607CVP+xOuAz8pFKJUeIzDlw
IcUNTYLs4S0nPLp9AGGYQBjkfXj1v6BBf42TLadjt5aEdnA0IUDhbr52LV4Tu1Y2
g+dyZ0DB6ER9xVJZkoWi7rg33Hw4dCjSREv9na6ASAqwC/5ncrmekB+8t7ZWqWCz
VqashKfkghJqFBZk+sUV0GmVqi0vzM+sDI440zekR48OhhKJVd57ofrztg1lWGD7
gIWZqKB24ez1Dc7ilkY+A261yotHxbszaoBiG7y0aNttpWz76COnG2VXEeokRMer
4m6LJWaTs2OP9jpZ8Hi1sUfKBu6mna9cCYtg9C0akCQQTZIn57pTy+KoLtPh0Ytn
KJV0Iog2pWXgceKm3KTRipD6RQTkePri3UdHH/kMsAa7fM7iE8bm6iK9xKTMUe+T
9ie4v0BgmoLWclrQKPq5eCHn71mPNSFqsWjc2FC8FXUwqxTyvvRMpMeCOt16sV8c
OptyXVB/NLlh01Wtgol3rHiRGJPYM+Xd9OJsI27E8VmElKoDay1dQA6oYqKCE7Kj
9SmtkRho242HnD/kkP1luCZfjfVRpmKR5Hd7WcaIkJNWUpJfuuow6/tSoFiRsCdn
bMW+ZSD0BzaeQu9tHx6egSm3/gC5gcEOVrRv+E5awawXfnaDqODGSOenNXWy73ll
KjhgP8ldNGNydryyPa3YiEOAhVU0niUvBO6hosADFlW2Il+jAM7vOptkPS4uGRso
2+f1+JIrfEgNWNXwxuDWS1OmJWQGTg7RXKxgKYTQKilmP0fqqX+P+MZTCy2trGVk
b50kJiCaUIGmx/QoysrnVR/1fq84tNhidr6rna9qswRLJpQx+i4WWwDN6MzFsgZ4
De4RZu4HFoqafyIcHcVq8jWHMDQoy4VbOE53gUA0FE3jIA86DiPPm5wYD+HuF1Xe
XFEyn3VulGASn1gMv1KJy5rtC7HIA3oj4jTb7yG68Up3hDQe1aQ2zUKatjEeorY/
CKA2LPXDvU3zQerZBIRXXz14yrtm9GIIJ0/CxaTPRvJxFA7JrQaMEaBUxcry4xya
9x8FgnChTISoSyMfwzL//Sc44oY+YcAruruEI9MunUkNQL43hRxd2AIx0NQ7QBDU
chJStaDYtdpY3yOc4zICio8uKRqxDRYWt01jo1cLJZ6MkWL/ugcRLfOgaoC7+Tfi
F+Xr3SjpX4Ajkwol5y1fVagpvDwiZDRn0jGfBIHhY5ONprD0XP1QVPsfxIVry+ta
sE4km5vCx1Cn1z62xfsqolNYf0brk56lssG0cVqb4DrcZBWwI2069H8i4/SRq3QN
USg+63hCNO0AcO8GuWrt/LEW705gDjsPJvIcjGn0NdPIDrtXGwhALvsXctWElPhP
GoMVa9DP8tcEAIk1Trs8z+WXfjxOab9as6iJY+tSSYAwJyBpNPcbv9bi8JHJ3rbs
nfN6Ji+7tDiceMwE14rqIh89Jyn3QEt0AmLy4OKOBhK9POqsr2gTMio6fCUa0W0M
xnzNEfjk3oPMwrn5Bkq2C4bsIZmPA0m2W6DMZ6VE4TGbC2CRq+OIa+o3GbDz9znx
mNFc7QXj+bBFsmIXLN1y88/Xvk1o60+5xX7BJ1SGufvAuaCx3JTqLFt6ByQeMHRf
KKy5u7CuhSh+OcwdRKWiFEddy7GsYXJ+KQnXTMw35+1tJIHekpQfYaUqY16akAX7
mViMpuFXA2S/+J5yFvbnbdIIJZsQObEZYrf1d4bq0GKNDj0wGbiKU7PoPg1EmbUh
FyyWl6EfNG7U7NTcHUMwySWO18dGcb54NXqk76bVvDp5fhGjw8rGBgiWiaNW0KSx
xf7UL3tGWtRLP4CEf/QU0mFcsMUKHrGb+8J7xjjMN3TDdh9E4umpd6WVgHOH9w1y
rF/LocUzsR51RbPXo6bz3wiOfnN7imJZ9BztOCxwQ6MB+KLJ6xhMAqAUa6zD5nS+
Ix14LwmriGPf7V1zHMbJMVbcisfpfPsKYGnJHNFeNfxjT6WT62yFWtm3nosx2VYD
OlcYHp9j3ZHh0QrFB7mcaDxfXWC7BQyxIa089QYgMeADsRSxAuOorhi+74IqwXCB
4EgKDA7/qQhOTYnJMftIS3Ooy7YkjKQ5OkHHLkk2HOFegEqysfktB5YpnAdE7W92
aZIMyV4QOLSsonm+4WyOh/mamWosQ52N72dV18JjcSsFKsbLfziJlAfhEoF1EiXQ
2HXqshu5d1aASPy8RWgeOL7Qeua/BUPUrLQNoS1Mh7c3eNFeiIaIwhKeJpTTfpr6
3hRqdlN2OU8v2PL+lT6hAzNzoz3g4zZ0VhGgHbTXGaGGGoIhWkUqn63iM0V+rC3i
JdJbxQczIxxQU+m26jQPFJjeJyFkbBeo8d63EnB/4zMUX0Ol1mzBC45JW47p6aBV
T13TC7+HKArafoldm3Y/uRmUW7t5bNpwIygBlcSrYRkS260++/r46fkddPTJm86d
FkkP4L2ParVIGRm6dLJsA5KSwfb3ZM6EtNuGOjNYaCQBLo3oTLOERE/7kjHuqY4X
r+TNqUU9opWB7PiXVnoChNxZidGk4HzFrUSu/w0od/3wfKWWwxWAmso/yVRvLNFh
uLWFH7cTGNYvL3BliGyc/9aDqN0AdzzcFVpW52gVfAvpImGhr4zfqNx3lG/rjK+9
d5naHuBa1aF1KYhePhE7FLTHnzBS5Y9Ef3GTE2pM5ckESMOQOxUy7d5K8uOISx33
k+Oj7wrW/TjNQhaJeND4DyVZn0xM/e40Qv13TY0Z6BjbAhBYKrpSHSmwQ1blvYMh
JJ4jLPvR4GmufUW7xc9WCwLkiiGX2OE3LPVeON4fcPNjEzxD4A2h4OgIb0KcSTKt
OvD1Ks4VtIipWsHKD/JUn+Hhq9SIRfBnPIYRqBDNw5Cf34jKbPZcwK10UByutb30
DP0LQ1sRRKK++5nSwBLtNUrKN7KSfZ2kpmTlZ8ZgU3TqT/t4+lKf70OQw64yvsBv
m2pJ0TxPdI3uouA5zHdTK8wVNNh1CPhnqNRWPO8t349yHMQZhqsP6LeiGEQ8QSvu
kuQ97OKn3dwBmJhtkn0agTtQioUveBP6C442Lw6q3nOS68NIPE9zfEaxMfvlrf/6
I22yYaR3GAp+ZFf+MbXk+3hDW8G6eajYKXMktFGxTcokWyToFGFY60XSfQmxMLnR
h+trxFfzoLQYCnKJlx43sw9W4mN/LxGC9HPT2tn/y01bgJOM1H9l000WNxidDCZn
ofgg0QOPKpct4CcaGbp4L8BicOix6SoGCBzzDt+WxomRdY+K2vEPen+uyEx4D1NU
BlvqF8fXsWOvIhnDeq+qNx1pISui0ikZ2quFTSUGOgy66QacftWWTW7ycgZTe9MB
GaiibVj9u3C+XYyvnjTFj+lYupQc/+vPLwGSP0v3srJ7FHH6n57K5tTldFG9Z1QU
/4q+XNJATnlKDLnMUq/okOGpWQjJMuN99UJAXppyZNXEc1MOe85SetSfHdNTQu6K
44oZ25j431+W9rFiRwgYK7pYZzerbTHX1n+iixhjNsajXS5OHHgE7sLSgtEUVdOZ
P9cgpnrMC78B3mfPHzDdG13UI0aRzBM1a2OREgIGc0fJzdW5hZUXjlw8uzsse6bS
jes0zxMkzM2rnMPd04TOVntg9ut5nezFkB+jm3gleHKPky0zOGQuVCVJ80DNlZMp
Pz27WUr2dA3XWsFIx80FjElLrqR7h8BuYxumT3qERjvuJ+JZppc19vd5t4HOSfGt
Mee73wm68g+L1WlK55s82UUBxsz7IfWkm9T6HLjIaPzNzmdWXKt8OQUdMkmsmZeM
NbrTZo551nYw6sOLsAoeq3XkQYPT6i42JGc4cJJUpvSFG6RaljGKmwKDfGq73Vtr
6bu0jtEOJz6e48h3nRqy5kj4Dt/b5iBlSnGxK7SUk2JmfWuyN+0YLIbPfzoNRkNW
NSCOp06sKzqo/PS+kWPNQMAU2pWwYkB/Fw7g15RaDsHpBV0M/l7PNgmxo+7YFN4d
I4StdeAluHY7YJw64f/DNfjBnD8RUP7iz6i4FosHecaCWcP7zyxPYb1GeAci9unR
gUqmJkJnYX1ckh3LY91pmi1jYvAdhT+wkJjLhgcWDB1oqs2LlYM7EPh3RQzUFpBv
rGa8Oru3otDdC5OTI5gJcNolgafDhqsfK1GG+UBAZwsYCtOlrkFOVRJ6FikvDQP7
YnnzE1zBV7LZnvg+ZQMJ4vMHmek8wc5DnpuAkclKwtzbNSl7Bw2FsTYtw6lDga64
b7uC9WFm0LGWB6JnkSENRdtGfcMkgXESxV4BmVHXIrsGJoZoOV79n+iHuvmqNzXw
8iGmk7ZWjdIg1HtmRstKv+IUCSo1NF4N9RUDxQTbtDoXobJEdZyWFkKPiqydzMK5
u77pHwskMh++WhSraD34LXxZ8TYw79YFBBW+ApmlmCPJU0cUsUOrO6EraV+mrDNY
0VQ5yR6gSgfl21VKajz2m73gU8X7zEtXjkkhSaMREvFljbW/ni9I0Eo+EzjtGDI0
ER4v1ktJXFjiLnVqUctdnvlEWVd1KL/89yKNVspcFJzcr58VmcGFCEdYhBKT57kh
RYO9bxdaGkXD8xqSyGxZHXbVIvxZ7O5IY+Y0W5Nu9jrVhFSknDc2mlJ729tO3Yc2
tSGXo6fHLX5D1IXWmE0T/MXlgmpUG5z9taTISL45VS3T2VdOuC+FuKLeL24niKz2
intGIBnC/8simfgL1ecZUT5tI7kAA9htItAG54bUfKAzXgxOPN500llYLeBAVIIq
lLheVoxNRxCy4soimBP0RqLBOqA96vi8778BZWXpz+wm4N8TmxU+qGhjkL7r0paV
17/nV8PN17D1r8ueSd+TJKoJsT1G4+nOIn3zD0bUs+Cz/YroQmevoFCCngYKuD0d
TN3cPkyIsbH1CMGvFGlKT3d/0y4JpC++nBKhsRcWm2J6ocDYxyNTBRrn5+ndBRs2
5uQFxGaxzr/qONVIMbMhtM4blH9GLvF+FSZnK12i3hB7xprR9nRVgEAsLJVSg7+A
+SqH7njDSqrVGgR8wFJJRQzZcHgEuEJi0QPv1k5Ka8K7m8DElYtOFIeX5IqO/YHD
EmvMjcvR/zYy0P2doh9slPFrcQwA7eKzeRRB7HZfJepSAvCa6foHMVwUBpeaY0qI
gmxtLboWwCV9zesWeSifJ8/SVAb9o7hokUjO7Lb5tNVaCg2lGxuk9X+T8ajLLPik
Xi0iMxApZsbaOUiNL/3sk16UtoAIa3HXTQoCiZjF9FCgw1IlQTnYcw1ZCsSvz3bB
cJ47Z/1lnkZ0RBDI7bWI1O2q63k86snbzD7SVDGZHrp6qZcvDkeXNfDm0ayRzwjn
zC1n1w0NRy6uPeS29TFbwfEqIuzGeNf217FcO79nwoV6xeMaWkER9pzypEKkHwHe
JmzrBa3ZwLwJXcziTdwyXlv4HiopWJWUx2SaQeWHC81uSOvO5LKuswujVV2LRLWV
nRObCb63a27Ic0kWqTkyP3xiEAb3R3CSR9nKbUxjfK0AAUJ9jKN6yo3nGbG9ESWm
MNQOH3yvCi9Q+gzpJMWS2zOnUuImu13VQXOZcj4WWSNKsDAIUDaJN85SFtPz4X0S
bNfKh3sk45+lNpuz45/8ckR8kpQiSdFiIgu7lTpWeRod4BU5IDmbswR1I7GEVu1w
O4+ZMNZ9mK+8GsXHimQM2sZwQRunTIsRGrKmBJn73j59fsRA+FQ/FfabqspdwUJ1
1pNdHYnns5NXY8sJSTUWJR0V8Sg/G0YPwWDSmP7fr7rz0hrk4V60depdCidPeHnM
21Cn3SB2WO+U12W1KGPl/0jQAk+afZnoC5fV4wHtYExlsBuhHHSEn1T6/sf3CR+w
94L1Gq/zAn3YsXRdzVYITNdNElF0V6IQAau18Ge74am7xRis2113DjCBB45xCDEK
25aJa8V754oMYAzsCT4+9MIT451jMuMQ/Um4CIrrMDvcds04oi7m/3zqlMFDqjMn
m0O4y3rzINL90TQFTJ/ulBes/LsjYYXb5Y96zeHDMnvCFXKsBZ7sjIV7DLSCMRH5
QRB3X0dK5ZEug/lZ1mHHSQ==
`pragma protect end_protected
