��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�@�w�4c^ �[M��d�#��������C3=��ؾdb �Āb��q�������)UZ�^���#�#�vubw�I���fo�T��t"�BZ��
�[-Oq���O/K�0]�G=z���f�֦�LhU�x��i�d�o��AkE�$�,D�QA�e�+�?��%}Hg�����m���l�*�BR�.!U��D��}���T,����2��F��"BHO�`��ֈ�2~Jq���*f�{�|����,����@�4^\;4�{1u�|�
�8Gm\-�TϩHᐈ�����N>O�'�O\'^�dR���I����EO�Ԓ���א�2�},��u9m,���`��&z���`p��Zf��u�8[_�Uag?e����k|�͉���l���Ե�
�vҭ�92t�>�V})55�+��k��'���!,Y�1�]~��̪N�Ѥv$�%��vn�6�M��>��[�zO�ag�t5�2�>6ɔ��(�נ]*��¬n��y~ƒ��-o�{�k��b~<�|k��0�1����Qݕ��=�g�t��V7�����='h+�P��˦ȉ��}���#�B�l�����9�/�S�g"/��Ou��c�7Nt����5$���X��A!��'\i5+_����A�w�DL��p�g�7p�RL���p��*]�$;r�J�bD1�,~�����OG��������ћ��;&#/��Ǥ--DQ�ω�?������M��ǂ���Z��/���)-�c�Zc�"qP��J���e��t��n]M�[��!lo���SP���>\S��R\�FWH-�����F��è�p�6Y�,�2���$�n]�|Ŗ��#c��Y���QfA��r�Wb�^ϹMS�n|O���&��ƒ���)��O�Vۚ�,?5,}���P�'ڼ��vH��ޯ����1�k���j�Ny�}9��<3� �ĳQ�%�`�M��s���VUf�Ƣ"7�jh�M��v�n�,�M%�z�'�h׷�c��L�Rq�z���P��u�][������O�n9	d ��R�M5�v�ߪ�1�y&�0uW�mFB�!�AM�C���$�h�8�a��A1e��Q��/e`�Et��j��T�>���b5�׫�ٲ�������ҖWL@����������D��=ݳ��'�Ƽ[ՔL������y�$E3�گ��	�9q�\�#�I�k��`J�4_µ`s��i
&	��i����ZҒKz
7��=�#e�*�t�f�Ǎ~�6���A�9V�P&��]e�^�Xy?X�*'���6��U��$���r
��6?JJ�*�j�֔P{e�H�W4�,�2��qr{e ��O,���3{")�t^�6����GOy]���!j�E�fB-���n9J�Ba�+.1�����K�
�#�ϣ.ɣhn�ŎG�˭�_Z��U=�.�>% �`�;sxDA��{�Q��EW8@#
֌3��e����	��LEnaN��ܸ�ۛ5�H�{p��a�~_��*��`;E�[��h��n]��F�AZp"�3F6��)�t��,��[�{�L�n��#���)�n����_���a�r�3���e���m�@��e\���>��3B�^��*fT4g��F�U��62f#XL�FZ���Oe�gl��N�{��7��\a�T�(�q�zJF� �g�ܴ�=�Y{Ll饍�?{q��,�UCr�f+�IO�u�6�m�O_Q٣_�oeZ2~J%������m�S�;����kG��SP-@��㼁2M�\�2Uժ>%o�hT��?���Hb���z
�試�l��n��m,��s~���"��P�y_X�\���}�����:CN���VʅZ�@����;y͢D$�_^$=M�d>��#�,�Ȩ�����"y`�a�{f� <�zX����@s�,O{��L���cG��y��(+
ORm���Z-8�P�jڎ�j�<[�1>�!��u�����c�c ;����ë}4m���Q�tZt�	9��0n��M�K�60��g P!,��Hk������z���f�xq�I?�=2�"��a&��_QbV�/:y9Pr`G�<M�R�����ذJ�R4�f�4����w��oՍ����G��.>���o�ϼ�,��D{�y/I���BW������R"o��"���h�e����^�@nQ�"��M��~�1�:���seu�<�	�
(��-kѧ���xB��Ìf�[ k́6��K�����DX<P��]��\���V�-�f�/�$���<�I�cg������J��{�z@���4	G,����7?�޲��`A�,�Aβ���Xbբ>�"�)��Χ������ej���2J�R�t��'���p�R�Ƞ�E��+�QB������U�vb��)\��c��l�q�N����E�K尻+����zi`�N�e4�5��Q�o`���˩���Oy�Gs��a{ܮh��6hQ�<���n����=
��&�%m���׷sSڛr���v��ޚ�󺙺Q�����2�,Dì�@a�Y"�	'R���B���z7�)�M��l��`ӃoK�z*V��:&s��^1�{�^&�N��:<����g�u�QS�$���v�X�����ǟ|Ca,���Cx��R��Z��?Su1,�qwJ`V}�Uت꼏)��e[�k!_!P�sP�NϨ]����R+:���fz��K�nw��6���BK!��ջ~_f��՗c��-1�I�2��OT'委�/�io&�w}A�Pun+T�-�uW�C�-Z�#���֙N�̸��%�����H՜�ۊ����r:��2��^<g A4��Y����@�K��#��|+k����^�+|�p]=�h,�Y{N�Nm�s�G�y�ҥ�"\�}��¤��������!�y&^��|Ų�)$��-"��c�a&������v�C��j� �N�J��h�m]��'�
�޷w73g���wZ	�C��O6j�e*o���9
ܴ������m���ڈ��x�@�B�&�k�Y��6�!6XN���BG[�9`��S�h��d��!�d��Ha:�H)%�:U����x�-?��نc��4�g0��*���B�9VnÒ�\����`"*�Q2��(��c�$�=/�Ϻ��nɬ܄�@�����f�� ���J�̕,.�}Α�VZ@A��+�S��H����r�C^��b̆�8���P✽�}ۿ�{r)CEP���`da�����/ʻ�)v��v/�U ����2k�U^�/�!{�+�Z�Uʔ�kHb���2d���p��V騳e�]÷���_��߀��l-ق�4sTSj��M4��ˀ��5�!�Ak�KJs��^���d�u����K坌m��8=����x�HU�;��4��L���R�Vd^�zq�г�b	
XaۏjJG����C#������m�%:IF��P��pJ�1#�,ӄ�!��~��~m[���/�k�z�;�A�_,����Z��� �v|�42s��;[~,�H|�_s��u�Ex��ʺC����$���BH�:^*ilQ�n��.؎>;i�l�-	����~~6��~�� çL+d���e�sI5��dwmo{�ſ/!�|9� N�US�l�?�J��=P<aV�������(ǰ]��_:��EB�!��M�JML/2$�Q��/��@}UO�p� bY�N�<nʃ�Qa���7���|�ܝ��n������&A��P5�͉��N��9p^�?1�%K��)��6�%2֓N}U�h�r�{?�ov���b�(�JO��7�žh^ݝ�2������>'W�px53ߗa ��e�PR���N�ӕ�=��
�YQ�i�vO��� �fY��/ș`N4��S�쬁CI�_L�N@ ȹ��pp�c�w�����Wg���AF�����c�{T�#�oNʀ�]L{z�{*��j@Tw���;'�T�l�R��?v%; Z�Δ����a���JH������Ƅ.�_�+�Ou��5<�ɬG,q��Ȕa���׋,�׬�A�&/G@M����|,���V��uْ�íz�5F2N�h~�G�Ɛ�6�0�ꭂ�pa�	�zE[��.�]�&A��lI�E���5�o8��J���?l���5��d�z�Lo�gNQ��c�ߨl�p~곧���H�ABM�$��g�Z��6�iw_���7~撯T7����}�
C'%R���+��x�Z���m?n:���z;gD!��ͮC?��?A��Y�ʁ�����,p�5]-� ��s+5�����.�����#ngY&<3gY��>���6����n]�����ji���?�7t�y)�Ǧ�����z�?4��įZ(qUӌ��ւ�|r��O��A������ý���{�s+������M��-��Y�l�^HR�lZ
�_�G	�V���v|"�8�-�g�]̎�E1� �z����7��0̑�5�v}{]� �0!4��`�4s���{ˤ�D�m�7��({NF������:V��|*��Q�PY]6��+Ňm��}W�8��`�7��x{��/���Y�����7�{�f�Q�d�R�i�`�z �#\�f���
F�/�'k>2#�{Go��2[9�Փ����(c��p�ȥՀ�#况�#(�1�Y `ܗ������C�;#|-�V����27�.E���h����;׫����:8��+�L=4���XIh$� r�D����n���42�tެ1,H&��5dd��9�I�� S�`���Qt��#D�z�T�6k��ٜo���]����ʞ���ϟW뗄ZI�MVGKLx�����
��Ci���3�ia�|��f`#��Ԉ\������-��_hd�γh�s�L7g~�ޫ�Jh�P��2����B
WJ�ѺZd�*n���w(NGw�q����/&cء�U����vݷD�7$��&��@P��I�M���!��;2�]���'��tV ���Y!�`���kw��L,Q���T�]zĨ��x��l�P �x�#��V?�PX�ҥ���z<n��
|6ME�Q�Q~�v y����D�VMI�"ǺE��-�:_�ɴ8a�Oe2�:�e����i����ه�)_K�\4�o]�"���z�%G�t>�l�������3w��C��_�﹓|�����{���$�$�$�x_�GΏ
��Xd�&G�^��2n�I��5���0� �̇��K�9�h��oE��a�R�m���R����>�x����u����}
�^B,��aV'����d��ߧ�9�O�͡D+f�I"��ݒpM�E���¡*.7������`�� <o]!;���@dMIw4�����Wс͏�km�q��X��˃=g`ز0�Kx([��(��w�˧>b�y�J�U��>o"C�����4g����xR�\i0r�mXҖN�̯��[�e�f�8c���W����}u���m�Chui���F���g)��*;{��y g"\,��[r�('�t8�k��ģ�1&��7`�L���,�(T��N�(��*�$SZ�q�>ط�@n~̌�x���B�ô�X	Od	��p�4&�0��1���P����U���h'E�@H�w!�X���T��%���Q^����	4��d�Pm� 9��n(}m���9vfl����(~��Fe|�E��+d\��~bA:���D����.����)��YR-{	�W1 |H��!]�zB�&Gh���w/�?�����\��1���}%�-�FwhY#�<`C��P���EF�O��,�u���:��ԟ�7�=TNM�s`�9p�Q���ߨT��#���|]�޹uRU1����5ށ)E�^<P�)���0=��QqMl��*��$gc55�[�>S��n�1'���#z���Y��n�W�s� ;|�bX�.��u��(�^Qʬˡaxd:\%Sx��q������^TT� $��e��C����qX�1��n"�vKU=y�+K!��kJ舱����2�&� [Q#\��"ȃ�i?����� \�Q�����m&G\�M1����Tv�r���&���X�#˷����m����8�V��CR���!��0�lZ1;�ù�o�I������&�Fcɹ�T�|�/Lg�{n���ޙPX�r���1W7
K)�!�sqU���Y���")��MV��a(���KX5Oڎ[a�s�LM��R�b�Q[&��"��U���=�+"��%��T#FS�Zc���!H��o�Yԑ�ӏt���I'QW���Y���B� ���O"ru��\�j�d=an����#�F�Ml��u�MÐl�]���=#ct|>b���(#�''X�GѲ�T^����8�7������6���2!DeN'��A%en�0�k���^d!u18ǡq����)��b�@�d��D�{m�*� e��:[�9B���R�e�G��엤�Ƅ� �)���p�,�ږ�T�!��𽪺�X;.������UU�(��\
%��a,��<S��P�w�D �jtIW��/�2 k�Z�I]4s�p�<�V�Da��1��B�)�|V1l�~�R}8�Y��+"�����6�h/�U�qy�@�rږZ�N��Rjr�H�zؑ�'�o�βM��~��	��O�,�D�J����#�����'���#�q
�/���:	��߱�B��)�F�.���C�v���z+T���s]�@��R7��S[�y1�^q�&����w	�B��.,�u�z��ۉ=���J�YWe"�(3�;�1��j���$S���3���dx\�T?߉�{�C�\O�(�IҼXk؛�{�Q���q���ս1G��&Z��3��&���AmIw%K�v���|�4��9��D\���02��?�<,���,Pz`�I�8W���J� �X�:ٱ�9���5�PV!
��5���%��X���q���&1(	����ˋ�ʭ�X��g:@0|�W�V��m?ܘ��s�:�U�Z�.�R�&�_e]��\ɻ~����ǃ��Z�����H���k�+S��~֚����a��88l�^��80��'�T(��b�u�_���ū$���8Y�7_�]g$�ʬ=q
>o=PS�6؅^���2�Y����E��&�A��/�T�k��z�q+0D`��KW�}.!Xi�d�Khv��Vb������M�Ζ��n�$����=?��islu����<*TE�||�i��(�pgV
����y9؀�t���o.Ԅ���2�e�߉��DC��!�Mu�j��m
�]G��~�C\9�H�d�m��ٛ�Ӑz{@��O��D����>8�;�s2���i���/U`�6^�t��U i�\��{r���2W��մu��!�����k�o&7ue44��h|?�+ݵ�6���N����'�7f�8�x�{����q���xWt��
�誓�Y��}np	����F��,��BəCA��wf��LFϯ����-�3�蛣�#J,F<RӼ����Cvu���J��=��)-k6FE$���	ySyb
<�0{lP�]����PV�h���xsh�H�B���L��$f���1��Ъ���:�ց��~�>!'�u)�8�#n��1��+�8���H�K5��(�lr:��7��T}T��*�+�AI�ܢ�9�;�n��e�f ����o���w |�rߒ(��@L�����u�+,�
\#�eD	u��m'x� �ӄ���$[��̔�y��m��5v��VOdaVTv<��b�F�9m�`�ӓ%�����>��i���Cb'M�J[���e�g�N�sJZb�y�)�<$�b��� ^�7��]~T�@�}^����㡮10��`[oZw;�PL�p@���'	V/a�s�=ޞ�R�R����n�H�_pJa�(���4Ο�;^~h���Z9x��EK��i�9��шg83�H�x�Fؽ�z����tiIUx��"�2�F�>��uk}>�N=�{ȽKC	x����/��`�����E���!^A�tI����U���%m��������a��X~��D~�%˵`�G�y�8K�+6� ��g�	qYe͋f�ETL�)�Fp�"[�`5G%�CR�;����t��	�J�n��ln`#�ۂ�/w(0 �Q�H
̘/Y��7>�
\��{��-xg:]ݲ኏�r[h�?��@�a�/�3��Z�bў+Ԩ��\{�(ػ�P�5͸;�y�W,\��i.0�+��*V�3�m7�I�aze��9�Ca+��6-��w�~���^�5Vy�N<�F�?�%����4L����t�C�%����83<��cE>�����[C}~�\`6ӎ�ķ�0_������O�mF�S~�:�y�Vf�,O��xpP�K���虌�j��@f�Y��T�Υ��<�o�����F��������|N$b6w;�¡�� �亘M�����f�����u��7-y1�rf�DE�����"sP��*U^A3�X��9���d7�z�J������RT���}PE��۞��[2?ľKI�V��]�9�|P�eiy�V�kuފ̍dp'Š�OXi[��{؅�<F?���|z���-��ם�X��_�c~�q��8�b��J��]�,��k�C��s��v�M�M�+,b�y~�X��,IN�	a�X�%�S2��`��1f;5��(th��A�_wb!Ŝ	U0��8�ﵹʁݒ�j���\rv����q���g�чyJb���Dsm���l~TX���PI���y�?&8\m�쓇7��[d��F�6z}�t�_&����#Q��On^R��?X_A��4����gT�����q�&xD�@i
�`3�~%�ˎ�7�Mb��]*����6��)멸h6�	>s0�>�Yo	�����*�늿���|�uZ���vԁ���́�T��֚~\T9�R)V=t���2@��� Ӛ��s��t$L�>�M�VU��WE��C���fYK�;�C�X�W�	V:*AS����]�1�ܚ�h/f���د_�p �'(1M�Fq�\�j�嗪�/&�N�x�T����ry�������;�cӮ�1�Yn4?��忆nM��"1�Ź���]��Vٻ;��e��/<�M΃k���^�b��f�١>�[���'�RO5���֘.Rc
�5/;��T�GCm�}��%��d��m�ݜ��7������§���-J��QL�,#�.�I#�x�0a9��-�fo���H|�2�c��.��
b��v��%���zm�j%��_�z��Յ��(�NڦN�
���|���\�n- ���U�v���h����Wy��Ѿ�c
���b�nS��\��%��cp�����|����f��"`���dO��C6	�����-M�ו��@�.��_���壃���a��Z�Q(̂c.�!e=ӡ���Iw`����ý���$x�Б��Y�,1|��Q_܊�ȹ7{�����O׸�H�G�Xj� �=�j���t[�@�A�)50�R'\B䛦�U���޳ˡ�F��j\��m%���ߩ��6+*����������QM��v��"�Pc�U�+��G��턧��2���!��S~���5R(��3�v�����f��W�L�Ӏ��p|$˙�����*5�Ȱ�U;A�f^� 
4���cp���j����ETAD���3e�|�ޝ�!�`�786�������Tm����A���+�Ö�X�H�g�����s'� �T�N��G�]E'?�N���ѿ�u$���]�*���/O;���'���эId��\ mVں�c3,�(�z7���MOX�,�'S�YL�w�>��dy��P_�mMxÊv��ͧi��e��6��b��>��C�^*���g����pbgb=OҺ{��0,�_l�����~\���7��a7˩�<<�[ɼG�_���,�|�������'M�;�������1H-0�����%Rgr贘�����o��i-L����v���D�i������ˎ�:�=NS�3BЗ�{�֍��M�-�`�w<Ö��2�I�9�.�Xp]�uV�>"3?�2����ìY1�ܠ ��o�R�z��~�rqd�9�t\p8&IǤ<e�֑3a'�|��$��_�k�!�����|���������d���=����Ѓ<�:�Pw��D��7O��p}�I왢��B�֢|A��Jx�c���ʺCa���Z
�0��w�U����[D�	_>vC�Xm�1�Xs1��Vv�K��۩����R�E��a�T���<����yDؾ���m� ��B~j\߬�(ڄ�ff�kl䆦�]�0�KKݬ8����/e��A�f|�&�&{p������e���:�p�f^W=��GU
��xKQ�����xr�^8��f6�D$|�8�ɨ�|�S�i�	�)ac9�Q�:O������X<Zb����3u����lku�Fs5����I�E��PH��m|v��cw��$ж����
���2Q�_�Ab��7C A��DRU���<P����J��/݀���%lՎnfP}��2�v�U�6�j��s�0Xg���1#��5u��P�_`~��/�Z(vʃ��w�g�Ћ,�3e�/��[��X7ݬ)��|c���^v�gzS4����̤���������2�u��[�A�r�������gIO�oC��J�x���8���t�w'=�~к�U�` �	�㹰�ʺ!��fs��UJ3��;� �z�w_o�^R?-��Pp^t*g|p,|�r�Z`#���}M��7okrj�Z`���#��e".���z�R��2 �<����������ʠ��_�𫆅 ����T�d�e
��vT|3#���Џ��O�Y�db��������޹���3��ؔ,��Z[�))蓨��%(R��_<�f�t��@��l쨭��׏�=̢�&�5+� o-R�^K]/\�4���V�IyUL��2���
g@_�-���oŽ:�ѐ���N�P47����6}61�\SD l-j�:M��v	l�P8�S�1��5S�U������� ��.P�"�<H�)��خ9�#J��4�&Fh��ևh6�js��p�Q�Q����?H��Gw�����I:����E�L�p���꼏��m+N��{��ݭř�"ts�O��)�Ts��?d�0���Ѓ��r���ah�������g�atV��Ǹ";���N��`	=�ǈ�A��?�t_\�%�j�e7����H��C¶VC��YViX"{�7���Cpt'?���s�_��+��C���OUPɖ*Qʝ1z�S�~��!v�,�P �Y���b����5p�E"��K�9�3�2͔�M�6�xj\�*Wmc����w�6���!i�˨.J���� �Ox��n;?��b���u��$�)��\������
�;�����_��b�� �QHqMkn��0g{4ő/8N9f+l|wq������`_N�Ob�lz�|�����U���eDP[B�Z���5ߐ�� �0��`}Hǽ�CՄ](~�8@�/���X63���̩�~�U���!�W1r��-�3�ޖi��w �&׎'�')���H���2���48Ҹx�ɥX{�3t��sr�`���R*j'�k��7T�9�@���(��*���'��h�UUO"pQ(��Y(���"�y��e�d���]'p6��"P�'�r]A���P8{��	�X�],!<MMH��ʢ�7H�BU�D.��1�RoT���E�"��b��#j��4�7�cƟ�x���~�I%��jz�g[��c��4
�{w�-�:�k��i(Ў�4�.�98�	H�@�m�70n�wT�v4�u_oFDX0��49�p��j���> �3"�p����53�i -�	K�@�n�������QN`��WHN��}!�@���Om�����EE%ޜ���:��z���M��LW1�����'�1XĞ"�9Q@��+�N�q��Y���^�}�W��1�� ����۾�3�3M����ϑ~M�o�N��#�?l�f�Ɣ�!�J]��E�޳s��<y,�����_�Zn;bM�0<�C�����-�����$�e���$�3���v���{{&qlb?.�v,3�����0Iݣf��2n�(�<x�36�z d|���Kz~&��ǖ�k�z�8G*uq�b�"�0lm�ʞYSi��\�&�]����MT��?�bl@g �{� Z���]��R�;/N��^038@��̋t���>�>�c#�@w�2�nb���@dtpڡ�X����ы��V��>���4�$2����J�`E�uܥ��v���kx��+*���L1�
 ���5�����uS̑�i�:�h�^\���!��Nr����n�4��Q�c-f�?��/H���YIT�@�;���2�sa�?��J �)�RG��X��AT�O=H[���\�j��8���W,z�׽O�M������"/�ұځ�Sp�̢H3�V���n�@Z`"H�́ a/F:gƬ�hO
U���<'"o`RvӡI�h�o��|��ZC���.�*["uYw-��9ƀ]���g��`�	7�h�A��V�:� \3�`Av�N���2V �ߖ�#����j�G����:m7}�2Jd����9���f����􌅠\�|n�7����kgf��d��v�K&���T��k3���oY7V��(.�)�s#� �SRC�9��G�܎H��nM/�}@�o�V�1��p��Hޕ�"��bU���:��${�>�1m�J�u�V��m��1}�HխR��W$ؾ�l�BzOQV�w����)�ʣ���y '�Gݠd��'W�ؠP�O~�d���P��!h�_G���[L�X�\��xƂ <x�5��'1*��>2 �������sΦ���8��<����l�6��d��3�mv�7�fG�.��ȤD���i9׮����BpB�~jH�?qs&��ѷ��2[��NAja�b��l^od�T�Lqwf}n���.�%�3��O�C��5L��2Bd���Nc98aD2���C��Y�RW_�9+�Z �L�e0���m� yK4^[�4dK+��I�>G��O�6b�a�Mo|�ٻ0@gԡ�������I�J�2헻2*^8���9�x�|T�,W<_b�n�t�D+Lq�@�m�&��|u����1e :9v�)��nE�[��,�|�t(^�\v��DG��s!��%N��Z@/������[;h�,���G��!�?5�(KѮ��7���	D=�ј�fE8�;'r�P��Z�K��7�A����':�*������
��"y�!ŮS2#ؚ�z����b�ypҐ��@�z��:�Q���YcU5*9i����@��v��z�	�9mr�v�Z�({�M܅�:x	��~f�����2Tqro1�`��g�C��G���	4-�4Ả�d�T��xZ��BL9{̉�JK��������!s�̊=Ӝ�|���}z�l��V�m�m�L�P[�Ɵ�<fc�GH��bϺE>���,z����yCU�'.�����XT�f��t�[�C�?H�7mqK]� !�m��5?Ȧ0�׷��S�����:#���V2����!�6��&yYu�]����,q���g�u��������.�! x���2`�[�<������c6P�W�o����=CZ���.�72k���ŕ4�ڼ&���"���9�%�R��T]M�8��6Q�%�5��@�Ųr
��q����,�N@;|2e�p���,�h+�����~��� [���>W�̠�W��i�����`�5���U�#�f ��j����cT0�'�M[1�dw52�H���=�j9���=��pD�����iZ��^/=�G�AtȰz#�z�v���x�܈���JT_��o4�C�Qa~C�����o�姿�ϸw����uTL]_�R�B���
���$�-f�Bc9��4n�#����Z��=�#$�ԙ�h�ZJ�hq-��9ی3h�;Ng�F`�����$�!�����z�w�VB�_$w �௘�#&�����>�:�!�bU���(�J�����;*��7�M"�����G�>�"7Q�;Ot����?}��qV�aEK�������a1����ft�������Fx��~R�����;P��4���3�C%���ty�������:�ed�3��9�Ԫh���o�I2�w�]�Q|m�VP�9A�>���&�=�nc
��3 ���0�����YV���g�ځ!|B�6/�����z#:7P
a�,��=����@���NG�{ʓ��$���r�ψ����9�Ei[.l���w�������D׮�M�b/�Z�����ܳ��B�	�;���6mYGR�w�x�#~Vb��
/�w9�\->��[y/t�e�SÉ$�*������|!Զe�l�j�!�G�D&��<:M�s�g ����uom�i�B�F?͏����PM��G��9�;�����0�
��v�q����7�EB�i��`-$秿n�ʡ.D��-��B�V���N`gnC$���KuP{MC%jnok����b]�_�k��"�9&��V�,��;�Bf�"������lat�jڊ)���i���Y!4�7~�6S��0-һ�S��Xkb����
���-8$��i���ok�6��]��бy���@�/لpk�G�"/�#�c����_�����q �����ܻ��Z�k (!:~B�[O�WZzʫ�W4������1r�1�N3����Ҭ�[VM�M���u�T�b
Q�ZOf
�����ǈ�ct)�R���q���r��W�D�b h�(^�d@�gb��^�f��ɳ|����70�-đ�"��׶&jj�Mlw�^hn�cC3�"=L������}��v$�?��"��mْlCV��j��Ç��"7���`��K6O�\ �����(|���8C>��3<�G���̒���+E�z�a�IdEPn9Q��r(� ��+A���JX&I��� �u����4���>�BjH�>f�6����M_tI%O.��%��Ж�F 3�4��D�A�`I����;zՍ����*U�mb4��������p�4�����XhT	'��'~y	��v�y6��k����1j3[�=�<8�x����� �&EX��P2;U���!��4�oÛ�3��)�٪	��E6�@ !�e/��9ze��3R��RG�.�u�![�?���N'V���TN�n��l���=����pҴ
wʲ�г�"/�d��#^	P��K<�5L�_Ţt�|;��o�7g���x�ҫ-�%+��a�ֆ?ߌ^�痍2586����ʫ
�u@Lq�$�˃�g0�M�
�gW����0aA#���Y-2�񺙡f"F���z8�&��l��Y���f��1Ƌ������wο�}�.T-R��S3�0�qS�i�+E�Gg�h��}����ܘ���o��س�4f�ܪHY)�)OZqrD��q$�w�eء��{���~��a�#���i�ܣrG��g	׷���kfY��Q
=���[��?�@������j�+���ӷ l����g��g(z �of�IY���0��3Q��1MymV��o�iq�X��w���QG]�檑/r��y
;�<},6{U�.t^��*� ��O6o5%H.Y\�rB>�۶��X��O�@ڽ�acP���C��������\(V�׃���l��5�B>WV%�8�u�g≭3u��^�cn(I�"m���0k�2���"z]@㈺Ż�����p[��Sh�vhGw/��| z.�i膓D�T�C��|t�p$���-��P��[=@�Cc�֦`S��h�I'�¡���AoK/��m�g��~�[ ORi�UD�����%`��Z�6�.��C�+��qN\�2�X��b�-5? ��X��(/�c�B��?P
�ɼS����d�l���Zdr�����[�O��5WvZz�׀y��&��-�|�FlCJD�쇛*Ċ5����7GFt�%�q�K��!�ұ�� `8�צ#��&ŲA���+�V�x�0�P�q����x%���\�,�T���P2�L�T	�N��;�g�6�_B�o�-V�_����J0���M2���?�����L:������l���D�C��z¥���Iz��o�x0�/),а$��G:Y��8}�Vp(g�/���ת����������7�J^��4�$���n"b��&�WT Z�c;NF�N؝י���g��: �e⋚,��XKy3�cu�q3>:����v%��F��FTxh�I�����i���qQ��ȷ}�vP��쬱�P��%�Ps�'���u��Sm$��ag���-�Ȭ�������A�Yn�$�-��+��N��&��ZR�/���� 5���Pm�<+�)�-�Ẉ���.��i�U�����\�"'�C<�����8g�	�#����ΙlO�*WX���#��|Z�Д�Om�2y�(,�RMAM���L6)<:��2���7E-���O�JўX~��#��ӛ���I�]�ב�OR��\�����B�q`��a7�J����e�Ů�q����iv4L_m��������%�-��O��i�gȜ,���a�E	ME.�49�׭�8Uc�M\LIB�j�N�R�-H��-?6���������n4`x^-�M�mdv1�� ����}w�WU�B�}���j�7�Y}�2�x�D�����f�c�,|�6B4r��_�������O3:�i2���'Tŗ�W_��r��]d����G��!�9<���)}�LZ���������԰Z0������B�Q��`9�x]�Sٚ�_�����GOZ���0�u#���N�0Ă�V�������#�?Wk\KK���r����V��<p��P\�lz5U����t�(c=�,P=��`ʎ?"U��\̱g�>�4I�;ӌ2���ʢ�좲��I=q�<B�B��aN�����L8��>��?��e_�˦��a� EP�C��A�[���0ne��W�U$��=U�ה#4Gi���?EG��/k<�0�u�0���p
�Zp�%[�y5�tm#*ӧ��~��B��#�V����/j���g�&��h�4��8j;5�f I� �h��.D7Ē��s=�؜:,�l�V��սt��y���@u�u^!XF0/��u줘��8������������Gfx5D-�����r�����2Q'�2�oQ</8�:�V�Bj��[���Ң�R 9 d�����͖T7P���qS���_v�J�5�L���M
�:�滪�v�pl�G���?jxTl�)�s��<:���*Yg��S��+m��M,����|����`��-񂣢q��a&�Q��������cQ��IF"��y�eB0��v�3�񸢜a�L*6F��,�@9uw�$l��nIT�z�LrK�*����h��s���:������G���a�# ����8����g���br"����V�ڙ��T�do0*�ۼ�H�7k!z�xI����N$�l=Yf���_`.�Fͣ�v�x�hM�mc���m��u�vp�HY��[+���ٹB�D�3�㕥�@��]��n(��!!S�w�},�1'K׎-�h0����/�Yi���/N�1����X�\6� ,`��o܇6H��J���q���P��j�V�C� �����:=wk6gwy>��d���Ţl�R3�����}��n.��d{�����jjP4[�R�I��
�+����M(|8 �� ���))�*�������5�G��Es}挹i��9��d�yN����w�H��2-���劾:_fZm��Aj��-��ꛍu#�
Rt�m���pːVq���Q`�2k�}��Տ�JX����b� j���5[n6��άb�B�"`�N9_b��|��M{��]-B�dak�(l���Y���qw�*�ܢ�$�%z��*C]������*�r���S'��������paE��m+`z3�W����n�kP�5l��w�$��1���a5JG��U�2�1^%�����IXI㵸��S�0\3�4},���:����y��-��4����?$�����Z����� �ɰ�4n{4
K���:m�;k(Ǩͬ�R�GV���a�eό2��C�suLh�{�������6��($�a�)��&���S���&�q�PU�{>�:	�j��R&��ߠ���Yݭ��E�.� 6(M�'����p4[2md��0(7h���)-&�Hp$�]ݑk�;/#.�N�Zs<���=��� o���6sG�$��i��E��1�}��I�pr���*Z��%�T�Q%n�%��	�$���h���ܷ��f�D�JJ�u�FN���^ s��	�]Y�ҋ�|�r(�Ÿ��G���0IG��P(�3ӽk��e)��U=�̤�Q�0���.�����	�q�=}�H��{=C��-t�J3��mr�V=Cs�9�у�y���Sk:H=��e����+s:DVq�m�Y��X�|�^`	{I�A:�Lq�]r�#!�l�M�u���D���]eQ�#ߥU��+:P��k�`��\{��+@Q0�a#�֖F!W^�eP�7�f7K��|Ӄ���O�=�~'�L��~��*1A��@<5�`�Q��4سz�la
<�H�+gDm�X "�%������w,�,�4���֢�a�S&X.�����qr���g�YK�(?Q�"�.�������޵LsjA���#$��*T ��N��\#����g S������� e-��7Ԇ"�&+�M(K�z��6b�7��$Ǣw��A9���+���8��(y�hBȧ�l��	< ?B}B�$9���|^?�!����@8�"q�s�,w�Πm�_��������)~��ʿ�7�T��o��&�UC�O��J���^Gf��b�k��<�E+ҋ`����i��T�7Q?]�P�X�(�42�0�(�U:�}���|�J4�*s�^@�oW�ឺSD��U(��(~hʶvx�!B�H>Z���7�;�Rx���.��� ��)���Wf��=W����Thz��J�� ���?�6���<�X�虡n���KȂ������q��.V@��F!��Xiӵ�Y�-�0G��\��,�˨,�~�j��Y.1'���dS����g�wܘ8W�Gx��k��ڄ�[�V��K������WPs���MĒ�哌W�������ha�폓QC���*l6�0fN�&���m�d���v��7k%�X�W��4��+����p��̚��R��bz�x��昱#�a����M�������e'�g�*+C4�nC���ի�<g�I���V=>����l��Ez���ڠ��;��1� n�Q��hEOF�a���$M5~M�����h�f*Mf�m�����Ë@��w��u���
[�!\n���/�H!���D,�Ã��&#�U"Ū���z�`^��鼢���I6C����&M�Ux�,�C,c��<0��F��IUx��T0�[�;VV�AI�v�n�K�O�;��`�}�dwܔ��P�H�b��4�!E��t����
[�8 Mz'����>�mK�(mi3��s�{�
]�bN;�i�bbo���>P��i:�����[n� �Iר�i����{d�h�`1��xtl.��: o~��I���a[wPo2�`	�_^�c��a����p��9�{c,N
}����9c1���HQ�?nb=�=��=��VT��'-���|������G�F�,z�Y_+�wL�wD���,�l�~����~� .�V/��(>%�А�;}��
�a������kz��=���O.>�x3��P��Z�a�+��鶣&�5�3�T����,�|�m��&����J��f~/�ǽ��:X
�Jm8���־cJ��!xD�
���&a��ᤂ��[1��"��T�i7\������ؿ��?/n7Rչ{4��h�QB#�eL:��E��Ӷ��R_v�~oǖ7��\�S~�!�qs�n3$=)�2g�?�P&S���Py� q�?�KY����~릭I�x��#�z{�`��Ud��u{��Rr:�ё�Я�d	:<���z9	�u�w�7���E�;`��!��T�r�`���/(Ǽ�����
�\-�������*Z_�rں� V��)�A=|@���e6���U�G:����|�qr}A����̖���	Em�*�Â�^��gL�}�MN{>)I����2�����"���1���Ie�E�V4��+ ����
mjx&礂��TSƁ���#����j�by����h�>��i��_(0U�����a�C?�����}&����g����� �2$?0!�M��L��XI3��� A�����a-�|�*E,U���mx��;��^8s=���m�w��8)y�HqXK�ˈȖ�* �&8u��غ�&�Ĕ����|r����3d=~TNzȼ�=G=������D�w��46y��arb���3d)+DeRf����D�-�2�UX�۪f"+��<��Q�|b{kx_8C��#�R��rto���5/e�ڌ�x\KmBY�'�KX�b��sZ�����HAG暵�5IX�����'�8w+��[^��F�/fCOd����-���u0����\%ƁY��J<�d(���1*ѱSD�0\�"��tn�8�.p�/�!0�یG(C;j1����N-���g��|� �J�	y{X���9�"lL���bφX������3u@x��5���5w�4,O�v^�hC�Z=���$c5��vD\��3� n|Ƭ�%�^���樭��oS����vFp�r~�C&����q=�� ^�e3ϑ�q�c��mf-a��*�3��6�Sa:���9��h~���H�HF��]��x��:�~�"�A��7A�������Ks��!���-z�1�ɞI�����FKoRQ֚A�X���:+��z��6k�e��2�\A}�յ�\����ΰ�M���8���j�F��8�}
@.�����!RQlng�+�pQ���.�PJ]D.��[�Z�t�W�e�r�&��l������ZqF�.Ѯy������5M�m@�V�D����^B~�$��V�E����mѠ)�
�!��v$z.#��,!Q���KMR���R�{�%�M�a$�r):R����"�����Z,Ŵv�k{�#ԫ��5�K�p��v�P6ġ��>����q_N�
�O�1�����'>�m~��ʟ�%�Fq-����z<" ���l���f�(sRjL��p�D_(1/{%"�Z	18=WH��%�<��.ĝ��:���>���+C�]Y���S��PhJ����Oڭ�cZb�F_Ni�x�V�ղ!�A�o}�{���~�� *c�щ���G!8P8`4��e��^��{���'�0L�	\{`��p�B����\�@��B0�)�zn_��x3�ƕp>d��_��["���X�b�,=B���3	暚jC���r��p��/<�*�Xj�`��Kk�2)�i?e��NP1A���1����6{D��*����7�az�ۃ��.����[<��%HiAt��|�>��̝���`��v0��$�{��L��</������,r'W>j��x�����]���^���F~B"�I��A節.� ����� ��C=L�f��y�������6��v�b�H�	F�t�ޥ���w��BN��$ Kҷkȼ�bݬy�.�?�j�=e��p��wE��F�֧ٮ��d�so;�������mA��a|>x-��j���A�vH�C��>�����r�����J=Xt�a��(�����o�+N�޿���{,���^�H�rXy�D��ٴM���{�׮Ł)���Y�=�TK�^����~�a��T��@@����nP�JaW��v��ms��u����)]i��]���w3��"�ʊ����F�����̵o��G ������J���|)��v��L ��BIm���\ؤ�
����:H9��m%	�@��,��M�(m��墨6ߥaܞ+"@A,��mi��Yw�0s��E��EB���`n��$�^�z���2PQާ� 7��A:����_���m�W/7�8�q�6��́l��<�󢌖c�>�Bl���p��ӕ��=��ꇷ/����]��a�Inȼ�ah�bup �"8��dČ�cf|������/G�`z `T��-��r�e�'�̾��Ŏ�J�z�B-��4=w��8����˓�����[�~����S�m���^�j���P��Ң�����!*�x���_ �߹H�����臃m�YVx���skH�W�2�_^K*����kR>d�(����3}��Qh���>�؆�j8ĬBw�"���pv�1��4��������4�A�ø�Y���[��G��_���j�5ѵԎ�%�W?�ݍ7.�u
�k�<㞱���L���=���"�./(�����a�WP$���|���kQG�d���Z���ژ�Ԓ�&Fk������Cّ�L�e��Hm�pt�U8�t������`ڍ&z'T͎r�� ���&�k9Гh�����T.x�l
^������I��.�d����~yЧ'�
;�f��pU3�>30���y��C��Z��d5&���YU��F���#`�i��;`l@F%�����PRҺ{b"����	QE*N��ƞôX_ �q�P��rq C�6J�73.,6T��y<s�5.�	��SU	RwI�8�JJ�M#�,��3�p���*��)����G��7�q\R頑X?2-�g��f�a7ډv$_ě@i�~x�y�0M.�U����+ ������Z��~��͕��>!W#�k�qys^ё��35�`�2Y>6L���&�4d�5����Yh{y����^4w �����p1c���k�� ����b�)iO�Δ�j
�O��:�$9'�����>�9̣��0@U�|�By�Ai�=lY�n��	�ڍ���j�`��`Sn|�R�A�G��Ō�h�dZ: Pl��$/BQ�d�޵dFa/62��.����R�������ʶ��Ȟ*�o6}К$[��iŊIᎋ�Rɏ̩	�,H���Pz5��oz��+�R;�zJ��R&��ټ�J}��io�o�g�׀K}E6�a\19PxK��tE��s�#�k��0@�x�hoNډ��:��&���D��g M6��x��r�×��b�?7��).X�f��Ɉ�rf,m m�4����Rp ����$,5� S��o�v.%.�B}�8��~~k�����1ʲ����=���[�d�U�#��r�ro�s��w���r���R� m.�PӮtW�c��냳�9c�w�׾�q����1>O0�7 �s��1�s�n�+�s�К�i��O�8�d�?bu�%g9�����KFE8Փ�r!�)@�\�RbFv�����c���m�;d���Ě`���� '��ޏ\�bLvX�R�Jy|~@wv��Dl#4��'�q|$'h����
��P�e����g�j�um�y�'�);5�����Pz�lx%Ǩ�G�|�<M"������2^E=،�|ދL"G��5&��k���1���֘r^t<��5=��Z	�u��=�/�;�������#�j�������0�r�I�h1A�jPW8$�̗�l�8���J_�D��d��3�lv�+��dR�r�HB�T��OE�X�܈���C�L(�ۍfh�q߾o�T)�~㱑�B,m�f��A���PU��]��$r���1 �:u�:4�uaY���s�>���w�4���R�r��"pFi��kwe0Ҹ�_�����)h�x:q�[C=���V��,�u�3��hWw�����a��P.S���ж,�Q���O���|l���-��D=6v���{[�EhI�iwIM���g�<'f�[��I|��'�Ľ���'�w��F٥2��mާ�CB�E�Q�޻�;����6s!���=Bz-
�����F>z=����u�hf�	=����[r����6�]P�s%�KY�$خ&�(rOYT�H��Xk�wä�s�8��s��9�RR��y�Zf���+�dϱ&f��bwJ��:�ly	�m�9�½H�JS�(��(����Rya�=�
���䓛 .4Of��]f}�8�W��g/k���?�j�*a�E�,i>���p��B`���_��ѝOy����8��7���O}��z����4��G曱x(�ݥ�.0f��5IK0"+zߒl�Х�\KI�i���Ⱥ��_�����~3�?5=n._��=�r&Q�R�vW7���
Wjd��.�����`=��u�>M�_�� ] ��@�l��\
�C�R%D3�\?���,�E
s�T�x�V�������Ó�a�T�#��%���E�y����I��O�sԋ	�_��A����U
�=��	Z��ž�6L�ƽ�v�e���1@@UY�Kd��8&@��� {=����2��./��������KO�.Be�9Y��ɋ�,M�žcZ�Y9�k@<�TW�߀F}UU�fi`�K�6���sq3A
��ׅ������C��W�M�O(�h�W���^s"7�2	�Œ���M��E���u��٠ ��I�{�?
�]Ǒy69)
U���:��L��O��cCP�ԔƱb���.z �AU��& 3Kb�H�0l�3����殍G+�Ũ���PS>ޓ �G�O�	�� ���a��veA;� ������Ql'a#P���I��	�7���5�R�r����!<G�ɯ�/�"k*f��*����g�W�B�˯��I����B��M��_��G1�l�f���`U��k�FX�7� 	9\�]�e�+�8�=��m֌��"�H X���5�J�/��N���{8��*��s��eN[��<٢��������U�~��T
Ő�2�f�;�JXy�x��I�Ԃ~�7��q{ɔ�]0gay���*a`k#h��Zu%�4Ǩ��y��8�y9j��Ն�� 6�-
�����}�t��Q�y���%���`)�)�Hp�������Gv�~�Z�k|�����~&z(���)�2x[�Ֆ��n��+�>�B������G�j<��̠Ku0��_�Df�IsBt��s�8<k`5�X�?���|/�qo����^S-]G�Av��`b�vQI
�l5�ES�Dd7�#��Q?�[�ޢ�M�h
��VnQ��T���2f�&am�z��u�}�bG1�ߟ��1%ϴ\6���f���tN����U�t&��i_Hi�h5��Ab7 ��S�5�ܺ�\������!��=]�z6����r�G�5�?_B�C��Nzǭo�_���9-���x�C��(���Hy�,�U>H/-u\-�(��b�_ӏxG�Q�>#o/�q�I�\�ձ끟�\1�����8��LR�'�%��_)d|%��1?c9x��>��q���M���w`ޅ`��ID޳]W�1�}���?�Sa�T�]b��s��@>�r�{��#�툈N�~k�|	��� =��P�׹c`1Xx�N���KMa�\�mh�`�d7�x�������%��J�U�n�BN�6�9�vG�K�S�T!��]��:ؾ��a+�T%6Pȉ�5{��)U�e-��G��a6d�)[��
"��u��
I=�h������wy���b���:�q}J�H�͒��I�}$`8�(� u@�b�$������AJlo)�U�c�3���
u�h\C��g/5�Z��X���'ˣ���o���`2nn�<rL�*2��8wc1�Y[��"�������c�V'u$o%�͜r�"�0H����
���0̦��S��h+�]/�q�م�$tjP������<d/8�y�[���ڱ7�Z.41���j>���$m���_}�T����}��"�L�jR����A'��h��S��~�O�����F�n���E��]�t�Iۊ�*��%�XC �Z�/�=����|�^�RO0EM��c�/" �#4��]Y[.sj���I� �I.��yj]������ա?�\}���O>%͸'������t�-�e�-��
ARj��>��P������!);�32~����0Wc��
�����w�\'����9o1hS�)BC>f�#�Y�*�z����u]�I�5$@��u�i��*H���h�1 �/s��ͳ������q�O��̾���͂v�Qy����g�_)z���}{-�������M�B�DPd��y41u��� �tE໣����]r:~��#�+���~�0C��X�?��V	�wM�xz��v�iP�	�c��t��aS���t��?e�1`�jP�#Yt(w"����z�R.��d�ʻ���������O�% W)"�/��À��V���Q��0 ���2Ζ;���u��@s��=X���Rі��6 6Ӹoڽ�X���_d`�8�N3b'M�u/���B��:+l���y��i�O�L���OH2���;ς.��� |��"��m�n��䶛.����5!���ݪm�J�ӝJ`
����<��C?i*���Wu8 ��li�|���mƃ=��,��5Vd��J�����+h��l!Үg�ۜ��O�����p���QHfdl�E��lU��x��:��H��x�Bu!y�=�����>ǚfе0�X�fG��A0Bs�p�]�J��g��8�Wb�w�_aD��*���Ԅ�D`
���
X�9�BʕL��#i�Q>C��͝�IA"x�lN�e��4e1��,�LC���n��2 (��g	Y�:�FvkZ?�G ��􇙡� �]ʻb�5cw�ej'����o�Хb�h�N��X�&�����;��D�^(�1��d�V��}
l�b[�A)�ѡ�<E|�<�%�R��R.��L/!`����7;��.�+:K7/�=C��li�$k�2�}؇���K��WA��
�y�����b#Z�}���z�Q��kɅ���a�[ �|��C� �OC��Ĕ���?`�[3�,<�	?��J��=T76���S�R��
�8W�)�9�e!�������t���)u
}z5�K)ظ�Tx_|���ٟ� B�s�~����h㘉�Cx_kMx�a%��ӝ�?�}2�k���K�my23��_&��G-e\���`&=���
A����W�3��[x�F� �.�>���=��`R7+�>��A�ؙ�.Q�6$�Z�L����v��?\�^�����I���l㏭A4�+@�:v�$���.hpp�m��ica��O��L����"���nE�w�+/�3���w~$�|�����e�N��P��z]\V�&�xɷ
��e�;G�Mt,<S��� �����/ʽ�!UlO����-b�Rk�C�x��e.a����\�@�\=��.J鼁X�a魖�s`J��O�x8�U�P���g�/l���8���<%N��}&���*��$�[�cao´����������+��)��I̗
�\� �l�����t7�y=9�c1���[��j=����-��G�>!<;��Q���,���7z���W}0EԄ�Y�Fi���z15@���5.������WS4��r���qEI��u����]M��C��7��
���op58�u�D���ʱ�Z�䥗����e���G�Wx�Ne�~�<a���~�$h qIetr8X	�=�����%٦���)���5�ޱK��:'�ȧ끫��3��FK�"�@�ߏq�О���c�8Ţ~���M����VҒ9�Q6�<���
5�A�vz�6@҄�^�)�2���!�����7k��}��ڶk��U���e�앺��1�E��m�^[>���:�b�d�2ƘS�N��SE`� ���\TZ�BKS�v%�������N��Mmϗ�3'?���M�͕G#(�:D-1Y����L���9F�����_v�b*+�˅GK[ ��ڛ}ɠ�`���O�y��s�@%-
�,U��)�Y����"�<������d�\�n�X�l�g�
��zsy\�g����{h�y���xD$W�̭�lʲi�Ǿ��E�[�]�}���٤-F�Ջ�jjا,0;S�QJo#�<���\�:l*�b� ��R �3%r	��	��12Ƀ���2W�m�_��<�2��-��I�����S���*j��a=4����ŝ����$���5�`��5웴�l-l��0��L�m�4@�֮�)�h��j6�S�O�TU�@�?�݊ގQKL��b�_3�T��`��3�h<���u�f��*@��GD�5�ʉ��'	��;$�'����!�nW����� !, d~e\Yn�g��an����~͝j��d7����t��II(�O�'�FvaE}�H���re���nT����ڿ��NG�O�֒V������Ȗ#V0���ci�O��$��O�r�O:�I�"��]��Ϸ��2"��7L4A0r�������u�+����T�ǹH�ƒ�3=+�|�1:<��XԊ��r(e
Q?�^n�`��F|V42�Ǒ�U��N�#@�I�P�ٵ*�7� a��iu�ew�
�2@��Z�3���kaD.�d�B�wxlH�q7��e���Oh�������"�C����1g��v�;�*�
�+_�4��r�׼������Ƞ�K~ʞ5�9-���D����)$��e�-}�%$�;�����5﵄s�Ir�*�(&2:f�����vluG�sR��|0�f��K�F+ZN�[��s).}or�0���FDlV;Dk$~��Tm�i���q��{�Qjá�)�^YF8��o��&�İ��E��+?�ap�W�һI;��
�|��La�4�j�
pתn�z�v���;64�N֓�ľ@��)Ư�oL(��1��x��2���Ow߿�R*�SäM�Wt�Q*�x-v�òp
�ي���'�?�voO��FI���e�V�\�q�:C�7d�goB����cu�s<o!��L�*{iv�YHR(�z�uiZ��vWG�<�ꟊe�Tu6t*��:#t.�N�N�!]�n<���[oF�&XW���VI�)���5`��xV e�69�@Cb��Gaa`u��X�-v��θ�����^N��-z���9|O�ݚ�coZ��hV�*��$I;���At ����C�;"I賍d$�2�Jk橐��#��FWA������`kZ���٩"����2�R��MB5
,�X:q�I�P�_׼H<�]d�*iR?хk�޷}�L,(�p^S4�����rJN=O1���X#X._����P�.��a��EF��%b�#��~�
t �cFٔ��҃M�DE�-D0 �{�U)��i���)�a0�{rZ�F�N�/�aQ%�Z�%?�F")���9.J�ڒ�Ck�j�$�qH,���*��Z6��l��EG�h5��j�g
N�������p�O����$�r�R�x������>I�u���`�@{����wjC;6�X�c�1���c3��rC*�I�h ����w�>cg��PV�'�ŕ�Q�Zp����F���̒C���"��):އ�?��YX�������r�����i���܆8�&�����ܶï���2�뮇�2{�XB�A���𥫭�d��9o�jI��8x�S�h���tv�z�K}�3�epE��^]�x��J)�\�tχo�0��Lc���c�gv?�����@�Q�%v{sS�Wa���uE�b�W�0߂,�2,��~ �OǬ1��vnQ|4^e��	����&��`wk�l�$M��_��;#�}r��W�"n��ɉc�\��I<�G�ޡ2��D����Ba"n�خz��5�����M������uRk�(?-������/%L���>0��Ձ���Qi��}��Ֆ��,�q��t��?	�!i@�q��<�&m5��^�.�"b���}���zOD���
,$�� ���@���_�F�Ɓ��;X����T�y�^sʊN"�q�*�&<ң���#r��I��;��H֩|���EU��&MʠZXm��qy�����j#6m��﬉,⼉|�j��Qt�=�h��G�J`�Xn���� _�6�ɈY'se蓢�B�%p���ğ�4�uPbd��c�Fi�[�}A�3B�z��S,�5^EX9ėb3�5�42�:�AG�חy��dO�`�VID��������H�[3�|�y,`;��ZuQL3�V�5���ϩ�����`Ĉ�⃌�¥�ϵט\=:/&Kնi�\,p=��ͪ�闏F���8�f�����2�ߡ�)�Ѡ����MH��ʘJ捲�?��&��ۺ�D�U�b�L\=�_�i'��Ŝ�[v������	��sO~�����_�iG�eC�8�~l��m��@7c���5��=�Z�)]�O�A�)t����zt��a$��#��� �n���Utw��$~�����}["�w�X�l�Ȃ�L�}ڠ/R�(��o��+��Q�ɠ#��|g1�>���2e���c��K���o]g����,��J1tf7�@�١�\�Vhҡ`7׮�SՈ�z�,�@D�n�A�r�,<8 @�|y��Qש��x�}�Rz���\��C��l��|��C=�jb%|P�3���i��6�{{����.Z7�A���ڿ��>A"�a6hB�K�O�B������e�"�H�z�QG6���x���D�8H����+e�3�1E�m���ݿO�7e��N��s(�7�ɶ�B�9����0�p̩�1�����8�:�8��O���@����k�c���U��L�'�8��֪h��h�߲a�_D�\�z���G���(iǲs�l�)��o�v��֜b�j]at<Q2g�����o�U�����t	�aԩZ���{��y�/뜒��&�ÿ��o��+D�it&�%�~ZIF��xwE]e@�Kfg�+��p_Z�E5"bm��ڙ�M')��	Q�Q+"i%�6H��b>4\�p�':Ui?���x��{��ĵƘ��eZ{�Z��'`N�.M`1:��N$����H�bA����F-�R��$V�LiW��ܻ�t�����& ���6x��X���!SAΐy��_F	��<�����x
���g�B���dj�yW N�q"s.����S�琱�!��k2H>Kxˠ���Ξ?�x_��5��-���5�d ��͒Ǻ���F��61#o7��C+�|���Q>��߬>	���Lh�K]J������9�o�[B�X��S( �K�2�
��Y����4�7t�mÒT%��*�r��vE�Ҏ��ϡ�f��i���k9N�Ǫ#cRp�@vy�P�Xe`:��P�i�8��a�^�n#�K ��{ұ]�Nk��m��V)&Bqv������m�F�N�W���Ղ�%�8��mf�=VH�����q��|�jl����5��GEg�w1� ,�������>ρ��O����Z:�P��m7��'3B������\�.��+F��*-(�2�Gu�����=*4]"�I��.4���)c���ۮH�R�,���o&�ϗ�ml��we�;�v��+bD������>T��x=�Nw��|���0�U����q^V��O��$t���ȡ�z�s��mD�_^sHa�F�.��TP:k���֡�"�J�4tV� Q��S|�����e9�uj�]�}�f�ֹ y�2�N&�/]@�����xU�Ր��Qt�f�%�A
��� ��KVaj����R�ƚw�B���$�&,�l���ݯ8rz���0�Z�g)o���^��0�k;«�q!��k�[]"hNv��Fw�]0,�7�d2��C�����"����L�l�l������(��$~�혙�B�rj�1���j&�x�F�����q~j���/۔���ܮH̤�N�$��,s��!��N��d��������UEaf�7Q�*���=�pY[QD#�:%�o+��V%N���zȎ6�x+v6<׿�`r�K����)��v�cCh���5�0���Ο�vxB1_�8�gn�o7�]�̌U`g��7�+:R��D��0Z��=�^����@Kʚ!eY�T�D���,�)z�ǒ9a.�,"�x���5��Q���@���#������X�@�ΔY���;��L��-k{vV�A��<*�v�A�T%�(`�қ,qz)�[~��$ݜV���Gn�0K{�mY�����7GA���Dk�QZ�*U����qüd&�N	]�#"�� �Fe�Ǔ��O\~�Q%�=N��m�t��2��NR,�����9:�/�L�nDE,U&���K�2y�e�=u�`6��I��z��z,��2��w���?�Lm�~
r��k>�'�ǿ�Cee�w�x��Ra��a��L�72B�����g7-M	"�Q�����o��Utr��<?N@A`ku�"`���^?��R�w![�7:�j[��F���T����S	��W��JXNW�R=.{GIg����H��PƋ�\�Hv��A�0��~��Рt��u2�k�̡9���s�1�"�Ǌ&&5�B��r)�G��_�� ���Cf���;B�{�����ߗvuSvy�=���b층\˻[���c�Ĕ�#���^��nɋ��V�}�8D]BT��	����-���=SJ��WG�/&����c��=V���(OB^�	Ui{��Fo���D/�(�z%��V�ұ�u|�'ӊ��k�SF�ʧ2��j'=p�U�Br����'lN�Z��x-G�yqt�N{�.�6z�!i�˴@��$�'T��T����f��["KPiǙ'���@�f����SC2tS���T�&�4����%>�����ʼa}߁ņ�S=[(�nJ
�n���@��o��XJp����~�{�gE!�#nz���|C��)�~3K9��ֱ����]f2d�L:i�M|#R�˭'q`�7�k�C�94���@U^�)��ӊ쯨+Q��zH򽓳�l���s4�"5��?F���"�k���u�Ip�v�!^���q�p{6���b�S�j��>�:|ťh"ַL�I�9�y�ǅ�w�\��L|�����w������7ω��\��jxI��V���E	�ҦIJ/w=�0 Qɪ�0{� \6����a ���_Ńt�(7˶7~*v-ĥ+ǫ�9�-��R}4e�֘���|�(���=�~ᐨv�k�6-�1�,~f85)r�Bz�q3�U����$�ww)�)'w�/o���o�ak=+Yq{NWs�����}Ĕ��˟ڬ��P��R7,ML�����8,���ORu["
�g�l�_0��e����F���|6�W�[�0���>�
.�*S��㗲���L�%�4����@N��C3�#>*�>�6w���V�=��Ɯ*8p�5l�p�O�isR�m4�dP�t/����׌��(ggY����l�jZz7�w��v��5V�:Y�K����Qʬ���L5%{����gq��t���h�Zh����t�<�K����E{e<��^_j���܇�(��}x�^ʕ��pj]"�RK�<��2�	�@$mӾC=��Y#${�U[2�s�����ҟQ^�GQ)$�>z����*=�p�=�َ��+��Q��o��^��4�O�ч��3l���씄��v�o^��v�c��6�G-��j��8�� At��0z� �;��<��� ���M ��a�K�j-�,��]E:���H�����Q ZdOcsZýۍ��|����u�N���-kx��.��H�ůk�8Nl%�����i�,�bc��R�ӟ&\$��5�
��`�4ݝ
�ni`{И�&��9dB�L�.#ܺ��W���C�/�^�.�r(�E^�]�8�f���;a��V��ae�n��,�kU$��A)k��"@]�B�� ;�w� �9H��z�g��Aي�\#�%{S�1�
�k�eƂ�F4qX��V��?�3�f"�
Ǯ�]Z��.D��#ܡ��3�y��5ɟ�
�:�`{/�s��ɑ>�"VYņ`��G��ތ2�mt�Rו���x{�핈���bW ��$[����F,�ۻ�e��6tB��7�lXpZ�-�m(�D%܀��3�`c�zHf`�t���X�ޠ	RC+�GX����>c�BT�{�)Vbt�%�k[:�ۘh���#zw��uzn7ZP%V�F�=���/�A��V����X)Ӳ�����	/ӓ|�f����ҝ9A�h�<���M��N?~z�U?+?@�G�����&G��i6�P!���U���2��L�6~�m���eWv�2��N�G�?Z~�;8�T�����nO�ݰQ��UC���}��8\�`]
�Z��f^Rn�{��*�\�e�j�w��-� � <�p�Yڛ�[�`FAZX�J�3[�[�w�Dt��U�`���g�*�i�Z��?���Y�y� ��D�Lh�1� t��E��[�4��I.SJ��nm�"���en�G?�o<�(�cI��ο�1'n�	<D��s�q/4����n߰ �qdVO�M](�]p���9BC�d�j��닂<�5���1��D�������	�v�="���J�蕨��J�R��M��n�B�-�vo�Z�H,bO�2�и��P�����C�\U��r������Y��/���~�:N����?�v��Ynv�դUIӂѻG��3���i�\�h1J=��qn���I�q���T7%v�QU�� ��©�^�vNlS����0�ѩ��i����&��b�{Z�K��BB��*��*��'�����ik�\0�]Ӈ+��6_�xn�y�-R�&ǡ񬗆�ɟ����j��Q5�RBо ��xy�Jg\�L4��o�&�E�i��v�"ɉN!���0s�fu_�"449&��|�k�Fi�^ny�+����Z�+���J�7���yv;��9��&W_� 3����%�
�W�;���&T���x8^��B�kM:�dF�v9���y��Z��-XԱ�Fu�h9d�)���@IxT�<���էw[�1(F_#�{��j�7O<`U_�aRJ'��4�>��n%g�d�+���"�%yn�����tã	�f��j�"U���������I��Ki�����'�H6���ߌ��C<�v��;m�9bx�wvt�����9�$�/8`[�v�bu�w�����3?�B���>}a3�m�k��3%u��9�-��|��t�Kĥ��x]��I�%K����1��I�Z�ȴ��iO�Yb�bMwI��mNu�(�ž[�DE#:�ˋd�5H47&�$��X�Z �R�ѫ��8�Sk=�`\�T��{�[i�QK����|��l�(5����)t*�g�F㏤���;�Q��Cо��[�C�����:2:Q���^<����n�����z��:����P�F.����<��:_����(\����1��.uX��M8�c$�ժ
�s�N%?�(����[�FZ "	b
a�ȇ�C�-`]a(��~?�fq����.L:q��m�U�lO�|C��,����J7�؋�����.�die�z��#)t�ע�d����������
�\3�&#�?L�ke�?P�w͒�	F��M@XT������B�\��F�Fc�AN�ΥXϫi�K���zh;q�9+��B �5�6� �d�	��B
�A8���B��� (�JLs^01���ڵ�%H3�zN���Æ�4��1[
L���GKM0�EXώS�ɒ���gG���Z`��!�E���o�UM0<�2��#��+�b�*��T`{?�s��7�^�i�Sk,}�	*����v|���ׯ? Jq��4skb5�j?r���w����b����)y�VG���rYc1�\���L;xO���џ�;�'|qc	Ly���b���Rp����wj�W,�����C�'�;1i�-�u5��M)D���ȫ>T��D��������-W����{�u8M��zV���=A"6h"(><;Pƹe�,�h!�Iپ7A�@�����������ۣ����h~7�霏W�fs{�n�L�4i��O[����3�?�+ E��� #:|_��g����bj?�G�Pa�𪢶N9���I%s�1�g�5�ѷ�80�s�<R����G�������b_=O.)�9�͉��\�%M(R�{�֟W����(t���q�(a�?��;�23�c'BG�,1C7��:��o�~�l�B%H�T�رr5`跳>Q~pi�@+[�}��[컑�!��m�t�v4#��eס���f���`8���R��Gh��|E	�LZ<ޏg2�76¨(ĭ�����[��֯��h��*���S�&r�����;7F�bT)�'r�"p�%g������4�U'�F��㙤%`��y�;C@K����f�n1�����^��/ ���ʩd�Mm���9'�S����� A�l0������,��-
̶�X�"�m>�3��`N��?�b?C��i�V�)�yER���^���G^���0��>{���u~�1
�iX��9%h^5_�L.��PG=������>L�b����7��k�drݮ��Ί����t��r����1��m�p�\�$�V�6��V�9۫�F�>����2 �\�������wU�lz�\�v��h���	��p"����U�R�њ�a�k���z��M`Р�$�c���e�Z�B�-�L�Gp�.RlɛC���΋�h�R	S 4��Aح����N��OfyfBF#��t�BZvF�Y3���W%1`��w�:��{>ԍ)�>Jn�;{4ͼby�q��5cZ�M�?�L��m7y�v�����r�l[>fŉ�<�.k8-m�����r��"Ym�}�Z����]�8aw�Gw���d�)���Ґ���9�3�S�[��C���h'��Sە�TР�^d3s�m����y�P,���
ԣL��}6���#K����7|+I0>�����0X�����pL,�*�m��*�D��̾.xO�Tڱu�6c���>	��"��M���V����J�I�2�&���rYg�-���M�W{������<���A5M��r���f9nd��+�G���5�CF�Fi����^V=��-ǂ�M�Kv����7�Mے�C���