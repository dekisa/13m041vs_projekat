// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:26 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aLiDXAZX5HZ0mTneiX3nnZ/K299idM9nQyFX4v3ptYzoVBopfvEDcZhEXQCKVCek
IXNn0bAzAr2ILj2pMHp753QBWThlfYFJHHd2RpFzCXGpawNXKplUPfTMYwYxib+x
duYio2zoNJDAm1KAkKtK63r2JtumhVDmJtHo9Y9f9UM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6576)
iNW75ew4mDHZMtESEOwPaLruBLEqEDhfuZcdGCTnthTytmStLaShaevTGh3AmMCv
a7KxIz+3gjTxuBUlchMoJQaPvDJ6UWk0sbx2IsYKs1bGyqcewh4qEKj8TGZtR7JG
4QTU84dWyTg4ff72sLEOfyp9lRiAr08A4UcLAda1BlnYDUg2l3F/TWrNcR1pvz7j
59imrY1AF+1Myge3awhywIduu5vYOXRa9CTTryyhxyMM64Wvo3UYkfOLqEpvU47i
RnLl/+FaG0lmJPs0YLMfyGBTylFvcYICo9/apMx7hHFYKRe/aKjviyfgYnMO3LZA
yAa63cOWXqHWNehmyPKVqrOQQMIyi5ikUp9L+MTgi9yw54g0c4uJa9B8FpxxyOZS
5C7CKkwUekTiIjzOj9ctvEhB4bj9rICMY6QkV92f4KPsM58zVyMMT96ve/ibRdt8
xaYlRH+BiW8Mzg6suHtBpKUC6Kilo8BK07Cb9vwzuHX7G5OWSQRwLeEH2YIgEqAp
lsh1Cdy2jUJiYcoLuw7CqRi8fFQXZSWOo7IhG30XoFApe7dvgmY6zYMSiZnZFDub
ryl2d6S8Wu/zqBv+TlWWLMAPfApe1xck6aDw2hg5dk1Zh0e9VSUlAvWrdAYxSGJD
4/dpXZGoos9FFai8Fw/BbzUsMfNRo2DWnTFt0EhYoOU2S8pWqDq104EbO1lC8dg7
TNZEJbe7ZMidFhWuIkkKKvsTUkWScLVhqnjCBP/0tcrXOLGbIBcHRXh0RBnB8ev5
b1Kp7f7exRO84xBPP3k37a3M+ZlAxpGdQkGKMAJoGIiqDIWsChfjNozA7gUYHuk5
L/E5UpEBGsCt/+E8W3GjoBU5iLa/nS1ImC3zxIwh10qgkAoDfcUEKHPS+er01QXy
oqU1GEewPOBJd00tqGJhu3xibmmNMqu+BxXlm2qrfnkljNUKZaSilnrP7pT3zpP1
JTuZcXhGW6lpJTE2N1M32DyQL1ZvdU2W2Fz64MUUM0Hrhd1ZhQADICRgUG9Hdcqn
e41Kc3YxL6Q9CbTPKmHaCwhW3ebtwb7b5xqabIzq4ZCwBigRi/NJf2PFuQ5dBNeA
i4uxgLHShOqhiXrqQBuRhYVGmfTbPvu1+Ch0meJ/7+qTU8jW/JjYpxKOtGBHk+2u
3FZJw3an0dcDnN3yJxXjg7g9Ji322hF9wyJgYYam9KTtdLj/VA9ACHwjU/k/h76Z
nAHZknBS1Meb1gJ0PtSIVsKkSkp0FPskXo5g+43m05zGqxoie8XQXww/KAw+cSOp
aNdkmMJPbSJMJ3Z0Dbt7iMDTHCW2MUR8TDLCcNh9pmsiKtDswq3Xlgw5whwetmJy
CF1h6625j5PiNxuKhECZ/qM+YQ5q0U66h82wiCKN7YDCVB4FXz7nhkKjCpaBrAM0
K2ODTTWirPWnn2GjjBT3hpCoz65smhqByQq6k24MCUbg4EtxDgu2YGs8NH6xCusH
0KoQT9oOwM86l2SKNkf1qQfqoXla1Yk+jnn2gimePFsUA+LYByqsPuSW24o5BGQ/
yZ307sddrNxC7YF6u5wCW2yZRKOVrLTeZuqXmbLcngbjLTFSPV7pQ8YxyBQCeBIS
zuut0qsTarT/RRjUOCE6lhYTxT68nWaO3gfqfAxgGydFRN5pEPy4EQKq54AKTd82
b4JGABVhu0b8X4zWtzQ6uCmAN4bA+zxvUzBec6PSbV8Qi0IUcmaKgRj0MpbC8M/3
+sHqsG1tER+V8mtD0BmimwpaUCUkU41wb7JpwR7XWVM4kJZl2Wc9it1oOQ+HX9Kx
goCv61Rj3masU5uGUjYRljD8QP02bk05SOiCNZcFCTFW1Oj3EsEd1GjEM0sWBlsg
WUKQFFPQPG95KJxv8pbHpkf5Xt8tfQt2j/rvB1+/2aWWafTKHG0Ninp1WmeevCEO
LN67wgDnaVIH55XkGw0btuftFKqd/fnWChmrcRVCNfrSYXnbIEy04MH4EWL8Cx4s
frik3Te+fJNRzLxReqDYl6hppXJ9BaEMxiQKcuBhQPSq3fOhYCxHKCEXeZyIpHDl
ROU3mgQcUIzR3xQxDJ+H2pyLcTttoOTpEyj1Vbd+yQdcB44YkCmTa2KqLKvYZeLQ
PG/BNC+jAjuQkM2/13rXmMm+k7jNIiqOy/x+5V78DObVw2OEUHNaYGumh1IrBMXa
7/8cphz3drv/yLrZ1SLk3T4BVZEMVb9XrXp23fifsGO8uRvU7YKRZgSwBKO8WzEp
mQTnwf7Fgg2LI5dZKf9JDqXeJ2bcD4K73hHXMhOhQ/a3aKHbOnfbRO12xqqkQIxG
Ze+5NridWIRW1KH6RUzTr2RaUuiqVXcdFhqcZ0W9NOZJqGvdikSmVvbT3YLRfw1S
y3kVKXNm8o+ML1v/fg3MqtqvFvW5GT9a+y8p7jDx9LFllcfdh74FtFb/eIzYHwj+
pDDOQ6FlrbQPc6vJbf43j9Ic9fh1w4gMLh4Z1TwS9BMksfhM9bcK7l6as1ObnEF1
eb9jy3cZQvGcJgxWjSqiq17Rp2Zi6RpwxRxBKAqyQPoI75Dgxii5xqCEr/jxrAPy
Cp21coaQCMtpXvw16oQBjSlHOv1sUgaOQJGh1Cg+KsdLghjxgDvZDrMQ02DXRFsc
6X4UuJFRra7nGDbwuvAhzjd28+XxLpAgZysU9VNMxdplApPYyRNX6Rt2iS6RYg5o
S3fE/f3tAJcg9MJtmUzsPy2sFgTJcXEPjsgFcjHHEEKxgqx5/eA+OLHyfhUCYUve
bla0i7kmQ8dSTGI9UONEFJmSgxnOiQcfcyjtP9w9BkBbJsCM0NPsN3C5mBJvSbih
VqHzLS1MOyomr0Gwj4+J7+mSIr9IcFncY12ojbapVcmg6xZMWjDOFDIzUJHVoNMM
hxCLr9CQvw9LWtF7DZWMaZimj58JGCOAkOYNmG0nF1ZH9pnhH9aTPaYL+XXVLvQ8
UTl4QOXm+SoA4BbX8bglVmhCJbD5K/vDS4XuQuFQfwY2n62zsBs2zMx2ZbG3tqH+
DqqaWlRLQYa+MXWFEP/lx9l2dwQmJBCcI6Vg36faMLDrjEHKKVnC8cal5ly5iqLy
2NXkNVN5GsTOOwZTgn/YiQNzbcOO9aXcWa3lvSZatLZUdcR2mvS6U8v4uUtHIx6n
XY3FZec8EHSGYvsJ2Z9oY6yJUGSdoA2e/Adav48CQ1kGh9YdeNN6neU/V/xix5f3
JRtdbrTfsN3+2yeiZQpNeMKZGro3juDjxPjrW5LjkM5aJkLcsEReNIVfq3TgY1bT
0au7BUbOzuQ9BLwJXnIVpRZ9fiHHuWbnuM09QKupcPGdd6rx5h3VpJlmJ+0vjGhG
2t4nimjRjqxTWed7TUvmw+mjcI6Qf2D1H+aKffV8pwTQO2nM/J1berbKWXAoSSvu
1XfZNrCkxQG9SygrUCwv7NAajwB57+t0GEFpj5Bk9lLDHia3LPl1rTflrkJvia6R
yQqkXul3HE4UHqfGO2/ErxL4Gp9pdB7BIh1ckaZ8BmE0HgTfWXTv+C04A06YcZi1
l46O1U/g6mFTZ9oM220CMHYqBFztZxiYZw1oHZ3PBul2CmQ9ZjMF/WV2QfC642hm
uekv2++nK+8J2utI5GYRkNZ1RCm+SR+k7VL1y258Ps3InjaT3US6n2ChyrHekmZa
dyiKsd9aBCNGd8NhG5+DXekehfjxjrokWgSl4NORrEhSoLljEhUndaOe0JlkQCv7
2MaYWIBM8zVm7bs2Qy763M5iYYNuIdRpeLc+ufptCwg/YEmxgAx5KnZlAf3j+Dos
WcVK+fVG5PvevRFPlY72nVUO846uULYymf3TZmtechWyTmvwD/1zJDRGljgLVCte
+4enZqhrlGilWNmJd5OQFCWBvA1Vng752LTiQGmx7NPTa+sXbH4cSQUjjelBVFDh
CG8wi/tU7kYc/7Ka6tNG9q7PV+74ZW7uZjXezaiiboIr1ODg6YSQt/5CxuEHXQZI
B7wl8tDmgqIsbal7OLGZewbmv3XakGEd8a/xR+8RWoEG1UGPEqU7iFgzupl9jGb0
JubawnS+J8y2QTP8C0zpkFhz3tW17Dm+y1sQKxai1EhUgq7ry/4xfHvQYKoE1SAP
bTzOEQ01S6Gfdcsinjt+Bpbq67P6D/A1wbO7m4jrOjY8LcJd5zg9LVWABEzOUAUs
/zGH6AmvykisGxygVva0WHa4xdVsenEsLR6b3WDNWzpxk5rdU+7t8NzgsZzlG0jX
Eg68AJNd3CUhxF1Q1Tf2SkeT3nC434HQMcFu6VBJcOQbBaxn4Gc6rt71i/v0a+mv
r41VPic0kEi87mAih/8ka/0NcD7JYXkvNpF4vqVF2Fkg4H00x+hHeOuzNvLq4MXU
M+0gGubeMr3hPTQQQh34NWKre5Xz7htj2qKL48wsXrPI1mZZ9E+aLAHH0kA2c6W9
6Fwp3yevilryBmtL3Gn28pQq5pVNZ/Umk9zkCTLDUcMDQhI+Tinji5KaUchfzh5E
rHk2uVHcChcIUfPxhl5PuxPGPZtGXRnjfQzYHGVMEIIAa1t+zVxGtogBC7o2ZyDQ
MZZK+Cu+KD7fJGBrtxzFB89frxFUN69dGrqtMZKVBKOite7DZu4AJo9l01cZ8J9w
AAqXpz4MgKVxnZf3AO+vTK1pP3aBzygtzJHiCBD1XAM2IMin9AT+aXZKByia4fZ/
sNe6w8OuGKBzmF4p7WTDJ69FQ7RZTA21ZxUw01EOghqQQSzgmGLK2mpbkRM2Jr8v
SdgJFrGM3sYDS3abPetQ60oQQfGf8NSaeMypnthoGYU16LVlgwV+o3MdJpd03hVr
diYGgtpUXecc7DXgkzlxlUvrTiCdiEC4GSIvAG6OXe95jU4laX/y7fDpSEdyoZle
1OsGyXnc+FyhsXFgDnqvShEHlBanklz0AwZXJuDifMgDhvywFyBrHzQW1X70E7mA
lF42ImcIyiF2AsfOFReXtEV7Y49m/oQCj6eNUjWvpIH8ahRxzLbTB9KDOHYvXos5
HYF1rP9OFyMTAdmoBmJHsz9fR8AJiH3tILdziWMFFn2B7b8t1TVfN7dGNXXlU9Ea
nldnrnc6mOyj0vuT3ayM6l0WiF5iX9xLN2QQf6undglhBGNMRbV8SMiz215g5lCB
aK3lmr3kLMjShn4ozfdVXwVZz/RWKP6/O/TG9cbfA0f3Wb+rZ+/0xvPiWCVLCdCi
kggmrz1oFMBDw7rVyUXfleQCqFN4x4gbVDft5LdqUMmGqCez33VQ/xv4WvBovHAP
GtWEqSgI5HR+dyGkNtuQCx/jHWjHUxHG2gXuTa1+voF81phms194rWkHkt8t/jkL
pb2oQdz+PZdvkI9JFv5SyqKSz4SlwnOA0fySUeZuvntRlYwOOQ3GPyh7sMGlPaWT
Slpgn9bMUwxhZ9RF7arP/UBI9biPidnBYiASoT3RQdMwmQGoTqyu5Sxytq6DUPAW
IQ0xgnHowOT2U1hhfn+h4PS9YEZ4szCHCF9WQvHAHk/puRDTCkP5jditMnGabndm
J6KV268LY8bvwbaxjkDGnPRW/BggVNrbRD2agiahx0o5NJRwLXJZDkel/JrSin3f
fZZOGzwg6dTvAC9iYclBRL6matcMrvCawOTWkO24V29IOR9+HnnmkytccX+L7hfi
+wQ2Wn8b3MHaBohY+h/MnYZapal4OYtZ384B282ZYtp6OvWBHnYVJZ23hURiBgOv
YjrkVczxLzqZ+3Kz9Te0d3xCH3zZ5b8niAxMH5Jdfe3/3fzATKfekjaOMGj6lSMt
mcRBicTh8swO7WwS+JdsDcuz0UzMBxuQCmSeARcejVwTXwEk7FjCsTbuXMQQCk03
a2IpeB/+ose+zKMaIAbWNYh7Fz8zstDkUG3nL/9EZDniEaeOLIUgk4X94DXMt845
wVCrP/MoJX97u+dGSIzKUQnxDkqh/BsPuQ83V/vAxTGYR2hPGMUha+BJfqHpt/ql
AVTXU7XxvI+01OY7Glsld7tYfe0LKCBkRk/ZtWOqeUNw0kXhV6tTcPhjf4YMzXA2
Zo9MbLyqGw88DGmmLInWoQvdEhUanR2goIPK+1a8EHAjZuaeOaC8nJ/3+Crw8m3d
SWjvrCWqHEpdflA2B2/zcugm1FuFN5BPwTs4lbqzsINoR/0AhnIo3u1DO5AyV9dw
6eOMcAxII2fcre1LIKSRnmZAHoRlRjixNN7YvqJg+IkQEW3y33nra5Tp6G4lSZN1
AmsJSuA1jI5Qr+9m9x3Z48GrxbU5W6ZnNbPmGUdDYCXgXZxs0LZDXWtNHJ7izAqK
L9I4vfWHQf/iwKQUUDfoese1fQT+v5ZoXPh6cU+sKgEPkIA6m53CgYbLTIDdNjD5
0Y1TR2C/Y3n9GLk6EcxR3ixRj5WxsFEY3UAS1Ph/1stnAt3dYELKGjBbtW31y0oO
3HWb0I535KiiMwPQ0aHDsXK2XcT2lKkuiSTtDbqSvjQCj32H8PMx+GicwdvAjgDA
95yl0sQu3tR++aqoQTxNYVwCivkK3ATXs7YUC2IFBAhJi1/qdEz+kozwi5lFZMAM
zOhr1W3wnkHfn3bFPfYeANitRXCwRv8mZfYLk5eGEIHYTHR/QJFOFSqsX+wuX+ke
t9pqNXC5mtyCPg+NKxK79+7dKH09kUPUNpgU7vp7QeCYzo1v+dR3J/J52Zuk6Uvm
d8NmE/cCjUtnvuixkhhMnCV88Eo8zW7gxHnGRdohxgJ2joKbr+P0FnKrbre0uvAK
y+qG0CdKiekf2DIFWYRKxhC1ZbG83qa8dgdLd6CH0UZHwgcvIitkM6OewO1L77Tt
p0x57upGjZX1wP3jFWa/lWR3H8ZN1YHq7YxOY+MoFj9F+5bMuE1kuEnHhmwng7we
gDyQf+QaoejnmWwvV6EpSmrNvfoZHzOnWIZDYdAQEt9rkjWDY/CnSt5jV2ufE1qj
x7i19ePDbiz/3dt3y+LLEDwKh0eE7eQxZIWSq4uj2wwS5jzh4Z0ZR+45GI+BEF7a
W6Y0L+hfbp4bKRopJ6NnIt7ddMhfNXNL+uKY8DG51kk5m78FoeLdllFhRxSzAVWF
UzLPWUPjS3wlgNiCM0Y6Sz8SqNCdqyCjDxBoFkFdMp47mffayxU56kxeosdl2yz6
Bqa8eITYy3/o0FyYUe/+3hTx3KFzwenpYPhAIXNiXZjlJ8QSFOalGJ9D1cDaJyno
oQtVdfNuSxb7Q4WtgI/EllzZhJYIjj95YEfMe9h4sPFLbqYcXlPr22cShnTSbCvQ
ziaUv0mm/NOMV+wopZyPMkQjnmGUJss+6QC6KlHefbFMrW7mZBm6wL212hW0V4Vy
17bd2EooMSKm8ArfmTjuTkNNO/ZulkJtvsWOVz4f3fub3OzJQvvZ6+ImLRJF1WCG
PSmFykhBAxH344s6LOWrpRUnpleTYA0o1w5o9FXxAt/lserFWRzHJ7iRdldGmogr
li8aJM42xiPcbG30NrhSnLnpSqYaklJlPCJuKSXEzLFFs0r0l4eWz8NR6koMudN3
Yg/QM3w2wEYDz3yBGHnCviGcVVZoX1jJJoef+aAeX8AaIrPTR1PhL9iO0Ap3Xj0u
Us2MwFHC8/FuOAT/CptL0BssCWuLOFnbeQzHZxmClZkPODgeNZdzi5+6G/OTU56M
YmlrpB40faVCwrz5au78/+KP8xK2a86M2clSLUBcAwMVD9ixd3iC3VWG4BzLFTKv
xiLkpDEDyJNlIo86ikqCWe+6zOzWhN81qctqjUGmnc3wjNsXdddap+pUNAa4s3gg
o5hyVCP+Ks9uh9XZijMF0F3/yUTGDuzmZmr1t7he0Vheufcdt2rcTRHK5i5LaPnS
b+5dVEgE+iIHxUABFGG0jJNKoT3TsKoRxDWyXNdBqknkDW+WBdwXl2Hi0n8cV7zb
R26eKjtrzQ5b5Rp5x7uhpQvOg9CTtyGkH1szBGolJhWDhtiqrwLbHMkCvZ1zmW2V
a4jB0yFvtTWWJKMTkLhQomxMJDSeasqBgZ0T9KZgT+Zadb8LfJY8ONWwd0AQ9PTG
KXigBhh96LEbl3KFSWoM7Ntmpe5bfMxjZoZY8E/DobinrdDFHOnM5IHDcgRsvkzV
iJlcG0Tx8HE1L3zhkZ8GV1kfNZxGR0L/GCgw8zhfdxZwWUrk6hSsxKv1UnsPonsq
Z5NCmD/VRg5peakOKXQa+VXCpSUFbIr2yXYSthye2q6UAAAvBecp2XuSM2jESJly
JB8kZETQyU7pb+HRqors1oOwOVqMm97/oWnBolWlrnaNBC5qTR4WfYd5In8rvw/g
wAuL8pOVD3hAuION4bNEiNb+PLwStL8PZcpFwZogWUWBIcUmNk2TtI5dr2+lXhD/
sYR5n2VrT/+vBMG/OiDMSaF97/VzSEl/2t53DVtpkCxnha0qvBM9lindYlvN2+Kg
KF5Uf19OmLEVi0jODISJh3s0B5P43VmG87qSYxVNRkhtZqgG3GPisc+yvfmtjJ/w
qkK/x3xkiOpThSKAS/Cn/pdvOakmcwJFBX1O3VTcnYU7TNh0UPhZdqXmViHHInXv
haa7Gg9bWrmhP4RDzbbzlDIFUsVhZkgGKCU2JX7KtcdgOTHl0NJvAf9/XwO94z4S
b68PIo4l6otQlCJPemJxEE2CP7/rNYhGZ/cHSCi+D2Z69Z2zWJim1+C/SvrvwroY
DxByDI8Pyjrdqg5HsnqaWgD/2rBOpUP9TtVqGtfLivwxZaS6RE2rk9k2ECGhXIGS
1hWTN3PGlOvpHeORyPUQ3NHuUBMc+dx/LSaJ4EO7718EnzS/UnRjEgR3nXPzcPlN
`pragma protect end_protected
