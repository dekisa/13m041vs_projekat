// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:56 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dBF364sWMDbYJBUXuKM4QhfJMdcVpcd4YxOpOHUxrK7pX7dAI+h6SHnDHWaLgWTg
ngy2l+BqpYglXyEnh+ThVPFWgpwUiq65zpjpUO9yWTCmTnOTZaMMI/zmXWjEIXM1
7iO7jUwjT2LZf9gRw9kbP15fS8r+76CQ/FVoWq/ci1o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3216)
rMVpBTXw3xkBC/d5jwRee0TwFQlb942v08dVhE9Ln32paKC/r+e27w61a9vGdz/t
1BcE/SlhyXZz+MQfVS7EZFA9dIg+mKRuaXg1xTjBT8TLw5mWeqp78HW2Vvmy25Vn
M5P01DSN70P+MPDAoZggYv+Y5R0AM9GuDR2OgY1phpe+RzVOB6K02nqLtG5YuqCm
LW2/YvYOzAgxlfdW4GEXJuDjj24198kXSU614CGss7XjP7t/tGKym64jWVcN+0dj
WRuU4BguST6HOR8IeX2dU7WP+vLBto+C+ZwU8u+ll8mLy2mlWKZiCd95OcTt3OIx
jJGX1Q4dNaZsmROmdA73YKJbal11cuYnBLJDYEEf2h/MOsF94sk+2lHExDhMBy9n
gvG8bW5CtqQSUe9e+V5pUEqB0SgeP0N2p29AlALSJH3pwjAeDIoJnVoa7sfq91Bc
cH/J1irmRBmeEXkF/wv6CvfzTTdWAvI/UZUs5qMFQnU1VK3pBp3tg+Q69wklcNey
R+SqeqW61bK/aV3JpFlvmL62rUUQ5bSNGB+m6WbUy5fG6wt9+Gzi7Hoe6QDDN7SI
f1+S/a5xchmo3x/uIFbmQjNjeQAjFoht5bkZ3PFI4LikCq1EVI/KldVjXbq/t36Y
k2jlPkJ3lzcVGN9uq0m68lSVS6GQ3BF4sR3Qze5q+Gs78soX5EM9hsKhexJPiXs/
/grNtm+0THUr34UBF2JXU1N++bkaXYm5c7E0Gz2/D77YZqQSnLncFqfQFdtWG+sf
lP4lzFIaSSBgDakqGTsj9i9i2RfAyxd27dXiEmNgvd6Kb3g/VU2X615x86n3npwA
WbxFYBGx+lYLk3xHZyPJvvQPoBTCV8TEfxpfWrjkjiq0BQ0ne0VEhp1YyoUKm+Wj
ZMTgwWFv8Ts8249nh9PiwMqAFOds4J40ckkeD1k6ig8uIfurgtwZp5aRf1lcmFPO
OjCPob6cs/XZs1PVI5a4kjx++XvILnubcxueEZSdAuQb5h1JEEGFnlmQXIEbIppU
ZANUEGBA7WKKM0KygflMyOAYsr7Z1JP2nr/Olfdxc2QOeUj1M94srshfcgoBe3jd
zscBXA30Jmp6rH4H/3/hzORwc1tQ/UGEzmSUIXXsUEgb1cd7cXY3ceAb6ZiaKApP
UwIHkelX2DOga5BnfwVCqcpl+lQTTt9zdZwLe5CJWY8TJay+yPPG/glhUP1Qwrzt
4rTucOwLgO1uToz8UCAkPNQupeNBuV/tlDYkMaRLC4ghegS0DE3N45bWsnSX0wgz
YHtOPsTzk10WH0FYt75pwFQ17rSoDUO3LPGPDduCfhmzhz9FgF+TlFZRtoI3E9HE
d+XLG69A/Fd01mLOVrYZFXnXJXMH6v5MQU0R9bcRa9TbwtfDUkGdlrjNaJdaJVf+
0S2qtpdwFcOg01HHhSNFkqwAuBn2+EdVMiltXLDY2sNKuX3Zh1BxSRirbjLz+pcb
HJsgQUGK5IRR3gTAKLp19cEPvux12xH77Rfyeu1y69lIb6dkEze3SjRPTRQFkGHh
OWJ8drHX9B0X+kxsiowP9v360f+8XV7IZeb37HKONXMQPe2LOpWNquQvf6XR0XbK
bBZ0nE/gRfuqQgEzP4nmIDYluzUKkrI70X3KNH5v0hvGPaPTTrhr5pUlGpPBn5nr
QMxjEPgZOmcBDbQa5ECtFxj+YhfYkFlGy13lhEFfmbeExBYLDBvuYwxdeV5E1cS2
9THRPOzg6xFhDjhruIhuahWUzp8nXeyzPe77pVC0MfXdekv3r8syIusA2xsibUqc
HQ+n+cHZUyU0SwKYiT4MAUj/8y3KMXmIRwrBSg3qPQ0ndLsILJreOOnvwg2M47RM
aOA+c7HUAU4PRTlCA9sNkZ05itlc4T/7tz2bpz7zVqlCnfw0H3r6VA+kgdInWsUk
9XG76qgJ5/L4HMGfdHjw/ls/Pbt0fXSv+WBJF+zT4PWJmmiRrYZ166zqFaE8SB1E
iXSwv61X+phkdtqx0PyDqUBLwNbDmBYS0HiiJj0wdPgFjNaPRuaoXKNJk+wTIWG/
UssMCXcoPffFNLaPp/eLOLgsBu8fkWO/VKlNZwzDvEX99lCKxbfmHeqdiAdqr/7B
KqnT69/y9rA69iisXPiUwY3vggl9eX6NspFNhShWR4G9nbCqclpGfpHi/7GSDcEg
m2OUMj+EgruI1wOEHF6JbwtwZuf71Oq0I59ZHLdyhNcqNH+qRbxEZfp3WOHho6FW
xJicSyAVDqkfH2T/GYDMIKnlPZj8Km8d3Sat7IxsOpnVnwOmwXHAvayqd17SdFvC
DVzgbZiYoBns4gYXHt0B8DG7DAP47Ny97ST6PWzIlo9o5JCF++OJ/bRColnYpjSV
QjyrZ1eCRL8BhxAApXvAY+Z+7i+VkxEHVEqjZ5Kqzwj15IPLgiJDa+aSusji6s2t
32dvXpWpIDkviBrMnBxmzKLS3CuBOz2jkOIoWMD1LFEG4HqlRB2YaVJf4OKEU3jG
hI/Ru4rlQHdL4iH6HY7PK710no6TmHyl0CMnhUylw2BOvVO7nx4R8co/goIc+QAb
5X7ePDTjowcSj16k/CZa3jfwjArSFyJaCWkIKahd2C2q07W8bUibHuDo0jWpYoHm
Z0jLKEBDfUn2aVGEnZlORTTW+sf+tXFQAYI2ghLHDp+k5c8h1Jp2FYSBPgkF59Ns
+vD7yR5AuiPEWXMMFd1V80CzPO3C79GUFqdtoUXAzm2AtLTEUMFDQWoYgnNuiU+G
yu8gkbkIsi1TdnPEauBvk9IDjK1ggqCNTo08g9tqurm2BuLlaV3tV1KzHdpG0jIQ
znXfArRxtIlaBbtnZPoHy5e/N/apx43H0nmW7aHof8e6PZVh3JtGiF9IA0Hvq/Ua
X9mnW9q31iHK5O4F/YRJ4BweM1qUeyUU1fp9LnLEZkAs4v6HkQAovq/SO/lneYVw
/JYSWb+eUhoXEq3lQN1fi328HpqGoL5LccotjZb01hauNmNyksyGBAFLnYntac0l
wslrRi1ILW8OXiHMVcOg0eKpGbuH3bySWvbbCKQ1333nHjLRN+LMTfSZxfqm6Lc/
W5ZZyC3neiBL4WqnjWCTj3AZg2g7G5m8bIOzCj3Vz/41it5z8UQw5vKFis4nvRtY
8KLJ5YftenyE7XNS4DeNezyCJ5Fu48BRQ8Y/E7kZBZDzzRgUK0LfsJjF+u/kIYZY
7RrAhDQIMXu6UCSdgwG1qXQZQoRKfI3Nv8mrVF4D5F8yrqQYJrdcfgR1/PV2Q+Cq
81Wpm3ejIkqlKBX/VcwK2bsUelAMySuqQxe/G1AKnz4E+5rBnkfTfCNnLxK5fPF9
gnz2W/IGh8J/NBJitctyUzo39bNao6CD2T+2V/fRjZgrR5dTSAxcQdleoPkJmJC0
2wCgK42F6azjv/TkVgJJqIknoAjJt+b5BMZhRiWn2J6RsnrZad9RRUZ6HM75jcnZ
YfycCoBw137W04OLqFqaSwT0nbRMjrb9ecKWfUDZ1k5/aCOJkBDVX4bzRQA6tXlU
8AO/+Nbq129OfPVvQADSCRPsAH6hweVApGQSYegoXk37NVjhAVkbiQ3YX2BAauBW
5zFl+bEt7/JkyNQNojhMJIqCk+wuIyPMAMnhAxfHtVQITPNVBTJTAVIWBo619Q/B
DTK3Qww4+mBU2nIRMlsW4htI5pSIhDlPNsBXQbErqMzb5jc4fwEBwdxpBfN33gpJ
qsT6J/r374sJcE519TO8cEaGL/cFpNr1WISJC6JR39JQWz6vap7BWiQ0QbWjKj7K
uhbQj/ewZcKkDG+L2CtiUyZhfxqNr8d+bY8cbjMtDOGkuGwkxX9/GDXPEsMqt/Md
yTITGtCNBWptBGQaGJsPGxgUjGiybWSXCAN4E22rzBEGxFbnUmZiT916aBxhYWJL
K+w4+EbFC5KNo9bDOllW/zneD3vhQkO034LxhB2Oo2zoU9sU9d8teZsC7DTNSSVk
kuP84bY99NW2g2d7WojhhcN438evGBmhOCvHmXszR10A8pyzu5oSYgJl5EPbRekN
ODXDPgY9J21siR8ruqwKibROS8UrcA4i4ADKMmj+EM1A8yvycTAD9NvKBOB5qxvi
uvJ+Dejjm2gtG0gnhsEK2a7KDvijweR4aarWqyG2zT51+ApVsvNgFmO+rxw+2BZM
gF8cIjtPEWEl03m4ObohqIvjpk2OsuW2AuBgzL3W+Yza8mtmJhDEx0COLQ7VIKh2
sUHX51v+BdzjdfGWUrDRhKR++o0t8oTaIacOamurXgNCfoHm/X/BtL2QvGG0lRIb
`pragma protect end_protected
