-- system.vhd

-- Generated using ACDS version 17.0 602

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		clk_clk       : in std_logic := '0'; --    clk.clk
		reset_reset_n : in std_logic := '0'; --  reset.reset_n
		select_export : in std_logic := '0'  -- select.export
	);
end entity system;

architecture rtl of system is
	component system_client0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(14 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(14 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_client0;

	component system_client0_jtag is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_client0_jtag;

	component system_client0_ocm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component system_client0_ocm;

	component system_client1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(14 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(14 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_client1;

	component system_client1_ocm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component system_client1_ocm;

	component system_client2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(14 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(14 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_client2;

	component system_client2_ocm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component system_client2_ocm;

	component system_fifo_client0 is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			wrreset_n                        : in  std_logic                     := 'X';             -- reset_n
			rdclock                          : in  std_logic                     := 'X';             -- clk
			rdreset_n                        : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonmm_read_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read         : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_waitrequest  : out std_logic;                                        -- waitrequest
			rdclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			rdclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			rdclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			rdclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			rdclk_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			rdclk_control_slave_irq          : out std_logic;                                        -- irq
			wrclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			wrclk_control_slave_irq          : out std_logic                                         -- irq
		);
	end component system_fifo_client0;

	component altera_avalon_mailbox is
		generic (
			DWIDTH : integer := 32;
			AWIDTH : integer := 2
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			rst_n                : in  std_logic                     := 'X';             -- reset_n
			avmm_snd_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avmm_snd_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_snd_write       : in  std_logic                     := 'X';             -- write
			avmm_snd_read        : in  std_logic                     := 'X';             -- read
			avmm_snd_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_snd_waitrequest : out std_logic;                                        -- waitrequest
			irq_msg              : out std_logic;                                        -- irq
			avmm_rcv_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avmm_rcv_read        : in  std_logic                     := 'X';             -- read
			avmm_rcv_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_rcv_write       : in  std_logic                     := 'X';             -- write
			avmm_rcv_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq_space            : out std_logic                                         -- irq
		);
	end component altera_avalon_mailbox;

	component system_perfmon is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component system_perfmon;

	component system_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component system_pio;

	component system_pll_100MHz is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component system_pll_100MHz;

	component system_server is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(16 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(16 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_server;

	component system_server_ocm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component system_server_ocm;

	component system_mm_interconnect_0 is
		port (
			pll_100MHz_outclk0_clk                    : in  std_logic                     := 'X';             -- clk
			perfmon_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			server_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			server_data_master_address                : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			server_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			server_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			server_data_master_read                   : in  std_logic                     := 'X';             -- read
			server_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			server_data_master_readdatavalid          : out std_logic;                                        -- readdatavalid
			server_data_master_write                  : in  std_logic                     := 'X';             -- write
			server_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			server_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			server_instruction_master_address         : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			server_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			server_instruction_master_read            : in  std_logic                     := 'X';             -- read
			server_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			server_instruction_master_readdatavalid   : out std_logic;                                        -- readdatavalid
			fifo_client0_out_read                     : out std_logic;                                        -- read
			fifo_client0_out_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client0_out_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			fifo_client0_out_csr_address              : out std_logic_vector(2 downto 0);                     -- address
			fifo_client0_out_csr_write                : out std_logic;                                        -- write
			fifo_client0_out_csr_read                 : out std_logic;                                        -- read
			fifo_client0_out_csr_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client0_out_csr_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_client1_out_read                     : out std_logic;                                        -- read
			fifo_client1_out_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client1_out_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			fifo_client1_out_csr_address              : out std_logic_vector(2 downto 0);                     -- address
			fifo_client1_out_csr_write                : out std_logic;                                        -- write
			fifo_client1_out_csr_read                 : out std_logic;                                        -- read
			fifo_client1_out_csr_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client1_out_csr_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_client2_out_read                     : out std_logic;                                        -- read
			fifo_client2_out_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client2_out_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			fifo_client2_out_csr_address              : out std_logic_vector(2 downto 0);                     -- address
			fifo_client2_out_csr_write                : out std_logic;                                        -- write
			fifo_client2_out_csr_read                 : out std_logic;                                        -- read
			fifo_client2_out_csr_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client2_out_csr_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_client0_avmm_msg_sender_address      : out std_logic_vector(1 downto 0);                     -- address
			mbox_client0_avmm_msg_sender_write        : out std_logic;                                        -- write
			mbox_client0_avmm_msg_sender_read         : out std_logic;                                        -- read
			mbox_client0_avmm_msg_sender_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_client0_avmm_msg_sender_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_client0_avmm_msg_sender_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			mbox_client1_avmm_msg_sender_address      : out std_logic_vector(1 downto 0);                     -- address
			mbox_client1_avmm_msg_sender_write        : out std_logic;                                        -- write
			mbox_client1_avmm_msg_sender_read         : out std_logic;                                        -- read
			mbox_client1_avmm_msg_sender_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_client1_avmm_msg_sender_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_client1_avmm_msg_sender_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			mbox_client2_avmm_msg_sender_address      : out std_logic_vector(1 downto 0);                     -- address
			mbox_client2_avmm_msg_sender_write        : out std_logic;                                        -- write
			mbox_client2_avmm_msg_sender_read         : out std_logic;                                        -- read
			mbox_client2_avmm_msg_sender_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_client2_avmm_msg_sender_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_client2_avmm_msg_sender_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			perfmon_control_slave_address             : out std_logic_vector(3 downto 0);                     -- address
			perfmon_control_slave_write               : out std_logic;                                        -- write
			perfmon_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			perfmon_control_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			perfmon_control_slave_begintransfer       : out std_logic;                                        -- begintransfer
			pio_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			pio_s1_write                              : out std_logic;                                        -- write
			pio_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			pio_s1_chipselect                         : out std_logic;                                        -- chipselect
			server_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			server_debug_mem_slave_write              : out std_logic;                                        -- write
			server_debug_mem_slave_read               : out std_logic;                                        -- read
			server_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			server_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			server_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			server_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			server_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			server_jtag_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			server_jtag_avalon_jtag_slave_write       : out std_logic;                                        -- write
			server_jtag_avalon_jtag_slave_read        : out std_logic;                                        -- read
			server_jtag_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			server_jtag_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			server_jtag_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			server_jtag_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			server_ocm_s1_address                     : out std_logic_vector(12 downto 0);                    -- address
			server_ocm_s1_write                       : out std_logic;                                        -- write
			server_ocm_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			server_ocm_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			server_ocm_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			server_ocm_s1_chipselect                  : out std_logic;                                        -- chipselect
			server_ocm_s1_clken                       : out std_logic                                         -- clken
		);
	end component system_mm_interconnect_0;

	component system_mm_interconnect_1 is
		port (
			pll_100MHz_outclk0_clk                     : in  std_logic                     := 'X';             -- clk
			client0_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			client0_data_master_address                : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			client0_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			client0_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			client0_data_master_read                   : in  std_logic                     := 'X';             -- read
			client0_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			client0_data_master_readdatavalid          : out std_logic;                                        -- readdatavalid
			client0_data_master_write                  : in  std_logic                     := 'X';             -- write
			client0_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			client0_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			client0_instruction_master_address         : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			client0_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			client0_instruction_master_read            : in  std_logic                     := 'X';             -- read
			client0_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			client0_instruction_master_readdatavalid   : out std_logic;                                        -- readdatavalid
			client0_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			client0_debug_mem_slave_write              : out std_logic;                                        -- write
			client0_debug_mem_slave_read               : out std_logic;                                        -- read
			client0_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client0_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			client0_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			client0_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			client0_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			client0_jtag_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			client0_jtag_avalon_jtag_slave_write       : out std_logic;                                        -- write
			client0_jtag_avalon_jtag_slave_read        : out std_logic;                                        -- read
			client0_jtag_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client0_jtag_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			client0_jtag_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			client0_jtag_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			client0_ocm_s1_address                     : out std_logic_vector(10 downto 0);                    -- address
			client0_ocm_s1_write                       : out std_logic;                                        -- write
			client0_ocm_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client0_ocm_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			client0_ocm_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			client0_ocm_s1_chipselect                  : out std_logic;                                        -- chipselect
			client0_ocm_s1_clken                       : out std_logic;                                        -- clken
			fifo_client0_in_write                      : out std_logic;                                        -- write
			fifo_client0_in_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_client0_in_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			fifo_client0_in_csr_address                : out std_logic_vector(2 downto 0);                     -- address
			fifo_client0_in_csr_write                  : out std_logic;                                        -- write
			fifo_client0_in_csr_read                   : out std_logic;                                        -- read
			fifo_client0_in_csr_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client0_in_csr_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_client0_avmm_msg_receiver_address     : out std_logic_vector(1 downto 0);                     -- address
			mbox_client0_avmm_msg_receiver_write       : out std_logic;                                        -- write
			mbox_client0_avmm_msg_receiver_read        : out std_logic;                                        -- read
			mbox_client0_avmm_msg_receiver_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_client0_avmm_msg_receiver_writedata   : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component system_mm_interconnect_1;

	component system_mm_interconnect_2 is
		port (
			pll_100MHz_outclk0_clk                     : in  std_logic                     := 'X';             -- clk
			client1_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			client1_data_master_address                : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			client1_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			client1_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			client1_data_master_read                   : in  std_logic                     := 'X';             -- read
			client1_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			client1_data_master_readdatavalid          : out std_logic;                                        -- readdatavalid
			client1_data_master_write                  : in  std_logic                     := 'X';             -- write
			client1_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			client1_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			client1_instruction_master_address         : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			client1_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			client1_instruction_master_read            : in  std_logic                     := 'X';             -- read
			client1_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			client1_instruction_master_readdatavalid   : out std_logic;                                        -- readdatavalid
			client1_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			client1_debug_mem_slave_write              : out std_logic;                                        -- write
			client1_debug_mem_slave_read               : out std_logic;                                        -- read
			client1_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client1_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			client1_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			client1_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			client1_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			client1_jtag_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			client1_jtag_avalon_jtag_slave_write       : out std_logic;                                        -- write
			client1_jtag_avalon_jtag_slave_read        : out std_logic;                                        -- read
			client1_jtag_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client1_jtag_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			client1_jtag_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			client1_jtag_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			client1_ocm_s1_address                     : out std_logic_vector(10 downto 0);                    -- address
			client1_ocm_s1_write                       : out std_logic;                                        -- write
			client1_ocm_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client1_ocm_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			client1_ocm_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			client1_ocm_s1_chipselect                  : out std_logic;                                        -- chipselect
			client1_ocm_s1_clken                       : out std_logic;                                        -- clken
			fifo_client1_in_write                      : out std_logic;                                        -- write
			fifo_client1_in_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_client1_in_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			fifo_client1_in_csr_address                : out std_logic_vector(2 downto 0);                     -- address
			fifo_client1_in_csr_write                  : out std_logic;                                        -- write
			fifo_client1_in_csr_read                   : out std_logic;                                        -- read
			fifo_client1_in_csr_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client1_in_csr_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_client1_avmm_msg_receiver_address     : out std_logic_vector(1 downto 0);                     -- address
			mbox_client1_avmm_msg_receiver_write       : out std_logic;                                        -- write
			mbox_client1_avmm_msg_receiver_read        : out std_logic;                                        -- read
			mbox_client1_avmm_msg_receiver_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_client1_avmm_msg_receiver_writedata   : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component system_mm_interconnect_2;

	component system_mm_interconnect_3 is
		port (
			pll_100MHz_outclk0_clk                     : in  std_logic                     := 'X';             -- clk
			client2_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			client2_data_master_address                : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			client2_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			client2_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			client2_data_master_read                   : in  std_logic                     := 'X';             -- read
			client2_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			client2_data_master_readdatavalid          : out std_logic;                                        -- readdatavalid
			client2_data_master_write                  : in  std_logic                     := 'X';             -- write
			client2_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			client2_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			client2_instruction_master_address         : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			client2_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			client2_instruction_master_read            : in  std_logic                     := 'X';             -- read
			client2_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			client2_instruction_master_readdatavalid   : out std_logic;                                        -- readdatavalid
			client2_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			client2_debug_mem_slave_write              : out std_logic;                                        -- write
			client2_debug_mem_slave_read               : out std_logic;                                        -- read
			client2_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client2_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			client2_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			client2_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			client2_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			client2_jtag_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			client2_jtag_avalon_jtag_slave_write       : out std_logic;                                        -- write
			client2_jtag_avalon_jtag_slave_read        : out std_logic;                                        -- read
			client2_jtag_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client2_jtag_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			client2_jtag_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			client2_jtag_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			client2_ocm_s1_address                     : out std_logic_vector(10 downto 0);                    -- address
			client2_ocm_s1_write                       : out std_logic;                                        -- write
			client2_ocm_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			client2_ocm_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			client2_ocm_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			client2_ocm_s1_chipselect                  : out std_logic;                                        -- chipselect
			client2_ocm_s1_clken                       : out std_logic;                                        -- clken
			fifo_client2_in_write                      : out std_logic;                                        -- write
			fifo_client2_in_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_client2_in_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			fifo_client2_in_csr_address                : out std_logic_vector(2 downto 0);                     -- address
			fifo_client2_in_csr_write                  : out std_logic;                                        -- write
			fifo_client2_in_csr_read                   : out std_logic;                                        -- read
			fifo_client2_in_csr_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_client2_in_csr_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_client2_avmm_msg_receiver_address     : out std_logic_vector(1 downto 0);                     -- address
			mbox_client2_avmm_msg_receiver_write       : out std_logic;                                        -- write
			mbox_client2_avmm_msg_receiver_read        : out std_logic;                                        -- read
			mbox_client2_avmm_msg_receiver_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_client2_avmm_msg_receiver_writedata   : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component system_mm_interconnect_3;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component system_irq_mapper_003 is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper_003;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			reset_in3      : in  std_logic := 'X'; -- reset_in3.reset
			reset_in4      : in  std_logic := 'X'; -- reset_in4.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_001;

	component system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			reset_in3      : in  std_logic := 'X'; -- reset_in3.reset
			reset_in4      : in  std_logic := 'X'; -- reset_in4.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_002;

	signal pll_100mhz_outclk0_clk                                           : std_logic;                     -- pll_100MHz:outclk_0 -> [client0:clk, client0_jtag:clk, client0_ocm:clk, client1:clk, client1_jtag:clk, client1_ocm:clk, client2:clk, client2_jtag:clk, client2_ocm:clk, fifo_client0:rdclock, fifo_client0:wrclock, fifo_client1:rdclock, fifo_client1:wrclock, fifo_client2:rdclock, fifo_client2:wrclock, irq_mapper:clk, irq_mapper_001:clk, irq_mapper_002:clk, irq_mapper_003:clk, mbox_client0:clk, mbox_client1:clk, mbox_client2:clk, mm_interconnect_0:pll_100MHz_outclk0_clk, mm_interconnect_1:pll_100MHz_outclk0_clk, mm_interconnect_2:pll_100MHz_outclk0_clk, mm_interconnect_3:pll_100MHz_outclk0_clk, perfmon:clk, pio:clk, rst_controller:clk, rst_controller_001:clk, server:clk, server_jtag:clk, server_ocm:clk]
	signal server_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:server_data_master_readdata -> server:d_readdata
	signal server_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:server_data_master_waitrequest -> server:d_waitrequest
	signal server_data_master_debugaccess                                   : std_logic;                     -- server:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:server_data_master_debugaccess
	signal server_data_master_address                                       : std_logic_vector(16 downto 0); -- server:d_address -> mm_interconnect_0:server_data_master_address
	signal server_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- server:d_byteenable -> mm_interconnect_0:server_data_master_byteenable
	signal server_data_master_read                                          : std_logic;                     -- server:d_read -> mm_interconnect_0:server_data_master_read
	signal server_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:server_data_master_readdatavalid -> server:d_readdatavalid
	signal server_data_master_write                                         : std_logic;                     -- server:d_write -> mm_interconnect_0:server_data_master_write
	signal server_data_master_writedata                                     : std_logic_vector(31 downto 0); -- server:d_writedata -> mm_interconnect_0:server_data_master_writedata
	signal server_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:server_instruction_master_readdata -> server:i_readdata
	signal server_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:server_instruction_master_waitrequest -> server:i_waitrequest
	signal server_instruction_master_address                                : std_logic_vector(16 downto 0); -- server:i_address -> mm_interconnect_0:server_instruction_master_address
	signal server_instruction_master_read                                   : std_logic;                     -- server:i_read -> mm_interconnect_0:server_instruction_master_read
	signal server_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:server_instruction_master_readdatavalid -> server:i_readdatavalid
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_chipselect       : std_logic;                     -- mm_interconnect_0:server_jtag_avalon_jtag_slave_chipselect -> server_jtag:av_chipselect
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_readdata         : std_logic_vector(31 downto 0); -- server_jtag:av_readdata -> mm_interconnect_0:server_jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_waitrequest      : std_logic;                     -- server_jtag:av_waitrequest -> mm_interconnect_0:server_jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:server_jtag_avalon_jtag_slave_address -> server_jtag:av_address
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_read             : std_logic;                     -- mm_interconnect_0:server_jtag_avalon_jtag_slave_read -> mm_interconnect_0_server_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_write            : std_logic;                     -- mm_interconnect_0:server_jtag_avalon_jtag_slave_write -> mm_interconnect_0_server_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:server_jtag_avalon_jtag_slave_writedata -> server_jtag:av_writedata
	signal mm_interconnect_0_mbox_client1_avmm_msg_sender_readdata          : std_logic_vector(31 downto 0); -- mbox_client1:avmm_snd_readdata -> mm_interconnect_0:mbox_client1_avmm_msg_sender_readdata
	signal mm_interconnect_0_mbox_client1_avmm_msg_sender_waitrequest       : std_logic;                     -- mbox_client1:avmm_snd_waitrequest -> mm_interconnect_0:mbox_client1_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mbox_client1_avmm_msg_sender_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_client1_avmm_msg_sender_address -> mbox_client1:avmm_snd_address
	signal mm_interconnect_0_mbox_client1_avmm_msg_sender_read              : std_logic;                     -- mm_interconnect_0:mbox_client1_avmm_msg_sender_read -> mbox_client1:avmm_snd_read
	signal mm_interconnect_0_mbox_client1_avmm_msg_sender_write             : std_logic;                     -- mm_interconnect_0:mbox_client1_avmm_msg_sender_write -> mbox_client1:avmm_snd_write
	signal mm_interconnect_0_mbox_client1_avmm_msg_sender_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_client1_avmm_msg_sender_writedata -> mbox_client1:avmm_snd_writedata
	signal mm_interconnect_0_mbox_client0_avmm_msg_sender_readdata          : std_logic_vector(31 downto 0); -- mbox_client0:avmm_snd_readdata -> mm_interconnect_0:mbox_client0_avmm_msg_sender_readdata
	signal mm_interconnect_0_mbox_client0_avmm_msg_sender_waitrequest       : std_logic;                     -- mbox_client0:avmm_snd_waitrequest -> mm_interconnect_0:mbox_client0_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mbox_client0_avmm_msg_sender_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_client0_avmm_msg_sender_address -> mbox_client0:avmm_snd_address
	signal mm_interconnect_0_mbox_client0_avmm_msg_sender_read              : std_logic;                     -- mm_interconnect_0:mbox_client0_avmm_msg_sender_read -> mbox_client0:avmm_snd_read
	signal mm_interconnect_0_mbox_client0_avmm_msg_sender_write             : std_logic;                     -- mm_interconnect_0:mbox_client0_avmm_msg_sender_write -> mbox_client0:avmm_snd_write
	signal mm_interconnect_0_mbox_client0_avmm_msg_sender_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_client0_avmm_msg_sender_writedata -> mbox_client0:avmm_snd_writedata
	signal mm_interconnect_0_mbox_client2_avmm_msg_sender_readdata          : std_logic_vector(31 downto 0); -- mbox_client2:avmm_snd_readdata -> mm_interconnect_0:mbox_client2_avmm_msg_sender_readdata
	signal mm_interconnect_0_mbox_client2_avmm_msg_sender_waitrequest       : std_logic;                     -- mbox_client2:avmm_snd_waitrequest -> mm_interconnect_0:mbox_client2_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mbox_client2_avmm_msg_sender_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_client2_avmm_msg_sender_address -> mbox_client2:avmm_snd_address
	signal mm_interconnect_0_mbox_client2_avmm_msg_sender_read              : std_logic;                     -- mm_interconnect_0:mbox_client2_avmm_msg_sender_read -> mbox_client2:avmm_snd_read
	signal mm_interconnect_0_mbox_client2_avmm_msg_sender_write             : std_logic;                     -- mm_interconnect_0:mbox_client2_avmm_msg_sender_write -> mbox_client2:avmm_snd_write
	signal mm_interconnect_0_mbox_client2_avmm_msg_sender_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_client2_avmm_msg_sender_writedata -> mbox_client2:avmm_snd_writedata
	signal mm_interconnect_0_perfmon_control_slave_readdata                 : std_logic_vector(31 downto 0); -- perfmon:readdata -> mm_interconnect_0:perfmon_control_slave_readdata
	signal mm_interconnect_0_perfmon_control_slave_address                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:perfmon_control_slave_address -> perfmon:address
	signal mm_interconnect_0_perfmon_control_slave_begintransfer            : std_logic;                     -- mm_interconnect_0:perfmon_control_slave_begintransfer -> perfmon:begintransfer
	signal mm_interconnect_0_perfmon_control_slave_write                    : std_logic;                     -- mm_interconnect_0:perfmon_control_slave_write -> perfmon:write
	signal mm_interconnect_0_perfmon_control_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:perfmon_control_slave_writedata -> perfmon:writedata
	signal mm_interconnect_0_server_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- server:debug_mem_slave_readdata -> mm_interconnect_0:server_debug_mem_slave_readdata
	signal mm_interconnect_0_server_debug_mem_slave_waitrequest             : std_logic;                     -- server:debug_mem_slave_waitrequest -> mm_interconnect_0:server_debug_mem_slave_waitrequest
	signal mm_interconnect_0_server_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:server_debug_mem_slave_debugaccess -> server:debug_mem_slave_debugaccess
	signal mm_interconnect_0_server_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:server_debug_mem_slave_address -> server:debug_mem_slave_address
	signal mm_interconnect_0_server_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:server_debug_mem_slave_read -> server:debug_mem_slave_read
	signal mm_interconnect_0_server_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:server_debug_mem_slave_byteenable -> server:debug_mem_slave_byteenable
	signal mm_interconnect_0_server_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:server_debug_mem_slave_write -> server:debug_mem_slave_write
	signal mm_interconnect_0_server_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:server_debug_mem_slave_writedata -> server:debug_mem_slave_writedata
	signal mm_interconnect_0_fifo_client0_out_readdata                      : std_logic_vector(31 downto 0); -- fifo_client0:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_client0_out_readdata
	signal mm_interconnect_0_fifo_client0_out_waitrequest                   : std_logic;                     -- fifo_client0:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_client0_out_waitrequest
	signal mm_interconnect_0_fifo_client0_out_read                          : std_logic;                     -- mm_interconnect_0:fifo_client0_out_read -> fifo_client0:avalonmm_read_slave_read
	signal mm_interconnect_0_fifo_client1_out_readdata                      : std_logic_vector(31 downto 0); -- fifo_client1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_client1_out_readdata
	signal mm_interconnect_0_fifo_client1_out_waitrequest                   : std_logic;                     -- fifo_client1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_client1_out_waitrequest
	signal mm_interconnect_0_fifo_client1_out_read                          : std_logic;                     -- mm_interconnect_0:fifo_client1_out_read -> fifo_client1:avalonmm_read_slave_read
	signal mm_interconnect_0_fifo_client2_out_readdata                      : std_logic_vector(31 downto 0); -- fifo_client2:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_client2_out_readdata
	signal mm_interconnect_0_fifo_client2_out_waitrequest                   : std_logic;                     -- fifo_client2:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_client2_out_waitrequest
	signal mm_interconnect_0_fifo_client2_out_read                          : std_logic;                     -- mm_interconnect_0:fifo_client2_out_read -> fifo_client2:avalonmm_read_slave_read
	signal mm_interconnect_0_fifo_client0_out_csr_readdata                  : std_logic_vector(31 downto 0); -- fifo_client0:rdclk_control_slave_readdata -> mm_interconnect_0:fifo_client0_out_csr_readdata
	signal mm_interconnect_0_fifo_client0_out_csr_address                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:fifo_client0_out_csr_address -> fifo_client0:rdclk_control_slave_address
	signal mm_interconnect_0_fifo_client0_out_csr_read                      : std_logic;                     -- mm_interconnect_0:fifo_client0_out_csr_read -> fifo_client0:rdclk_control_slave_read
	signal mm_interconnect_0_fifo_client0_out_csr_write                     : std_logic;                     -- mm_interconnect_0:fifo_client0_out_csr_write -> fifo_client0:rdclk_control_slave_write
	signal mm_interconnect_0_fifo_client0_out_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:fifo_client0_out_csr_writedata -> fifo_client0:rdclk_control_slave_writedata
	signal mm_interconnect_0_fifo_client1_out_csr_readdata                  : std_logic_vector(31 downto 0); -- fifo_client1:rdclk_control_slave_readdata -> mm_interconnect_0:fifo_client1_out_csr_readdata
	signal mm_interconnect_0_fifo_client1_out_csr_address                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:fifo_client1_out_csr_address -> fifo_client1:rdclk_control_slave_address
	signal mm_interconnect_0_fifo_client1_out_csr_read                      : std_logic;                     -- mm_interconnect_0:fifo_client1_out_csr_read -> fifo_client1:rdclk_control_slave_read
	signal mm_interconnect_0_fifo_client1_out_csr_write                     : std_logic;                     -- mm_interconnect_0:fifo_client1_out_csr_write -> fifo_client1:rdclk_control_slave_write
	signal mm_interconnect_0_fifo_client1_out_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:fifo_client1_out_csr_writedata -> fifo_client1:rdclk_control_slave_writedata
	signal mm_interconnect_0_fifo_client2_out_csr_readdata                  : std_logic_vector(31 downto 0); -- fifo_client2:rdclk_control_slave_readdata -> mm_interconnect_0:fifo_client2_out_csr_readdata
	signal mm_interconnect_0_fifo_client2_out_csr_address                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:fifo_client2_out_csr_address -> fifo_client2:rdclk_control_slave_address
	signal mm_interconnect_0_fifo_client2_out_csr_read                      : std_logic;                     -- mm_interconnect_0:fifo_client2_out_csr_read -> fifo_client2:rdclk_control_slave_read
	signal mm_interconnect_0_fifo_client2_out_csr_write                     : std_logic;                     -- mm_interconnect_0:fifo_client2_out_csr_write -> fifo_client2:rdclk_control_slave_write
	signal mm_interconnect_0_fifo_client2_out_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:fifo_client2_out_csr_writedata -> fifo_client2:rdclk_control_slave_writedata
	signal mm_interconnect_0_server_ocm_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:server_ocm_s1_chipselect -> server_ocm:chipselect
	signal mm_interconnect_0_server_ocm_s1_readdata                         : std_logic_vector(31 downto 0); -- server_ocm:readdata -> mm_interconnect_0:server_ocm_s1_readdata
	signal mm_interconnect_0_server_ocm_s1_address                          : std_logic_vector(12 downto 0); -- mm_interconnect_0:server_ocm_s1_address -> server_ocm:address
	signal mm_interconnect_0_server_ocm_s1_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:server_ocm_s1_byteenable -> server_ocm:byteenable
	signal mm_interconnect_0_server_ocm_s1_write                            : std_logic;                     -- mm_interconnect_0:server_ocm_s1_write -> server_ocm:write
	signal mm_interconnect_0_server_ocm_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:server_ocm_s1_writedata -> server_ocm:writedata
	signal mm_interconnect_0_server_ocm_s1_clken                            : std_logic;                     -- mm_interconnect_0:server_ocm_s1_clken -> server_ocm:clken
	signal mm_interconnect_0_pio_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:pio_s1_chipselect -> pio:chipselect
	signal mm_interconnect_0_pio_s1_readdata                                : std_logic_vector(31 downto 0); -- pio:readdata -> mm_interconnect_0:pio_s1_readdata
	signal mm_interconnect_0_pio_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_s1_address -> pio:address
	signal mm_interconnect_0_pio_s1_write                                   : std_logic;                     -- mm_interconnect_0:pio_s1_write -> mm_interconnect_0_pio_s1_write:in
	signal mm_interconnect_0_pio_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_s1_writedata -> pio:writedata
	signal client0_data_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_1:client0_data_master_readdata -> client0:d_readdata
	signal client0_data_master_waitrequest                                  : std_logic;                     -- mm_interconnect_1:client0_data_master_waitrequest -> client0:d_waitrequest
	signal client0_data_master_debugaccess                                  : std_logic;                     -- client0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:client0_data_master_debugaccess
	signal client0_data_master_address                                      : std_logic_vector(14 downto 0); -- client0:d_address -> mm_interconnect_1:client0_data_master_address
	signal client0_data_master_byteenable                                   : std_logic_vector(3 downto 0);  -- client0:d_byteenable -> mm_interconnect_1:client0_data_master_byteenable
	signal client0_data_master_read                                         : std_logic;                     -- client0:d_read -> mm_interconnect_1:client0_data_master_read
	signal client0_data_master_readdatavalid                                : std_logic;                     -- mm_interconnect_1:client0_data_master_readdatavalid -> client0:d_readdatavalid
	signal client0_data_master_write                                        : std_logic;                     -- client0:d_write -> mm_interconnect_1:client0_data_master_write
	signal client0_data_master_writedata                                    : std_logic_vector(31 downto 0); -- client0:d_writedata -> mm_interconnect_1:client0_data_master_writedata
	signal client0_instruction_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_1:client0_instruction_master_readdata -> client0:i_readdata
	signal client0_instruction_master_waitrequest                           : std_logic;                     -- mm_interconnect_1:client0_instruction_master_waitrequest -> client0:i_waitrequest
	signal client0_instruction_master_address                               : std_logic_vector(14 downto 0); -- client0:i_address -> mm_interconnect_1:client0_instruction_master_address
	signal client0_instruction_master_read                                  : std_logic;                     -- client0:i_read -> mm_interconnect_1:client0_instruction_master_read
	signal client0_instruction_master_readdatavalid                         : std_logic;                     -- mm_interconnect_1:client0_instruction_master_readdatavalid -> client0:i_readdatavalid
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_1:client0_jtag_avalon_jtag_slave_chipselect -> client0_jtag:av_chipselect
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- client0_jtag:av_readdata -> mm_interconnect_1:client0_jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- client0_jtag:av_waitrequest -> mm_interconnect_1:client0_jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_1:client0_jtag_avalon_jtag_slave_address -> client0_jtag:av_address
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_1:client0_jtag_avalon_jtag_slave_read -> mm_interconnect_1_client0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_1:client0_jtag_avalon_jtag_slave_write -> mm_interconnect_1_client0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:client0_jtag_avalon_jtag_slave_writedata -> client0_jtag:av_writedata
	signal mm_interconnect_1_mbox_client0_avmm_msg_receiver_readdata        : std_logic_vector(31 downto 0); -- mbox_client0:avmm_rcv_readdata -> mm_interconnect_1:mbox_client0_avmm_msg_receiver_readdata
	signal mm_interconnect_1_mbox_client0_avmm_msg_receiver_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_1:mbox_client0_avmm_msg_receiver_address -> mbox_client0:avmm_rcv_address
	signal mm_interconnect_1_mbox_client0_avmm_msg_receiver_read            : std_logic;                     -- mm_interconnect_1:mbox_client0_avmm_msg_receiver_read -> mbox_client0:avmm_rcv_read
	signal mm_interconnect_1_mbox_client0_avmm_msg_receiver_write           : std_logic;                     -- mm_interconnect_1:mbox_client0_avmm_msg_receiver_write -> mbox_client0:avmm_rcv_write
	signal mm_interconnect_1_mbox_client0_avmm_msg_receiver_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:mbox_client0_avmm_msg_receiver_writedata -> mbox_client0:avmm_rcv_writedata
	signal mm_interconnect_1_client0_debug_mem_slave_readdata               : std_logic_vector(31 downto 0); -- client0:debug_mem_slave_readdata -> mm_interconnect_1:client0_debug_mem_slave_readdata
	signal mm_interconnect_1_client0_debug_mem_slave_waitrequest            : std_logic;                     -- client0:debug_mem_slave_waitrequest -> mm_interconnect_1:client0_debug_mem_slave_waitrequest
	signal mm_interconnect_1_client0_debug_mem_slave_debugaccess            : std_logic;                     -- mm_interconnect_1:client0_debug_mem_slave_debugaccess -> client0:debug_mem_slave_debugaccess
	signal mm_interconnect_1_client0_debug_mem_slave_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_1:client0_debug_mem_slave_address -> client0:debug_mem_slave_address
	signal mm_interconnect_1_client0_debug_mem_slave_read                   : std_logic;                     -- mm_interconnect_1:client0_debug_mem_slave_read -> client0:debug_mem_slave_read
	signal mm_interconnect_1_client0_debug_mem_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_1:client0_debug_mem_slave_byteenable -> client0:debug_mem_slave_byteenable
	signal mm_interconnect_1_client0_debug_mem_slave_write                  : std_logic;                     -- mm_interconnect_1:client0_debug_mem_slave_write -> client0:debug_mem_slave_write
	signal mm_interconnect_1_client0_debug_mem_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_1:client0_debug_mem_slave_writedata -> client0:debug_mem_slave_writedata
	signal mm_interconnect_1_fifo_client0_in_waitrequest                    : std_logic;                     -- fifo_client0:avalonmm_write_slave_waitrequest -> mm_interconnect_1:fifo_client0_in_waitrequest
	signal mm_interconnect_1_fifo_client0_in_write                          : std_logic;                     -- mm_interconnect_1:fifo_client0_in_write -> fifo_client0:avalonmm_write_slave_write
	signal mm_interconnect_1_fifo_client0_in_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:fifo_client0_in_writedata -> fifo_client0:avalonmm_write_slave_writedata
	signal mm_interconnect_1_fifo_client0_in_csr_readdata                   : std_logic_vector(31 downto 0); -- fifo_client0:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_client0_in_csr_readdata
	signal mm_interconnect_1_fifo_client0_in_csr_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_1:fifo_client0_in_csr_address -> fifo_client0:wrclk_control_slave_address
	signal mm_interconnect_1_fifo_client0_in_csr_read                       : std_logic;                     -- mm_interconnect_1:fifo_client0_in_csr_read -> fifo_client0:wrclk_control_slave_read
	signal mm_interconnect_1_fifo_client0_in_csr_write                      : std_logic;                     -- mm_interconnect_1:fifo_client0_in_csr_write -> fifo_client0:wrclk_control_slave_write
	signal mm_interconnect_1_fifo_client0_in_csr_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_1:fifo_client0_in_csr_writedata -> fifo_client0:wrclk_control_slave_writedata
	signal mm_interconnect_1_client0_ocm_s1_chipselect                      : std_logic;                     -- mm_interconnect_1:client0_ocm_s1_chipselect -> client0_ocm:chipselect
	signal mm_interconnect_1_client0_ocm_s1_readdata                        : std_logic_vector(31 downto 0); -- client0_ocm:readdata -> mm_interconnect_1:client0_ocm_s1_readdata
	signal mm_interconnect_1_client0_ocm_s1_address                         : std_logic_vector(10 downto 0); -- mm_interconnect_1:client0_ocm_s1_address -> client0_ocm:address
	signal mm_interconnect_1_client0_ocm_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_1:client0_ocm_s1_byteenable -> client0_ocm:byteenable
	signal mm_interconnect_1_client0_ocm_s1_write                           : std_logic;                     -- mm_interconnect_1:client0_ocm_s1_write -> client0_ocm:write
	signal mm_interconnect_1_client0_ocm_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:client0_ocm_s1_writedata -> client0_ocm:writedata
	signal mm_interconnect_1_client0_ocm_s1_clken                           : std_logic;                     -- mm_interconnect_1:client0_ocm_s1_clken -> client0_ocm:clken
	signal client1_data_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_2:client1_data_master_readdata -> client1:d_readdata
	signal client1_data_master_waitrequest                                  : std_logic;                     -- mm_interconnect_2:client1_data_master_waitrequest -> client1:d_waitrequest
	signal client1_data_master_debugaccess                                  : std_logic;                     -- client1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_2:client1_data_master_debugaccess
	signal client1_data_master_address                                      : std_logic_vector(14 downto 0); -- client1:d_address -> mm_interconnect_2:client1_data_master_address
	signal client1_data_master_byteenable                                   : std_logic_vector(3 downto 0);  -- client1:d_byteenable -> mm_interconnect_2:client1_data_master_byteenable
	signal client1_data_master_read                                         : std_logic;                     -- client1:d_read -> mm_interconnect_2:client1_data_master_read
	signal client1_data_master_readdatavalid                                : std_logic;                     -- mm_interconnect_2:client1_data_master_readdatavalid -> client1:d_readdatavalid
	signal client1_data_master_write                                        : std_logic;                     -- client1:d_write -> mm_interconnect_2:client1_data_master_write
	signal client1_data_master_writedata                                    : std_logic_vector(31 downto 0); -- client1:d_writedata -> mm_interconnect_2:client1_data_master_writedata
	signal client1_instruction_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_2:client1_instruction_master_readdata -> client1:i_readdata
	signal client1_instruction_master_waitrequest                           : std_logic;                     -- mm_interconnect_2:client1_instruction_master_waitrequest -> client1:i_waitrequest
	signal client1_instruction_master_address                               : std_logic_vector(14 downto 0); -- client1:i_address -> mm_interconnect_2:client1_instruction_master_address
	signal client1_instruction_master_read                                  : std_logic;                     -- client1:i_read -> mm_interconnect_2:client1_instruction_master_read
	signal client1_instruction_master_readdatavalid                         : std_logic;                     -- mm_interconnect_2:client1_instruction_master_readdatavalid -> client1:i_readdatavalid
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_2:client1_jtag_avalon_jtag_slave_chipselect -> client1_jtag:av_chipselect
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- client1_jtag:av_readdata -> mm_interconnect_2:client1_jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- client1_jtag:av_waitrequest -> mm_interconnect_2:client1_jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_2:client1_jtag_avalon_jtag_slave_address -> client1_jtag:av_address
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_2:client1_jtag_avalon_jtag_slave_read -> mm_interconnect_2_client1_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_2:client1_jtag_avalon_jtag_slave_write -> mm_interconnect_2_client1_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_2:client1_jtag_avalon_jtag_slave_writedata -> client1_jtag:av_writedata
	signal mm_interconnect_2_mbox_client1_avmm_msg_receiver_readdata        : std_logic_vector(31 downto 0); -- mbox_client1:avmm_rcv_readdata -> mm_interconnect_2:mbox_client1_avmm_msg_receiver_readdata
	signal mm_interconnect_2_mbox_client1_avmm_msg_receiver_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_2:mbox_client1_avmm_msg_receiver_address -> mbox_client1:avmm_rcv_address
	signal mm_interconnect_2_mbox_client1_avmm_msg_receiver_read            : std_logic;                     -- mm_interconnect_2:mbox_client1_avmm_msg_receiver_read -> mbox_client1:avmm_rcv_read
	signal mm_interconnect_2_mbox_client1_avmm_msg_receiver_write           : std_logic;                     -- mm_interconnect_2:mbox_client1_avmm_msg_receiver_write -> mbox_client1:avmm_rcv_write
	signal mm_interconnect_2_mbox_client1_avmm_msg_receiver_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_2:mbox_client1_avmm_msg_receiver_writedata -> mbox_client1:avmm_rcv_writedata
	signal mm_interconnect_2_client1_debug_mem_slave_readdata               : std_logic_vector(31 downto 0); -- client1:debug_mem_slave_readdata -> mm_interconnect_2:client1_debug_mem_slave_readdata
	signal mm_interconnect_2_client1_debug_mem_slave_waitrequest            : std_logic;                     -- client1:debug_mem_slave_waitrequest -> mm_interconnect_2:client1_debug_mem_slave_waitrequest
	signal mm_interconnect_2_client1_debug_mem_slave_debugaccess            : std_logic;                     -- mm_interconnect_2:client1_debug_mem_slave_debugaccess -> client1:debug_mem_slave_debugaccess
	signal mm_interconnect_2_client1_debug_mem_slave_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_2:client1_debug_mem_slave_address -> client1:debug_mem_slave_address
	signal mm_interconnect_2_client1_debug_mem_slave_read                   : std_logic;                     -- mm_interconnect_2:client1_debug_mem_slave_read -> client1:debug_mem_slave_read
	signal mm_interconnect_2_client1_debug_mem_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_2:client1_debug_mem_slave_byteenable -> client1:debug_mem_slave_byteenable
	signal mm_interconnect_2_client1_debug_mem_slave_write                  : std_logic;                     -- mm_interconnect_2:client1_debug_mem_slave_write -> client1:debug_mem_slave_write
	signal mm_interconnect_2_client1_debug_mem_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_2:client1_debug_mem_slave_writedata -> client1:debug_mem_slave_writedata
	signal mm_interconnect_2_fifo_client1_in_waitrequest                    : std_logic;                     -- fifo_client1:avalonmm_write_slave_waitrequest -> mm_interconnect_2:fifo_client1_in_waitrequest
	signal mm_interconnect_2_fifo_client1_in_write                          : std_logic;                     -- mm_interconnect_2:fifo_client1_in_write -> fifo_client1:avalonmm_write_slave_write
	signal mm_interconnect_2_fifo_client1_in_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_2:fifo_client1_in_writedata -> fifo_client1:avalonmm_write_slave_writedata
	signal mm_interconnect_2_fifo_client1_in_csr_readdata                   : std_logic_vector(31 downto 0); -- fifo_client1:wrclk_control_slave_readdata -> mm_interconnect_2:fifo_client1_in_csr_readdata
	signal mm_interconnect_2_fifo_client1_in_csr_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_2:fifo_client1_in_csr_address -> fifo_client1:wrclk_control_slave_address
	signal mm_interconnect_2_fifo_client1_in_csr_read                       : std_logic;                     -- mm_interconnect_2:fifo_client1_in_csr_read -> fifo_client1:wrclk_control_slave_read
	signal mm_interconnect_2_fifo_client1_in_csr_write                      : std_logic;                     -- mm_interconnect_2:fifo_client1_in_csr_write -> fifo_client1:wrclk_control_slave_write
	signal mm_interconnect_2_fifo_client1_in_csr_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_2:fifo_client1_in_csr_writedata -> fifo_client1:wrclk_control_slave_writedata
	signal mm_interconnect_2_client1_ocm_s1_chipselect                      : std_logic;                     -- mm_interconnect_2:client1_ocm_s1_chipselect -> client1_ocm:chipselect
	signal mm_interconnect_2_client1_ocm_s1_readdata                        : std_logic_vector(31 downto 0); -- client1_ocm:readdata -> mm_interconnect_2:client1_ocm_s1_readdata
	signal mm_interconnect_2_client1_ocm_s1_address                         : std_logic_vector(10 downto 0); -- mm_interconnect_2:client1_ocm_s1_address -> client1_ocm:address
	signal mm_interconnect_2_client1_ocm_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_2:client1_ocm_s1_byteenable -> client1_ocm:byteenable
	signal mm_interconnect_2_client1_ocm_s1_write                           : std_logic;                     -- mm_interconnect_2:client1_ocm_s1_write -> client1_ocm:write
	signal mm_interconnect_2_client1_ocm_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_2:client1_ocm_s1_writedata -> client1_ocm:writedata
	signal mm_interconnect_2_client1_ocm_s1_clken                           : std_logic;                     -- mm_interconnect_2:client1_ocm_s1_clken -> client1_ocm:clken
	signal client2_data_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_3:client2_data_master_readdata -> client2:d_readdata
	signal client2_data_master_waitrequest                                  : std_logic;                     -- mm_interconnect_3:client2_data_master_waitrequest -> client2:d_waitrequest
	signal client2_data_master_debugaccess                                  : std_logic;                     -- client2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_3:client2_data_master_debugaccess
	signal client2_data_master_address                                      : std_logic_vector(14 downto 0); -- client2:d_address -> mm_interconnect_3:client2_data_master_address
	signal client2_data_master_byteenable                                   : std_logic_vector(3 downto 0);  -- client2:d_byteenable -> mm_interconnect_3:client2_data_master_byteenable
	signal client2_data_master_read                                         : std_logic;                     -- client2:d_read -> mm_interconnect_3:client2_data_master_read
	signal client2_data_master_readdatavalid                                : std_logic;                     -- mm_interconnect_3:client2_data_master_readdatavalid -> client2:d_readdatavalid
	signal client2_data_master_write                                        : std_logic;                     -- client2:d_write -> mm_interconnect_3:client2_data_master_write
	signal client2_data_master_writedata                                    : std_logic_vector(31 downto 0); -- client2:d_writedata -> mm_interconnect_3:client2_data_master_writedata
	signal client2_instruction_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_3:client2_instruction_master_readdata -> client2:i_readdata
	signal client2_instruction_master_waitrequest                           : std_logic;                     -- mm_interconnect_3:client2_instruction_master_waitrequest -> client2:i_waitrequest
	signal client2_instruction_master_address                               : std_logic_vector(14 downto 0); -- client2:i_address -> mm_interconnect_3:client2_instruction_master_address
	signal client2_instruction_master_read                                  : std_logic;                     -- client2:i_read -> mm_interconnect_3:client2_instruction_master_read
	signal client2_instruction_master_readdatavalid                         : std_logic;                     -- mm_interconnect_3:client2_instruction_master_readdatavalid -> client2:i_readdatavalid
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_3:client2_jtag_avalon_jtag_slave_chipselect -> client2_jtag:av_chipselect
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- client2_jtag:av_readdata -> mm_interconnect_3:client2_jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- client2_jtag:av_waitrequest -> mm_interconnect_3:client2_jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_3:client2_jtag_avalon_jtag_slave_address -> client2_jtag:av_address
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_3:client2_jtag_avalon_jtag_slave_read -> mm_interconnect_3_client2_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_3:client2_jtag_avalon_jtag_slave_write -> mm_interconnect_3_client2_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_3:client2_jtag_avalon_jtag_slave_writedata -> client2_jtag:av_writedata
	signal mm_interconnect_3_mbox_client2_avmm_msg_receiver_readdata        : std_logic_vector(31 downto 0); -- mbox_client2:avmm_rcv_readdata -> mm_interconnect_3:mbox_client2_avmm_msg_receiver_readdata
	signal mm_interconnect_3_mbox_client2_avmm_msg_receiver_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_3:mbox_client2_avmm_msg_receiver_address -> mbox_client2:avmm_rcv_address
	signal mm_interconnect_3_mbox_client2_avmm_msg_receiver_read            : std_logic;                     -- mm_interconnect_3:mbox_client2_avmm_msg_receiver_read -> mbox_client2:avmm_rcv_read
	signal mm_interconnect_3_mbox_client2_avmm_msg_receiver_write           : std_logic;                     -- mm_interconnect_3:mbox_client2_avmm_msg_receiver_write -> mbox_client2:avmm_rcv_write
	signal mm_interconnect_3_mbox_client2_avmm_msg_receiver_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_3:mbox_client2_avmm_msg_receiver_writedata -> mbox_client2:avmm_rcv_writedata
	signal mm_interconnect_3_client2_debug_mem_slave_readdata               : std_logic_vector(31 downto 0); -- client2:debug_mem_slave_readdata -> mm_interconnect_3:client2_debug_mem_slave_readdata
	signal mm_interconnect_3_client2_debug_mem_slave_waitrequest            : std_logic;                     -- client2:debug_mem_slave_waitrequest -> mm_interconnect_3:client2_debug_mem_slave_waitrequest
	signal mm_interconnect_3_client2_debug_mem_slave_debugaccess            : std_logic;                     -- mm_interconnect_3:client2_debug_mem_slave_debugaccess -> client2:debug_mem_slave_debugaccess
	signal mm_interconnect_3_client2_debug_mem_slave_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_3:client2_debug_mem_slave_address -> client2:debug_mem_slave_address
	signal mm_interconnect_3_client2_debug_mem_slave_read                   : std_logic;                     -- mm_interconnect_3:client2_debug_mem_slave_read -> client2:debug_mem_slave_read
	signal mm_interconnect_3_client2_debug_mem_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_3:client2_debug_mem_slave_byteenable -> client2:debug_mem_slave_byteenable
	signal mm_interconnect_3_client2_debug_mem_slave_write                  : std_logic;                     -- mm_interconnect_3:client2_debug_mem_slave_write -> client2:debug_mem_slave_write
	signal mm_interconnect_3_client2_debug_mem_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_3:client2_debug_mem_slave_writedata -> client2:debug_mem_slave_writedata
	signal mm_interconnect_3_fifo_client2_in_waitrequest                    : std_logic;                     -- fifo_client2:avalonmm_write_slave_waitrequest -> mm_interconnect_3:fifo_client2_in_waitrequest
	signal mm_interconnect_3_fifo_client2_in_write                          : std_logic;                     -- mm_interconnect_3:fifo_client2_in_write -> fifo_client2:avalonmm_write_slave_write
	signal mm_interconnect_3_fifo_client2_in_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_3:fifo_client2_in_writedata -> fifo_client2:avalonmm_write_slave_writedata
	signal mm_interconnect_3_fifo_client2_in_csr_readdata                   : std_logic_vector(31 downto 0); -- fifo_client2:wrclk_control_slave_readdata -> mm_interconnect_3:fifo_client2_in_csr_readdata
	signal mm_interconnect_3_fifo_client2_in_csr_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_3:fifo_client2_in_csr_address -> fifo_client2:wrclk_control_slave_address
	signal mm_interconnect_3_fifo_client2_in_csr_read                       : std_logic;                     -- mm_interconnect_3:fifo_client2_in_csr_read -> fifo_client2:wrclk_control_slave_read
	signal mm_interconnect_3_fifo_client2_in_csr_write                      : std_logic;                     -- mm_interconnect_3:fifo_client2_in_csr_write -> fifo_client2:wrclk_control_slave_write
	signal mm_interconnect_3_fifo_client2_in_csr_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_3:fifo_client2_in_csr_writedata -> fifo_client2:wrclk_control_slave_writedata
	signal mm_interconnect_3_client2_ocm_s1_chipselect                      : std_logic;                     -- mm_interconnect_3:client2_ocm_s1_chipselect -> client2_ocm:chipselect
	signal mm_interconnect_3_client2_ocm_s1_readdata                        : std_logic_vector(31 downto 0); -- client2_ocm:readdata -> mm_interconnect_3:client2_ocm_s1_readdata
	signal mm_interconnect_3_client2_ocm_s1_address                         : std_logic_vector(10 downto 0); -- mm_interconnect_3:client2_ocm_s1_address -> client2_ocm:address
	signal mm_interconnect_3_client2_ocm_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_3:client2_ocm_s1_byteenable -> client2_ocm:byteenable
	signal mm_interconnect_3_client2_ocm_s1_write                           : std_logic;                     -- mm_interconnect_3:client2_ocm_s1_write -> client2_ocm:write
	signal mm_interconnect_3_client2_ocm_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_3:client2_ocm_s1_writedata -> client2_ocm:writedata
	signal mm_interconnect_3_client2_ocm_s1_clken                           : std_logic;                     -- mm_interconnect_3:client2_ocm_s1_clken -> client2_ocm:clken
	signal irq_mapper_receiver0_irq                                         : std_logic;                     -- fifo_client0:wrclk_control_slave_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                         : std_logic;                     -- mbox_client0:irq_msg -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                         : std_logic;                     -- client0_jtag:av_irq -> irq_mapper:receiver2_irq
	signal client0_irq_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> client0:irq
	signal irq_mapper_001_receiver0_irq                                     : std_logic;                     -- fifo_client1:wrclk_control_slave_irq -> irq_mapper_001:receiver0_irq
	signal irq_mapper_001_receiver1_irq                                     : std_logic;                     -- mbox_client1:irq_msg -> irq_mapper_001:receiver1_irq
	signal irq_mapper_001_receiver2_irq                                     : std_logic;                     -- client1_jtag:av_irq -> irq_mapper_001:receiver2_irq
	signal client1_irq_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> client1:irq
	signal irq_mapper_002_receiver0_irq                                     : std_logic;                     -- fifo_client2:wrclk_control_slave_irq -> irq_mapper_002:receiver0_irq
	signal irq_mapper_002_receiver1_irq                                     : std_logic;                     -- mbox_client2:irq_msg -> irq_mapper_002:receiver1_irq
	signal irq_mapper_002_receiver2_irq                                     : std_logic;                     -- client2_jtag:av_irq -> irq_mapper_002:receiver2_irq
	signal client2_irq_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper_002:sender_irq -> client2:irq
	signal irq_mapper_003_receiver0_irq                                     : std_logic;                     -- server_jtag:av_irq -> irq_mapper_003:receiver0_irq
	signal irq_mapper_003_receiver1_irq                                     : std_logic;                     -- pio:irq -> irq_mapper_003:receiver1_irq
	signal irq_mapper_003_receiver2_irq                                     : std_logic;                     -- fifo_client0:rdclk_control_slave_irq -> irq_mapper_003:receiver2_irq
	signal irq_mapper_003_receiver3_irq                                     : std_logic;                     -- fifo_client1:rdclk_control_slave_irq -> irq_mapper_003:receiver3_irq
	signal irq_mapper_003_receiver4_irq                                     : std_logic;                     -- fifo_client2:rdclk_control_slave_irq -> irq_mapper_003:receiver4_irq
	signal server_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper_003:sender_irq -> server:irq
	signal rst_controller_reset_out_reset                                   : std_logic;                     -- rst_controller:reset_out -> [client0_ocm:reset, client1_ocm:reset, client2_ocm:reset, irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, mm_interconnect_0:server_reset_reset_bridge_in_reset_reset, mm_interconnect_1:client0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:client1_reset_reset_bridge_in_reset_reset, mm_interconnect_3:client2_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, server_ocm:reset]
	signal rst_controller_reset_out_reset_req                               : std_logic;                     -- rst_controller:reset_req -> [client0:reset_req, client0_ocm:reset_req, client1:reset_req, client1_ocm:reset_req, client2:reset_req, client2_ocm:reset_req, rst_translator:reset_req_in, server:reset_req, server_ocm:reset_req]
	signal client0_debug_reset_request_reset                                : std_logic;                     -- client0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in2]
	signal client1_debug_reset_request_reset                                : std_logic;                     -- client1:debug_reset_request -> [rst_controller:reset_in2, rst_controller_002:reset_in3]
	signal client2_debug_reset_request_reset                                : std_logic;                     -- client2:debug_reset_request -> [rst_controller:reset_in3, rst_controller_002:reset_in4]
	signal server_debug_reset_request_reset                                 : std_logic;                     -- server:debug_reset_request -> [rst_controller:reset_in4, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                               : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:perfmon_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                               : std_logic;                     -- rst_controller_002:reset_out -> pll_100MHz:rst
	signal reset_reset_n_ports_inv                                          : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_read_ports_inv   : std_logic;                     -- mm_interconnect_0_server_jtag_avalon_jtag_slave_read:inv -> server_jtag:av_read_n
	signal mm_interconnect_0_server_jtag_avalon_jtag_slave_write_ports_inv  : std_logic;                     -- mm_interconnect_0_server_jtag_avalon_jtag_slave_write:inv -> server_jtag:av_write_n
	signal mm_interconnect_0_pio_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_pio_s1_write:inv -> pio:write_n
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_1_client0_jtag_avalon_jtag_slave_read:inv -> client0_jtag:av_read_n
	signal mm_interconnect_1_client0_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_1_client0_jtag_avalon_jtag_slave_write:inv -> client0_jtag:av_write_n
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_2_client1_jtag_avalon_jtag_slave_read:inv -> client1_jtag:av_read_n
	signal mm_interconnect_2_client1_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_2_client1_jtag_avalon_jtag_slave_write:inv -> client1_jtag:av_write_n
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_3_client2_jtag_avalon_jtag_slave_read:inv -> client2_jtag:av_read_n
	signal mm_interconnect_3_client2_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_3_client2_jtag_avalon_jtag_slave_write:inv -> client2_jtag:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                         : std_logic;                     -- rst_controller_reset_out_reset:inv -> [client0:reset_n, client0_jtag:rst_n, client1:reset_n, client1_jtag:rst_n, client2:reset_n, client2_jtag:rst_n, fifo_client0:rdreset_n, fifo_client0:wrreset_n, fifo_client1:rdreset_n, fifo_client1:wrreset_n, fifo_client2:rdreset_n, fifo_client2:wrreset_n, mbox_client0:rst_n, mbox_client1:rst_n, mbox_client2:rst_n, pio:reset_n, server:reset_n, server_jtag:rst_n]
	signal rst_controller_001_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> perfmon:reset_n

begin

	client0 : component system_client0
		port map (
			clk                                 => pll_100mhz_outclk0_clk,                                --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,              --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                           => client0_data_master_address,                           --               data_master.address
			d_byteenable                        => client0_data_master_byteenable,                        --                          .byteenable
			d_read                              => client0_data_master_read,                              --                          .read
			d_readdata                          => client0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => client0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => client0_data_master_write,                             --                          .write
			d_writedata                         => client0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => client0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => client0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => client0_instruction_master_address,                    --        instruction_master.address
			i_read                              => client0_instruction_master_read,                       --                          .read
			i_readdata                          => client0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => client0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => client0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => client0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => client0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_1_client0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_1_client0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_1_client0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_1_client0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_1_client0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_1_client0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_1_client0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_1_client0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	client0_jtag : component system_client0_jtag
		port map (
			clk            => pll_100mhz_outclk0_clk,                                           --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                         --             reset.reset_n
			av_chipselect  => mm_interconnect_1_client0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_client0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_client0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_client0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_client0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_client0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_client0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                          --               irq.irq
		);

	client0_ocm : component system_client0_ocm
		port map (
			clk        => pll_100mhz_outclk0_clk,                      --   clk1.clk
			address    => mm_interconnect_1_client0_ocm_s1_address,    --     s1.address
			clken      => mm_interconnect_1_client0_ocm_s1_clken,      --       .clken
			chipselect => mm_interconnect_1_client0_ocm_s1_chipselect, --       .chipselect
			write      => mm_interconnect_1_client0_ocm_s1_write,      --       .write
			readdata   => mm_interconnect_1_client0_ocm_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_1_client0_ocm_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_1_client0_ocm_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze     => '0'                                          -- (terminated)
		);

	client1 : component system_client1
		port map (
			clk                                 => pll_100mhz_outclk0_clk,                                --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,              --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                           => client1_data_master_address,                           --               data_master.address
			d_byteenable                        => client1_data_master_byteenable,                        --                          .byteenable
			d_read                              => client1_data_master_read,                              --                          .read
			d_readdata                          => client1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => client1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => client1_data_master_write,                             --                          .write
			d_writedata                         => client1_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => client1_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => client1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => client1_instruction_master_address,                    --        instruction_master.address
			i_read                              => client1_instruction_master_read,                       --                          .read
			i_readdata                          => client1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => client1_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => client1_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => client1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => client1_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_2_client1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_2_client1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_2_client1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_2_client1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_2_client1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_2_client1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_2_client1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_2_client1_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	client1_jtag : component system_client0_jtag
		port map (
			clk            => pll_100mhz_outclk0_clk,                                           --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                         --             reset.reset_n
			av_chipselect  => mm_interconnect_2_client1_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_2_client1_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_2_client1_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_2_client1_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_2_client1_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_2_client1_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_2_client1_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver2_irq                                      --               irq.irq
		);

	client1_ocm : component system_client1_ocm
		port map (
			clk        => pll_100mhz_outclk0_clk,                      --   clk1.clk
			address    => mm_interconnect_2_client1_ocm_s1_address,    --     s1.address
			clken      => mm_interconnect_2_client1_ocm_s1_clken,      --       .clken
			chipselect => mm_interconnect_2_client1_ocm_s1_chipselect, --       .chipselect
			write      => mm_interconnect_2_client1_ocm_s1_write,      --       .write
			readdata   => mm_interconnect_2_client1_ocm_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_2_client1_ocm_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_2_client1_ocm_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze     => '0'                                          -- (terminated)
		);

	client2 : component system_client2
		port map (
			clk                                 => pll_100mhz_outclk0_clk,                                --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,              --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                           => client2_data_master_address,                           --               data_master.address
			d_byteenable                        => client2_data_master_byteenable,                        --                          .byteenable
			d_read                              => client2_data_master_read,                              --                          .read
			d_readdata                          => client2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => client2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => client2_data_master_write,                             --                          .write
			d_writedata                         => client2_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => client2_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => client2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => client2_instruction_master_address,                    --        instruction_master.address
			i_read                              => client2_instruction_master_read,                       --                          .read
			i_readdata                          => client2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => client2_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => client2_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => client2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => client2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_3_client2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_3_client2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_3_client2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_3_client2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_3_client2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_3_client2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_3_client2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_3_client2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	client2_jtag : component system_client0_jtag
		port map (
			clk            => pll_100mhz_outclk0_clk,                                           --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                         --             reset.reset_n
			av_chipselect  => mm_interconnect_3_client2_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_3_client2_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_3_client2_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_3_client2_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_3_client2_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_3_client2_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_3_client2_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_002_receiver2_irq                                      --               irq.irq
		);

	client2_ocm : component system_client2_ocm
		port map (
			clk        => pll_100mhz_outclk0_clk,                      --   clk1.clk
			address    => mm_interconnect_3_client2_ocm_s1_address,    --     s1.address
			clken      => mm_interconnect_3_client2_ocm_s1_clken,      --       .clken
			chipselect => mm_interconnect_3_client2_ocm_s1_chipselect, --       .chipselect
			write      => mm_interconnect_3_client2_ocm_s1_write,      --       .write
			readdata   => mm_interconnect_3_client2_ocm_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_3_client2_ocm_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_3_client2_ocm_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze     => '0'                                          -- (terminated)
		);

	fifo_client0 : component system_fifo_client0
		port map (
			wrclock                          => pll_100mhz_outclk0_clk,                           --    clk_in.clk
			wrreset_n                        => rst_controller_reset_out_reset_ports_inv,         --  reset_in.reset_n
			rdclock                          => pll_100mhz_outclk0_clk,                           --   clk_out.clk
			rdreset_n                        => rst_controller_reset_out_reset_ports_inv,         -- reset_out.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_1_fifo_client0_in_writedata,      --        in.writedata
			avalonmm_write_slave_write       => mm_interconnect_1_fifo_client0_in_write,          --          .write
			avalonmm_write_slave_waitrequest => mm_interconnect_1_fifo_client0_in_waitrequest,    --          .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_0_fifo_client0_out_readdata,      --       out.readdata
			avalonmm_read_slave_read         => mm_interconnect_0_fifo_client0_out_read,          --          .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_0_fifo_client0_out_waitrequest,   --          .waitrequest
			rdclk_control_slave_address      => mm_interconnect_0_fifo_client0_out_csr_address,   --   out_csr.address
			rdclk_control_slave_read         => mm_interconnect_0_fifo_client0_out_csr_read,      --          .read
			rdclk_control_slave_writedata    => mm_interconnect_0_fifo_client0_out_csr_writedata, --          .writedata
			rdclk_control_slave_write        => mm_interconnect_0_fifo_client0_out_csr_write,     --          .write
			rdclk_control_slave_readdata     => mm_interconnect_0_fifo_client0_out_csr_readdata,  --          .readdata
			rdclk_control_slave_irq          => irq_mapper_003_receiver2_irq,                     --   out_irq.irq
			wrclk_control_slave_address      => mm_interconnect_1_fifo_client0_in_csr_address,    --    in_csr.address
			wrclk_control_slave_read         => mm_interconnect_1_fifo_client0_in_csr_read,       --          .read
			wrclk_control_slave_writedata    => mm_interconnect_1_fifo_client0_in_csr_writedata,  --          .writedata
			wrclk_control_slave_write        => mm_interconnect_1_fifo_client0_in_csr_write,      --          .write
			wrclk_control_slave_readdata     => mm_interconnect_1_fifo_client0_in_csr_readdata,   --          .readdata
			wrclk_control_slave_irq          => irq_mapper_receiver0_irq                          --    in_irq.irq
		);

	fifo_client1 : component system_fifo_client0
		port map (
			wrclock                          => pll_100mhz_outclk0_clk,                           --    clk_in.clk
			wrreset_n                        => rst_controller_reset_out_reset_ports_inv,         --  reset_in.reset_n
			rdclock                          => pll_100mhz_outclk0_clk,                           --   clk_out.clk
			rdreset_n                        => rst_controller_reset_out_reset_ports_inv,         -- reset_out.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_2_fifo_client1_in_writedata,      --        in.writedata
			avalonmm_write_slave_write       => mm_interconnect_2_fifo_client1_in_write,          --          .write
			avalonmm_write_slave_waitrequest => mm_interconnect_2_fifo_client1_in_waitrequest,    --          .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_0_fifo_client1_out_readdata,      --       out.readdata
			avalonmm_read_slave_read         => mm_interconnect_0_fifo_client1_out_read,          --          .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_0_fifo_client1_out_waitrequest,   --          .waitrequest
			rdclk_control_slave_address      => mm_interconnect_0_fifo_client1_out_csr_address,   --   out_csr.address
			rdclk_control_slave_read         => mm_interconnect_0_fifo_client1_out_csr_read,      --          .read
			rdclk_control_slave_writedata    => mm_interconnect_0_fifo_client1_out_csr_writedata, --          .writedata
			rdclk_control_slave_write        => mm_interconnect_0_fifo_client1_out_csr_write,     --          .write
			rdclk_control_slave_readdata     => mm_interconnect_0_fifo_client1_out_csr_readdata,  --          .readdata
			rdclk_control_slave_irq          => irq_mapper_003_receiver3_irq,                     --   out_irq.irq
			wrclk_control_slave_address      => mm_interconnect_2_fifo_client1_in_csr_address,    --    in_csr.address
			wrclk_control_slave_read         => mm_interconnect_2_fifo_client1_in_csr_read,       --          .read
			wrclk_control_slave_writedata    => mm_interconnect_2_fifo_client1_in_csr_writedata,  --          .writedata
			wrclk_control_slave_write        => mm_interconnect_2_fifo_client1_in_csr_write,      --          .write
			wrclk_control_slave_readdata     => mm_interconnect_2_fifo_client1_in_csr_readdata,   --          .readdata
			wrclk_control_slave_irq          => irq_mapper_001_receiver0_irq                      --    in_irq.irq
		);

	fifo_client2 : component system_fifo_client0
		port map (
			wrclock                          => pll_100mhz_outclk0_clk,                           --    clk_in.clk
			wrreset_n                        => rst_controller_reset_out_reset_ports_inv,         --  reset_in.reset_n
			rdclock                          => pll_100mhz_outclk0_clk,                           --   clk_out.clk
			rdreset_n                        => rst_controller_reset_out_reset_ports_inv,         -- reset_out.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_3_fifo_client2_in_writedata,      --        in.writedata
			avalonmm_write_slave_write       => mm_interconnect_3_fifo_client2_in_write,          --          .write
			avalonmm_write_slave_waitrequest => mm_interconnect_3_fifo_client2_in_waitrequest,    --          .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_0_fifo_client2_out_readdata,      --       out.readdata
			avalonmm_read_slave_read         => mm_interconnect_0_fifo_client2_out_read,          --          .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_0_fifo_client2_out_waitrequest,   --          .waitrequest
			rdclk_control_slave_address      => mm_interconnect_0_fifo_client2_out_csr_address,   --   out_csr.address
			rdclk_control_slave_read         => mm_interconnect_0_fifo_client2_out_csr_read,      --          .read
			rdclk_control_slave_writedata    => mm_interconnect_0_fifo_client2_out_csr_writedata, --          .writedata
			rdclk_control_slave_write        => mm_interconnect_0_fifo_client2_out_csr_write,     --          .write
			rdclk_control_slave_readdata     => mm_interconnect_0_fifo_client2_out_csr_readdata,  --          .readdata
			rdclk_control_slave_irq          => irq_mapper_003_receiver4_irq,                     --   out_irq.irq
			wrclk_control_slave_address      => mm_interconnect_3_fifo_client2_in_csr_address,    --    in_csr.address
			wrclk_control_slave_read         => mm_interconnect_3_fifo_client2_in_csr_read,       --          .read
			wrclk_control_slave_writedata    => mm_interconnect_3_fifo_client2_in_csr_writedata,  --          .writedata
			wrclk_control_slave_write        => mm_interconnect_3_fifo_client2_in_csr_write,      --          .write
			wrclk_control_slave_readdata     => mm_interconnect_3_fifo_client2_in_csr_readdata,   --          .readdata
			wrclk_control_slave_irq          => irq_mapper_002_receiver0_irq                      --    in_irq.irq
		);

	mbox_client0 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => pll_100mhz_outclk0_clk,                                     --                   clk.clk
			rst_n                => rst_controller_reset_out_reset_ports_inv,                   --                 rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mbox_client0_avmm_msg_sender_address,     --       avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mbox_client0_avmm_msg_sender_writedata,   --                      .writedata
			avmm_snd_write       => mm_interconnect_0_mbox_client0_avmm_msg_sender_write,       --                      .write
			avmm_snd_read        => mm_interconnect_0_mbox_client0_avmm_msg_sender_read,        --                      .read
			avmm_snd_readdata    => mm_interconnect_0_mbox_client0_avmm_msg_sender_readdata,    --                      .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mbox_client0_avmm_msg_sender_waitrequest, --                      .waitrequest
			irq_msg              => irq_mapper_receiver1_irq,                                   -- interrupt_msg_pending.irq
			avmm_rcv_address     => mm_interconnect_1_mbox_client0_avmm_msg_receiver_address,   --     avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_1_mbox_client0_avmm_msg_receiver_read,      --                      .read
			avmm_rcv_writedata   => mm_interconnect_1_mbox_client0_avmm_msg_receiver_writedata, --                      .writedata
			avmm_rcv_write       => mm_interconnect_1_mbox_client0_avmm_msg_receiver_write,     --                      .write
			avmm_rcv_readdata    => mm_interconnect_1_mbox_client0_avmm_msg_receiver_readdata,  --                      .readdata
			irq_space            => open                                                        --           (terminated)
		);

	mbox_client1 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => pll_100mhz_outclk0_clk,                                     --                   clk.clk
			rst_n                => rst_controller_reset_out_reset_ports_inv,                   --                 rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mbox_client1_avmm_msg_sender_address,     --       avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mbox_client1_avmm_msg_sender_writedata,   --                      .writedata
			avmm_snd_write       => mm_interconnect_0_mbox_client1_avmm_msg_sender_write,       --                      .write
			avmm_snd_read        => mm_interconnect_0_mbox_client1_avmm_msg_sender_read,        --                      .read
			avmm_snd_readdata    => mm_interconnect_0_mbox_client1_avmm_msg_sender_readdata,    --                      .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mbox_client1_avmm_msg_sender_waitrequest, --                      .waitrequest
			irq_msg              => irq_mapper_001_receiver1_irq,                               -- interrupt_msg_pending.irq
			avmm_rcv_address     => mm_interconnect_2_mbox_client1_avmm_msg_receiver_address,   --     avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_2_mbox_client1_avmm_msg_receiver_read,      --                      .read
			avmm_rcv_writedata   => mm_interconnect_2_mbox_client1_avmm_msg_receiver_writedata, --                      .writedata
			avmm_rcv_write       => mm_interconnect_2_mbox_client1_avmm_msg_receiver_write,     --                      .write
			avmm_rcv_readdata    => mm_interconnect_2_mbox_client1_avmm_msg_receiver_readdata,  --                      .readdata
			irq_space            => open                                                        --           (terminated)
		);

	mbox_client2 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => pll_100mhz_outclk0_clk,                                     --                   clk.clk
			rst_n                => rst_controller_reset_out_reset_ports_inv,                   --                 rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mbox_client2_avmm_msg_sender_address,     --       avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mbox_client2_avmm_msg_sender_writedata,   --                      .writedata
			avmm_snd_write       => mm_interconnect_0_mbox_client2_avmm_msg_sender_write,       --                      .write
			avmm_snd_read        => mm_interconnect_0_mbox_client2_avmm_msg_sender_read,        --                      .read
			avmm_snd_readdata    => mm_interconnect_0_mbox_client2_avmm_msg_sender_readdata,    --                      .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mbox_client2_avmm_msg_sender_waitrequest, --                      .waitrequest
			irq_msg              => irq_mapper_002_receiver1_irq,                               -- interrupt_msg_pending.irq
			avmm_rcv_address     => mm_interconnect_3_mbox_client2_avmm_msg_receiver_address,   --     avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_3_mbox_client2_avmm_msg_receiver_read,      --                      .read
			avmm_rcv_writedata   => mm_interconnect_3_mbox_client2_avmm_msg_receiver_writedata, --                      .writedata
			avmm_rcv_write       => mm_interconnect_3_mbox_client2_avmm_msg_receiver_write,     --                      .write
			avmm_rcv_readdata    => mm_interconnect_3_mbox_client2_avmm_msg_receiver_readdata,  --                      .readdata
			irq_space            => open                                                        --           (terminated)
		);

	perfmon : component system_perfmon
		port map (
			clk           => pll_100mhz_outclk0_clk,                                --           clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,          --         reset.reset_n
			address       => mm_interconnect_0_perfmon_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_perfmon_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_perfmon_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_perfmon_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_perfmon_control_slave_writedata      --              .writedata
		);

	pio : component system_pio
		port map (
			clk        => pll_100mhz_outclk0_clk,                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_s1_readdata,        --                    .readdata
			in_port    => select_export,                            -- external_connection.export
			irq        => irq_mapper_003_receiver1_irq              --                 irq.irq
		);

	pll_100mhz : component system_pll_100MHz
		port map (
			refclk   => clk_clk,                            --  refclk.clk
			rst      => rst_controller_002_reset_out_reset, --   reset.reset
			outclk_0 => pll_100mhz_outclk0_clk,             -- outclk0.clk
			locked   => open                                -- (terminated)
		);

	server : component system_server
		port map (
			clk                                 => pll_100mhz_outclk0_clk,                               --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                           => server_data_master_address,                           --               data_master.address
			d_byteenable                        => server_data_master_byteenable,                        --                          .byteenable
			d_read                              => server_data_master_read,                              --                          .read
			d_readdata                          => server_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => server_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => server_data_master_write,                             --                          .write
			d_writedata                         => server_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => server_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => server_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => server_instruction_master_address,                    --        instruction_master.address
			i_read                              => server_instruction_master_read,                       --                          .read
			i_readdata                          => server_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => server_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => server_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => server_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => server_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_server_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_server_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_server_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_server_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_server_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_server_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_server_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_server_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                  -- custom_instruction_master.readra
		);

	server_jtag : component system_client0_jtag
		port map (
			clk            => pll_100mhz_outclk0_clk,                                          --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_server_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_server_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_server_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_server_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_server_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_server_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_server_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_003_receiver0_irq                                     --               irq.irq
		);

	server_ocm : component system_server_ocm
		port map (
			clk        => pll_100mhz_outclk0_clk,                     --   clk1.clk
			address    => mm_interconnect_0_server_ocm_s1_address,    --     s1.address
			clken      => mm_interconnect_0_server_ocm_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_server_ocm_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_server_ocm_s1_write,      --       .write
			readdata   => mm_interconnect_0_server_ocm_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_server_ocm_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_server_ocm_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			pll_100MHz_outclk0_clk                    => pll_100mhz_outclk0_clk,                                      --                  pll_100MHz_outclk0.clk
			perfmon_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                          -- perfmon_reset_reset_bridge_in_reset.reset
			server_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                              --  server_reset_reset_bridge_in_reset.reset
			server_data_master_address                => server_data_master_address,                                  --                  server_data_master.address
			server_data_master_waitrequest            => server_data_master_waitrequest,                              --                                    .waitrequest
			server_data_master_byteenable             => server_data_master_byteenable,                               --                                    .byteenable
			server_data_master_read                   => server_data_master_read,                                     --                                    .read
			server_data_master_readdata               => server_data_master_readdata,                                 --                                    .readdata
			server_data_master_readdatavalid          => server_data_master_readdatavalid,                            --                                    .readdatavalid
			server_data_master_write                  => server_data_master_write,                                    --                                    .write
			server_data_master_writedata              => server_data_master_writedata,                                --                                    .writedata
			server_data_master_debugaccess            => server_data_master_debugaccess,                              --                                    .debugaccess
			server_instruction_master_address         => server_instruction_master_address,                           --           server_instruction_master.address
			server_instruction_master_waitrequest     => server_instruction_master_waitrequest,                       --                                    .waitrequest
			server_instruction_master_read            => server_instruction_master_read,                              --                                    .read
			server_instruction_master_readdata        => server_instruction_master_readdata,                          --                                    .readdata
			server_instruction_master_readdatavalid   => server_instruction_master_readdatavalid,                     --                                    .readdatavalid
			fifo_client0_out_read                     => mm_interconnect_0_fifo_client0_out_read,                     --                    fifo_client0_out.read
			fifo_client0_out_readdata                 => mm_interconnect_0_fifo_client0_out_readdata,                 --                                    .readdata
			fifo_client0_out_waitrequest              => mm_interconnect_0_fifo_client0_out_waitrequest,              --                                    .waitrequest
			fifo_client0_out_csr_address              => mm_interconnect_0_fifo_client0_out_csr_address,              --                fifo_client0_out_csr.address
			fifo_client0_out_csr_write                => mm_interconnect_0_fifo_client0_out_csr_write,                --                                    .write
			fifo_client0_out_csr_read                 => mm_interconnect_0_fifo_client0_out_csr_read,                 --                                    .read
			fifo_client0_out_csr_readdata             => mm_interconnect_0_fifo_client0_out_csr_readdata,             --                                    .readdata
			fifo_client0_out_csr_writedata            => mm_interconnect_0_fifo_client0_out_csr_writedata,            --                                    .writedata
			fifo_client1_out_read                     => mm_interconnect_0_fifo_client1_out_read,                     --                    fifo_client1_out.read
			fifo_client1_out_readdata                 => mm_interconnect_0_fifo_client1_out_readdata,                 --                                    .readdata
			fifo_client1_out_waitrequest              => mm_interconnect_0_fifo_client1_out_waitrequest,              --                                    .waitrequest
			fifo_client1_out_csr_address              => mm_interconnect_0_fifo_client1_out_csr_address,              --                fifo_client1_out_csr.address
			fifo_client1_out_csr_write                => mm_interconnect_0_fifo_client1_out_csr_write,                --                                    .write
			fifo_client1_out_csr_read                 => mm_interconnect_0_fifo_client1_out_csr_read,                 --                                    .read
			fifo_client1_out_csr_readdata             => mm_interconnect_0_fifo_client1_out_csr_readdata,             --                                    .readdata
			fifo_client1_out_csr_writedata            => mm_interconnect_0_fifo_client1_out_csr_writedata,            --                                    .writedata
			fifo_client2_out_read                     => mm_interconnect_0_fifo_client2_out_read,                     --                    fifo_client2_out.read
			fifo_client2_out_readdata                 => mm_interconnect_0_fifo_client2_out_readdata,                 --                                    .readdata
			fifo_client2_out_waitrequest              => mm_interconnect_0_fifo_client2_out_waitrequest,              --                                    .waitrequest
			fifo_client2_out_csr_address              => mm_interconnect_0_fifo_client2_out_csr_address,              --                fifo_client2_out_csr.address
			fifo_client2_out_csr_write                => mm_interconnect_0_fifo_client2_out_csr_write,                --                                    .write
			fifo_client2_out_csr_read                 => mm_interconnect_0_fifo_client2_out_csr_read,                 --                                    .read
			fifo_client2_out_csr_readdata             => mm_interconnect_0_fifo_client2_out_csr_readdata,             --                                    .readdata
			fifo_client2_out_csr_writedata            => mm_interconnect_0_fifo_client2_out_csr_writedata,            --                                    .writedata
			mbox_client0_avmm_msg_sender_address      => mm_interconnect_0_mbox_client0_avmm_msg_sender_address,      --        mbox_client0_avmm_msg_sender.address
			mbox_client0_avmm_msg_sender_write        => mm_interconnect_0_mbox_client0_avmm_msg_sender_write,        --                                    .write
			mbox_client0_avmm_msg_sender_read         => mm_interconnect_0_mbox_client0_avmm_msg_sender_read,         --                                    .read
			mbox_client0_avmm_msg_sender_readdata     => mm_interconnect_0_mbox_client0_avmm_msg_sender_readdata,     --                                    .readdata
			mbox_client0_avmm_msg_sender_writedata    => mm_interconnect_0_mbox_client0_avmm_msg_sender_writedata,    --                                    .writedata
			mbox_client0_avmm_msg_sender_waitrequest  => mm_interconnect_0_mbox_client0_avmm_msg_sender_waitrequest,  --                                    .waitrequest
			mbox_client1_avmm_msg_sender_address      => mm_interconnect_0_mbox_client1_avmm_msg_sender_address,      --        mbox_client1_avmm_msg_sender.address
			mbox_client1_avmm_msg_sender_write        => mm_interconnect_0_mbox_client1_avmm_msg_sender_write,        --                                    .write
			mbox_client1_avmm_msg_sender_read         => mm_interconnect_0_mbox_client1_avmm_msg_sender_read,         --                                    .read
			mbox_client1_avmm_msg_sender_readdata     => mm_interconnect_0_mbox_client1_avmm_msg_sender_readdata,     --                                    .readdata
			mbox_client1_avmm_msg_sender_writedata    => mm_interconnect_0_mbox_client1_avmm_msg_sender_writedata,    --                                    .writedata
			mbox_client1_avmm_msg_sender_waitrequest  => mm_interconnect_0_mbox_client1_avmm_msg_sender_waitrequest,  --                                    .waitrequest
			mbox_client2_avmm_msg_sender_address      => mm_interconnect_0_mbox_client2_avmm_msg_sender_address,      --        mbox_client2_avmm_msg_sender.address
			mbox_client2_avmm_msg_sender_write        => mm_interconnect_0_mbox_client2_avmm_msg_sender_write,        --                                    .write
			mbox_client2_avmm_msg_sender_read         => mm_interconnect_0_mbox_client2_avmm_msg_sender_read,         --                                    .read
			mbox_client2_avmm_msg_sender_readdata     => mm_interconnect_0_mbox_client2_avmm_msg_sender_readdata,     --                                    .readdata
			mbox_client2_avmm_msg_sender_writedata    => mm_interconnect_0_mbox_client2_avmm_msg_sender_writedata,    --                                    .writedata
			mbox_client2_avmm_msg_sender_waitrequest  => mm_interconnect_0_mbox_client2_avmm_msg_sender_waitrequest,  --                                    .waitrequest
			perfmon_control_slave_address             => mm_interconnect_0_perfmon_control_slave_address,             --               perfmon_control_slave.address
			perfmon_control_slave_write               => mm_interconnect_0_perfmon_control_slave_write,               --                                    .write
			perfmon_control_slave_readdata            => mm_interconnect_0_perfmon_control_slave_readdata,            --                                    .readdata
			perfmon_control_slave_writedata           => mm_interconnect_0_perfmon_control_slave_writedata,           --                                    .writedata
			perfmon_control_slave_begintransfer       => mm_interconnect_0_perfmon_control_slave_begintransfer,       --                                    .begintransfer
			pio_s1_address                            => mm_interconnect_0_pio_s1_address,                            --                              pio_s1.address
			pio_s1_write                              => mm_interconnect_0_pio_s1_write,                              --                                    .write
			pio_s1_readdata                           => mm_interconnect_0_pio_s1_readdata,                           --                                    .readdata
			pio_s1_writedata                          => mm_interconnect_0_pio_s1_writedata,                          --                                    .writedata
			pio_s1_chipselect                         => mm_interconnect_0_pio_s1_chipselect,                         --                                    .chipselect
			server_debug_mem_slave_address            => mm_interconnect_0_server_debug_mem_slave_address,            --              server_debug_mem_slave.address
			server_debug_mem_slave_write              => mm_interconnect_0_server_debug_mem_slave_write,              --                                    .write
			server_debug_mem_slave_read               => mm_interconnect_0_server_debug_mem_slave_read,               --                                    .read
			server_debug_mem_slave_readdata           => mm_interconnect_0_server_debug_mem_slave_readdata,           --                                    .readdata
			server_debug_mem_slave_writedata          => mm_interconnect_0_server_debug_mem_slave_writedata,          --                                    .writedata
			server_debug_mem_slave_byteenable         => mm_interconnect_0_server_debug_mem_slave_byteenable,         --                                    .byteenable
			server_debug_mem_slave_waitrequest        => mm_interconnect_0_server_debug_mem_slave_waitrequest,        --                                    .waitrequest
			server_debug_mem_slave_debugaccess        => mm_interconnect_0_server_debug_mem_slave_debugaccess,        --                                    .debugaccess
			server_jtag_avalon_jtag_slave_address     => mm_interconnect_0_server_jtag_avalon_jtag_slave_address,     --       server_jtag_avalon_jtag_slave.address
			server_jtag_avalon_jtag_slave_write       => mm_interconnect_0_server_jtag_avalon_jtag_slave_write,       --                                    .write
			server_jtag_avalon_jtag_slave_read        => mm_interconnect_0_server_jtag_avalon_jtag_slave_read,        --                                    .read
			server_jtag_avalon_jtag_slave_readdata    => mm_interconnect_0_server_jtag_avalon_jtag_slave_readdata,    --                                    .readdata
			server_jtag_avalon_jtag_slave_writedata   => mm_interconnect_0_server_jtag_avalon_jtag_slave_writedata,   --                                    .writedata
			server_jtag_avalon_jtag_slave_waitrequest => mm_interconnect_0_server_jtag_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			server_jtag_avalon_jtag_slave_chipselect  => mm_interconnect_0_server_jtag_avalon_jtag_slave_chipselect,  --                                    .chipselect
			server_ocm_s1_address                     => mm_interconnect_0_server_ocm_s1_address,                     --                       server_ocm_s1.address
			server_ocm_s1_write                       => mm_interconnect_0_server_ocm_s1_write,                       --                                    .write
			server_ocm_s1_readdata                    => mm_interconnect_0_server_ocm_s1_readdata,                    --                                    .readdata
			server_ocm_s1_writedata                   => mm_interconnect_0_server_ocm_s1_writedata,                   --                                    .writedata
			server_ocm_s1_byteenable                  => mm_interconnect_0_server_ocm_s1_byteenable,                  --                                    .byteenable
			server_ocm_s1_chipselect                  => mm_interconnect_0_server_ocm_s1_chipselect,                  --                                    .chipselect
			server_ocm_s1_clken                       => mm_interconnect_0_server_ocm_s1_clken                        --                                    .clken
		);

	mm_interconnect_1 : component system_mm_interconnect_1
		port map (
			pll_100MHz_outclk0_clk                     => pll_100mhz_outclk0_clk,                                       --                  pll_100MHz_outclk0.clk
			client0_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                               -- client0_reset_reset_bridge_in_reset.reset
			client0_data_master_address                => client0_data_master_address,                                  --                 client0_data_master.address
			client0_data_master_waitrequest            => client0_data_master_waitrequest,                              --                                    .waitrequest
			client0_data_master_byteenable             => client0_data_master_byteenable,                               --                                    .byteenable
			client0_data_master_read                   => client0_data_master_read,                                     --                                    .read
			client0_data_master_readdata               => client0_data_master_readdata,                                 --                                    .readdata
			client0_data_master_readdatavalid          => client0_data_master_readdatavalid,                            --                                    .readdatavalid
			client0_data_master_write                  => client0_data_master_write,                                    --                                    .write
			client0_data_master_writedata              => client0_data_master_writedata,                                --                                    .writedata
			client0_data_master_debugaccess            => client0_data_master_debugaccess,                              --                                    .debugaccess
			client0_instruction_master_address         => client0_instruction_master_address,                           --          client0_instruction_master.address
			client0_instruction_master_waitrequest     => client0_instruction_master_waitrequest,                       --                                    .waitrequest
			client0_instruction_master_read            => client0_instruction_master_read,                              --                                    .read
			client0_instruction_master_readdata        => client0_instruction_master_readdata,                          --                                    .readdata
			client0_instruction_master_readdatavalid   => client0_instruction_master_readdatavalid,                     --                                    .readdatavalid
			client0_debug_mem_slave_address            => mm_interconnect_1_client0_debug_mem_slave_address,            --             client0_debug_mem_slave.address
			client0_debug_mem_slave_write              => mm_interconnect_1_client0_debug_mem_slave_write,              --                                    .write
			client0_debug_mem_slave_read               => mm_interconnect_1_client0_debug_mem_slave_read,               --                                    .read
			client0_debug_mem_slave_readdata           => mm_interconnect_1_client0_debug_mem_slave_readdata,           --                                    .readdata
			client0_debug_mem_slave_writedata          => mm_interconnect_1_client0_debug_mem_slave_writedata,          --                                    .writedata
			client0_debug_mem_slave_byteenable         => mm_interconnect_1_client0_debug_mem_slave_byteenable,         --                                    .byteenable
			client0_debug_mem_slave_waitrequest        => mm_interconnect_1_client0_debug_mem_slave_waitrequest,        --                                    .waitrequest
			client0_debug_mem_slave_debugaccess        => mm_interconnect_1_client0_debug_mem_slave_debugaccess,        --                                    .debugaccess
			client0_jtag_avalon_jtag_slave_address     => mm_interconnect_1_client0_jtag_avalon_jtag_slave_address,     --      client0_jtag_avalon_jtag_slave.address
			client0_jtag_avalon_jtag_slave_write       => mm_interconnect_1_client0_jtag_avalon_jtag_slave_write,       --                                    .write
			client0_jtag_avalon_jtag_slave_read        => mm_interconnect_1_client0_jtag_avalon_jtag_slave_read,        --                                    .read
			client0_jtag_avalon_jtag_slave_readdata    => mm_interconnect_1_client0_jtag_avalon_jtag_slave_readdata,    --                                    .readdata
			client0_jtag_avalon_jtag_slave_writedata   => mm_interconnect_1_client0_jtag_avalon_jtag_slave_writedata,   --                                    .writedata
			client0_jtag_avalon_jtag_slave_waitrequest => mm_interconnect_1_client0_jtag_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			client0_jtag_avalon_jtag_slave_chipselect  => mm_interconnect_1_client0_jtag_avalon_jtag_slave_chipselect,  --                                    .chipselect
			client0_ocm_s1_address                     => mm_interconnect_1_client0_ocm_s1_address,                     --                      client0_ocm_s1.address
			client0_ocm_s1_write                       => mm_interconnect_1_client0_ocm_s1_write,                       --                                    .write
			client0_ocm_s1_readdata                    => mm_interconnect_1_client0_ocm_s1_readdata,                    --                                    .readdata
			client0_ocm_s1_writedata                   => mm_interconnect_1_client0_ocm_s1_writedata,                   --                                    .writedata
			client0_ocm_s1_byteenable                  => mm_interconnect_1_client0_ocm_s1_byteenable,                  --                                    .byteenable
			client0_ocm_s1_chipselect                  => mm_interconnect_1_client0_ocm_s1_chipselect,                  --                                    .chipselect
			client0_ocm_s1_clken                       => mm_interconnect_1_client0_ocm_s1_clken,                       --                                    .clken
			fifo_client0_in_write                      => mm_interconnect_1_fifo_client0_in_write,                      --                     fifo_client0_in.write
			fifo_client0_in_writedata                  => mm_interconnect_1_fifo_client0_in_writedata,                  --                                    .writedata
			fifo_client0_in_waitrequest                => mm_interconnect_1_fifo_client0_in_waitrequest,                --                                    .waitrequest
			fifo_client0_in_csr_address                => mm_interconnect_1_fifo_client0_in_csr_address,                --                 fifo_client0_in_csr.address
			fifo_client0_in_csr_write                  => mm_interconnect_1_fifo_client0_in_csr_write,                  --                                    .write
			fifo_client0_in_csr_read                   => mm_interconnect_1_fifo_client0_in_csr_read,                   --                                    .read
			fifo_client0_in_csr_readdata               => mm_interconnect_1_fifo_client0_in_csr_readdata,               --                                    .readdata
			fifo_client0_in_csr_writedata              => mm_interconnect_1_fifo_client0_in_csr_writedata,              --                                    .writedata
			mbox_client0_avmm_msg_receiver_address     => mm_interconnect_1_mbox_client0_avmm_msg_receiver_address,     --      mbox_client0_avmm_msg_receiver.address
			mbox_client0_avmm_msg_receiver_write       => mm_interconnect_1_mbox_client0_avmm_msg_receiver_write,       --                                    .write
			mbox_client0_avmm_msg_receiver_read        => mm_interconnect_1_mbox_client0_avmm_msg_receiver_read,        --                                    .read
			mbox_client0_avmm_msg_receiver_readdata    => mm_interconnect_1_mbox_client0_avmm_msg_receiver_readdata,    --                                    .readdata
			mbox_client0_avmm_msg_receiver_writedata   => mm_interconnect_1_mbox_client0_avmm_msg_receiver_writedata    --                                    .writedata
		);

	mm_interconnect_2 : component system_mm_interconnect_2
		port map (
			pll_100MHz_outclk0_clk                     => pll_100mhz_outclk0_clk,                                       --                  pll_100MHz_outclk0.clk
			client1_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                               -- client1_reset_reset_bridge_in_reset.reset
			client1_data_master_address                => client1_data_master_address,                                  --                 client1_data_master.address
			client1_data_master_waitrequest            => client1_data_master_waitrequest,                              --                                    .waitrequest
			client1_data_master_byteenable             => client1_data_master_byteenable,                               --                                    .byteenable
			client1_data_master_read                   => client1_data_master_read,                                     --                                    .read
			client1_data_master_readdata               => client1_data_master_readdata,                                 --                                    .readdata
			client1_data_master_readdatavalid          => client1_data_master_readdatavalid,                            --                                    .readdatavalid
			client1_data_master_write                  => client1_data_master_write,                                    --                                    .write
			client1_data_master_writedata              => client1_data_master_writedata,                                --                                    .writedata
			client1_data_master_debugaccess            => client1_data_master_debugaccess,                              --                                    .debugaccess
			client1_instruction_master_address         => client1_instruction_master_address,                           --          client1_instruction_master.address
			client1_instruction_master_waitrequest     => client1_instruction_master_waitrequest,                       --                                    .waitrequest
			client1_instruction_master_read            => client1_instruction_master_read,                              --                                    .read
			client1_instruction_master_readdata        => client1_instruction_master_readdata,                          --                                    .readdata
			client1_instruction_master_readdatavalid   => client1_instruction_master_readdatavalid,                     --                                    .readdatavalid
			client1_debug_mem_slave_address            => mm_interconnect_2_client1_debug_mem_slave_address,            --             client1_debug_mem_slave.address
			client1_debug_mem_slave_write              => mm_interconnect_2_client1_debug_mem_slave_write,              --                                    .write
			client1_debug_mem_slave_read               => mm_interconnect_2_client1_debug_mem_slave_read,               --                                    .read
			client1_debug_mem_slave_readdata           => mm_interconnect_2_client1_debug_mem_slave_readdata,           --                                    .readdata
			client1_debug_mem_slave_writedata          => mm_interconnect_2_client1_debug_mem_slave_writedata,          --                                    .writedata
			client1_debug_mem_slave_byteenable         => mm_interconnect_2_client1_debug_mem_slave_byteenable,         --                                    .byteenable
			client1_debug_mem_slave_waitrequest        => mm_interconnect_2_client1_debug_mem_slave_waitrequest,        --                                    .waitrequest
			client1_debug_mem_slave_debugaccess        => mm_interconnect_2_client1_debug_mem_slave_debugaccess,        --                                    .debugaccess
			client1_jtag_avalon_jtag_slave_address     => mm_interconnect_2_client1_jtag_avalon_jtag_slave_address,     --      client1_jtag_avalon_jtag_slave.address
			client1_jtag_avalon_jtag_slave_write       => mm_interconnect_2_client1_jtag_avalon_jtag_slave_write,       --                                    .write
			client1_jtag_avalon_jtag_slave_read        => mm_interconnect_2_client1_jtag_avalon_jtag_slave_read,        --                                    .read
			client1_jtag_avalon_jtag_slave_readdata    => mm_interconnect_2_client1_jtag_avalon_jtag_slave_readdata,    --                                    .readdata
			client1_jtag_avalon_jtag_slave_writedata   => mm_interconnect_2_client1_jtag_avalon_jtag_slave_writedata,   --                                    .writedata
			client1_jtag_avalon_jtag_slave_waitrequest => mm_interconnect_2_client1_jtag_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			client1_jtag_avalon_jtag_slave_chipselect  => mm_interconnect_2_client1_jtag_avalon_jtag_slave_chipselect,  --                                    .chipselect
			client1_ocm_s1_address                     => mm_interconnect_2_client1_ocm_s1_address,                     --                      client1_ocm_s1.address
			client1_ocm_s1_write                       => mm_interconnect_2_client1_ocm_s1_write,                       --                                    .write
			client1_ocm_s1_readdata                    => mm_interconnect_2_client1_ocm_s1_readdata,                    --                                    .readdata
			client1_ocm_s1_writedata                   => mm_interconnect_2_client1_ocm_s1_writedata,                   --                                    .writedata
			client1_ocm_s1_byteenable                  => mm_interconnect_2_client1_ocm_s1_byteenable,                  --                                    .byteenable
			client1_ocm_s1_chipselect                  => mm_interconnect_2_client1_ocm_s1_chipselect,                  --                                    .chipselect
			client1_ocm_s1_clken                       => mm_interconnect_2_client1_ocm_s1_clken,                       --                                    .clken
			fifo_client1_in_write                      => mm_interconnect_2_fifo_client1_in_write,                      --                     fifo_client1_in.write
			fifo_client1_in_writedata                  => mm_interconnect_2_fifo_client1_in_writedata,                  --                                    .writedata
			fifo_client1_in_waitrequest                => mm_interconnect_2_fifo_client1_in_waitrequest,                --                                    .waitrequest
			fifo_client1_in_csr_address                => mm_interconnect_2_fifo_client1_in_csr_address,                --                 fifo_client1_in_csr.address
			fifo_client1_in_csr_write                  => mm_interconnect_2_fifo_client1_in_csr_write,                  --                                    .write
			fifo_client1_in_csr_read                   => mm_interconnect_2_fifo_client1_in_csr_read,                   --                                    .read
			fifo_client1_in_csr_readdata               => mm_interconnect_2_fifo_client1_in_csr_readdata,               --                                    .readdata
			fifo_client1_in_csr_writedata              => mm_interconnect_2_fifo_client1_in_csr_writedata,              --                                    .writedata
			mbox_client1_avmm_msg_receiver_address     => mm_interconnect_2_mbox_client1_avmm_msg_receiver_address,     --      mbox_client1_avmm_msg_receiver.address
			mbox_client1_avmm_msg_receiver_write       => mm_interconnect_2_mbox_client1_avmm_msg_receiver_write,       --                                    .write
			mbox_client1_avmm_msg_receiver_read        => mm_interconnect_2_mbox_client1_avmm_msg_receiver_read,        --                                    .read
			mbox_client1_avmm_msg_receiver_readdata    => mm_interconnect_2_mbox_client1_avmm_msg_receiver_readdata,    --                                    .readdata
			mbox_client1_avmm_msg_receiver_writedata   => mm_interconnect_2_mbox_client1_avmm_msg_receiver_writedata    --                                    .writedata
		);

	mm_interconnect_3 : component system_mm_interconnect_3
		port map (
			pll_100MHz_outclk0_clk                     => pll_100mhz_outclk0_clk,                                       --                  pll_100MHz_outclk0.clk
			client2_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                               -- client2_reset_reset_bridge_in_reset.reset
			client2_data_master_address                => client2_data_master_address,                                  --                 client2_data_master.address
			client2_data_master_waitrequest            => client2_data_master_waitrequest,                              --                                    .waitrequest
			client2_data_master_byteenable             => client2_data_master_byteenable,                               --                                    .byteenable
			client2_data_master_read                   => client2_data_master_read,                                     --                                    .read
			client2_data_master_readdata               => client2_data_master_readdata,                                 --                                    .readdata
			client2_data_master_readdatavalid          => client2_data_master_readdatavalid,                            --                                    .readdatavalid
			client2_data_master_write                  => client2_data_master_write,                                    --                                    .write
			client2_data_master_writedata              => client2_data_master_writedata,                                --                                    .writedata
			client2_data_master_debugaccess            => client2_data_master_debugaccess,                              --                                    .debugaccess
			client2_instruction_master_address         => client2_instruction_master_address,                           --          client2_instruction_master.address
			client2_instruction_master_waitrequest     => client2_instruction_master_waitrequest,                       --                                    .waitrequest
			client2_instruction_master_read            => client2_instruction_master_read,                              --                                    .read
			client2_instruction_master_readdata        => client2_instruction_master_readdata,                          --                                    .readdata
			client2_instruction_master_readdatavalid   => client2_instruction_master_readdatavalid,                     --                                    .readdatavalid
			client2_debug_mem_slave_address            => mm_interconnect_3_client2_debug_mem_slave_address,            --             client2_debug_mem_slave.address
			client2_debug_mem_slave_write              => mm_interconnect_3_client2_debug_mem_slave_write,              --                                    .write
			client2_debug_mem_slave_read               => mm_interconnect_3_client2_debug_mem_slave_read,               --                                    .read
			client2_debug_mem_slave_readdata           => mm_interconnect_3_client2_debug_mem_slave_readdata,           --                                    .readdata
			client2_debug_mem_slave_writedata          => mm_interconnect_3_client2_debug_mem_slave_writedata,          --                                    .writedata
			client2_debug_mem_slave_byteenable         => mm_interconnect_3_client2_debug_mem_slave_byteenable,         --                                    .byteenable
			client2_debug_mem_slave_waitrequest        => mm_interconnect_3_client2_debug_mem_slave_waitrequest,        --                                    .waitrequest
			client2_debug_mem_slave_debugaccess        => mm_interconnect_3_client2_debug_mem_slave_debugaccess,        --                                    .debugaccess
			client2_jtag_avalon_jtag_slave_address     => mm_interconnect_3_client2_jtag_avalon_jtag_slave_address,     --      client2_jtag_avalon_jtag_slave.address
			client2_jtag_avalon_jtag_slave_write       => mm_interconnect_3_client2_jtag_avalon_jtag_slave_write,       --                                    .write
			client2_jtag_avalon_jtag_slave_read        => mm_interconnect_3_client2_jtag_avalon_jtag_slave_read,        --                                    .read
			client2_jtag_avalon_jtag_slave_readdata    => mm_interconnect_3_client2_jtag_avalon_jtag_slave_readdata,    --                                    .readdata
			client2_jtag_avalon_jtag_slave_writedata   => mm_interconnect_3_client2_jtag_avalon_jtag_slave_writedata,   --                                    .writedata
			client2_jtag_avalon_jtag_slave_waitrequest => mm_interconnect_3_client2_jtag_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			client2_jtag_avalon_jtag_slave_chipselect  => mm_interconnect_3_client2_jtag_avalon_jtag_slave_chipselect,  --                                    .chipselect
			client2_ocm_s1_address                     => mm_interconnect_3_client2_ocm_s1_address,                     --                      client2_ocm_s1.address
			client2_ocm_s1_write                       => mm_interconnect_3_client2_ocm_s1_write,                       --                                    .write
			client2_ocm_s1_readdata                    => mm_interconnect_3_client2_ocm_s1_readdata,                    --                                    .readdata
			client2_ocm_s1_writedata                   => mm_interconnect_3_client2_ocm_s1_writedata,                   --                                    .writedata
			client2_ocm_s1_byteenable                  => mm_interconnect_3_client2_ocm_s1_byteenable,                  --                                    .byteenable
			client2_ocm_s1_chipselect                  => mm_interconnect_3_client2_ocm_s1_chipselect,                  --                                    .chipselect
			client2_ocm_s1_clken                       => mm_interconnect_3_client2_ocm_s1_clken,                       --                                    .clken
			fifo_client2_in_write                      => mm_interconnect_3_fifo_client2_in_write,                      --                     fifo_client2_in.write
			fifo_client2_in_writedata                  => mm_interconnect_3_fifo_client2_in_writedata,                  --                                    .writedata
			fifo_client2_in_waitrequest                => mm_interconnect_3_fifo_client2_in_waitrequest,                --                                    .waitrequest
			fifo_client2_in_csr_address                => mm_interconnect_3_fifo_client2_in_csr_address,                --                 fifo_client2_in_csr.address
			fifo_client2_in_csr_write                  => mm_interconnect_3_fifo_client2_in_csr_write,                  --                                    .write
			fifo_client2_in_csr_read                   => mm_interconnect_3_fifo_client2_in_csr_read,                   --                                    .read
			fifo_client2_in_csr_readdata               => mm_interconnect_3_fifo_client2_in_csr_readdata,               --                                    .readdata
			fifo_client2_in_csr_writedata              => mm_interconnect_3_fifo_client2_in_csr_writedata,              --                                    .writedata
			mbox_client2_avmm_msg_receiver_address     => mm_interconnect_3_mbox_client2_avmm_msg_receiver_address,     --      mbox_client2_avmm_msg_receiver.address
			mbox_client2_avmm_msg_receiver_write       => mm_interconnect_3_mbox_client2_avmm_msg_receiver_write,       --                                    .write
			mbox_client2_avmm_msg_receiver_read        => mm_interconnect_3_mbox_client2_avmm_msg_receiver_read,        --                                    .read
			mbox_client2_avmm_msg_receiver_readdata    => mm_interconnect_3_mbox_client2_avmm_msg_receiver_readdata,    --                                    .readdata
			mbox_client2_avmm_msg_receiver_writedata   => mm_interconnect_3_mbox_client2_avmm_msg_receiver_writedata    --                                    .writedata
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => pll_100mhz_outclk0_clk,         --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => client0_irq_irq                 --    sender.irq
		);

	irq_mapper_001 : component system_irq_mapper
		port map (
			clk           => pll_100mhz_outclk0_clk,         --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,   -- receiver0.irq
			receiver1_irq => irq_mapper_001_receiver1_irq,   -- receiver1.irq
			receiver2_irq => irq_mapper_001_receiver2_irq,   -- receiver2.irq
			sender_irq    => client1_irq_irq                 --    sender.irq
		);

	irq_mapper_002 : component system_irq_mapper
		port map (
			clk           => pll_100mhz_outclk0_clk,         --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_002_receiver0_irq,   -- receiver0.irq
			receiver1_irq => irq_mapper_002_receiver1_irq,   -- receiver1.irq
			receiver2_irq => irq_mapper_002_receiver2_irq,   -- receiver2.irq
			sender_irq    => client2_irq_irq                 --    sender.irq
		);

	irq_mapper_003 : component system_irq_mapper_003
		port map (
			clk           => pll_100mhz_outclk0_clk,         --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_003_receiver0_irq,   -- receiver0.irq
			receiver1_irq => irq_mapper_003_receiver1_irq,   -- receiver1.irq
			receiver2_irq => irq_mapper_003_receiver2_irq,   -- receiver2.irq
			receiver3_irq => irq_mapper_003_receiver3_irq,   -- receiver3.irq
			receiver4_irq => irq_mapper_003_receiver4_irq,   -- receiver4.irq
			sender_irq    => server_irq_irq                  --    sender.irq
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 5,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => client0_debug_reset_request_reset,  -- reset_in1.reset
			reset_in2      => client1_debug_reset_request_reset,  -- reset_in2.reset
			reset_in3      => client2_debug_reset_request_reset,  -- reset_in3.reset
			reset_in4      => server_debug_reset_request_reset,   -- reset_in4.reset
			clk            => pll_100mhz_outclk0_clk,             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => server_debug_reset_request_reset,   -- reset_in1.reset
			clk            => pll_100mhz_outclk0_clk,             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 5,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => server_debug_reset_request_reset,   -- reset_in1.reset
			reset_in2      => client0_debug_reset_request_reset,  -- reset_in2.reset
			reset_in3      => client1_debug_reset_request_reset,  -- reset_in3.reset
			reset_in4      => client2_debug_reset_request_reset,  -- reset_in4.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_server_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_server_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_server_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_server_jtag_avalon_jtag_slave_write;

	mm_interconnect_0_pio_s1_write_ports_inv <= not mm_interconnect_0_pio_s1_write;

	mm_interconnect_1_client0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_client0_jtag_avalon_jtag_slave_read;

	mm_interconnect_1_client0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_client0_jtag_avalon_jtag_slave_write;

	mm_interconnect_2_client1_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_2_client1_jtag_avalon_jtag_slave_read;

	mm_interconnect_2_client1_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_2_client1_jtag_avalon_jtag_slave_write;

	mm_interconnect_3_client2_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_3_client2_jtag_avalon_jtag_slave_read;

	mm_interconnect_3_client2_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_3_client2_jtag_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of system
