// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pSSMoMzqWpKKxMZVWVGwLsTgr2Z7z28yUH72qWShzIqEEjX0sct+P7kbmCr9XU9uPYqPTzoB9yMb
8+VsLni53AmSzT1dVN6XqT2wtZ1xFgk1VXY6yOSiyD7F5PhZE9I6K4pVS8E7Acj7jC+LqvXdx2P+
qF5Z/5uB8OCuQxWsUGWUzgTJwd0oICAgw+947I9fF3rduUPlA4X4wnY4rU6eaDCX7gewU3oNv8Kn
PPAHQAY8emE1A8bnEi2kncku+c2wxUZ7i6q72/sdgpAjsvUOe4o3Q05r8kJQlIubW0beIanAQM9W
B3rE6VH5vYyGi9vn68E6GFBf+IN1/ZYK2swwTQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12880)
ZlVC8irAbxUq+6gwsw15PAsBMfUYTmQepWdaRVLh4AW2teruNBXMvtt+cX1JWnA94yIH/y/kss/z
ItgaHumCKK5pGDHvhO/xxRfG8AfqnvucQNNXRzC1zRHKV5ZbcGVWwV+UPXA/Yzw94JdsiLxU8x86
VmEDsUclz70rsTK2tW6zXXuzJTknky4L4Ht7gmzhCnyZnC/tEP3/daeD2QrpW62l2+zF81Bj+HTt
wmmkdri8GdDCLMX3a93id7Dxj/qpJDCtS3j1JwKDKbrTZWi5ZKFZz99K5NdI0Y3D/ozoUtrV9lfl
hspDlXRLMrLkfNrEZQ3u5VZ+ml0tiaa9SmIoCG+BXeuFTEeKTc6kYD7Oiz7Bg1tbU+lgkUwN/9Ni
C6SwXQ1rUxoBcd+kuEMPrETt3r9iHMkw35jprVPqBm0DOAyXB9zv2alZJXqzjb90TjEAmBdrNXbz
MygElB1ZJRx7UyK7rH1nYrzpWNVOiD9eV8phsIM2SU5LrasfRBy3Q6WTG7jsC5Hgi3NDI45r/zqY
LCoXBnZN33Idj6Ap6mOIZQsweRCWJ9OjPIIHuoKojxLvj8e+lzOwDrZYNSdaiExmV4rMQp07UJO8
EG1DvTSy85KZw1yXWB4BGDZaJQ/IlmsGBhpokG+rXgwjPzWiRh2QeyXEQ5A/3ZI5wMPFBBqsYGAi
OUsDfItN004pNeiZ3gPT4nkZWSXaWdlI9jx3WvskmRbpy+nbbNIZFkjFLPsl/NJVC8iyGFL0lAvP
bLkpbFxq8CVc2kPtj2YY1XZBNM9mq4RlWLbp83ILxX//bhc1o5GvbzSFHJQ+BnK8eC31pnbqmY0x
qfqYsAoC3JyFvzXv6UW3TFzp6N7aRzloj5sy19Egkk3YkitZ9chOzEmcAuoYEyerf/wqEn0QycG3
/JZl2NL3JAp6/Rl2c8sPXgy0aqb1RTlLYJCJtWjy6fmSoku9RpDINo3NLljzs0+SCMaDdbjAMelk
9XInDRLyNgpDO/H3ZSBufk3Eo3FM7Wb8EAu4DIduR+YUVApix8t77mWjGbO6WnhdRc+MhI32TFIC
buSgxDeqwhBBybi0KStEhHMrr26SJqt4c8wHXYHyD2QCV93tqRLLGTd+HYFbFNDwFtPSL6eGBGMX
JCLKI35KP6c8fS965doToJ86XoBIc6go2mg63DRLDHLeriKdTR+pY7mUgS7nMBPMd6EdHpkUmSI3
ZGFaAG5ZEuGQKXy2o4/HPgBB64UpRrax8RcFQzt9whBaR+RwGC1IO+4a7t/P1aqE/R5MUIYAZkFY
mHHS6U1kXZzSYHJYls9Hmmu+86/OZQCgpSpME7713DoLof6kI5ug76b2CwGTZd+N19hHTrPOibdv
Oj31XB7MD9m8mKcsneLKN3gDvwPed3I2VfErR0kinGemY6o1PWFJaB3IJcqA3c0zW4+ThzT9At2a
hb89CFlKQsA5BnM8xovRzxjyBGXRWz3yl4Bx80uSwmdfV6og+L93X4m1sPk7jdmGb5fVoiSakF1U
pTr32Qo60SZNnVldjnIlIganPy2XKPwztQ0OCHZGSoFyEVKIFgTTCDyK25J8EJcfx34q0gOkK211
dNQdEbrmWBuQn2T/exuHQ6CByJQpJLPcSPX/m9TRPmMr63SM9DdbjMufcGwkGm50IogBaH7Ur+am
bXEQZmOEoHg7SoDyHi90ITxmFEPBrAUAR8zXgo5vmzzhqPfIuuCksVLE9XpWODKV/HEXnkjL4YSW
zoVJ6X1m/B2fYkHY5kWI81XKDwl2IxRqan/FRXzNB7BS3aB4btiHfnJhI4e1YhDu/MQM05f6gFZp
6gSahJiNmxnsODaPJuCiKavWhiv3tvx1/kvuOVwD0IaHVd/hIz9jqotPoaelWaTH+KRYzcGC/Mts
+HyW55ovVNJbAQerq717hrRZe/taUxyQNMweWIFcUYoG8WtPtuid0DxWI2U3wgJ4HXX1AkUbVcRO
wS4GjVvtHLAuKuV5uvHGZZadV4cBF+W+cvdMHhkT4HuSUqvXGm+lMAkJKXmKGJ5ajmwyA6zyBcFN
6HJ7Wb53/UGwSqWogs8ghXEOeB/sqNfMEIGF4EYdWrLIorjxXkfzh7LcITuajVwHYs1vRDF6T70Q
qxptGvjcJqZe67JzdvDbqKJeN8y37dVuhvQOjnkGv79YaeObWb9rjmrqnxplFYqrfqiy4pghnpWi
UQm33Gz/4g8GmjxSTrWE3u/pZGfZHjhcxDISeVLgqg/NbfFgJuK8xqDVXukKsZp34uZCZ/rOpVjH
uKKi0ZX2IW0Ve7U1J1PvfItfzWJDvx9z2THl5Az2xhkBjTjBHGaT6tnR6pHLKPPZv3W8lSNeoMgj
pq4V2Yk2SQw6dmwDHMioyvtBG7DyRRyPYTfC95RKC4CmORS8+VeheHhapCbcUNUldx35OaOWEWOb
5rv8c83tnzk0ouZvEmJelNBgr5A3RcEKW0bUtv8p7+/UzbNOkO+xfs3JOfrEKpCJipQYcsEriUUW
JkeKHXzxB1KIOBk1aykuQQQ2CnuBaBqkto4HAWp1iInAgW3TRMHyY81sv0d9WgMSA6Az8Ju46PML
dtUt3m23Pn8JHo4EbbgJo140FHBGNFER1IbEbf7tyMCBL+osBmjTJzOSa3wU598oULFcAXOL/GR2
3wR7M1RKmLMfVWRWKQ25mCq8sFDEwHKMnxdbM8rlk2g2Lwb/ipMWnnmXKQgRQVFVdK862toBWlyA
zDgwNryJLPSqV2abYu61P03ieHE8TPP1BIDRq6hREZLC55vbpK/dYOjec6L9jaU8BmUsqD3TwI/o
W5nsRgMxHDDGZw88S/cyylRpjoU+1V7zDFPOBrX0+qr3ZRtXdanSeTGjaoMADXJ7FXjFXKXYtH4j
LgPxXdOHQHt39wnFHgcicS9I3kcvHHsAac0erbFfXPbbvF9ZcvwE6b7Wz08FVke4pL851zSxKu2I
BmbhpMpxkoR8Za1q7lamGZLGjYm8JpHy7kC3Ywn5+r75DKNi4mMvGNHakoYXg0PfEn28UJp3z0lg
d1XJqhlAMxEtb8dAP3eq830U0wlyg8u+rq+JRL5ydZkXccwoFUS4HKQOUgQeXBnu3F5kYnOjw3Ih
6xX3stogKsq1evB0+B3nFYfJh4eFB7CwSrYQHG/gtL7vXzzp2ePBVpEcDuChsRfJNY4jcxhoW6qn
YknmHhunv1mm+lOcL4zFXQxDFfcOU7dm7GCn+zDDXi1yf35aWwD6WMfnUZ3HJeUijBI4VrLvA9pz
i2zLDU01O02MIZX0Txq+mPd5m9yYf+8TnZ9+7CevxHML4vfVds7sAV7hhekFNRQ7i3g86QvkO0dx
I9xIvGKM70bOhKBqsubpAMJqA75zEAjefTYOD/U0zWZjeH01Otcv3of8VCQ0QmBakuycjWn+0ckL
0PWBb+aalFz/LSKXl29GdexPCPXnwCa4UOB7WJpi1SyJQKcNUGvBiGm7DXNdsTtdsl3WSIJGD8qE
mYvH9PW+cBbNA+H1ooVqLSUAa+2Tk4BZ7OHUv6iNQ+UWc0sVYtmnMvvjUH7eTEjxbNWxh/q9FOW4
g11Mo8YHuE15O2VEf2tFxXaKv37HVONOjWNSGW4NIMVwk/3GFyNWzUU5HBsTMnFzFqckK7WUdIQ4
k4BfT1e7cxxnaFEk3gFGOIzsXBl1EpxflXLKOmA3QlUb0d8KP6I/iAWSdIDGflnjF4JoVyP1YTVe
R+89Hwv+X2gzTVDafg3xL6rwwXoMuyVxW3f8s4avPqYfGnNPZzEYEdZUnSHUBeI7PEiyIY0OcFB+
Gw0BVSmY2jhPxwnQpT2W1hsjeMiv87LU1FkW2WLeGPSliHcBpZSOIN6o2lyJy1xLzmItXXZZW0Dr
RjD0YUSR2GsyvZYk1KLXyvAzfC9eIL4yFSpqmtRV6m6tsstiP81QWk2E+vh4FOF6xoaGluuROD9W
obKwn3pHhse4jH9ee5cWjYjGCDEjuxJduuPkc5bd99sabDlM+hKapmcy3rtmsZdqQyzcsx4/NJCe
zBydLUNdHrSVFzvcEfbX3DDvnqyqTEZik2KKcPeiFHfmO1I/fpP9eu8616+4Cplnf6vAbO174/1j
96goiMQ37yu4xMfLO50G2qF/jb2sR9mVX5vdg2pvk/ZZj7Ccdc63gYcu76wM9LL0uxj7z/J0icsH
fpBbTp3OQJeK00cOiS6uiv0CYop09zSz1EGE4T+PgKCYxG8pGBnq/smvwHg07cnogkhxCMZp6QGx
j3HVXy9+zPXb0DeUC7TCOp+KcJlm4x2AvASbpgJd+KI1pODxWr3dxjneadZJ1WhmrJeA2sJZ2Awi
ntU+nyhbnLvPMBJRcEgGlZfiBMnr84flNgV1M+CtvhCaoxBHWnDF2PrjUa0kXxjP5X+VRSKxzcpg
1Z1JK97z8rmBd4UKW8Ba5JhErGC44iEZQfPPR4j10y/3qoJYQbrlazwY3aD99fkz1wGcz0Rw4XI5
1RCZXenAYd0t4X7xnCS1PPbPtdXIuC8w8JN+HU49jvHnaH4h0u42YcWKzg6znJOGfwtXQbLe6hET
S7Txr/mG+AM56MBjjs7/O3PXJdqloIef/X05kphYa3TxnYF6cO8zrFrwFdc2NJA4f8vxcSfg/Arg
pVy2kgAt3O1UWD2qzOhgS/l8OjPkvhd9y9ogn/fk4cGqHAi0gHYW/SwTEQEjSNPtPoqRpR916bOt
1s2/6ivAi7l1LJDaWZsBoJjOxXSAjp8S5GLpEQnwlikXPP8flz+bksBCY13hDkO8a1yVNRxdoUYJ
B97tcfNB+3gNv5OauboMsg12PqyDV2XUhbqe906NtjeRadFMayFXn25U4nQSZt+VX4p/5O48Y/B0
zeFCZzzLDNUDDZGFLZnt8NvdcSOZE1bgxTSPZomXyaRT+zq/Dbb0ONmPzAJK3EVxy8oVCstrd0uJ
MImMupfCoGW/jeZsFMw1ZyZNFGWcXcgL71ka31kHDLvh9wa3AhMqVgbb0HjQD9uIBFMkJGmtu23m
vUUBtWg4waU7/W3InqyT7oWpowVVeFi8N8dh8fGkF5qFDZvyQKbCAGw7wAxzd76yH6AGUCg+pLdj
nekkzIKZkgzyvZas+Pl3xu2QFERNa7kwpDKvbedlICRXo23hZYQMm7/oDm+v3bzXYU8i+glMti+c
2bnwzoOai5qPbVaGM9Qba6NMdLo5WAsDU6uEg1gQMfbPW1QCEaC8Djjd+ETe79CgqAYEhF7AAODx
q7k7aclZx+jCMqdBpHCxf5NfSHzzt/u5p0hYjChm83pgHtuAmuDUJ6nCkZK31L1u7HGge60oet/X
WeOlg1x9mjBtlC6JaPvTuYgf97TCERuFBpTEbLoP2bUamb3l6i4wSC5oqjLiAv4r1mdJKkVQzWul
nAPGn3sEGZgHWVxB+lqkgyww87hpM8DfAnJ+wN+yNfzYV97LB+EsnT4/do1t9dFtIDAUJQHrRX3O
tSinl+gVMELF9KcqX9EAJHNCtxwVJhL10Uep0mFB1K032x64JPt+bfCc2mqeOY192882nov4EiX9
NA9EU2DjDSCoXBkkJTRqlq2WRede4ARLYSQ0E/S+uddZTq5/cw89P3FkY6KYXVhOX3RTFL+6gNrt
WVaVRsiSb9B4Qrea4cvdBx4ZArSs/AYzWJngaOxJqU9FJvL6gBQCzC63Z5Fytxtu1nh7gn1PCih5
OJ5bosgohiOEX+uMryg0lDfcwvJcoPMpJ6byLciTmWT3kQcsMkqR/RP/xT1kk3rmxq4uymGL1ujC
cp0jVoyTmt4pWZYZJPg6GFMkVYp2q1Nn8vfoT5XWV/gvtR4DFaN+7YhWY8ZUb9ij4mcEDNYIpLlL
VIXTyqYPEfzAv1y+s3OkwocPud/HoaAZhFrMO2IX/EmhjPXAsYJMJlJ0Pqcxx7O3b5QaoBnBff0g
IuI2CCVDqfNLUXEDkg4u3lb0iUBQ6dqITj+e2n3RfCJR40eQwkWXIfn88mvtyxdyiLfeGqOynRcB
c1oYRQFC/cQJJtBlJRVaij2jWHkvvhKgpwK5sEIIb0p6nhIsTKVu/T93x6ZV9oSgCuYwXV1rXM3f
65p6Vt+jyQkjXuu18zCHjbK8wp0XaBUaR8mejjfVvdRI1yjptF2Mc0Pt90rWAydkoAq+T8/LWn2Y
igXWJc1GZMTvCfPeUK9oC5lkabfM6xJjbljJ2yy/aa0OhS3Pg2soB75zojsyWpW9Cao0xcZB9YMF
7SqUAvjf+lFAF+vi0JUHGICCEVBCAVZKykXDhG/yJK3sUx9Agr/MnI9IjOKSq2Owo1FKuF8sru+T
DFdhHs1cRysfDsXbqkRnx1VYi7qT8wIaebgkXQXPu3yoUQ3d0V0AcZ3V6xRk7zDN/dXYZw6HUGyw
L2hJF7bJkR7xI/klDoAmnngRR2rw+MHcH7Mhw8o/C4Sd+F7rAq5hZsBDubyAGuuG+ttZnfIjNOZS
aH6LDserU8fqCHe6aDsx/+4fXo1nxNTlDIe2lx87vzO5j7vyvfRgmlMPTATx0uDjSR/MbGLJUbrK
csSz59+ycFHBz12WAukV+VQ9MvC6qJUkhrocgm3CGvi6yhRuyacisXWugR5sj4PPKybP5sAKZahV
Uyo6dd4bcaEF0f5MvIXhAPyLubJSMA+F4+PBlRFScazLXz663wRQKcg2kzFQYQCRgQr+xw7a6CT1
MZ0nw6w46a1qEqXZMA3bTvq10+UZQ+WLv+QuKmeYvFmSQyMXP0l7fRkx3cbfXcsvvtDbtOCeATCg
jnNHRxO69lqgGvlfSzJUXK+wogzPhoINowM4UXLTQhiiP3vj+rdvmjV+dETl9voS4rcluaPB3BnY
JEawcTg6fShWc0L75n33QFgCKvEhem5O2ajQUQYlUUA5WV8/FtsfKYBM3V5rpxnzVWX989CgsTH8
5FNGdwEvGZ8Q4aqA3zpZ85MXYFyO2siEtNZkOn0fYh41MB92Itc8zodWp5+Z1w4q2jWeWO8YnH5D
2Cr/F1/4fOOlAeihW2nD+79eUNRr/Qw++VoWbfHdof51Lnt9cNekca2qyqJ1AXtvqu8AHg1Pezxd
ZrpcauUuCVV0XAqSHLEP8/JWBLLPlOjW6UIQ7Yce6/Mtz09VGupCDBOP+S0zW3MdzFmWFZuWu/CC
OtcfjPasiFc23RAHceCiUQYn+N9LKi88MAV1QFjsJf1KMB0empjws2kQeD+Zo6D/SOSKRz9EGxUR
GRo/YHUBNVe2CktXJCiHlTF60mdg5WSgYONYDxz4NtpMj9PeZGskyBL0Q5751ekDkZkJMdpePKqa
YF1yAJuWSOxUGESH9C3qxgrRHsRzJP2JaaLpXpHf0o2EXUiEpoGNFzpe/PeI5jbdZfEsocP3XWNl
6GdP6BBQzOwpbnJ0KSCYEZmn2TTz01lZYrkBtIAIQbf0Y3wl5H1JYW+4nZGss8ksT1irtlrhMs1D
lnHzS/q5SR1EuBIHn+b15BZ2/kcsY0U9dxwcK9ZLsA3s6phlGr3Uxh1GBA6r/LjDUHURFh/2I2Ww
RkJvHJ8vN8ZlBtOHCPiHW0f61J5SSU7thHSI4txV0qV8CsnebguBavizIV+TuiNaeIAuVQhlCyr/
Dznb7Z+FyZ8dLVejNHtu6jRYqf+eYxP6nMh2UzIbockTvJUYGvRAqjzO0NewjDIgnIpDlTRBVl2d
lpVxE9Pku5nI3i5B8ebuGIhJkjM4XM0gYcfCVF8N5c7MS5DAx1oWxBNeSyxcfxTvx7MQnnkcT2N3
tZrBVtzkny3Di5m3EjvJtv4BrGyHZx6aUeV2UryoBmEHPSOsYmGqY6NplLSE1DFaOMD4s50zplwG
f7uU2Kf6mw8LOt2fQrrTfW7+XuQtEH/OLcvfZtDYMBVJZuGOhfbvTC7o61bgBWi6G1IlAOSn8ZoT
iVyb7fe8lfYMuiSPcFxnSNgPS+AvnXFSNqLP4wDrToz4V3nIQwH/HjKYO3BNCHLQn8iBkHG48p+L
XC5B7SDvXKYQexR4kRx5cnvYsGEGU8KYUIsg7IabcPdT8p/RcyEI0HDLofihAPigPkyBgv+KW672
QM+UYrPZJFsi+XMz2cI0JkOcTJ2V//XI+U7vBjPs4Iu/PuO9KjWXuF5Fko4jnLRygDUMhtK8xHmA
MOvVTju3YCmjPJklhyBmVHwhQTYzCFOUWcWRnQURYPbTkbWLtuRJuMZ+8xFoccwsarCbIkU0DelU
pZvSyZpjszW4DGKjlAm/vfC28J2iA0lPDcEj78j15FvjitAO+tTBBdzYdoXhxFZAjPe7WqI6OwMH
qmJdBs9d2ypQaGPpTIhaYOCBVprcrAzjkPW56VJ+rEWOZ9DrlQcFPiKypR1VMU/8xEQ9dt1yS0RS
mT5GSWpS4WRel/+NEmpqtWQfViSDw2BQdoJvjGVMAjiNEqx8lwcIrsausvR1U71U+K7gfYYxSsC/
rEfJh8boKuHl/TX+nJnL412EcBdfMUDmhNTxGcnC1Kv6BKtswxqi6r0YbtoN16sjDOQfzzH4vCJM
fkfOQrzeOnyjm7fsOMs6m0NYIpx4gCBFCE2gVp8Lv/1ny/bXez25M3GGEW4YlL+pxwhMHrck/LGB
p9+L/l+fttXkots4E0sXXRUGDuBMmpMhKTUAnyeCYTLsuUokVK3MOjVYNqvWzE6td3LR9ZX9x2mg
KVfGay95mIXyEbR955Z+tPhHgeleP3l3HThcsC3O2MsTqvoyUZ1sPSV0EPsDx0XMwloBbf93tasd
OsknhuD001wJCA14g1RoSceNdU1Egkr/57WSoUu6kKA3FaV9Nziz21otQhgnV6YL1qtPG8tMLHKb
WxyfcxqZABQtOo6tWiCQUwTMgD+kpcP1d4+JoMgygqaYnFhWYnL63oXzkSvQJsIL12fzwPAs9w1s
5RyWGsQeUceGKZL+LG1sK+SQOVraYrJ9rMpKjZzCbyRi15cLENYmeVMZBq06WNOF+kRtBMLFVJJi
/xykQjp85hBr4Dmm3eytnFJ2P7TdV8FG+qlipCFyv4cppwldS4vpwY09h60haBgaI8u7rwreGmY6
GHNbWGIB8Z9+ySUgsv3zZ50mvUe3bvHyIrD9SAqNZOK8xUx1eMgtoT+wk2oaUeMmLHDVm6Vo+Xc5
zGjJwoMTg4j/BFpzoXIM73E2IY57BcSmligtmSJ3V8L4r4GmajPO6ovRBER12dj7J/OjAUusyZA/
WTw7ZseqjpXI70ivJo00aqa00m5JmsjtITsi1qiPfrrO6G8OyfOElMn3zHBlYeHYXhdXaaKCWcm2
6cM3eraJGWEa5+wkqCxFqSzmw/fJZse7mkO4alLEsi+EjQ5bEMk2z4zu5B5MPv8XeSu5gBtLu2If
cRy54/i4xdsAjwu/PGZXY7Wg2v3RRh3V0vcE/wXOy0zfo5WTL5bHvV/lI6o6/g0Ecg1oN3MmVyVE
ypgSBgJeEj+DolQ0V9GnxKa5T6TMv4KbY8o1JsXJWzNAQfJE7zzoHhaVXNXTE2Kn8U/I2pQPMiwr
mD9Rg3tte7ldMqyyyjyN4YjjjeBfp5v4KjkyA5XanlbVjzkIrHAG5bSaViw8SsWWAEGedDf17HPL
YGFb8Om3UUBQDrGjpxZ3ZtJM47kcj+OilyJSQrbSNQ8a1CJqx6T9TFWArjViaQD6oOD0lVTKYV8V
/c6nbaOd0o/8kU3q/hBNq3xDQfS/cokgDzZgw7OSi2muc6LcHQmPhBRVbt5wUssR9eSZar1AvsuW
Ab1IF+d0Bg4K3snSKLcV7g9wj0tvWI4QgStqPREm20VLLHEapqiLu/ELHcn62Hvi0NWgH9NerdPL
a34KaL1OtedfaISWz6OLDRPAO20qSJr+sfvWL/Fnt+QEYMJ2ywttVBbbH8UygM8fd5vAU79XEnzz
AuHWUWpfK66VcOTj9KeD8n27iM5tcUKDblmDzzRTwME6g+nQ8IrXnxgEGkJXLisc43a8NwnDkABq
Yio95tZMsp/X0XnfbgFwR9Ll72UYAl1mt6x4Ac5L6D01jHbfm3kNFLKunp3nH6DTQ3/Mn4nQAZj6
b8ZoSYWIjtfIPqsyYWxyltQlqJJXsZyGDEefRHH32hfWoetq816YqkZaMuYoX/JlPqPT+4FIVisd
f1Hrz+Ea9vASkioRsOVkXDBWSNHLY8cV4c8kOW+L7jti57GFZ137eBN2RqywsqXx9BP4vBpo0rik
G21ElXNZ4HugXmj0J9UEpUzTFNX5+7anUb0olMXdAp8fPSLJb5hNujmyB/LBkmXwgxaaZdrYvlgS
vPcUfRJPbv+y4QrKIS96objL0vKKt+e/0N8TpJxnYwETiYNpcRzSHyrXtYLntv7TEOxmpEjyDnjz
FMIitjW2XUW7A8Rvh+FWqjnYaZoYrw08nkE8HNRol7oVhc9jOHnfHc5JLRzbVksXr8R4rU7WDctr
kB+31dQ+V4xi4alLr3VcQZjpa0gRmf2YQYnEn0ikfU0j8LwDMtN3ajUrBAae6sQFX6J7yIW1LM74
AS3X+MpesulbpOSVsBP3nininHr1t7eiv2NlKrbrC5imKaLKES8hIlezvkWiDIMja4PCXoozBLR3
TwKYL1eCBn+x69QqBPTTy7GriBS0mkG/VbHCZoVYrCXgh+jWAdCtCykMMGGMFbu4u/y/nNf/U0Lz
fgVfuthQZ5TJhL0jhULpSTaeCMQ00MS9sOHC2CeuFpc16vdSqvMxko0nc1fpfkobOyAinx/EELqW
wB3W3AfzUIXFoPfKWqPhvqn8vUPcdWad0fHzBX498lz0RZKhUNVxkelVWqBqI37KHumMmLZvVZsD
yA0RLxuZ1Ex+HRDAe3cuuzIqy65VFGnD30i8S6290OwN/HJU98yyWbQoPS9fUR+NvYG0PlKPtM2v
mgNttr06xrJbcvmnVGo2oR868DIhFLYSMZpE5ZvcJ2BHkcgosJBhth2/qtNEGy3JC3E+wIFE5iyy
Z/IzWzzGrT421BLpuEj8N3KxHOzwUeP4TU7iKetPiyKaYCfELkIHSJWYEii36VlWqURheO9qXIei
NH5p59jhXaI05awGvf4Awi3u+jKpBQS4ozC4t8P8YgS6WPy7CaS43Y+WFhme+0iJFiQAXSSUgVnD
q1PmyBxNBR4VVJ9OJfM8xDugxnCR/hYlUmHZv5DzyfaorNXJ0fnPLbc3BXpIR30TfxgnoGbC4OZw
NQ8sgthmwqD+uZ1JIXGyYDSgN4CynnYZXgI5DIWmfSs1G7fT2CZh71229dIiG/JqbhBRphM6y/o2
VakxejK1DsrCAEw1zGYUCX4PFHxz+XtAo23DLpskWzaYuCT7h1TdxlmEajEF2AxHTEoaoSWUAC+f
JMDZKuSlwKBDDNkFkzr2Is2SOPDZHtnbcL2rPLSaZIJF+GfBGol0ZQ/+WVylL5iuRGRwfFSsMfhs
xa1wp323yfxP+QvyH5NxOhUIAYuj+A1I26LB0dyCXw+eHDpqrwfLfF2jhe1ArliPaBRcsVuEQRL6
l8DbfOdbCV8zbmc+VhJ2r/GXG+z2rIgoVCfhgpMje0iOdZhy56QlCzMLW3I7xzbF48/EsA3kg/zl
LaKX1yx/jL2LdKN6Tn6eVNeUTomvz+vIHJR6ggGwSu6tVwmokpImcdIdDrYSae/QBw1o3ZnPTbvE
mHdaYQP73PtkGqe7yUpQp3jTdLlQGrX/65hSRWQUuhyNAgwHFgScBgJyfpl+Kis8UFlg6yvcxP0S
kt7Ot1dsICKZ628pqDWJQFLTGSIpQaHAhDWARbcX17+EfF4ZXLWjoybbVtNdDh4OCx5lzHap9vRv
jgxDwBF5/0SmzHq2mgCL4hX/INfhLyPCzdxOAFYL/bjeREdtwj3QbKXS20xJT617x9cocpoXsnT5
dRPP1IGgsAR6Phrs4kHmnkBKlA2LLfaYiOWGSzne+XeYK4EKC2iF7tQYELX7UNu1wdVV6uSZNICO
+BJ5/11Lwugo2WrHA0OpPJN+SSRvULEqYdqNhog8Z+4rti3pU+aVCQGHkstQIJ1KqUlmC5FrP2Ap
/kz2Jx9oTBxThQDKGSmtS4t6QCqU/RryrHUDMCJolVw83bgJpLo9/GA+rEcNuTClU3nvKxjw4gwQ
T2hi7dUIW6Co9frHo/C5UBeGiYUKtcYgr9vWVv5Fx2WmpqM+DpFxYfASxpY3V2cRlgYLV/bKw5Xy
AbsSFeYiRVs/I+KmmJH92QAUOEOo1HWwvzBM7bonZWTxxzNbMrcZ/nrGigIxf90tuRu7D8arToDV
nShrNYvQ0mQJZJH5Zy2Xa8bSPDm3P9sf1FMbE1H9+2ZSJr/y4DHn7evRqRUTH9KXh/aN9AFRb9Rz
QjjC/rF9kxjgxJuxVUpfI8xQ+IKpZHrE7FCMFW3WHD88QCiqjUGBg3EDjmNbCsEbDjJxfphrd38V
EtgRJrFF5w/3vepvZAlf2fIEm81Kv+gWcu7nhTqlq0U5Ok8nA8j3KsYhUh4cru2ogIPquPYvKmqP
PVMbPt9QrsLIge3NVRpNsHDBjreJeQUC6LwrNPMJcKYSH3F32OlRI0+wExD1xmi5bY6hh+cqcHb1
A3AP+QgdQnHkD1rQ/WWpeJ6nbr6onNQ/LEjfBZNsvGkCgpTyWgpW13oH49Ye2/bxmmRZbBfo/gSz
HwPqq6izISANVF7toOalYgwgBaV0wzu1INYafQwRW4Veo5/X6Y/pm2Rtwov8GO/0vIQu2Aq3YN4C
gD3RXMo4trOhmWVapf5ke5caXzntOHrU4BkNMRBE+9Rzd5aDdlVq2ucTTlWmVQYK7gptdaFC6+Fy
ls8tzxzSjxRT+qc8f99QjEnwN7/5SfgMqx9kSVp9VnkIixw9OCJ8xeGSW66D4TNnep5G7SIe8E40
DiYXbiYiJgKLYZmKVfEgeRZu9HmOrVTk+8GzZefkspfTUyhfWg+lJX0mK/G4AEFed+RpIiGEak4f
KQYDOM8McwDAmRcOQGZFvkmu+ba03PLvqKsX8nQiLNifmuk11w6yPI4QuhjT0Msh+oGREJfsibzj
c1XEe602skmRTpvtogY1rshzWPu0SCcDTtgWRrODPFrT1VWZUIFQIfOvK5bv2FBZgazNrEvBllcJ
sWF88W0mkqEhYEeNC0A3AGm07fpU+WtR78B0fyPW6tNvUeCpoW0+eM2JpYUt6hDP3E1snu7dDWwe
ZjM0tPYDKv4hqxN4y9pkrlVeT3ZEa7Us0QiA+2azgTsUnom5wyZx37U5+HGj9/V4d3GREzm//r6f
8k62N+AfVPhuV6UaoIyB9ilNz9xyD8IuA7kJB2yFYvXZ9Yp0UM6P939RqkGFaNbjU3oaY0/W/X2K
PAmSfewZ1XxQenfUFXYh2nXmioFKE4QJ/klaDstfQ2yiqfQGORmp09jzii6/dBpwsYSHZuVEuQZ7
pofwzSPa8MYEDKgHRtBHrD9K7pz/XNSq+c2Z5jNYVRfxVZOHaTE326R8ZkpI8dep1ugK2gzP0xBo
jzprVnshlVFmNRFw7HVTkHHLWp2quo7nZUOx0lKt9ISnOmv8Kous+Trf2rR8mb2vouuwWbW2p4SG
zf7YWzAd/oKje+r76yDQDTOAloH862j1EMbZiZ5UWedG+1vDO+QLjIXttQ/oPBZ3n1DjNPDK+hTB
wHUiNpG1Ry4+StMG7I9q2RltBRN8H0jt5HhwfV3QUMNIxqJDXCp0dRIr0QqEH3i0Eeq4pp4GfYS+
UUYHCL3FS6JZT1dk6NSKrw++2j4WUa79PUIDfxrSYLAkF7MI8u8xgdc1iSyNbrvKtFrzRdK+Oa+u
9Oq9qogOePZeKyQO7QuxAr/opJvxezYPl1rvlONDa43YwEvUyBo0OOEktezXG5BPAv4QL1YQIgsQ
RjDfdphSJ3jHIuTfZLfSb1dyQ683M/Hr0LfM5oRTGEq8Yn8zPtbLoJySNKlrj64NP4F62KicUDia
skgN6JHIS3W/VqXGyRfgEcQfhwcPeXomrfnY0xg8REIUMIuAOmtZIQ70C5KvI9ufJ5EK4W1xqgBv
/6IhT9CbHHUwkACXqT9R3Md0FtAYYMzGKTASIBNtiJls8aEGxkARGqS3B2SfRoOyoOftTzyv/wZA
s/0fD3YwwuhJ9CoAxejDhtVLcknfeFOB31g3V81outHXZcbmbtzscjd3GO3GRvmi2SLS7bsiXc2q
i/qy8fsNmdqp2FQL0hnS30wLY5HKpuwNYfupq7GWEXuDdNWhUiv2O8DzSRBeGcQNLBWcRQ2lIbQO
9J2SqnrhsmFpOisWy6GjV3Rf2GJkDwhIpRAW/N+rlmH5BCCb970ErCEMX34dEvFP6IOu/DTIAMOE
lBMKUZorxXKZMD0HSPmGjXwxIc2rkZ+RQmBN0YFKIHT/EoNRmaT0cGgDSddIcTjqArMzz5TdNHbX
G+GtmWjV18tA7kSg/QoMRtpoB9GKpY+QF3cRpBYpjp2czDc8cZ53ksKXsZdbGFjVFbj4Mts7z5ni
Fjf8Xpc5Z99DNQmWnWd3VtNLnde0bvUT8NNlcnMYc8tpjhKPsm6/Y+AMO9rbg/80WhTj8qXQtuKS
xd2uPeuGVdkgdr9orfbCVB8TWkiiRuR7Fr9cKfBYv/BXzRwv10g0wjvpF74jFkUzVxQ6hsyM9CCu
KgK8N84FXKo9Wz+1f7zxNZcjckGEc/vBwKbPJ8Ze8ofSCJZAF5PL6C8vomr3fKOgKA1zUlnExL1i
tn0FeUJwmY2uW9QeXCo+dFP6rTxDL3M8S2yE0coB6WIP3teUi+mwmuK4mu56kvI9yRjQ+q/0kKYr
q7QELS78zoIRtHrmuh5kZp1iD4ms06qWnPmNeV45uQ2ISRi2gPJoK/cuB+/29NC1jvWFMIXBcA2X
+ZkXKB5vGIyEKn9aEwiJwOkEk1umRgTd08ln5kFLU/4fYTWxlkaK+IfNsq45gb3V4MgmTln41pG7
QQ96Zo1/6CIzoXP6IHgmwRIfDyjFOIjTmSlBgqccEP7LvGtmXKNU8/WJ0pyoOVK2lDiAPMeV30Be
2wsfZQ1dCKjWdQwDrP5qWgjyA94njSSSgOffHtQRHpD4zoKF/cqroQPg7EjBGxcFYjpdwjml0SGL
qkEq2/2WLpGKAe8pLd2kicA0RQn/OfQqmCpf6Hu0zNmkTFi684l1jVx8nqey+Z0R+PrGqaJy6P59
YXdm7joPMzjPGu8w8BQSxLQauvV+S74sWEbnQMYXVHUeG7JuPgn5emBLVErnaHBj3g9sgp7hd+kj
7g/fdA1HwQevUvYN3hEVylOhnHWfxCrMbggfjH8iug22fS0hHw/dNG5ZQU9QcbFDl5kB7nrSJKoY
b9I8GSlYC5QVAF4s03trCPPkJn9JswrVki0g5T7XCBNCwcnHCmRI9T2F0anEmS2HwTXzOvxzfVVP
8+704gpBAHnSrjI+lIEOcGMCfhajmdq2Bd/91vjWHGpgMx31jNTzjZmq89XmqLQ4fojFQ/1jcsLF
VsBDOlGDf16DO3dv5Ud/Ni1bGDnlCpBTMp+CFe1XsLwx9KVHlW76tolIKWlAP6af51f1cksZtAr6
FfjUqh1Pkbdk6lhntJCHS/Q+YG7vdEdt8iz2ysdQZf3Ov+AhZqPr82TNJ2ZcgK4bZRDTMsNU4YmX
52AWd13ajmOVn2oUnqo+t/04MdaLrwSg9recBv6zX/ZEgEKoHScybALye4HRwiGRpBU8T2zTqWb8
c94ZkFO/jSqS64/BgNLw8yaUZylECXetpbOF+CS3DvY5z2dycs0zcNnlo0oqLkEB9MqQNmtWNiuy
w14UJ02kt34tQmXc0b8Kj51Yp9+G4/kjbJ80w27NHAWCV0lR5+TtaawYI6xcM0p1kZtyDjGwbh9N
wx6RzGbADOIlLY9dHbV0X1ReTHIMrHUfbRYNVbXz9o4EaRAhWWiqIo3vhiN3+6E3XbfSGI9ZIbAz
tImTbBa1W5lZerXc+c1fygf3LSAc8UIzjpaamxaNHZe8M/7vIZ7hp1m+autUtPDF6fOHWXUmhrJD
oBLHR4BSQzYwdp8HN1cEIzp/Nr8maJxaXsygc5ENDUnO6UdVUcbWbCyW/NS56QdRldY9gUcY1Aw0
JDG+9XFmkjpZa9+WkDuyjdXWmmYdTfS6QQvRS0HgNV1NeJ74woxO4wIEmuOSX4CYHKYjCviGpNhT
cjoOnLPl1Hzu181M1q/UlCi1arl4GVuAVkK95qX7omi3MEHIIjNbS1/x7MAh8qI2jJHhBHYOAmDU
Kf2B8ZzHGPA872WqKzWv935wR9KcHzuMByNvS2ZuPMq9JUBYvK8Ot5yyJrXgwcAik5oOo0TVgvyD
ypiaNQNZfSVGzTyG8jDLULlHbt3zWaLdDXxYu0psY2nJrC1iXZdHIv/mkQ/RkbIXzR3sMsFyZmAq
+HNHwa41aiBaxqBQcDoJUF2hoX+HTrtcu0OL7Xo7yA8NYxtGJ98qrssGuMZMid7f9gykr4/zfrD7
AvfShV0DSXIMu0ZuVzYhkLJ7SBrk/vAnBxdH3O26TnhS1FoYAVQa/3zmiYz8nkWo2CHrHK5k3L2r
MwDZ04wpwV5k1daRaXJuoW5rRAULke/yX1Yzr9Kw6a52dcl5NTq21XrPBKQQxo3Z7AVE3NaxnbWK
0qbDqk5J9IXbmpqaQrjZp0eOnB1CCUoqj4HaJmtlOXhFZuLY4kgtnqDjUb86wSqQrsVbqJMTZ6bo
ZwjNpCo/0LO9mnONR2tLW5niqZq2+jCtWXIs2fRTnDqGC/aXn6cL8jSdI8tqJPUjg8En1e6NYBGa
llCzDNZt4H3KcUnEfzV9I1pSJlKWGmCmni3E7ECxaOAVJZvqjNA+K0TrPDd0ZUEyZ48fWlN6PhrF
xkZhRvLAYaX2cyDehMK10L0VxLnrrrrpCSlN6joRlzL/RCaD4ybpsmyzTM9Zr0M4Ks8UWWF5+ym5
MUD0T9qWygSccfDTJ6Gk86uXY2ZHC/zzdMpPjpgjE2zCTcnFz6dFbkjrwPsdXjTQo0+s47N0rDlp
BJ8D808xFpy1XO7ABLD2j3dLz7EGQjqCmTVunydv2P9QyodmWri+FC2W5OG9jj1UboMjCsE9uJC5
Yf6u7mFGai0g2zISByykSaN2xItuk+kOVEnp0LqLG1Y1lcB8HdWJwM8hR7Jg73lTGcPUI1PksuQm
jI2oF60Pl/1u8+AMqriyeRxOcYBuCeTgRnzZsUYCJ/QVBGllKO1KNiNxK84XitWP4KLIaVlYtA==
`pragma protect end_protected
