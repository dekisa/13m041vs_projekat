// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J61KimdMijQyhGzha9APTrZNWEnnoVyuYsD8O0M+IvYuub9YPxmgqmKonhtr3g1b
XEGWwnLdZs9SWBSnEk2G3u0PAeaDSgXc7HpmwuN+0jiWzepe+0ylnThe49Qpxc3Z
ObvLKyI3XJAGe1Bu9JZN3Hq2eyNWWNmMRLabcB0qHsI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11120)
JOMav7snktz1bawOC5JdCqISeBJtkjOfcqlyU8w1z75Xyao/AzFjKU8DRQXie019
jUNJrO78zMrUjoiLPbzgHr27EdEVxzUf/uL7Te8Z9C0HWuX7qrrHrc04LR/FzNpb
wz16FEFyJLn2Ccpag9KnU7dvPnIWyIDs+JiuUiUXWDv9kmyrqh5NOdQWXQEN5cBr
AwzXLocuTdiWz5TzBy80D3/hrfgZ2++H2Xtx+TS46lSiDSZe+n4uBAW4Asa/v9c9
+3lICAqAWbvV7RXPBT2SM1Kmy0mjO+etNeYNzOTHLHGYZV+HGZImhW1THitJn1sB
f+ycg6uE8mwW+V5ea3V6hoJXWOUhyTf7SF9VX1poQ++fPorpJWuulUihgSSot+0r
F1Sd+kJi7/bOos/ya9DX+GvNdUKo/Xzs2oxkseM6H5MpvJEZsYOM5FieS6UZHZUM
amrpS1hmMs0ESp/2IiPCBrTekGhZn3mnWl8QJOplOIROha9Ak4gnt6LBz8/uxFdg
uM89Ut+f+Z9HpH31nFAuVZdu2i3J+N5wTz6VR8hBB3WKrFsVhQuQB97TefUijxHF
VRkPlry+ovqyGregmBQxKveVy565NrPeqZMf5Gm1d5P9cqGAsFhKtoxhAR7Ft9hF
yKbumkLM6GabLsto7md2+ZoEbX7qEU3JfHXQ3usPKduLa6FeZ0/wHgtqvF56OsC8
KRJY+GkepqdkzejeB7ggFLahQFTxn2qaDBukpf1geVNNGrmvfTk5/AdvPfbGwhzE
lgS4tw+kwSlG2hGp1cqDQfchi75/ghuOEqmnjJJoGfkJ45QuQFVluTM7tZOPjVbG
IhodZcX1yRA2nXyf5VqiEiRCTtVOzpc7zKV3w75OOpnDVUqo5Pm7kbsC55/oiguB
EekdkXfD5nT7ZiQ62TvJR4bHBzjJxY5N/ABdmX8Yw+j9Fbr3IRVM9s04rmFTP8SS
s3kqINGite49bia9xBmvcuOA/qYrTdEm/zoLX7nIqBM9opEC1dPv3qLHs2rcByl1
2x9V0LsaJWX3SGn31MECpHO04RFSyM57v/y1LDLOAw+Y+DFr3s/c+jTn09rdzCUl
Uwmr1O9TEF8rV0HwfBNYMcGEfHOh3kpEIYvhXCWLs+6opsCXRndlFPFgwAKGYKML
dg5VwkNQyNHJiRhVJMk4NGkCrJWH4ejguulJ2LEeXJmhEDWg5YrUKfS6jBRKPgBz
4v3lG61jb280CIteuDsTGr6wYYc/+F4R5tq2QcY8nPJCc9idWCRmgZbPggQA0NiR
YnXsrBdgTNulLq+DGc4w4+AWFPOlV8hwu3tAUKue33DwuvUY+Cej5wGK6/9Rj5LN
bsoPRT0s+S011v/1XYtht6z8mOeL64QManz/E01NHdJ3Ki2qLDYcu3c4OZ45HP5M
msKDzHepm+3Ty2yKiRb2MtAF9ZU1zZtuCV4aqL76l3VkQRJ4Sb34cAtxWU1Um+V0
KdSrgbDNPp8JeUms8DQR+ocIuX4rC38GTPvXfzbaDUF9o+GeO97uB2n+IM9d1S+c
jNZnQEWhLkYO0kerBcl1G2cCSANqVxay0jk5Sun4W2tJwjvfxypDHStVAzGxr/gZ
sGoG2IhL1j2Apg/1MkTHTFbg/49uyO6OqFgD9POn5lI2cusGgKSUT5pgkryp1D26
v66XTC++MrZ6Ew4PTCckljKz7M+m6cn8ASjS/fQH7qUrWp3TUGFx5oHXwiIhjUDy
YQX3Z0qG6wwz/SwL78R8LJHk2V1U3r7Y+DAMYYYUeBI2vEhX9wKuAzndlBYsnIuw
y5jaFM3q60fS5QEZBRIm6ajw3VpAih878lkdEaseVr0hsgsTFRrR+krPX+dv7HQe
uEXV9ed/HefNDR4fqIa5VCHFgYnK7+2fPi3XYcDGNl27DOZFLOe9olix1LgGbnJH
ZtDGh0PunkXZSz2fOsKrgc0ej2H268bUlgRREv0KLYj8WL9bFRIEq0IdwCB/4jkT
DgmcU4o2KIjSdTrRl+9uAfkhF7Er2qUaTbrbqOsQvyH9rT/Z5hCEpGo9o0lLdoWO
TShbv2nxA7HltXoQul9DD0mTj1msPMvQpbI2zNHaMJLAaHvLEoN7/vf71WYcRmEi
pB2BWOsCm8nw4QRTEzyPHV0xtSoY7O0/j7HIiedSvmxU0ETbJM9k8N2atSOwIVPd
yl8ePqw4opDjMboUFQSD52aJQCQCvd4So1qrK+pVVLKLlE2ZKrecM7M3RgK1YMEJ
dIFyYgvdCq0GFrlBxEwdb06QM5HreOznaUl6eBlOXEqSZK0D3Dih9l6683TiRWwh
sYEzqDEw7a8FcM8FnUU/S2NZwW1Z+gqeqDaWEXutre2kcJhQwK/ewM4sp4NkuvIm
Ver2wGhqlN4KLK/8cuNncNkBE7paU5LWahNfeoDf1RWl0ujZ1yOx0/bxV7m2V6FU
YR0lK7M4Z9Td4WCi0afgD8miXMXmCHckbdm5HDbPcZAN3E+ant0JzUjBlLU/8gL2
xOHc97VrV20Ksrec8ewxXanRPpdgS2v2UxGdHJoVMUve5Bsgpt4Wg8flpJnqIdZD
Yi+ymp4jeXp4vGZ0Q7n+VdLr36IvXIurha9Z0nto3WEWQEmzbTpsGg6SuXcGEa/2
OCYFEFfRXAVl39bNk8hLWfQ7MHw1H536z3WIQ8/XOxVAnmISpAJwigdsXHC5kl/P
cV4PeJg3x7zXbKvg+h53itsX1Vm0mwZN19I7u56Fm3jUMpTI7AwAcVrvzuCxJnHb
L7K5/Z9Kb93JGo0G0PX7QWXlXTGHhkcH0zW6anwi+Pcg/PBVxAlrPZstvQhyGLNX
ER6BE51zpKROOoXZ3QrZqyFOK9jra6xru0sRJeN1f8/XpsNH31RDOq7NwNR2fPPo
R/s1qvp0mN6eyRfTb8w6dzQ0qVbSkTy/X97IBnPuCXxqM3YM15bnytYaYvKzzjGg
UHRvmM1TC0hJp2Yw5su4IfO/UKf0sg1lylB2dtIQvAbvVtx7hbQGTF+4JevRtdDA
AQtDZWGsYgZ9R2Qvjb8cgP7+OAecSL+IYgBEtHVuzcfTHSC9n97XYgPnPcf3yKe1
YdSTcbc97XbTXUcmcR1/xKBR128H0ymI8unpW7Xght29Ouxe6U503yULR9FSHBJ2
PxTdVtJPiidbzCgobYKG3V9eAPD3Nbh47VArzEmdt3H0QuaeNvAIo4xZxuj994al
f1l34iUwJuiC56J5ZcLBoz7BufyGBcDKErtijxZ4oFdXO+jNJqeFXH4T87Nvu78y
uGJidgWmtGMUmqTWb1AnZzP+fCI+JPfRbmP+WKUe0/lEmcm+XoqL+dpF63fOTs9b
Qli1IOyXg8ISXjxi6PRl+suRFCDwG/zd687pzifbHtQPF/B3es48bZTvwXJ73XBC
u04hMV+FbQ2JZAoqqFkVhtpw/vrHL6HmPQkg/s4G7Bl8mg7WlM/Ej7T/4OM/T2qs
S4lcoY0+FYO0fuGKvaO+xj/tXXQSAxuNC3Rh5dFq54eKVUwUzLX+tRTdzLHSiurA
pcZ6xHDuHNEb5/o9ClRQlXiBQvR6PmfmxW5kpSyk/QuAU5kxZO1nQn8LYn1n0mHZ
zbpOWGUB7vmD7P/XnaW4yhu2sdlf7FAG2sViARS+hS3abEbY52YEV59R+Wid/1yx
5CXJtEirhMu/Liq0D+9q7/wH4FvrppyGw9UqZ/gScsL7PeR44PC9tZhP7zFFCoD3
B1/oI7HC1BQLbmMBSvvrod3sMlm1LmjWXMj6bVv+AJQFk0CaP6uD/AKleKhvqhYO
bQGQHmegFYm6Eg84nMLS04ZkoGuQ8UwNicuQnhZfmuwBlOax7iyYFb4FpL1o7gpb
xwtnEXpwzo/DX7sJ8SiNQLI9RuKnlmKsNeIBA3buqaHdNZ4g5RJALxdkmOTUQN3s
NL2xBnWFeXTX6tfykhDz5LYFkm0Is7o1aJ0H3ImgIfSuffCCGbaB72Fv4HmB3mJB
DGsbGkPK0prfpiBnYR3u6jDbnYwW12SJuMrG8Vay9P2FO7+s2sb3wuHt+1vC7amq
8wWQ/xuBXPMiKo7+zoPXjmck2og8AvJkATxPN+QRTl985/desf2EfYFdwewhSWCG
QJx3yE7XFWZ+YDlIWCZ3DOXsA0A6xTJHKTCDNxTBvJQXSA9op51+TRNyeqXI15SG
SvDYCaBdbvbVBGgj4ngB5kOY+8BuYy1+2byZpGd0kkn3HRTnq1VSCgMCHab+slnt
Zmik6lZBrh+JF/9odoPFRBl/g4frmUyr6ahAML5+sphuPPUHKl/5D1do3h5q3tzV
DLXuHnbwCZbyiZ2tbNbBIJBy8tstdA4z4e+opz1etYYHqncugPAdj6zYawNxhbGA
NE3qh38hLIF+rDNdY9V7C7q9fTc9vlTwGtGdOnHTMGTSA6kEnSXRD3ndA/Lfebrp
eB+lHB/+faDz0jSWoPsiuFunmz/f4wGJQHB9/6JUD2Uvrym04SMc7FFDirtfaDXK
Zu5c4ssj6+RPwCYanOFFCPBKc6CFpJ0Bpfvo2rzCETE9fHeoKUnAX3FCJA2dMctK
wazUBh2NhC64IdnPBRb8LXZL6L9dG7rbGgIhIMm/uHREVARObLrS6u3UuZ4USYGT
usiyvZyrd5gJ0VXMsYfjeUlH5dzGNuPZIPiPFNyaUf2wDw6pE3ITSbBUo3MpnBxy
St7a88Sac8S4F6dBk6SCmlnpF0TpxkEUyQKMvnMxs7b5Azbh0+tjnVxyjP3R8SmQ
nH8USnI49Ec9eXxUHvTxP0GPkdlmgKyEXhMVV0V6Fn1QNkjwRA9Kc3AN3RALpGoP
zOaj57MsH1ghndhU9F4vr4Qf96Bsa3ww7dqTTinwo9duspE5QVUC9jpj0ONpAUN3
Xn69mcHy91Mn4nmyCDuMPpi63duftVBsQTV7PBWyJvWIU1bDWqJd/h0rzejYvAN0
ReH17IFVVV9jgxYmXwmSrwFDflEj+8H7V0SnmZyvn57qbNlsfXa3PWLI04+gAGF7
dtKpEs/h8oqpJp1iET0gHo+oV5h4EDQ6Knz+j+peicUvoiRMTL4V9DcGT34Zl36l
A7BK00vihpdIcxODWEi2QnPqdK6NhXOjXRsgMINS/wWr0TbKg9L2yh6ae3LX5Fyf
5NiCYAHThIlF2Pf+/xsUrZS5SkwlUGt3iDUc9tgoPmusiiyQZHQ1jVaviz9TL7J2
qL3aDAgnh4zJP74wacet/Vcwj5bOeAaaadEibSKTew9IS+opFPdfahns41bVdrUJ
oqK3JJWz0g4rEqQcBfoCDVIVntNOwAJhh3JO1y3IDNvWgBit9LYWsVc3/Tz1/Gou
2VqxnhL1dLQyGRkA72Hek8DDkuxnk8zxpRJm1hf4ri4/488709HTH+lu2HwgE2hy
TPsW7zJbQsvfhgzMb6re9FXF1PsSMwYptbZJXNlVtuhoiGxBsQvwNtlv6dXxqniS
qFw8QMPdg12MMS1vmFjj11+2P9itPMuA4w12TtrJ4IqMYq5ZSuch/8wjDpIVzsji
GYqXimYtds9GDTbJ6h1kSgRrZw+8bcPGp3xdkLiFaYxozm2XC/nmiVPQq+pBoILT
ZPLS1Hzr9vr0IYxYZLDXzdhw4VubwtUKEgoUvyxffJ+sG+x4FbBzPvTfzG1cDdsD
cNXEtiZO+vmjWLePMTp5/1++d1eNj3TAcAkyIA7tt0kISLABtXFkCS/QbC/XM8qy
dkqmfLujiIJhUhAh9tQpRSYmUO1d0dq5VJX7ySEVTE72+drykTR3qxEvhmgeNkPk
WSysgjSVhBPLDZM4/1la+36bPmtYxqv75qX2wzxvahct+Ii/Sw/w9D1gl82yxWpV
q6tJ5Sp6k4/d523f6Iv4uxXh4XTZa+XEQxd/hHF5WB9C2yA0QolZIgIhyvqE2n0N
yhn9PfyN2gHBFMliDGLzi0ifz5Aac6L97oXCwgdOeIIG6o4eWjHWtSCwHr9jX25S
BvlLT3dt+SOSkDcniwwADd7gAyJ2vIGNmPCAIUlLM5oqHfePP8maN0RuR6AshYG2
Q/1QkVJ4HecTe92b5AXU3eRkwykvT8V6rPuSvo2sSvI8dR+ifcI5anKYtNAr5KRQ
d09FbsBG/ldiBkN5g6Z3GYpNaDD8HKl87kT+4Plx+kjM841s/aZIn8KRLyAbraYd
TIqB15p1rUs+ir3UDRSOOG1cWGV9qauAXOu8fyuUkPHmUf0SrOFPh6hqumh9L3mu
WbnhlV6m73kw8ldEQ3y+j75dgekQrFr8BeAxyeTtsWfWxYmnr9hw+vXx3mS3bmBm
JQ1+PV6bbHCO1+UpH/RGHDKLiquOZeTXlIZYAZux1zdv2k8hz7B1qEW5FnU461ru
vMIMe9pROSI4afPLjtr/fbTY+Mv9Y1co5iPys96kDy+zRUuaNXdPytPU9hpVAAWx
ICFwQRBx94QvnwERDh6rF+VqKhHCAGIpfR401sbmIgi2SrpFtmHpLMlPuK932ezN
nI4bklQRjFZpIIe5Ll52cuDy2Wm4COe+h1MPrUETOajKFvHIgnVPR5u2n7POmhko
J2EQT5h9xR1cmqJxNYSS/cUs/Y5btq+YlcOIFvJG3sm51WTQPdYK0ZLDtRKVpcsq
xP/50w76CpRW6eU9ZgAVLQa24qvaS0kjPJ00papxRWPlRpTyI0JM7uY56DNDioLs
JiUH0bAq5xokvl+WcPjDATN0wuU6MZ8iHfw81R1RV9EmUe04lfExMIo8cVw8G2Av
qkuhF4bDilNikhJXWRr/6ir78ME01hCGnYpka5eAx37wuqg+6ZygMUTOg2BTOsXX
JVQ3va9pvghx4J0etFCAz2nZKPBxiWOPuUhZPD1kcv9puNvGlaX0Mf+bj7RttnqL
CC8Zalx/LFJlbY94MU8rNN5XZLknkOlEV7G37AdSb5OenRe6rfEDrCbDT0KUf8VJ
kQ/JAiIIcDw3DcpJTprVKsnr9CmINulxvP5iPGxGBLzYgpvDBA8psyx22Uc9HgMb
2fPFcq7OhMjbdQx1TePrLLT2gwkx0Xu+kvQhl6uaNMuc9GIdTOQPNfLIi9veCeca
pZ6VTZMyFckW97HPYy98QPgoG0qO+WT2LQWctuFqydGtI5gVFTtv8dGzNPKZc+Io
jaM65LMr/Oa1HOUebBKgvnT+7IJuEsriTVJj82/pz6FV9p76SZC/UvRahK0TKz0Q
6fQEpFMnKSjD84o2qVoa94p1Lw9soZebtjWBHnMZT+kgrW4XuwfRVNawznZoRM2h
9y2ih7DwnXmmnwGwALaqavVfCVHZT4xcxNkK2ctQ/BIa3NTT+mHNxf6/hAI7nDrS
DRg2GOAEhu6WuDm3WWe45+wdKiR9HbNEoQ/YPj93CTuEUb9FSwpuYziQPyHyBG4I
G9Ip2YvXNqlOpD2YGgfxAThNuzOXuhD7FGMppp4fnMrPzd2KaSGOclz5lhnJJjIH
0PI7pWLNxlRutBeCcllc063WTSQoSmNgxJci+4QHLQ+O7fiUkCopoblObwsDrXFg
NS0zbq9jQl60xUdBKM2WjG76uv0uVOzm1pR7BJUL/RZzhVXAZN97n1JvOJrpoZ8G
7xPrWcC6xZ4M4iOIX+jqDsH9eFcXrtS7lADSIaS+dD4uPMBCZGyyx+bYNkSQQbEE
hC9mYrRFoiyLxfgjWrIYx7CDzAG9gRlIYGhbXs6D0QLLnvw84B+iwAq2NzbCA+YJ
Xz1gO4yn9uAgvO9zFztQRoBxuC4SzWltHi9tezCmjehzBGAHivBYkc1StMK3b+WT
Fpjt3O/HZyP/FAu+CXnsBCECtn6Ws3I8sCpmit1nnl75LF9eJluvVt0HLU8urnCS
hGwsucMCOcNuIql15J6VYnqyn4Su3UCEywGwJ7OESgyANj34I0m3Y8MenN9JM8LB
sS/tPK/aXs+kmMZHxjo1ga7VsVLajprME6pZ2r1G8Y5+pCbz4np/Yh/a4rrYXVCa
S9RS+LJxLaD2e0VN7YN/zczywecu5iApRFJVfdye/fqzkCtpvb8Ihu9LJjfBZv3/
CgrukszS6F8a1cLjVjAfiSgkHO8oXBoWftX4D3fXbb3b/JOJLB705nvcIzKqY/5p
G95sDlAphLaRuCkcmI/nYXExPe5pf+5ZwJx7rEvOTEwcnfYsssirDIzh+9z7QA2F
Px5hcnPVyl7w2JZQTZifJP+7ZPxfXczmeYVo+F2uZzP9XrOl3DhfY/DQRuqtUVgz
1o0maThpCP4BLDhJSKbLfPAxWiTo4uHTxCzibzP3VqeEqXZ1kOuT4dm9w/Gzo/8Y
PpcWjwYVynySRAOZkFfJLZaoSD7oGw1+heu3DOHj+qBlB8JC0AekGwoBxdsqspXv
CuV/il4J/bKRlogo5Hc+OMAT04u+0OuhrXoNOCBivZayLsrb9eSqwlgFwwcw6nP3
eZdEJLZCF+hrvyktiUVU9T3MUrVl1RMCiegIC8HCusxEVA2MTbE3qOzuDP4eNmN9
SeZWLHP8Gw2QCwZK3gOvmDoxG9/SCVkHTMIgOrejWyfL48u8IKSK/g38n+PiSpir
LT2vCrT1cJD1LLs42WYkXzW2OMilMeAI5+Zc4Uz725rPYWKTl1Y4ySJ2Jyj2GpMr
yA+5I5ZAWtpI451LY5R1c+JGppHv5l5H+BIKon0rZL8XwtBUSgvgMy2zSyNAVnz2
AtI6NIys57vkpM7RkSE9ONrtIMgi7h8d7cvLn0N0rha1ogZkt5kISZZP2RyP8YCy
nlMr7qlSky3924gkQCNHzqGKDxaDgHOGk5q3MDRQl4x+5PQb4qYakuiSwuRgBVu9
1QrNX/YOIhy71ajPFBouf9QjegyxkFX9ADIzzqIaFwkZMCO41BMW3xFvhiXdq/tO
IBBIl034GeD6vU5auZLaH/V5kr4urhQUjCDsvQtuNh9mp6VFa0jYEGdGKXjz49yj
Wa864DJH0n4L9asagE0Y1rq2MZKe8eEbA/yHoMFkCUhuqynVF5eFcbjwfQ4xWpmF
QSBdpavzqI2beh/apOBalcg8K5NJp+wVl0pO7la54k/PEFPA61vcw3uq5dqA8FbS
9CkuKeccHpElnqmL/KZ1qexeJa+7wCVguzt6RvmL+CKIQfEArLLXbQ1K3NGXWpmZ
R8TRdhehxvlCjxV8ZHD5VcXD8pwZmL6iJsv35B2Ts5G2nE9wxBWaRoAZMmp02pOu
4c4HxKO00gEOjVkQKxxRmhwZo5wDnfESr7QdeGY46McWUm9GwdcjdnWYWn64KXrh
CYyKeuqGKuv8V65Fxmor/Ti5fKVn8qI4Ps5/KZZZ8dYO/5A+MAG4UiGyOaZ7k9c6
lmqMBzxuotbXP9Rn1wqxrz0iuQ+k2LXeGrdv5Wj+UB2X58f3dbobGJjf154bLURF
XGSRXY2j/KqGzG4b0pdv54NKk3r86W+ig2bPDlVxzzhyiR4A3CTbTRKg6ADBwxdL
Kb2liyvPsEjRfeyYqAVuJlAiOpS1joEw39XWbPOFvvw0LvjqhfMHz/j1sHJjFma3
S4FGUdIWGPmh8HOMuQ6AmxoQCmO+67XVjtg1QHCR/rwuyn7sCllfbBzQ1GNgN+yI
NDyqxFb7Tl4lEAk/J8jyct1WoFQPTNvIQfoSmqFfJHeIO+MWoHrDSx4YEd1dH8Ey
XSXW2x+dNRG1N6f5l0X3R4hMwGcWBA9FSuy7fCdj6urJ0q11MZGxBoGZQnOTrp/E
XN+uubrqXBZMY7oFhhdPpGXTi4bN5RNuvIi0HuSYLvQXKb6xEwi3tGpDV9jCnWq9
eBrCjeP+vaoy7sQXwS0eKPGlkOlVgk/WDt+LT6jEkBDOq2GvGXxbaThE1H3rRSEW
dHZaRKKu+VoAPZpGbjClCqhu+IFnzJ6CU0DHhJ+RSn5W3H7D+CmpQdymcCECNsqC
zYLqmoof0C1In6VBihXND39QAOhR5BA3K/mm2TR8vOvlRAnhwBo7XIroHaeGnXx9
Q3lV/TbPuS7oLZ6hV8q46prprpIIMc8UTonlr/hwOeFzx22mLSkIOo+BQ352dU7h
HKEZ23XDgiKS1dQne9OetYLYpi8BDdXzpr+46V2K6fjfudYtnJcW72s16o40++lq
Mum1D8X1m9kEwSKLtq+sTEQaamD/HIyz92ppQNy0EADa5UJbXkcYVjCA6uqmw+fI
v+6SghuCnDsWgSSnr9akdqnR1O+6ofI8X7ntj+9YOMgMQLpJqeBooevnaxhDlvrH
UnACKJw5MHbe1LnuCDzqwrbQ0KmhBNd15nkdrBGfMB1WVpcHXMJz5RsiSM9PmCUZ
ehG3p/7kMfJWE2P/TRcWagqOqIT+Pl0ATGn32k3cfNPo7S70R1adaS/DhXv1CyLi
5T+USiB3jIPFnhoAvF0en2c35aRQBcpLbT9o+a/cXWhvWtOty0yCgswgKeMEbNOR
HGexx0O7Ec6r3ygOQkx5k+UUd+Ga/h+vjOsVk4k9U/1RR5VEmCFeF91XWg6u4gok
pgF3Dr0zDWr9vyicOq3e2cO6IGUxOIjObpK90g+lp+Vqo8FAyTjP81ECuPIScswz
h1IXX+Gql0L0BlixWAvF6NiWSShx41rD0uDkLGVa1Qcye/pEguxglkKzjAqbjjXY
rrSvo6jE4HcoxgWqDuTA1xR2ZaaD6bLI9O4Hi+B7XjWfz/e6iYks6YhsO5uzYfdP
3FzI9DHWylzLaxmXRiovRgU0e/VFuUpWHPieMTVDVXiUCJq/+GzA2v5Xx3WxAtGm
59dOYq/ikoIWHr2IA941NXEkdpo0bAfmY9EX29XBgMUl9ulN9FvQrmzomozEXSEU
Wx0F+LcpoZt7KtBLyrzq+cRWFFKjKLT3SzpiGVKv69pAJc+JiBgSeDFln/IjOXJO
D1VgqRHgIYyEqnBStwYOr2a9SAVaTIMnTNPCoKSl/R4eYuffqjU9ysCr2QiurDvT
mhmdvK8gjQqzW9YJydJpm2hb/TxNZVHhhL6gDxMVuAxs2AAA/RPLv0TzxYPk8AsG
ZRrAOScqtCzRcLFMAAUFwaQXgBXFDuRg+vs3lAH1+hZZ7dtE4TioBUU8S43/5x4J
iEBFveq3QXz4gCI692Nj/96rxsXwVniVbD6EbRGItra2sgx/Or/gepzkJCxZ0WUe
T3bjZ/hh9qMMDTLuCCef2a6Fi3s0RuTHZJhcMXQRvUPam35OVJdnHV4GUQkYZO0A
OCarWGOtjuw7E5jLX3rBHzBzR4yzny4RiYWToA0NgE5ys8+cyRu1b6UCw8e0H/62
rpPHvC4OTFIVdQal5wslsbyLSiP1EX+Nw4xvKmCPRfMUbK1zivewFTKxaF+7uF5Y
Hbu85K1L8xOEw574/rihfmNI83vjwjeO49lnl8VqbEzHF/L+pW2+xRZEAlYb/258
z2wskRtpIYK5IwIHUE7c566nMY49ZgyZ8m2BK3JXpHEesvmyqPJSQqLDGgIYtmpj
zWLwMPvNs1WP8jMQaH0xFpprRmRXw+36llWu5eb6Y9JLVCSDURlxiivacP7tF007
0GQX2GTKx123MWKMhJX6gqq9x+OKcifrZNMXDqUQcpz5ct4jvNFheyx464URUpns
QI9LpQMjKzFMhe7dJvxHCawT6xderZj67VOx1JVZmu+vqxhCxIYNYEO13wD1Qg5b
67a8GTRb8Hxo74gwPelNtJ/ce/rlKNcZOJZEFr1D7nJbdev/wRjclnLxxJFXFVXA
Ah5Q9PKQPQf1WKrl9ieEzhka/OZ9ytUaosKNBNJiWTM24GGVSZb2muSvrzDDU9p8
noCCWJstG5pRBpxcc3RE6gWH8/lAwMSPkJLyEUdW9xOnEZHsKkke1+WBu/KuttHW
kBeMzuCetYXhgbROkq7j+F5Ds37R/qA9Tff4XRn7G4dx76+pRWWC39LE4thLSgBJ
oDjr9svwrrtaTeuBN8QHxxv3XKcM1UQJCOPxDUAo6nPQzGuN48ZyTt+9F+ntSVeY
4POhmXqr+TLp2yRn1XOyLXARGjwht2yrfzn+8Sbk1LIZFTfKpCkxlhzLxHLPoGqu
/KEQxaKto8aFdfFF2AZk8E2YDX35FmmZfC/PceioRiyc1Q5L90iAcXSu/Ns2fk7N
VXh0ys8xMATAXJj50Sz4eicEhMT1Qu28EpAvEI4Oi9T2GzSIizLBL/dPHvS7Fr0Y
+EywAttb6nksaVZ3SjFxqFVIVug7EzHpbZYaKXii1+XCBRVrnwI8ozud9a3PGXmi
yHrfHXDNMhhVR9X4qzsGB+xzAXpeTc71h2/Moi5t4GMOtyt3uAOgzrxiylswBAKA
iKcyxxjLgc/eKuHUZZ2w/isGpbHbgY2NJoJwmfYU4pjQVCY2rrAwPlcWhg4QpGCe
nLwd4VX7rhRe4/bnOKsOw97R9fsA6HUv+CTh/DvDoKcdHUZPUgy5HVFFivJd+i2P
j4HiYu8yltYWr/iWGDFGGMaOssNam8YT08RwjNEbUuxHa3OpcRq8zrxNnWzV8iG/
ZSqu6g5mz88xeKmwMNW7y4Y+1/2QJsKWpW92McLMfBv+4nyV01Eu+f1hlquDZ8nM
R8s1zPPp5/Tf/nLxAQT08BEEItDO7qF32j/CD21JNSgX64WBk9Dax8p+Vw62u4/Z
gs5WJsWg0LqNzy4aIqasKNcFAfPE3q6d2zMKvuAO077O1jaXLxCG08rn1ZhYkcXg
taRZ4bPT68Z76dEGZ5G6BCOkrIFOItXUDfx94p3j5tKXzNWxEH8tWwqwyNe37YFK
U75JaYq0S6cwxU3ecw34gCAU3KEz6zyFCSX3RQv4G4ziBc4Q/p+0VcSIpIbu5QU5
ozgnW4zDq0tGcrqHqkcGWan/bUagbzUNCV5gpWtUXAW+1OBwEUqjVHyhWgwnD2Eo
ZJEDSDp/1s36kl/3Tsw2Frz6Pzls1AqL+4ZT1CpcXiKJKgm2SFSpY+p3EjnBrvqr
GvDg4lvN6rGU9h974yhsnIdGyO4gW/ZDtaV/3TXKWqHsvgU3PBgpaHDet/dO1Xa5
Ol9TCQ7Gdp01lungw2T/2yddFTyNmBZkq6UD5Lc/WIcA68pppxNb8qFPqnJMtO60
Vj/XNLDIqeZ8n85JEYa6pOtMocYFZIWqB/E4VIhjGzZMuiHOMPBPFBzzlVpMSJkd
VTWmnboo+yMq4uUgFTnrIdOWI4vq0I13h5qjotUJdTX1ra51lWGniuVr2NCrG/4z
iP/9jVEwD9RNEV4TINxzzjfFuJuYh+/0rRRNUDKXIuP/b1hamQzxIgOkCOt7kMMU
Wd20FqvCi/+/nLO0abUvGA0i/l4htwwn2OztYHEggWCGGInIg6dLZJGkso6VCW3g
pOs2v8iOMfAlRco8r49JZs7fem82bqjfM4M3eVMnh9mWNC1NbQPXFgmvPeSRZES/
HamP0cUXg9k3X0plgJkHbEDjalrjnHf6+FTeyUZCDDCt85AXtFPT80OSUf28ntbB
48mo6r4Cd31SYIoezHq5E34Ifwaaij9hNKoGwCuzg1hZexe69ufDJFxWsNHeWkJ8
F/vhYGeR2BHdHcvIXyldmIJs01kNMGBBX9rFyvIgh1Vrnn5MaslYc8LXtTlnu8xE
fUkV+2R7YhETl3uE7ajscDOo4Zrr9v0sNzvgd4yx6h4VBoLRYmxwdapqkjW5bTrY
Ylq4uKEmDQ9FcSGMdNHzf2MAA2gjgV9H2wWTRbuliiITl269vdZoe78kz67VARMG
a7V04AUgeJbXNb1Jfm8VIKXmObPUhsUkmAzftbIuH/c6Dj+r4xX71BU+Jr1qeE3A
9GS/wWnzEfAkspg2GW8KGYqIMMsEhaZOA+iOyYzbDbQr/679bFkHeTfRiBkg6qGU
Vqxf3gC9jWhQWJOFlMzFA0xHLAmG79rwBWXca0WGD6W5EYYnK0RLSpJFSKsBWEAz
T8xECW2pU2qYsEpog/cKXw+TbN4IhQZ51mNyaibIb8Tm0zJJXbzjS/fgEbwuBLXv
6EfGIkZuBtKq00LjIFcSIwIzPT63C/ypgdDgCUW2+Hh6FsbrwSc5q1ZLBYCw7rPt
FoPaARZNPUxKSE0AqwFKbxw47O1OAPf8aKk0QP9SURbT+L8eTNSs7KwXNrON0PJt
e98IdWRHXQM2nyOV+2kl/DzkSBVld0TZ89B/xP1kIRgPph5FhoTAIQQUHCK7Ky4T
qcjj7MnAUz3PSu6Efol+piOg6f9R+j8vDZ7y0DGSMJT5m6y7MN6XoPDCogLkIdCu
1OIoawn6fqKUllVLARkTaMhwk25mecw6dmX6qA0WGAkXJPRG/79uZM2+3lfPzskc
U7XKNHBXA9iuHW4R2b51NIAMGraARgDaSvpBkaxFAYb1WBcMXI5diTMGYYOBKOqp
TjGh4U9kKzlDP7wqyiFigZyTx603NcVo9QOTDUolp2mRIkwvp09OUjsnt8ore90v
wTi8PcHgiiKILSuWbwiXepWY8Cx+Wf7scb4SAxQurr8zxtihEOFCvigS41XW7dWc
ORgJxWHpAWAIyqc8H9qLifpqk9vP5oStMLEL9IEYa2x/RXWo+dyswVxS+8C2vBaL
6B1EGi+oQU3oG2b1QnaQl2JBm3RfQr432s3n0tasskSAfQtgMxVGxgFCJIqLIw0R
wOyDnhIlN9RnogBhWPcshVk/LuaMHfZN1vqcqCzMphasLeTJrCqLflWKSXAZ4tFv
K76EjRy5n1xqb7WrGez3EvM/ZlSnJoaxE7/oV6gc1B8xnI+xXLycSfTHhheMYr//
zA5TH2MP0hAeeofhe827sztc/bfBnNlJqpmSi6sDdxk0G4/R1T4QW37dVoH0ilhO
b/tyyGDelmnx6pAU7pq9oqxyjTGi8Wbs9UHgchBBC7vha+CGkJxZvmlG5D697Fyx
8jJCSBZyJLkhdYlexoUApOOMtma7dQPeIx6FOduySa0=
`pragma protect end_protected
