// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1COpwNHueGGQjlnD8Lq2Z42OiG8V6iw7PH2djvoLT29LuDnxKnAq/FD5CI8nAs8tdG5RqX9VF4Ti
WPWtLp+Qdnr1WiZR643a5GeQ7j/4BYfbS78y6fNOW/HUptKBwAuR97BlCWr0/ZCIKAhMNYZjr1Fa
rBsAiDHadeIRSHoBC2Fj9VAm+RSdtm7QgcI7MID1dpSlOBSGiC9301a03QcRREvhQ3V8G7NKLIy5
pdhVbIQvFlH38N/W94o1UrM7uze/vG1HyxNrfCQmarrd3B8zOYVixbnQYY6iFKnnrpOhWM42qzoJ
zNaiH5WSlpo7TGsLNxu/ZAbwFuuoARwttSO+YQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 25104)
gys0RZjw7TceZekVyqSYjmPpjn4VIhNGRDkq/MM4oVBbf5XeeQBlWrlCWroV/T5fjmuHTL8g267Y
Mmhv9CmkKLJcgiJ8ws99j/sOqEP84Zd4aRY80mDdcfEAp7E17yF8qbX5JJ9+ZA7Ma3KcUQNE0Lnm
myH9IKTP0lvPi0aI2/dFZqK5ngsic32zyfTAwhCwr6wlodsH6iwdopUkjAXKPDYLWKtgnTPhx+N4
sc3sr2rwwaZz7EeDnEbWQJWE3/pihBcJAJ9+hIWWudqcqDhsrUaI7k6M8T1QyIXHPx9Uc0dmwhTP
riX38Haf3oQBFUYB+ZHDOAsX9xGY9J0WeeZSoVHHaz1pBlROEtbQZw6rwWyQP9DPe5g/37UmcygJ
rZtVmfo3CDV9ng5Je3bB1yc84SWe1CKv7e/VirWDq3aaT7F44pdVY2nB/qyp+Qmx32mRBWv/kAJ+
P2fyQXyHLlg3n2aMm/oSbRgtKFMJIMYmCGSEhA5IejZmlUKECbudZ57i7H++ntu7d9D1IDZ/9/G7
wRhiW/RgMIe8DBLufPp6QPoRLpsPWYq32iO/t5mc28iLPTRiI4TQS7G40HsW0tBWBXtuRbRkJDDQ
vq62IOGBUrMEkg6uEQG0dv7Kb1pbDrfO1rlunK5rFNydpiU20crnxt0HemZQkGaCsqA5iKFntd9Y
uWIbY1FDzG8fCvOiQVXmoIbUjfSXpKCvJwTINAKGj6h2/bG8yuC3te4ezXbYEH4pLViv3npV9OUH
s3OrUnS7Inizm32FUIHTgMrUeX/TuWUxecL6/+HlBQ+vWJ9aRXvAVSFG+Q1tsvDgjMApbNYTYkwF
3rsebpROUcOPdmQS7Ju4iIGglvSd93ct6I1Dp3+7IGcPC8mXvyFuHgUsCFCrsUrDeJH2EnJcmguT
KDLyufYNenGeiQxBJQlqZs666Ps77IJr3qYS+EkIXI/o1bugauMEME+i0O8NIGucAUKQVFawI1uD
7Nwr/zAS1P/c7thfwoQVzodYwYPprBhWcOwIya9VeH3stIQUqe3jWy6DWblQW/bgvTp1vs3RrEdX
p3KqhosfREf0A3GPodu/Bjmu2G5ISWONzVxXQ9v+NDdUmnVMumciMeddhH1/FLtegkA/JznyU4iO
z9YqhbxIOTQXc8zbbvXlMIDiQVimfWZHY6Wj/elCbvfT+x8QJe57rUxR44Iawy3zMrJb7Sm1H+TC
WKyj9aIEzmtklfTjQzPKVu2VaUXLJ2KSyDkDsCjWQ9bWmmepnDizoNoH6YCZADKqleY58uqFB6Qf
PZrE04Vaeh7XAQHHm1ZqY8NOqrCKkQHd+0nowbxnMBtqFqe7OKhO1CZ/heuM6gu/wShp3hgKXvAy
xuXI6zAMxukjoY8yx4/saNRXBjXluUPkN5rJt0R8plavW8QUAYkV0mKenGL87UE7xn8bGMv7k0iM
XNMrLs4hQM2aAqqYiFhxLTvHHTKABRurivZl31bMIeSUvmt8YGqXm17usWtJMYlaaNm0htzgPHrA
5Si3yyWoZp8w6uu4TSrHhx4rE/9OZszlQAMkjO5rjS+G1Voygw9oPlEUdick53korjpTOMCaIgww
MVjmyYOX9bJOkDiFEADiAUz13I4jAzcAnKyPtCTgElIkHPZcGw1jgwi9/A1UYGzJ/CAPnuqlElkH
l9aRkf5zcu0Qo6EB0OPWzt98fDGJUs0jAWnuoEsESN8y+GZvJybxh2H0TcPHmem1fLcfQvZiRtGX
ULXmd4JOqY1QF8hEUp+vY4QbalrMFH8TQBR26A8DvfysPX/C/DV6ty2X9nn/lYe6lZWuh3nM0zko
KTtMqvdiOCuoRWsFse9bB16hCeC++yPbe/Wl7oj+DXn1mq7dzm3zlOqHhTIZDq5WFVRzH5nE7DRP
hXbsWGjyP9pH7g5Q2baLN9inZkJt4vtHkJnreFQBfmngvNBhDlE5wqnjHkjp02CgwoB7ERhRbeX+
TsS4Dt+yYY75PAs1156mfqB3/R0Ygy6e9jI88zsWcL8zh2EodQmNcs6t+E3afbIBiDHD6U7b5DH4
fbIFarkeRMsoGEnrHoX7UDGq4Vc05mrmdFOqF9vkwXca4jE1ED2cv8k+ErLoFOET4edtTVozBeR5
DseJp4gD6kRZiagSH0WiyPh0VRDojkQjgfH0u2GG0ZY//sb31u2prsN3F0+Ad9fWaEuP8XYP4saO
5Pyk3NsGFcwFGmKIHW51vCCQ+q5HukeWycyPn3yZSYxNjdEbGNh0R57/LfuDJhRi8LydOxz1Y/xh
pKYuodrK3dQJOuOXlRWh/nvW4UGVnFpTSEbJ3PhkWjrJ6oy6WynhD3HaZgoZ33DzuM6VIdvZJcbe
3GnQHfkPmZvmqaq5UIrOX6fo71mZPOoiXs8kYpPsrHGLEyYU8nO+NEcUAn45lGl2XGJFLfXWIghj
pOp20awDpGZqN6p/OFnsH2j2cTEkUvKPDNA2qxRndbjOhnlIzx+o8V3ZyS1pGKRjrXo9myT8hexN
XKPQ3dPvZuvr+RS/sJpb+Nb6axCbB7oxVXzqLwP3efQbfsIhQznltwb4EZ8KfL0jodQREKyumqti
b9zTU7q80bwZXTTpHmFcaZ8jLJcypr8i7KTU8oksubXqbDyqdK4xUd+nmQwyquXVkbnvQe8AL6QP
FIlZtL738kZ+I4BioJeYII0XPkMgTw1al09UwVmDdszRDb0aGgwQVx1Td6TxHcKATXLAxL+gGH9D
+ioM3TRsZEnXMyFfAsqrxBVpmNdtjMqoJZ8iTaOZ9NGoQWOzGlajXtxLsX9LAuGp+LkWUzpvMHGf
aBv1j+uhgFgCVKo8SPhCakMcuBu9n3qPgK/0D1l9xWHPB82GRYf0ecR7BBStD2qsTqn0pXN5ObzG
TstMpziuZYKHEAtFZS0EVpY6mpewG3lsyWKr8V1E6UQTH24BVT8EnE3dEKQLGnADP7EJupGvr36x
Ck213yJ7LNMufkOTXhXPw+eeOAugHFAjfHP+f+9HH4oyFCWdcjAyxYvHtsSCZwZmVjR3SphO21Jp
4xq5Q/8llSQ6Uh1qm1sh+QUaY/LizsrzAJ9CrVJPVXf5HZzbkcphaERWV/XYIhJHRdKAGsEqApci
UG6n7l+zg6vJV5VMnyR3LAplP4igm0n/MElgJRxLlYEmre7B5T06SSKAjBp2ufndNFno2N4PfH6c
0uioec6iFEBndKAsVzOnezj13kRALi80yTDg45PwM3y1I+7RW1YMWF3SH1vC3oy1jXGO8pU+rfqV
MZkQfb7kjYzPndlvLr3cScqzI2wyJJgl4k7u5qo56SRtXYMHHrhGFiH6+/7UIjOjtJm37fDP0105
5cb6hqthP3fAZ66Sm/oOAGVKaPq8RkZ8cCibUvwaNibkN8SpD+W5DUyquvKR3iXwE0OTSEv4cCVt
iDuznG/jLF3trzX1iW7HOMKqgAkwf0PGOq3YLRmsVNbv/pHIopeHvA2ItDkI/HFuJ7OAbivHbWeT
3/+DGpfiGOnKEYZVKlYnVTZI1WBqVWepXYLupchnUxlvPShFniBwHzZJGDYsDPlYNPO/GTYUTR56
uDogDhu2Y2FSPP5aNJCqgJ9RBZN4kyWP8GFCK4YWa8VKM8x7uHJqKu+3DukYst9g/Xc/ZXoqc5/o
fR+LmmX7N4RmGPRdluwZcnooXXgQ6N2TJYk2eZYXc8CTr0KemjvEmiwRSYQvLj4iXJ/z6ZfOQg01
NOG6E7PIya+UaINRx/jGazE45vyrGf+UGuOmyCX/IOgndVgMezLrtFKKeNyLmz4Q34Fi0sTE9Z35
sTlAMq6FWqj/uWYOMPrar2u5RctUR7duF4XwbtpyQPJTv880F0Q3PXNBrb78suPIeOO4KKHvJ7TZ
hb0RVu8BQvpJE3jfc39JJpVkQ37EiDsL0U/Rlvg86Fa8MMjaVHWEsOI3QOE+rrZWanipzOS4RWUm
uTytTgHgZ854URAX16IiaLk3+I/VISBblmZDN7Ga3tZiQQRjK22+h0due7HEAZBzkCmYPAgRH00A
ZJlyB8PYXWSvcoLRz6FcSHPhTwtcSd0BGiSlvvyNvsk6nW9GfdSH/4HjG+NUQo5ZYgzGwcUWLcwq
k9+w0kf4MNc3i6tw9wQsJLleXHe4UlNLqK8vvDaWJO170J3aR53ruZ97cCRjfCw4AXNdsfA+SJCS
87DJqsM/5vfcS1/mkHFBkvRFU69mT124bEVxtWMD6OOGuMDXHbFNg0pCnzxTIU6z0G7P3+uFmPDG
Sok3BuvLl3iey4Xa9O7NbilMCQJtycY5pc1ELfMnQDSWDbsyjv1sCYaMWUBT20F1M0ktKn2yOfDR
aFgBcJUVBFiSqXTkO9wVMiizNq191f5NZKj9mgP8SVtZzm8xbX9HSw6s9L8MyqU5urLb4qZja5gD
EdsoY89TDBc5vb2K/bfz71eRFHiOGo0FShc4OTSGh+KkBlA1M6eKc5Fpsbo2B/lis7GbBAg8CSLg
nZT86a9HPCMcwOijU7L4HxLuFJyndYarHATFMVBt5A/j46ok255u2Zgy5swfiZq8GyatVwjwEgqu
CQIGmo401gx9TtzM083PIGSOfebyFYA376VBsXH7e49fcjwFMoWXZ7HDSv6EaAuwgrkWJl18tcuS
exmyK+7KXwY6jQKKhQU8xwfkY5lPQHgXEPXTQYsT8AEQhG5eMkFleTbUZ3PhySBLeS8zCBOMMJQu
0O8U838ySivuYinpyGyXJKglOGYPzUi5VCFuTP5FWsUWR3uc+hGR+FjyUXAnTn3V2GCdbn33SENq
m+wMmbFaxVvns56/4CxlUWz/9w5kQXFoWUsBYRST89d6uoQYmZcX3Dx7pU/7pCCLJossinCKp/NY
twUkBVOfWRCHXOSpC7ntJGPzJer8sLm0euYjEexKJzeYIk8zUKmm/AWhydEuRtRGu2ZpDLJwfShp
XLAAGJU/YcbQWqdtfXnzaS3dssUH3QWwH6KQ3oR3rMNeD44uXG41Jmd+W3AzWRd+iBM6+/v2LjDp
vTMysoTsaxtSbQvW+bYgjNUMdp8aBrIzdl5mF1+jTpmd9lw7RAWptJjVB/TPxh3M/lCit4jRugtM
bJtEbprCSGYDqoN6LoIk5thy/+JeLiVHk0MexgNJ0d1njvUEmKM01/h6/wMHtjGfH+8a/w6m7Wem
c0PP0ZHuEGoCyaM2FTnZszjxU3R49sxOp7mMST1eW5o9gIgzXYJgK6D20QONQVtzHhpWyTIdG0LJ
KrB353+4P/mGJEhxd2XScFCZ284kLn/1golM+pXMB/rF5MG84hxQhq3B3wEAlkyOw1QAediKvEvG
ZUXYr95HEE7CEoy53UsvtoAWhwwlDcmfzflkwriphdlPxGAMk7I9asmOZLHn7uutJCpYw2NU2MIb
HMqrrS4hGei5cTfTQ0sfGS5rZ0qWIC2MN+SW4jwgRM8TJ8Cs3+I1HDIsmp1WQ3wH1DzvOkNeXWzk
blE3nlbW95m0/BlWLfMjeVQ2J+azsYjL65szwBuE7S75hu28fmtnj4p+vCrSMFCafhtRa7KOSJZ4
ivCBrjf8aSoVyG7+N9LX/KvxciAJbC6tvuEx4Xkej7jmAGn9aDykRh4cxC45FWzZSHq4u2MQIhFf
jwal7YUEvSlx/fE4sg7yqPy6NZtztlDkeic9wbC7nTEDUnRAoMqLMLo/T5SSpc3AAJbmJWSa30B1
OtbH0gT7j8oMFS3pfEHHrmV8SzF3IqElF1QPddSLpPn8n35Orjjsh6yJlar8ligPesQ2WWZXao8q
zcbbaFByV0lr4LZOSRdApry1MWeQIYjTbhBFK/vHofLyn+t40uVEzt+WKUJ1nPE5m+vg0LwnjEJP
dmK7DV9yiWlM3Qf7FpX/NIc9ZFsdi0TENKNmbyIUIi58vj43hH5DyHFepKsdKvKGIgd17mU1yNL4
6wnQGXjFfoxur2e0nEE0FdYZz6pnO1X6r66tMjXTANmzPSWKixFsZFJn+tvJca6aEIGyGB5x55Ul
g1Au1xYx+nryGuS8szTsHXbO9Lwu+ZFlaTIVl3Bjd8CQYLP90C1/c2N/kOBH3gbq+GBYvoau84Rb
ezBkQaC589YEmb09JtKltFcNIlMwVNlIl7AImywmyAPDkQ27ddw0PXWSKYQicb2Hb8BzrPIaNQtR
bl/M93F5VXVRoBEDUPgrE57eGrGH6+wvTcfaOBzxsJEZnfkC/IyA1K9rTEDYZl0X/1JuK/XM8eEu
KjKLBbR9ujIrPlfR5M2LiItPp8mpfP5+0hdBevxDQx4BJ26nIIxfVnHFyHSm9xUOyBWerijDVO5A
tuwoBAtmwxqzSJFhtvfM2A6/zlzEbo+4eKJd5U20XzsOGQLz48LjoB7yZ4MFksizMqbfvXq+371E
0GREyNntJgS70lQCU9Z8+YN7075nDNbSKdoiL87WdcPTiT13l+TAq1b+OllW8qrj4htBPRxsiQe1
HmIfFWZYh0Ld7q0Ybw57k/rtvsuNWKffDaqnIPUacDHtjwDd+PDPXbmdATEdfM599cI9AQGx1ID0
qqVuEwny4XZhYAWjy4x3PQAtUR2vLjCjABsPz9WjWVFF6M2cW4kCPViiLcfxct+5ShuzvfDQ1qBc
2Mm2v0yCn7zkCHLBD6R2zIC8SZGUE+oUH8rUYNIThxTXnlmaBdoafq6sNxocAaZrQJkCAVkW3kCf
NCh8oft8Y8oemVYo5SudVoWnp0BKVbkThZ6arTWJvvjPOP5K9rAFYeK9CuzbqWwZG0reCAulyLrj
CzbMbTHlxemvJ7wtEjllNfxgSiwmGzZdqrjHaDttEH0/MuVx8zM5s6AhDpySjM520tXnvLzdVP+I
TY0k/clQUpfQYHET7+n+Nk93GJFrKlgm27n/2sdIuEl6MH0mzp9NOv8YjqsDTLeSGfJlRfhVdTRY
9QUSxtc6RN9f72KMn8/KY3m+fgZ+LD9MuVqHq/WmysVIiqxKzu9puIZhkVbFOpMlFX6m30uaGKNa
xTJXehjmqz/LMKs6CeYTOqGVlDIcsKjFVjHNNtSdFnqfroldfNtuKn/sogVp0gUCjl/cY1IIxpAZ
dxpGEAGZh+41AIbyyHj1O6qFtUYJWrOoEQY6w9u8XGCiy4QQk72CSzEqa+VI26nLXSnNMpgr/z+6
03xrLmWkQZZSpujFCn1IfuO929xqSzLcM/yU0W++rsZjc+JExMlnK5GGp21skbV76DevURXsfrAw
MaX7pWxN5yaJG9/p2TuRG5mgamYLzc3sSAyVqnoOs6W/zHVzZjaOlAOK3rYgGRK37tSiYOxuBM42
eJR/WUkUgwDqovgamyQmwHKjhvvKULDKmJFNz7ShPAz2EdnKx2y/GFXvuRazRX83ts59C0NPrhpl
bIWMEQQx+mlYwvsf5VLbZm6Mzp5jDwvcWFxXbFmQU5hqqJS5QdGZfGSCXYCO2C7DnaP3IV8wjfog
bBrFqQL6UogS3QyNlhP1hknsq+j36qbZTvH6qBJAXHKzmIGeIDzxizSMW4fqGfENLCHAMVUbJ2Dh
a8gzBhVaoqGN/GBPFjMI44h82pL4COAIgYGr7Qe/pTjScDNg9dA6oVmb0hVSA5cZ23IB32fDdq9W
a+qsRnzEHYzorai8vcoNz/oLQFUfKjIdTMHx+JquswFgD4k2kWQ9wC8xtTAvkHAEdwsuTXpT9CN+
aCfWM1rZn+RXD9OnHDGZW9lZiC5aEZYbKwaBBPaURqyFtDz2r+urHo7lPiCgsxgwsnbvYrUj6Z2J
tAHzjlOeoTq5PkaaWYi4HfBwf49oWW9sJr6PKmEGWdx3a4gu0X25gfvIdDdiixmlD5JEP5jUPmuk
nkd+pa1/w0GokoaysfbOqietkr2debXrUNQRtuJAcjWu70fz4INdsI1SsOYnq2mWuHKGK0PiTCBl
xRpWRiOyoeMwlz+euHJlgiPE5bxesU6hQan0nAt4jlNbuVdM8UieL5VAaW2BwLFVdi6uwaQ49w0K
6+ecWWy2CkI9eT9+PdB5TKUjECQvoYHagFBcj2C7jvGNiQwZvDfu0+LNuTRXKMtqRvmHpa7fQGvX
m70FKxvfrfzgINys8QUtCtAMjTbHyl+bWESs5FnChdrtpwlhYUavCJDi3HzXPc4IG/JOoY8yCVk/
n1oxV9xaAKTnpjXOfro6IgRoH/JcHSD0jAIz+kzNohBX1tFmtlBMUpRqRz3qkA7+SZu5oEFLhPXE
aL/Vv3gHMqIkLu4QHLGlUrTrSn1skba3J7Le7bGEingUzjA0mfTW7yMq9HEZqa6+3/s30nRuFqp9
Hs7b4xxoE+Hq27tPD6T5uGgEC1XuvxNRWHiQ54fje5WXlmuLVVZ892XVFRgZqrGEks/n2D3fBxqQ
d+Ssh6bzWbCqnzgWQkHn620kwR4nDRCqtbEHWaLDJJNI8A6egRteWe2gRoGk/FSq1vvABND9QTh0
ebcjzihLnzlL20GXKm+wFD2gq+iqwwhlqpyu9c89IS+GHMqz5Fg6JvPF6vxLDzrdYq2bsOS4frFk
+oOBo5yfRowf/FQls9G4TSjFKddwPVeOaeZ3r4ijv0r1ko0f/qi2GccQf4tgR60MqzHBdbH2IpKn
k5LVWb/ItZMisJhpJkhXaa25PDmnYiMlntEEZlyh1DzxukPUUB6Ep076uQoOUf6+9nMKZVOF0kIt
I5Y6p+r3PP6OKBqzeREIjSo7m4rgbSsx7bvTd95fLqaKrSloOtxkFVwBk3ES9LQ+nNg9sjgvDyez
60fuNMiguGM4yn6MLM5RkVaBsVWuB+mFCeft7UIovBq3Q82Y6Na7RoNMBTZlcFdX22K5weKL3TFd
voTWJciEhzMXVGHqn/7n8bNVGScUI6tczIjmfUbM0tYNxcdPcK6gzR4nkNAuDJFczNDHJ2R4j0AD
fHwDczr4hcEOrsfV21v+rSPQEzQ1gDnhB9moII6NlMw+KIrIyzCz4aRd7a8xtf4qSAjBFTH/P8qV
Z3NWMknfGxVuL0KkYfgfolKL3G93oIuQ2+00CMcTIVqgsNQOIdKuanPR0HhE5b88GQjLbVrOUdUn
1KedR28JCMuXyvTkZZW7+3DyIZCVPq/FiWw9N52prHp+gkt87DfAdZPMb1xlTojXb6OpRcaq3XaL
AuJouV3uxaq/bzSj6rEfmzaSvTpPFB94cCNB+22Z/v4dYnnzv9jJ5g7zUn+Vl/O9e1+XRbMUszlR
vjidVFsNv9E2JR7B9GtyELfHmkjh2yJrfAXNm9E0k5x+Jr0RFwjjVqw+VmgoxMjnG7XYoDP2Iakk
FFZRO6XHsVJCLLEEBii8zpeRYhxBN6cEMZ0TDyRHbZGSXUX2eUIGfFi2D48E0ParCCOuG5XsOa1Q
luOlZbLkOB5V8vImPY2uPRCG6B9lkojsZugdzjLTS2+rcBQDZ54L3SSaJMbbyBTvjWZvs5byTeO5
kNc/gR8bZ0wXZJUQkssZAWIB3odirhedHzxmKvs0UuCW4P6PbHh1bpRRCWDoiysPBUMgQzsNYXQE
86wn0lw7dFuf1QAG/8DB/FKh2K1bATwOa2X4WRU1OMQMsxmG7Xoh443XQ6UJzsyzbkeQh9Ttw++a
jUrUjDPqCbvQ3UPneQWAgBxrAbXAzi75ifacEZCf17NG6j18UT/+52GC/a475b9xVrbMzbVJWjUs
ykPHdqZU/2b11ySbPcSVT2o4CTE+qYcf3gs0PzKDi/s/J8iS9t4YS3pVWHcHDVkja/CYNa5F4I0H
slyCpruON5WTdbrOt0QP8iP6QCiXuZ7N2lRlhirm+ymxNPM9jBF/T+NX1zjTswIY+tCzM3LYyTZr
JL8777oThRXndvkhQugtZyIv63yENQNXeLmbHTXzk+YmLTvrSnNS7x16fyJ00vYIICRn/PrOoXK4
jyD8vJdMonJ/9RBnsp0bcOUGpQJTqLNgaTFwN/HJx7FAE9WksSXa9tbdJ7eOxDJJqETBYEbCi/Yf
lK+JvcwQiAXvaikOurkqGLvu6aCRY/cEJcLuFGmbiqXDpQj+13wa3ajdynFONVPAMgWOBz6HPGTg
40MbjCQwraIhPUa5f4EYoOGp8GybQ00lL7+MprbhZIwvxd+7Pdf+VlOtbbDuhe+P6OhHZuEWprc4
mJFYzm9x2pWcb0PH3ZJj4CWiLfAaJ785ZWluG8pBKNN+IEQGOdJTey2B9MF5ogaWvvK5c+V37HUH
zEW57jhh+ga3rHpgxyNKIJBIRhvYhA8SKr2jlWVzS10nYRgmvY2r5GE6CLTjis7iNTEEXcWpuWF7
FqRUap+6Gzhnh7L1C8mgNyTV4m0/OGO4j0oOdj+rvQ9S16l9XcdBARlnKTC8RnS7Mh4c0c/SE/xT
TWJssCnGOGFBXth0FKLEKcJ6657O+h5XxZFvrYKKHneeyUGCsA80vdk8bdLloCqaCh5bws8UX6YY
2ZUBd88sOaPT2qgUQcT05xWGv346AnYLLXSp35WLe9lGjneWuisxb8od80E+jTjQGi5zf6XQRbat
BXXnB2i9ONq9EQaDxxFnFLtOWO5rccGDj44fwOFMXsgBv9wqcJCSonNarY8SCmFvfvTiyc0MLGNv
Mzt8RPkkFkp8F8Cdx/qro0svmHeYEEQxM+3CLJCkmjWqSdqaIKwBVnXFI5u+LHEwGZdX76P9S7nf
wcfOiIkKla8tYp/9Js/GQjgkQu3b2xci3TFyax2cCWgVOTVNiyNEqRRDix0DL9UYB54pxuo8zQM6
RDauzFXcZMpGtTE2n/0Xr/oqybQcS0yc8WkZoeweCoPQ4lZWKirgJuwx+7kAMmq3GsbaGXSDWGX9
a9WmkgnqScltaDvlJLqck3nlb6p+bwZPIT1QQ8fk54p2lra6VC8f0A7sgtu8iZlZ8vl1VHua+6wR
u2d6Z289QPz0iPbMV6XLgUUF7aHErzNikky/3Zpz2QpK8jP28ttQlUg/hR1414HM+h6gvRN5pXtv
EAMcNFfuHHZvqgVjHNZu56je1AkI5HKdfIg1W1gZSAIK41/1PnpD9+Y0jnY16F57wy0FDiTQzWKi
MRnSaiw9oXkvoay3Lt5C1hKfcNUA6TYU6Rfi7Wh/xNGJBR65+uZ6wziK39IaRnL0Prm1eQcB/M0y
0c9tMJgHBHVMBLiygmy331BzKvgmBzRpGnAMfbOb9TPjkk8pU5acxBT9br4psZpo8c0F6jnWnznZ
mE9jTyuclEp+qMrg/Tjfjogjbp1JpJtThLacVkQoX5xiTtFDGJiH5iunwLN2MJRnjzyZfqOfTH2d
lbQWVDgj+gdM3owZhMv4QQOBkbW8UQnDBDNAnPArOJ99u2ql2OESSy44F5VrVEBsqU84xFPFtJE/
04HH+5Axh4TSIdlM2m1A1cLG1gvDnbEpJWIOGwVHPGatjsbo67IhhPVlyr0a2jGZS+NYc4jfUPuF
jH70PxOzGmpg7QEuWWVhf1vZSNlcQkhAt8cIMgwk5fZUVjjnu41LKQKkSVmwrwFv3J1QYrr23sy3
raXoKviwEMr1B5FNwJFSyeC4zHN1NM1uCQDEUrtNGy5eh68VAOhHMh5nr4vfl7brK4OslqLuBtTm
40sPuaCHqOCdovNa7eoj4ppEghAVfpSP87o+GEhKz0NZjV9zxEZb9/pTZoJVBcrXO+JOsa9jTaSz
keVz9VnRGAvQ5TQwbDGmzvpS5N+VBjvdphJIb76mKRe+1LKHMJh7sJZLwIQ4ueMaQYpYVuq5Mocv
yc9nrSQPltPW+EVPXChKsbtYgzCKIQd5DpMf/og5ofYvu4+FZQyYZK2KD3bh07pzoXO0gnk6NugW
TWXKRn/D2EuWMEgWWxGjW9sEHq4pZ/hqUeIaa4USyC6JfhTLISW7XcxHRncCXJTMPo4E/0lwbt0V
ckEZYJHcAEBvvg8jSBzubtb1eCGjNH2QU09F8Vue4vnI3Ep7XUIGwbJ9yJoTZ/Uat+LFFl2q0kOg
bUCLfgN/iawMZuaxvGIHtDCZJxJ5LK66BpLM6J1UaXxVEqEXryEII7u2JCS7WaSdeMVShYTPEGyu
i1L0B0qrE+BPAaPOxwrBo1EfEiyQG/0mQ03d54ot5yyC/zCV6b7iRPQ9L2F7Ic808NqswWLshMpK
GLFGkLiWReVMng/xvfUKQOUJkzqAtjE0Wjyum5RhDk7SS5NGblhngmod+eI37RUlPOUhfLqtWaMf
yQsqSs5v/tF39ipsFNuj6gsLm8/4muEo9Srez80yqgnBIZhZyCELSSjJEIg9/+v3Ts/kuuO/XExR
SrQt6ZRosR0KtTFic1lQ/jbE0O9bR9ijTNMhfbALONlV60hFlHFlfQVYVPhxugnwIp8toNIffRqm
ahUlQncijcZio5Ss/xSzAF3TpZUPLwq39ZKg6lY08L9UjVw0TzupNR82thMpeT/vGAnqZourGr5s
A/TbetO/N4ffu+j5TSPpJZ/9yPrIJaCOIrDv7y5jQ/twi0ygoQh3KnglH/YcPpqLy9o0vFCe1p3e
8GYr45lD3PeLF4bTBD9QsW+SKhuO+qiHmtwqnWxssFlTIcVzNolHED2vciq5YgBVnOH/c8xjG1BU
3AWZvl3lPQMi1cPXUhNTydY8GIn1hmchpmrW373v9WMELr5lFj0Of4cBH1wxIKmnwR+AUduGO/PP
rXL8b7ZyDk6U6j98iyOJsSmR3Yp8kXxZvGrFtYJSxu+7cfcuWF5pJFFQ5T2uewCtJAKjfdPyybRr
oCoFSjbpMM4Von/xiSGUU1pThMwO0N4QQt3JfnT0iO/ZyMFEgTxkQnS6ysPKQ+jhmmZK+wARHos9
cTd4VSXjIusjSlJ5NUlUjvFeNaY0V1go4uQn6QOdQgfMk8qNGSckE3HUPYbVcySIJFLNw4uctimL
kkwm/xqtoC/HmN6+y5UceNtydAp747u3GiMJ+OphbXa4T+LT4dVZfAViD1tvbk9Yju3g/fK0FT4b
09stLyqhmxfYL8oFw0CiKhh4UDSmLEubghD5NnJu4q51d+2Ov6Lo52IYY7KB1ohkFD6f2x7AJ+4F
U8tvzqkpTs0b/9dhp3aHOb9wq2isP27TwWzpnqGUi+7ih5KzecXIMh5NsmnGvexOhZca7xW2Onig
WJa0MB5pdbbfzhVGZ9aqJphfl9iddFI+dXz2r0dXszRGKvS5sTreg4uH/NTgQtF2XzkoDUkKHsYx
sT3Aazzxbz5k3l5BNV18CiXkJPTk3HOAnPqVKYHcxnZmJHHVypchydmmN0aOHWjo4tI3H/QBB0UH
v3UapcXo7LLmIJJ/Kk4ub4NN235sap2BmGKTWXhjZSbYCzcrDMQR87vwMiiGcsUu2TVhQgJGFgFH
KbruzAGsastgfZFGv9TqTcjCgXSIPpUwh3op6bM36FrHZoE56JGvTRcYztyHKqcBaApvck0eD2Wx
tfMC7Okc4freKXZz3m2kuLSMRJiys6htoNWQQ49n+d/VQ1G8oJuW7eyL3HmPABsgk644YcJPbq3F
pYl5qb16WciQLOl4IEuPUVYpVkYDbI6EOYAylA8taFxOWo/KNiIbMOmEVq2dGmzaBKdpSQcmn26B
Vs9yOUwW1xfNb2A1WAbDuM9dpUc8IOrgr+7zKB38GD9koHx4hDMAPoTgSX2zTkhh4jMyQrn/w8p0
XRGcxe/bWyPSoljLzE9HGIdmIGWJAyAAQ1BJfaQIaFlviThuUQKl4VAQ5I/h+Mv4ncA8kaq9MQ2+
YnmtB1zVW6oprBundHdkJXQfA4BsFMM0uXkp2rgVK3ZslnDIc8gTi4hsHRvb0+jIvorESpmylJ40
Tgur7t9xNui7HyqWEP7J2icp2kCW74IfnZb49oq/jhO550ypmWoJ4N4Ci8QHUZCe9YTfOZdCD/vS
O6frijsdBHG9lxpU4mGGJN5Qwytc91FZd1kv7uw524T6Zbb0/uDSAWBaWQO7Qig4thrNVd+X/iqB
/fpaVPEYulo/+HK2K8QJBS9tpF3o14WCBfV2UPJ88Dks0rZtr0hUsxi5KLvdKgPY/h8AdZhJ1gfq
eu1IF8LWTmMq1jlt6fm+ZkcQhPg1DTe+qyvUvLOf4GNE/rWSjsPKOHeVp5At1UAUSaGeeo1mtnZ5
oKWjfNfF36D9Pv4pT4cXyqLXHQyHgj/1rttTxi24uvG/WAtFPHSppSB/vlTC+viZV98uGol/VMyZ
YZxfRsyuI3wXTX7euK6fPP/7CYr+Y3qF3Ql6aOcc/A4z1zWHe0xTCk2w7ve22BOsOuSghSjXdQ+W
djtyc0zgzblCrhPCB/GROI7R5DETgcg74fXjfEAtAl9hDLuBr5luKk6V4IFZ4VRFQ8vcaHWK/tZW
qtCyHUbpex8TR8LaEvVQwgLRk5Z46E5VSPraufoIrCCp6AIPEbdedYzL6mpzUN6Oxwkl8Um/e9Kw
kO5CdLmUL/cZn/wG/po12SOWA4tmB2mj15IJ0PmrJ/FfldxHvXZ11J98Z8lPXoymMG7IPPN+Tc/L
EKMmEwe1F1I2/5Zcnw+rdsModCoaAcSnRSNFtNMB0GiLpFs7JRHhnRQsQGrl1QwQkMySBO8Fo2LG
3JIDioua/QExIZhFIR2omb+QnS97kG4F4K4GWbnJhByMr+9mULP3yX2iresz0ULyILWC1LHvOikR
U9FB4ltx5m2toDW7yW+iEdiytPFnq2vZ+4Zh4Y+qjhz9/eLa5YVmlG1bbNFc9hsKqGyHIizk+BQ+
ZsDzCexQzcSVtMA32sl0Ifp07rJyLbvly7ePYngrbeEjEjO0Wo5BMBSbCDYI7hjyob2m2h+6tK5N
YYtPxxblHUF2RbKxKSPSTAFNwHNYsizs/XD99Asz7+4AJ7W5rspwqqLOVSAoc52bx6krfu4WUW9u
fw2l4td1UWlIfIypwaZxlbKmrBsAjTHxzAcHlKBwmWYPGRntnLmK4SXKNlt9qf3erPAAO8juDRYr
wc9IApqI3V23btyaMlywXZtOziW0N/bzO1Cjktn6wjgQO38ZFGqYK7KoAj0lgujEu0WFHV0LEguQ
4W30jOzhzAh9GpKaB8LgcxChdFikuKJglGJFGF3ctzUxwQl9cDh8oQYlLtk3taMAMWYyTwaRBhhF
hAhTqH7pRkps8XmPtpS5C2eio7AVOptUe11sqeCB8/1NiObtDyGkRyvJFq4IfkaUV5NWWfvNta1A
WMEOSU6q8+G7Wb11zszedfknwTSdU9XlWW9Mbtne/ouklwunBLEfbyFJxf27sPpUawgcSlfe1Nyc
efSesodSNAOSubIJYkGAzhRhlYaU6g7Cr3fwXuwOdVczwqCKKlwE2sqHwAVBG7j1WdPfKZTYkVlE
mwdi7yUyZZq0y1JbEZ3ZZWRVLwVnKQf5i/HIOcgmyM21eisD4H9RuF9uN6zR1jbjgeAaspcfR6SI
pD8++OAIuqUOfMBD0n8T+US/TVLPTY9xlLc1by0MqWdvljFCB5LWwMhBpRRqt3/1tX9inRd1Kp+P
o00vFDkaU5SSfdrKEFcLn2ZF1jfhqpzKkTF0vYz7bRYseS70HK2kCX9TwxE579kmWm1VXzGjdEcd
CgwlBQFGDsUr4QwGWfjjAPVHYIbHeNu1mKOtUbW1o7UUIsHjRAqLhjegsRQT6T81K8L/d0kNAR2R
OivCOsyzZEP/nYV1LWqNiQfhnyVUXHBpyWA59VLo+OUojQxifT2SaGr3jlN28tdNQgGThlJfJRVy
oUXOfkTOLkSYgqX2Zurcu/8jIF9Z4OqLk+kiB0Ba2tf06P5OEpGFeWWaiWOCyh0N7CzrkJPS9r4U
yu0I+w6/NIi90a31fitDHjyxPeCDdIJCDsussxaKvFx9CbBEUIxhFiFR41GSEmW3FepV9p2SdRjR
LHSKeAE+aXn5HwaaLJzQHwU/mZu6armFCRAFhDZ2vIF4c11192uBM+rrO5dcv8rPZNKC6AxNOzkC
H+920A1RiYPkSlGLzp8bq6ibzCpHDWUlrQlXXLy/ti5WUD+q2o7l/1RsuCLkmOP1DW0Wdq7B7vzn
gNYqyXa+vg2FOehDC6VijInUB3XPKDtjB0/evvL+hwNh+bK+9KKuExyicFMqE+2zSuYIjl+ovpd6
0NX80YK6rBGLggoJcJFi4veE8UhWgsp2AED3741Fbmr/RfAwi2dlAD4/1gRsEGDTH1npj2LDhXZ7
SvTIIAMAC7ATNK8FA5qCAnkcrbj7ApsupvyI2lEQT2omfYAATCdm6EiIE8M+TGGMIlmHdvYdZ2Z5
56wCuvexvJ3hlz9jxIpcO4htPL2OpdC3/peZsyWA6JHtf1Qt7iAxqcSzI9P1fPoM7G3EPEIGqCk2
NsasFcBVQs8YwPsyfxpw11Bhj74mS22WAfq7SYuKKvtwwpwJ707LZccMExiX5enZrCWYcGVIH5Ib
KnvTOnl0XodQB7G53H60jMSmDL1J4eMQrBeU4WNky2E2cCayT9kxQkglChx/yeVQqh7ErxUg7dZq
i+WmZAnVpAYDunvHAQFbTAdvAg+xXx5p427c0hiNwV9h1GniOVGSRBo9xdXWBI7qGc0dknfvF8UR
C4FsV5ArLvkc2xZDTL05uU9yfnjBPvFOADUu0p1qC91WFKD5NqVe0XmDAcQaBWzu8hBaSAAsl/AV
EhTFP2rgoC4sv5dupoYQDE5aaDHBcTJctHLX9JvfqI46DgYQ/Q8ycIePOVyUiE8HVMmo6fZ+wW9F
TlNMLa67Mb+UyFetVCeNN38QI0V1PJmA1SXztCmVMv0gsnd9EFINTFoOCfCI/XpohHbjxh1p2gSe
ciPlqksFwxu7woYdHo/xtz9et1+VzsoQsjKMolfZ6q1tmxXwwqfGpg7xDgyx8BqnK8uxEAlAGRtV
L3AFtClAItQg2aemmFbtjBBh5mmWexpusyEN6MLQ37lzun4CK8/LeIg/CGb4o1WS59VdbWvF6FIP
GDUt8EZRyYsxpVXnOgapapXF5SuTXHL5f+toxOJ8iQ39o1B88WsKdi0XDOORHVuYk5Gg+V9gmsoQ
AxWYpye3xnoN2sxJjEV0CEYuDc3KaOXhTq9x9zXDteENfcORrsdMMs/+thjmgN69q/sBEwzCO8BM
kcXK33aEq9OgqW6GBiCfwK0Gs4OJWwkIdmMSdBnn4b8HVQaR3vAfUmdNViDVWINImAdPcWo+vUhT
6M25wmJbWNdU1cODMT+UDPOWwsBi89l9IM3wfK/Vs5cTPi0ucfAj1RUUbrZ1smVS8BYtFx4e6YEs
L3At0KccgeIcrzYyKkj/qHltdFDG0gZAF6HrwsTgGDfYD5nr5Mx9+LnEDgFlXALKNdlT/f66zXZY
3wr8wWA2Czf3sjABbEcSUrOtbweC23ZlowerR5sCp3BtiJdqz82+Ri4s/kb5xBa9DMzqn0VAbwRU
EnUwxqjxKdsJ25QIL2Q7Mx6d8prJf7UiMwICtWh+WIEKzaLGeSdacaJw2qMJMmoGbFeNqKq6DCor
TkjVTOQ4Kepq3t2M1QHVXRX29yx1eu8wqzF6hTa8X8hd+P/IJ+F+SlxbArgxirHvHp6875AIDcon
PE14kKnX1tMP7goNir75Gb7RbydpDtkF+34o0GwltmWOXPXlfsJAIAqnjBEGACM5UV0ooeHgBz4x
OaatjFYBb6mP0IQobq5EvWzm3YtmqKzpwi8XKacdnWHMDKQe+cq6GNJX8/KwkuS6b2764tz4lVhP
sNko1etdcaZFILsYcWeQqmF1dlgGSkUUk80MsXcxG79zxzNiYBUG1adk7Skw3qQ5z4tQWzOdylwU
U4bbguZy0DinaUfoJAJOj/pHLegB4uTN3hF5Yq2wyDcpSQrGM7GSaxf5dLfoeyAyFb3ighIXhErJ
JO6otpR672XZAn+pVvVrn8QD+pC9kchvsxx4oLr+tKAGo9f3lheBZ5+ngllaWgfmrCMrZOBErujF
eZrXZ12GcTw6yWH2zgFostuZho/HAPfBd0AaZ1nAtYljxnpFvCzOHU+Chp4+BvokTA1CyqW3ri+0
28fd7DiAB0k0udiUmMXz394U0KHdBSouIIF4Ku9CSah3r4L0CY7Ju3A2YmI1jYees5oMOZMRu5bs
BLguCxsg6UNs/QsFNd72zu3fptgHmma6JKqmdZrQCSnBm4jwwNo3hVTmOxLf1iXTjkXYiXq3Hgi5
pmpEI45dgvkDrI6uUqRyfW6IieRpCEwpUee4/SYDJftw7i0bF2P9AdGFXdAumBXG2ZNC/ergYzsS
+ccEpWfDdWiNZYymR4ln8zH4gEQvzcavtzmCVngm8sFyCOROUHy5SEi3WHH6oTFSHk5hJFrZX5od
NkVJwRixQjO+vSnS1mpUe30kX8wOWn1LSYqN2CKvbwL/URUT4HNMeEtjc7xhUstVjzrcp1X5AtgF
2d7G/+qxjfuaR1t7Qt3i16xS16OpAGrio8VWHESnsYKSCyrPDg8TTWaclX5K014x3bdUrcnlnKmF
v777F04TalNFS2lw0hMlNklTcKOMCjjnsHZ66scRH/1x2Gy1jARfNkP4oQ4Vr4v/pI+SVuew/aeI
tw7YBNgs7dOYjkJkOwQbFa7cQ9CoXQzaDyjGCwLF16D+TZllgZzA4BQrNWQqww4AADs6Hs570ELg
waUUL6TXQKh5pjwieGi16w4TEpjFCm0XfreVhJT3RyWrvbDDiCG+Ka3CAK5pG3jI0MPr/AYUcWQb
50r163jEd0hCxjDo5lNtw7VUQdhLxtUkLb1qhq/mhZC8E5Qbf5isUk8hosjDej+N3eUSSVI6trUI
v0hT+J9X8NBSTWsDgR+ndCngjJA46sKfM5pHS6+dwfHbU4A/30FF/ue3rM/EUkAI9GHNJFrEXoAh
6MXEEvupODtcN4RYQqjIyoaYurTvpg8fkLGY2OFQZzmf05dZtt62B53LmXxx1aPVwVn7ptpTYtl1
7QJkX5fyH4ICfhtCCTPN0/csx386fxCdgamSHQzPQTf7RtzQ8It5+d8Y4qjal4uFEQhqvRQHQO7H
y47BCNnaTkriSxdTQey6E81LpxJ81QcbGDV338PtSVHcyNHHrnBdRGZVHzvX+zwcO76UCx3wcToa
FonWzH1eWx+MQB7EkFrmieOojg2GGx7TFrJPsE+MBxY074znsHUPzJpzIMi+kIa7yrs42tIYQjfI
jBuBYxhvtFL96W5hovZi66DFuKCf4CvVdC9vPa3ljDqdg2syuFhx9xBMRwWptnYHvRz1Pt3PhDqC
7X6SNwcFcE+P11a9vaXEUuUIy4+vNwhqAWDNHhFpA9EvcfYHSOLTuFREFE12NVh7tp5Azsjkt8mf
Tz4POEiVdk0lsCToqLkvfcDmvk4rnrMV6t9I5heLfcVIIB78R/B/h6QBLoAfsV/3Pc8jvFovXvae
wl7pX7i1+xwXDHQvYqXLe+GkAeIZuSamxwA9dzvcw4HXtI8sIM6PEYhLn+jpBcTpzsLCReerSM8+
nxv9qD4Y83dDT394JguJmEkG6ekAFcG98z33rwAW0seL4D3lMkfjFXzvOZe2SXOSZi94+HcfpGm9
UsoNQLaYniEHlOxkkSOq8TrJyt/H3Qc1+0pEW6Kv1R/GaabGG4ERFvX/271MkfJNa6UpaJOkM/7G
ZQ7AY103WEODO7F3GSYbZukytkZlj7lSt+V+ydu30BDsQe8601ufwX7PeKJJpQMpH+O0kFwldJLD
CdYs6viXPHDRpMkmVAO7l6QkCgABATe0H7w37YcHaMZ26JBKj+3B2e/1hRYxYZW1eQau2jAq+va7
xJti16qx0YtbtN7V76uk2iOzqBMkK2f9yEPy9lqdixRv47j4h8EVIZwqndyEovjkCjX7v/EwiMFq
LsWmt4djHrxf0/49XyEvNAvUT4Q61CH43miXzz6S5aZaRtxtjwiBDHUwa6G0P/qNAQEoc0fe55lt
SDAUjoh1xfLrpieLRXeMe5C7HQmR93UMTPgIkxDcSiZhMqPcGMoNkHe0PhyLyJQmtFZlcMNSbVBi
imbh0JtmxtxBh546h5d2UGEL93ICor7+lxZ/JiE16op+YqlmEsCz1XcpY7bZgAamVZrQ2zjcbVKf
QHm7R8fG3v7gWiWTa6tniQCvSBw61lDAVkRA0K1e3EQewWfo6Xl6dZ9nceOyXg5V7Eso18LsgsL2
zVj1FEoM31LDLatC86z5XEpOu677jvBigDhO5DDCKuCT+dWl4zBXuhhPHD1jUwdv1bLgOZvPLoHz
MCaLPZWeciq0gs2alp69GqMJUNvcpwUbdxMVegozHO9ehnhV1O1n33PRVk5qAiCQJgYXC/00D35e
nsoA40A3gK/zfh6UDUXVr7j00GBgWsE+NbuV12l0UCji5IdbcPOJQei0CESQQo+bODHckRuSS5d2
l+3N9/12WFVeqIIW4UAH2tMfFI1qDyOeWogJdW5q8YA8OxtEBgquUFl0t15CnYq1rjjXrWvyQDMq
SERfOLZoG8UErHYmbIZiMNJbAlDR+CS6ihNAzyUzwsxuTdUrRc7ycjoXo5Mj3ZhJgyc3ouJRThpq
GI/t75TcVW+Jbep7Si7tFxpC5rX9YI8y/5uXsRDwntbleqfx3bAqNB6NvxJm8oOHbtOoofj2ib3t
YaVPeAPn7sWSjbqg4lcZeCxIr54pUf7Y5HPLVWkBmSTxuniAAvzh1Ew2S2Sxqey2srGUlh9u4DyJ
wut1wkoIC5Vdt/1o/WAPRVDEX9l1sYIwEIhw4sba/h2Z7IaV5QfP8P3gaJ5LJ6rOkFtMdpYNIJPf
kdKr7FLZRojrZ/EJmj+YYtASU6YcOfmrwZbsPilPBIRkYGjPWXIb7Llife1kJkF/bUlFwFjWQZUp
+QgNM1EPkga7Slz3Zc0dFaIjyZG4slnvf9PE6p/HTMtbHWMw8KLoZkTHWi3ZszXW8mGTYXu0p4MY
yi5ojIhjSIAvQ9eClTYwwvSJHqWieI3+wrn1o49nDlLSYbKVnnUGUsdRqp6Mrx8FkJUZ5Wss1j6A
k6f9mgHbPscahHTxEexaRCW1DIHFptcDTRPhgXqlkNaIKQXF+A+dBF3S0MkPPdab7C80hlhW47ZM
0lnfk7TyrGEFBtZXk1X3M59byUB4YjsUqktNTL2tLGOAfgqoDVrvpg/EmIYtb45mWHgeRVBKb2iH
pbCEjayhG8e9Mwlap2SpGT3v0U0t/mVeDTmKnS3NzGV12EPtcTOIp3ucZyHsc0FscO3qeuM9x96R
QA0AQdavr4oAzmSj6Uy86AZ2dKlI5LNLWcrVrydjxLASgSNV1orf3p0hKX8d4a2m7snccYrM1awi
5xdYhaDFdo24SZ+RcR2KXSO0r9pby/97HigDXQRdUhRUqW027y1GfPZcHqAR56foTnVEJl6S2713
LaID6YDejiyIwdoqXfC2ixsejbF370XCI6pIXpYugfOkLU03qbHied5qoFeIAhgyRz7HAs+SDzR7
cqlJhONvWvjvVuN8rULjdknAeAbUUNOPg0jg+2PnPSx6QpvgJ/zwWTZekVDgUBJj1CCzXoJjezr8
DiHr6UUbGF4yV/GaHjGsE3iQLOkz1xZYAWqVSpQnaRzU8B1XgSHuPByOZ7b9bsfvH8G+5r9W8Jc5
4C9utMIJOTC2UspmMcq/E9083J/DI5ttrsM/7iNHFUi9Ej/uKaEakGkqA3cyG5H96sBFQ7Xg0l59
l5vIuTgmxbbKJowl4sCF5njZC5HxQF/oAhTLrdFeUHeeYR2lnVoc1FjBB3eUwDh2EPOd7Re04mH9
HbQSF7H5KOJQVQJ5WtrwpNNq7/8k9cA/uLKTOMhptFtFoT6pc91KqwQ1eOdx6gFAgPRO+qCeMYA1
013rW5Y9lb9rrGAIx+olRl0HZxjTirjLTCCZta9MOrXIG6kH5yvHG6IS1UGqTOQbxyOYXOeVxMYr
Oo4qY9WOblaLkDE6CIZQpIzno77sQKYht0x+xrjxqkhrbkos3A/6hFq7i/Q3XtVmaYdx5F6IdFki
8dnVX7WnqjIbD/MnCBojJGIDDadGsnrXfz6B3mR8wUx9s5X7sSes2eSwZk/FuSrTMJ4uOLeKh2Pu
twSvAw9wiu8zvGivfrBPjgGh4hZ8+BgDw6ys+mZCvUewG/JDQiMxBVEFhR/K4nn26BatRqAiQbKB
fGAuyn1nqSIJwFCgjyyMGAiY1vUfGDXpWvEjfHMoEMveTgOZi4NQ5rpVbhhELldyI+4HevmZiw4+
2fADH6jtdPOCX5gcyJgpz1cwUgabKxr32TZ1UZyJOXFrAR1dI/dEUJTA7IArMZzXYDYScj43ham9
1wyusXTKJbgDiF143YdYnmtIkHVuf0sW4MH2LIHMMcSeKxIGZlpqVs/O5fwt6XyvTrhV/zsDaiNo
BWbZpmKhXLAnaq6Br2x2G+IGN+tOBmq0RMQ+wbuUcJOUeOl+/t+7dE7TGdo2hVoA+v2fFDqo4xjX
TbT6WjiNu1wDSaBI7DfdEhUoA2EIM3kUy7nOsBc1J9gYeDwIb02Bmap9xFGkiDDQ1ZicCNklaDKy
1DL7VWhtSqwz9Q0xuhKAciHijDr5Dw+YIMrQv9KVaKncYQtI6xt6OlBEZUj8SMLkPzJ8sUlNfCU1
WednSsMkmVo6HB5ti+FUkimLmMnesVox0hYLtLIzmNTEfScGj+mVZbyHLT6nr5ddYrotOo2TdCt1
ABPtfxhEGmoOjYS7+gK46lKdDc4BQt3l3j2o6jcBmvtlxPOu1sLCaA+PgmCrnY6rHXzXCX5DDy9M
tTLsmKZX0GmR4G3coEkI4tVK3gDJWj95ySOlxgCCRcKCQwtIS+QSCwyNbLTo1MqEOmco+LvZVBg0
e73rDBCdG70lsYZfS11kg5/a+ay8/pCSO1uTqlfZBNW2evR4TJwcbOcPfBAGT4i8y1igfHOKBPe6
71/kTfrPEAT44MQNyutxZyFzdemlz2u1Mr7omBMnhtilZRhHnrX6HCcp8Pel9h4b/6q6Pc14iX4s
D9jMioOjyJd1ARiJZvOWuqrlwZ29xLJrJip4Ce8NKq70CDPg1JA5YemEIQyu0EY6IuJbCeR2gMxd
J4eP5/6JaFsD9iAASuf2JGNz116LzgGQV9aBY6f2GZN1IO34Y4zd03QNJXbPoCzf4LwO9TIYuF67
PukmQNdzaRUXGbk+d2KF/Bp7OAI9AqyT/KfiS/RJgr5HXyyGr7eR5uzR2Pnjqtxlvvs86tqmGdbi
Z3EX7DQkVMQc274eHSWCet2y+e1hEKlG/mJ87aXTCWJa6Zpyc2sa20azy+Vb/cgPzNCOs7rIngyj
BvyTc3djNYrwp5IYN7sYu3HYTgzkkE0m1PYTAorXb2YrXiSslu/vb0inZRWALObW/v8/pJodop8r
pnIp3n2QqznvsCBm8/YSBGP5KFbzgD0PDANkIrk0qL9Z1l3xOMqokIGEZpwaEjpTa6FJyE7Tw4Jb
v7hQa9x5qCGt/RgdCu6Y0u4D1oLID8eO4sorPJaXPrHRglQyQEO+g60UxRGBLTkk2IKjKjHWZAaf
qBdhTmCRiPD4gDkv9M9VG5BaZL8VDkFtaxXLd0wtbD1kdfcjAnbS1O6RIydgT5bInihrJW76Ngye
WVU/QpKpqQM0KUvxkXKNIiJNfTfFJxIiD4R5Vo1ZBqe8aejVAp7RrXSPd4zrL1S6VK1Iaq08aC6s
hKHKrX6gE95YYi9+DZf0ITsyHEL/15w3ISHoQWFrFJYHJLP/Z93N+fDFUtm/94SJVqXCAhvpSEDL
flYbcHiMB/X/3jBIXDn3oeXTD/VOq65aH+fPa4gD0iTqnU+YhPVv5R7KgqKEMhG5OE9hcRQW1RzC
dhXPaetTFWM+jgR7Di6/5GgtOkJEKSkwqEQZfMa700GJNUWBklO3WvhisJKxRot42TSerWPlZ4s9
JzIkY0lMINMsCUD+ImfN1lnEI151vhy857kcTBjZOIEadWc3tAZPMIuxZs7pG7fLNxziSVwUbyYc
gmByqhmVuG7v0OzZLGL9Ke1lrojQk5Z5QWycugN6sNYcnqB5/YFzrMT0WjtNL/+wi7oCDcDbzb5Y
JlIFZOiLxT4DoeVPvCacTgSXtZ4fCcW+QrNeEk5kam8ak+EvsTPC0CiIIIvd2UUQ5uC7roPkJVfo
rmYYwi2e5bYe58WZr5DHPjg0gao9mYp01PgME8Hmfc92BXtesd/131zpfVerAn5zCxpG5ejHHfIg
UhfZa83DVfNAtE9qvcoCW7IzXotTiHwnNJiaBfLhujwfy4s5hrcGOY4exDvTEsZRcjWXCCVP+s/b
DKcZqqfJLsSOFskhJLCOEDBxgAET6ma2e2ntVIjlRyHgET/SosBsbhYrrwoRBjl74z8bi/81L03K
+skXGTiwWuuvpwB2V3h3nmlIcD9hLSREXWHTPXMQBebibVDMhmdpPxLHZin/ELLHloin+C9zhhoN
rbEXp81aPU4gMu+RMyuO7ILGYR8YMHxwrPK8Qa9R15Q0FqJOgSEh0FEnOfiigLA2L3JJpbKGbisM
V2rRckSfHe5hlhI5EPxu5a1NWJjO0u6k3vbJ8Sz10ZF//vG959rLlCotSc2iCMIbTOL8O6rG7m1/
UNavsxAG1iTWtUyvq97upsImozaXTfxbzibHuDpT05BvQq8Qzm78LnRxMC7O00N0WD77r/06JE6g
u2B/EH3ipFRXybNPkVgfUOizy6ifYFTXnNaKQcrJ3fDvFUzUHEOvGTu6gMOhfp4oJsGhwSvCL1aA
4eW5Q1TPANqJly9bQ29po10lWDLty2b/XYu6FY7TSlVaMcHGWHpoQE38lqur4nvXXPqNn2NK0qIW
Iu0uwOyEt/YocWVcAyj40OAUZHBu8dQaeqI95nGmOkeJL/PTApAX1/mFJbAktRx42QHy8Whey6tN
zlkYO8L1EISDU8okaDYUKQqoRLOer8cV+YnypAY1KQRwc9CB0tfiYm17jAFVNZnwH5NnM3trnoaI
ZFHoTlj4WRrOVjph0gNgNZQ+zjvPJ0H2IH2bXWRsceT4tk52mkzRWfDo3+l5uJ126EljBj29QaAa
2ZjN5SHSvVrJkNYvUrzu8JuTLdeI+GMFiEcC/Ir4DPGrgDeGKCLXnOg2msGuADVLMTgQHfY93RS9
4VPXZfpawhfujpIeQFTRtMDLLY6qNnaqCC4weNR4rVnH3vOuDasjk0WrnyHUaChsWZymEsz3ZIkc
AucX6QoV6KV2EbPORhCnVHUHnir34zSPaUZd3nvJel3MunHhxE+VpfEGqj6XXrZLMiwdUers5dbW
9NFvGymmKI6qvaWQhB8kjUpD38jC0RzamqNBQjf9pvtEjDNaO0GQFLGa/AfRZr3iSGpBUVgqyd10
W/QnpBVgF2fx/o7Rci+zYFcQ1I9xJafRv/JrZpZUhXIFyme8jLHU0wu9Bi4b/cZ6hbcNyPgIg2bZ
Eq3rFUY+To0F5frKEubzUii7qsM2vedLAtytiF8AEIfr2jzGyZCu9THyxbFpH5zTqGRyJd+PfPeY
EnA++zSwKq9qfCaGnwmklNufARHNRrxrtYMafzDsMmLAU3MTp7U4osFkNoKChpTN329kBOI7XbGD
DlRuztqoyMPSDOOZmmZU14iZLxWHNTTF3Y/phK0q6Je+74flmZ7BMZiZ7dF74Xh3z3zxLHWNhNTz
Q0biqeQ/yfkXn8PWWUaeOmMO60YPigF6hDD1T/zRB6UwyaNMcNz+EfvGXoRKxPzt3nhWdJvUsclg
Is2McmmbqFyhkjxHo/brneuRaQ77p6Y0MFKLsUdJcbQeXzo/V97ra3NkStQjxjFeF7/AKqc59+od
iqmMTOQ99gZaqS5ME1lqmYnzkrX/xlaeUIfrrLRq/urN36DqZkp0Zl9UEZtj+LK41XibEAN1k5Nd
dofnzyXMPiYC5fQJO1C/MZh8e3lIcAwhvjPSfFL+akGVPokrsnRYzcl5in73r2pJCQNUxGExLUh5
tmUskiOequHt7MdKm7ZMvIXHEa6RBfA+MK22QN7psliTn4c/Hoh/q4AjkLQnMHWJIAxcYr1e7j9+
PhkShM1BlbWmJSqGo1/XD2KblO4Fu0BLAKoBAgMRZa7VX776CREJL4hC193dPatkXC8p1IDq398B
9T/yquSQ/feW1HxMhiRdFEYuXRfw225milK7A36/+HV6R3XP+qdaNL3ODgESLsWWERX7A8xcmOEM
WVx33cMx7+OBECZlOkAgbk8gJQ7kn4FKmZSrMPlgV6coYd01uyeIZsqZT4jYr77/94RIzmq5Hfas
+wbPP1AkSORmn42LkRmHFp6OsZ8WTav1vBOyUtexBOAtMzlgr1j/G/yqEHTELqa+TdPw/3OeP4Ru
FCg4mkw7+ANRo4frNkX5QyzqhFWkNyRUZsdMIc5cYrkj78vNnnKib/EstxAv73XopGmCXWiSuH/O
yQ2XFzIBL8bqs/fmobf/If4pM+n8wuks4o6zQ/BoBQjdqN3IhCojvWYClMZ5pajNbHUqSHy4kHEP
F7Hbtf/08hj8brsKZoQI3aJnhSto9c24GRJdOXExJmvzexhlYoiYxdY8fw5FOdP0zyuEYN7cu884
mEAhquL3bTege8qYZwDs+onKFftyswek2F0h61fofMMp5Qqqy0wcCyGf2sDJ5UQEoOBejEz/42hi
e9SnzmqrTSRNe4YcXOXOOTv9P/Fhxv1kY4q0EfFy+mRnE1CPyoYxYs2mKoB/wqDo4v6HEBA5fGwd
9+PXrHxwt3AC3nbhGL/Xs2BD5nmpQAdfOL56OrhRisnCXWQb2mducfyLVLXLaPqZ+yDyUMqGdSa4
PAQO4scilONOkvGY95aup2YnluRC0rMOycoSbSVp/0n6PZfaWs1ju4UiRCZftu69JkA4epzIA90U
mY/XdOqhEg//wuHcEP54bTZv9UDeWsDaykPzuerYNHuExcpzHcto6KY1UuOAq7PQsb+ld2cA8aDu
Pd9L8ClaZwO08MxoIiGpbl3IZcO49sPkfht8pxKYbr7Wbc8NjNG0zjuMGaY9mF8lz9OQtBvc81my
B4TEAVwbhpm3cRTVVuT+RYti6Uf63LCNKdvuBhDsOdt0axG21niqoipTQRQNGeXoe7ybBiNtNgft
WiWuxf029F3hGD76I/qC4ghMse3Ajcbi7U+uUV08I77Dj072b5HMglbfxi5HticCAGB/ZhwsT4rH
vFgOVQzqrRew6MalVIgM9/1/kXaWQJF9T0fhptMz7BQNrxarMbBU6AIN4pGi1xV1+ryOmRkmDDPw
ASMh8edJluMJ9X07dqOQ+A7oNi5kP3i7KSIyuPRUXYthHsK7dQNhygjnVS0iIfsF10XIeYGmkbg/
2NgHI+B1yWySaxbtrDDoAqtMlu7KFRDOPjTp7AMkCOpzADRawyYvaeG6gV7nLNbwlOTxXHm1tQOg
Flb8s+cdoJmTJPd5ctm0oAVyasN7ExIZ6PWBE/pwqHtD3cMlglLlvlwmXWjX5DW65xPz3oHdbywM
X2Ix4kNx2W0L+OlOHKOUE9MKltSvwW0R5gaE6Pfpa1x3mx3AyPM5AKbc8i10X4zLfvw+JSj+GCIP
zp4mSZhlqTUjgsE6htLqQ2QtNxsz4QqueFyMNwPdnog58CSb1lvhc5SmT2DWCEIRWUMcaqW7WFpr
IwakToXSSOIhqLr7fdVPCjJrlX8zSx3ewrFE/fkcNYNEHWPRR6kBySoSdzEFHLUZUyI5dgeKWGs/
5WtkGZq59zLWNlvzKKzf+P/OqvsdRHqHWplQcheqDPsGG4Uu5c9Vl0IUOZkYbrc1K7ONUC1iehlZ
D5n3FfuiTqhZIDm6tvJ92VjvJL6JzYaVgeBVDvRnCrD3XWcMt5P1BjjR1AuPLBcZ115stkXh0kAr
Alq0Resj/ZlPkx3tqRyjyyRJWhtBslAuj3zOy+yGZh16PRZDeUaDafFPIvOebL3rsZ07F5iQptZi
zHYkEUojpvnAfV/0ik1YYa2P5OiRe7ovWxnITJ0oyqGGg/h/AmHipK7zfwJ+S/KRAjqUIQBJO8bT
00f/UHe8SDl57ikFUIA4Yv28p9axRh5fbCdzkilF950WVwKAFfL2b176rxHUL5fz3qb+fabS+cfr
7eVuQdpF/Fge2r+zzZiyQIi0w32mR1oMkN5QhPimd3n4hSqmfm7LhAXcBYHafEdjjCBVkw+nhB/L
uybSdKLs+lY/gfmEDNj+xG+uUqc+iAvn7XVIreaLnB0mmvg+hbR3oGhVCpX/xrBK9PH1BmUQG2A7
QGd3tw1r5O5hf9rwdUfFcxxOBhTF5v7la6P1WLAjHrmQ9e83KRnT87NneyTOqKcmNgNTNkVHvDMu
Td5sMDvOzuLV1ce8MAO4cAcCXa4oGwY1k+aMNJ54wOlaDhGjHXpbpS9E5To5xEiXQplRxSNvKV7V
96Ig3cBWNH8mBEZHY2kBEmpFDbYY6ziz62TyA0MTfWHxTMV5xN5zd3DeLDddOenQMxB620z9XEK2
VrqMJK5v/OGwdFKOEcQ5LzAr4BjerrviOdRm8KTfnPAE1BDyzKWFyVwMKRA9pBIQvOfwzbDM3+wa
C0jQnf8H5lK0lqC7w/rmm2okcJqv1yM08T+FmTI9c+k8eX3nBLvq5kQuoAfCKFejuWsJLKA4sCfh
BSJ6mHEbzcTmxHouF25PQkHPTIYNB8oKu4UcX3SyLLlV+7doZCLY6TFs4MQ+aM0Fo1vSjgija478
unmwuBKsz12dLpmGyUSAHNFkeJZn40Kxhy6mM4ZD8YPhKANKachLBK+8kSOkSKqlZbikLJJm6nDK
xQu14PxVGTXQE1wp2crVfihS7BzQUuLiGXPMCT9zAUsNXJa4cjN26A60NozG8NkKN0hN0Uw76e3c
QTrm7fPUCYIk2NwC42MJyeL53Gr4klDpLRf9pq2sgju/FFa/Q4RcwXYTXx71Luq5164Cj4Xn6EbZ
+stSVMPoSqgUc8JYlB0CoFbPMb62qPOTFNSaI1FWMxzat949VrLeWpvh5P5RIWQQVSk3jhaex35r
wAPCcuH0IRjfs1AE2GvnNd1GqX7YFEP8gBHusaB1d8AeZ5xDNlMK58xJ1ang5pYmUHUHvd9d4pRj
1Ra6uLMZaDYqafXM4QwFYKK1L9wVdCfK45NEyTrAhmTqdvWcSG11ePl8KR4ag++7BEH/nt86llLw
OPmIKGzd+4/WigRZhA9Di4dyDpeerQXJLz6hjfjS4qIkJ0OKljHnabrfrOrHlfuGpuKaSF4DLdPz
lkM0TAob31q2A4FDRJOUcaNXD3VLVmRmJB1eJ+m2O5QVPhe2XfdEt/xWvUgWcVHlykdPdw3eRiuz
fpDB7jBNVNdDfSTkzg4dcOKn1pVIvYeuku9o4lShPzfdcqniovz56fqv07ku+nEX9pxUDsFf7Pde
/kUi9CiXkK3QiNMsb6V1/Ar/3/AGia/Bnwg02RReZLaESolXZm3PjlM0aMhhkS3zVYAf12YZzgI0
Ee71v5WjPjSwXdIQhSHu36ZAk8GoUBT6H19t6aNEQOQy3oz+pVTRBpQhz7DdhS5OHp6DVrfB126h
5/V6KWt49nkGx2RvYMBbGZvsqEmrWaRZhHrspe+ivOrrgCp7Ux/DJS+fUlL9xu3ephAqTVPDUfbx
1X2lQdWSoeRUj/6HQ7Il15BgK1Cjb6/pjYX8fzQeyafdbRv3fL88h+UDF9jTy3g90sGj1dUA5Mux
4t2IpBiWSyqfg2rrmXfHDyRrPj2OBsHutCmBxCBXT9EDOgHT6ilm2/+QQBblsd3mD7k2s9uJswNX
9vBB+0qT+ppNBpcmA08C807C+HRrCoWEM5LwoPQHFxQT0Stc/bmvhsDgisqdcNEmtDhzpli4Aav9
jkJNj5Icir07+5luLBdCvYeM+VudU2RVGF0fPZTDuJ5uA1jWTLSQssCrjM3h2LenFdERt7VgocDz
XsqvohPQ/qxgBUmW8b4zKF3GziiNlGWunsGf1cftFdp+9IkufTCBmJ2W3mJ7yq/bdD70XSMJK2iM
voI0f9AqApwkVMP8+n7XXSVBXn/5/TB2wqWxeKhKBMUrhj0tQ3uRwU7Oxlvijk2z499Slo0s4cKa
IR4i9AKFZOvRyub15cdCTMoCH6J+h4cyZhqJFbgpbeuPH3iXQYV4GPZul4YFVP/pYyj+jsY1aNCm
metaxaXzcBXitg5klf5ZDiqkW9HmhtiKfiG4IvVWdeM+peIGPlQvotL1343Oq4iTNzmOGBWCuMg3
UpY6EWAH+hZ3rvT0UN37AH+HdL27Jspr53Vgge3mK4ZbrcoHyYfSG/zA0gv32SfC66T/17s/V819
QBw73YIbXrWK+F/k9XATaqhYb4HUHNcwsrCyOMWqFcq4hdBn9byLdIlPRM4RkiUF7G3mi5yLJo8M
Ts5jwESi08YVMMiQvQ7CZ4Rcxu2mLMwKnWKAYrjmcr9Aau/3g/odu7AQuAwpYIf+N6IlAfj93kJY
gugJr/sRaqtZ0tQYAkNA4Fh3bXXqOzO9qjz5zCQmbLBmSYKJ20W/2N6k+1gL5FFnyYW3wqYxFvif
4raMGeJIPnIqM8qwW4IfBJQG3/L0QxY8p94beNuDICUEq5VzgEYShfK6PUZX2AC07KmJxSJ0vvFB
fSWiSY9yqY/98/Glhu8h4V5E/8g1BPlHfmC9psciFYo4QEPgZ42kTOz7v0ciMJJODoGl4HFUyowW
kgWp7O/eGRg8RKwDaEKVn4lRghTLnxWZ29MtTJkAMMiwtFjYogiMQ9L1LG3evneBrFEp/ri3TE1e
pISBPZZEBJ9wCSj/AdyxmfmZ0NKeIuhdGZNZn+0ST12XGPXvzEFtaIqY7jr3ATJRonEfLw9Koz1P
IhZgYEUC2p327glNwOeZCdGSd9pBbdVr3ZHjVym7PiApdVWpcnQLdMivjwNHhttq2chhOB+1R3sW
dqxW6gdHsMEcODGXX2uITJzjMk7dzKsQIwzza3q4q4iXc8GK2Dt/QEunU3OXFSwfakmKOa3PP3np
6L+OeuXJD2QLdEci2aPE2ymQircMsbb5m64zhsbLFTzwMMUPuuRhg6X1sna8EmnJf1tZKnJfTkZF
mYKT12cxzJAMSSdSr1zTT+Jaon6M6fpMCKq5I9Hphd5F1/lnia3Gph/2eE0dPwhKuhsVdtYQ4zOl
W2veuq1Gsl9oRzNJq84bhcik++8RrxhJ2Ssb1VmlUwizT4xC/5Ni/B2QsKEjgu0C6i+GqPcvH2Qm
RtnluM05G90Lvm+tEnr2I9/D9VP/EK5fvqfyGmMjPb35+AD91QT2RtAtHABaf5aLj7I3IuGQYycE
psVrdp81UdIccuJbgZLcrIWomcjK4pNzhANTgmSEjYXR7LHf3hninnt8cX+o5aScPxnXZ0oLVORR
NsY8mfaQGYDbtgnz0bqnPoYPdGKUPyU8bnMzPCBWhjQ8iJKDNOcagKQYvoQi3dBsdnUtnkACZq4S
W470kdH+4LAtDg7xP/nwynZq16w27rMeI35TEjwZfJHQtUgY7jgKImoS/TMKKBY7hgIcdSoaoynW
tRnIp23peMtlxzkJHphYThTESmHjmAsEt6PYOZrTtfHH6B7cEUDUOgK9sWW3Mjg1irV/qfmnkMHg
xHnoBtmHcXLVZHR895W5z51rc3ZsjuJTM1tPiw8TTZFeUZrRhRUy0QFvEufHJLzkZd3NrjYHRnIt
mZ6ilUZqJ+LYYbm8VIsKQoTM4MyVYKpOPoCxXaKPVmdlRYjJwN5t9dOyhblTc9aRHQvkawO3BcFf
iD1EfEA9Xk0AZcGtYVKAmPJZI+w4ST3EzfVT+FF1GVvkhMSmt+KXdGU4zIdXWTnBFxKrHZkaJFZo
h1zaiUtViGoHuFnv4G83e0/pgkHtp3mUYuTNr2Pd+iWMO2rpbM7s+iEeL6ND4nTO6CR59EZtptnm
GB5q3b39dul8hpTku+/eM3EKd/8cZ3MhFFLNP8+RV15dOVJpm04nxpf/t7YrJBV1GbBeMSS+8bwn
KOvl3hsta+/2xWQtKNnZwawnCKJoaiZ2vZRYWlKIuroXM/EdLVR9ShKlR1Nx34pHoID0q4XtUDpr
v5L+QU89kdxXpAxNEN1Tu1Q1o+iIfHcBe8vVE0LdSlQNS3hKmSd2lo1ujcUIhUGlw90iUSeeji6S
yroMV1FXZRtpE2D3XcFeJ+21ZHoJh/HQU2b0DQPTKh6Ucz/p4RfVmvfYKOhW573uyySQqSGLx+gV
8fEBoy/Jm8Bzvt8UOS3XqyselnJh4wVcpXEuBpTrh21bHgbBkc4WJYJaXiIp3t/RY9EgFEB6LtgH
hojWlC/ZF7X2Ffve6jLHkNGEupppOVz4rXM+tW+2nWnjHTYyu4Q2VpVPE2Z9cDAQE7gnMA1vJXFb
SLMCMId0J19X2NhgiBi5Gl13G8lsFVV3nWZlUT7Ft4p1lv5Vpec2Kk6go3C0jbOFaJtDDSgXjdm2
Jc+CpQ/BqRFe+/ifKS9Qaao49UUcET8Py5MDtPOS+Y7t0Z0uER/Da0nMAenAbDuL6vBhx1ruNyza
7QGMSF8LdsjgQP2FZ0Qei/kQicU1HNRwAUxqgFjrel2p57ODX2dvcVxhwXD6nwdyTdmc2A7imkmJ
hyPkdPmxnkX8IJomzaU9U7X62Li4RmGEz7F85vCUE1l+oNj2ABQdaD9a3gFRwausZek9YCq9Sbya
9XR6gecjOuCYPZ5fI5HQcPou94uHIAbL5Stl/kpBBVtoYBh6AiEinUAGd8UnD36bK47mfriKag7g
ZGmr16AmbWufGU8sOxNDqFmKiXgro9OpVKh9hrJ80Li2glo0+uB+vd+sU3eHhBaiWoQrbACezy5m
kN9QwoRmhEMvKs0PPFShF5vpASBzfgybZZ+yBYjeA+Dv06PQIi0ysfGT8uVRW/WlzsnbM69aoot+
2+lDdoqhS4zHd8qfHCP2HGFiLr0Xhlbdp2TLhMfqJcbHBLnb5hwk07E2AaaJmJQc93Hk1UsPliLm
zJJwiRcTi8LAnAp0t7Cir+/wz3B3kEQHw/jjvTxS4VZQVvE6JybpE2DZ5mfvtpBlhbAHzJWLt6/2
Q8HCxYGxngwX0VvXfdMSmzfwRcAaJ/TVrh154YPiokuJnqY1ICC8sIbQjFQnr4JdQsqGWT58+sjU
BPVk+vpvdgQ7ao1bz1XGZ/GjFpGGiQKcjw6OmAU5lx3GZOTpj6tKXtNuSO0wK8MsKLoG7uv/wZ9q
tG1lK2BczW55EQI4cBIlSUfsGozs4XGiD1yrqL3UCsemJ5oEtfN/em0+tDQH1diTlhbb9G0Qzk+q
zHwQ5+rIvmwde2Ei1UgvBMwTH3FzBF1Eb3UNcigrZH59hIhtaj6k7KLhuqdj9jZK9TICkJMtSbUF
uvRRddo5eqeoYrp+swQ6xhF3BT0RtkF93OOSSEE/QMUJEnexscNDxZXj5MdWJJdzRusv9MyLLn7E
J/YPLqXc5WIUAvEzcFBV9pV598tsUFxLvKq+y0N5Ty4mkiFezdCylRmUMxpPpbXeC95Ucaf5Ehsj
BYjZtFVyXMDdxYHAH6fDCEDs1Zh2q/ZwBEjsFFAdzKIQpzMFb3yYjsa9KgHNDI+FjSrG/vxX5zBH
ZMCITi6nBvIRb4U40yP1y0JDxMCOYWv0
`pragma protect end_protected
