// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Wu/rcUHD+bV3EZquvSS9D9/07V1rvi76c3jxxP+6BWknBod3h1BXzzwzBprz4vdttbqokPjXuknd
h2bAxNw6sdR6A2Swq8l5GoGE9rQorAxRqA8lMwGZ8OqZ7TSz7Gq7OhcNXw2DohYXlhMioX5MxRa5
r7P/zJDC3hRWNoTVEt06PJpuugviTOkR4crqLIvO+VfJcYBAMH53r1iNpRa7EYKROyCsxXn66HII
Ja2WG/rLudZOfKZJb92BkQbq9tW+m7h2e7lGGyUNSW+3QoH3+y8SuNeEB/x8dkTkhEq3k+pkHRXh
tRj1LuIZoqBiEYYGvtn0tMMo3ODzs5t9ccN6gA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 77680)
Fh1EtBYrXBka/VG95An5IOyY016YJMRm3V9WeZPTQojYJOJzNTQIyX8QIOEcN0FcSNEWkDexm4qK
4bXwgSH4LZzqJT87+ZC6Zo2hdCfolT2YB9wmY8rlGqakeupELVK3DIxP9NKz9DfmEeslVeoU+d4o
Ph9aKCxUmJdUPj8/wREwLza9MWfg1IWuecKWlJdLPZ3EthMJKioytJwDCs6crVGHg4wFvOa+MKu2
u70DkMFqtQpcezIb8QhU3BtXN4AU76jgagVcIkiO2MvXd3j9Ux5g9kt13cD9/MCl5fV8nLqEs1mQ
DxZ3o03S6OAYyjfbTb4uqFPz5rWsOEoiqH5r6ieLF2tzngah3j2t6+TrQRpscl+3k+I4WuPGp9/9
p45AqiLysPtzgC8KAlDqQfpCzVGI4dGkK8Q91s2hh/CjpWS57H01Nla9DHrIBPf+VyhIWHcuUQMq
r/eM52wxElzremH1xPjtB6b2dgzqrUgajBLDcXPBGanocuU7FyUBkeLQbk13Kz1oePPTrZ2HcTdM
dqbdhgsAEa4aWz3vMi4i8bVC2LWrwltAGaGTrjV4B8ECgaAMz/znlBF/7UtrJ7fONMyFKxkxtdHe
oF7A8gvFnYVea9nhpo+2G5+recNnnxq3f7/JxniVRP32WOqvvF3mtJxUlVDrtXcHayJ223J4NN9w
O22LpEe5ZAf93TKw0zip3XqIYorA3Q7NP0r3Qn8JF1uvTpVLZeL1Ho+T508AkNs35CkjlF2cJXFn
KzK1QkBFMhpPLYbkNrD/xqGrljKuXACo8/WuPJ8KQb5qyfqbctj6v8iX6PiCBA1RDXqpRUB2mYVL
oklCWhUyRe4fIJBles4kKZAX+LSLh2AYt2QRJeX5qCVCW4j5lmsFnKv6wu0z2nO2uAtvWFp8ISh1
CbUkZs3+jWTu0VHl3pKwJ8A6xq+q6qScowKS8rCaoly/V9mlCczwOkW+SE572s7tzxQdihlGBPEW
NARhdL9IfGoMb+sR2/lTQvrZEaDB2jxOOjeEFa5JYzoTHG3nRML0vSaTYHXvptumJfmLMkXCBHef
A15/jKcLPebNLGsnSzSSie2GteMKr+VWXNU7lJ+AXuOl0l1Cfd7ExuyPqMO8Ovo1vqLUF0dIBeAt
EF0sViQcS7hE3XtBms+dTVEilttfdDcGu3URnPB1eStE9efMpkgVuYuSxDzawVlofC0z18+DAGna
gInNHBW0Z4yi1XF7n9zSaIuerXN7L2nPXjKaSEimsoWJppDuzJOp86PY6awbs3unp1CSGsM59ir1
koO9s9UmQWxt/rNSHBilBJmuu47ubxZ+B1p/fMINotA5Dz9Mu6IpE8hZcSmZt09WRj7rGDbBb/xg
rKPYVN7hqsfgijGBlH4f6YWSqnc2edbewZ12Mw8Z7Lxa641nh4NIA25TN1gRu/G5rK/MlSRcUPOn
OoT63XmBRKL/ElB4/aSo28TGj43VDnDh9jr2hciwT0kZKPYwDEXAEGScEmzNMaRmLJ+LPSyKYrjZ
rZWPamiwvuKTJU9VaOStRL8iJ7cPFC0KZaN7gM5VLKjwfT00aC6v8PAi/+OEBP0ui/Ck93KM/ZGr
jgayZnksFojjnXMm4U44WeQBxUFzjEsbLD3paR7kqhkou6hrL5X7XgeRbfIlr5d3GqVLwYzoH8s1
KWmQIpq9j3irXf02kDX8jZHK4V8wyekao+qvVptnA8jcItc5c3TrDBIFQpg8UJ3y1udMcrJ/DiaQ
AoxLC9YHP4OFwKUaUERtLqbCcjZIiG9phSsZl5oXlUrfIFXw13FmfN6arYwlBVO6SyhwSY913Hju
VaP+Uz3XTx7+RahMosela7g5WKCU8ZeJXclGfuPY1Oj+2whDjl8QUFJ0Lg3B9x04HnRtzqaDkAVz
qIeylkga/KkMEfUF/EiCAWzc9fisl05jNdmVbTZtHUthjvngYnFcHlZYefURFBcK1L9cOLwevpKQ
EhOOcz0eyQg5NnJYldqkbH745dvOTT/LAoGgeC8TtVDcQkziZ2mf4dzocPJNLoMH+6hFKD2x1Vox
T1pY6zaIjrGLF+CvK77xkkYrCQDU6gaoFR0TEEmD9x6gIrVbcWKtblNvS4Cq0lQbC9mCR7EpPMwO
QKoagiP/N9wtcJPbwhU6WSnx4VFzgdlpDiits2brI27mI7/VaUn23kdb91M08lPvNs7kNryYPOZd
+UZslMvBm7DsIj4nHg0HF8r7lv1zGA7cMEek4WJxLgpxoyJvfOtj+1YwNwgtU14GIMhGzgfrkyrc
bdjgHPMl/ChmDD5W2oq9Z1GwL9+klX4EhvFPDHxsfbWH1FGNjnEvUPRmpyeWvsKVmmx6Tir/s/T4
GPiEBlMMgP3hytzb0uQoyTn874QLdN7VvkYZQuC3H9454DxnsrczzsCysmMI5IdtD93RmEFG7Pak
PUg4zyt47NsDcKIM/uC4ypRbvva7JQ4mUYYEBMMvSY4HaAverkeNCAB9O+zBCgTZn+eTvql/YYuA
bE94e9VgZtzbIpPnm6RZKBmC7A8+v7GQlHsmakoHpzYxGzApf2FzbnaGiNlMxNUtaNeDcD/rk/ns
OnafuQd4ozeMNceK/7BPG8ewiCsI7TlYfU7QorMJAS2usSIzMgbAfsv5cNq3tpwJusa1fc/C+H4k
OfaOzpMzDz7Aoitnjkv8QQ9LqxtuAEk3LbMPSkyMkhiz+1vLq/xLzjibIdHBbsFuULusml41XMFr
svA32exfubJ3anPJj9ZWF1Ha/amAu4zDANJnEBLaJdj/fWzZqC5JpEpfakM/E1QBo633T4Fd9lhP
ZuBpavmSolJcV2p3+k1qTV4asSU26YGCiOWu7X4/L4C3geimvMFNKUVs2Uyi9X6fimAtNxzOeLHG
BfRu1Lv2XInA6tDJUgSmdVkO5ot3BeumqdkEFjKyGZ1kZQUj41c8C+o1FbERvZoY6Kk/DLZoHGea
3Z23Jx8E0La2zWrQ4w8jntKKDtV+bQbaQ9uxQKKqeVV37dXcuM56X247ErbaNZPdXgGOtlNYZgW4
zmMn6DXIu1WnKjUclOh6495iG4OQuEAj0ZQZ5HTJYEs7gF8q9N4oPu9wZ0rRRjs3nGax+Z8UEmPV
COky9BIpBxms6OeCKvU46wtnCkkOukOHQXelORVdJHpfXJv1BBRuEL9zDb36et3rb0iabRtlVPiJ
60N/Ny9hltfaLHIf9c8pBmA5IFPmewEAY6n71tjqCAy0gGl6UBynuJ5j4ccDzwQvPvrE57CDG116
nYTnzZvFapqzOG8wqjHuVzx7WNpydVR831HooaMR5Dckm9pr0eNrEljUtwKvTskpqSz04egr9IyL
W7LOtcg5/bS1SXhA+hzaOOobgYnDhxwguoueW+M/jQVx1X4EWMvzU7/K1Ga+Yl6StndaBjFE/vjQ
Uta1ScCsd1cusItC74ErMzYLY8MrtuURtCIS8GwpRMQ2e17PQFJ+AieS9nOWCvMlZUWKCwiQ53FO
7Up68pnBfVSCORD4VVj+mK8D2qaILnNsxOYW20h5n5RWz5F2ZXgzjkhJoPTRt8IqCaESCjzX+HnN
Ns3BRMwTtrNoxJY7n5MY9FXbk1cOiH6H5ZXq7wn7GgotpVvXGTPtSY5KykjMwR6EnyF72X4RmdDR
QFSr5/0Djc2hfZ19e0fQM+2Xst3fDHA1L7Weayl2npcrhLLjujq5hulJwVA1dJuE4Sq3eCu7SmNJ
Io27jmupEc4GADZdkF8MvCoSwxm6a7v3mrybWmtKJfp5XwGq9yh6RhlBMIR4pHfJawcP4kEcGWEQ
bO3l/cY24sFsoJnW1xCiJAmorfL50l26kT6x1iI9rBINYzIVdjCGuOylHYmIYJyHAFg8rb/IH+K8
YEfvPgAzn9bIed62jrzCBGtsNQ+E9a0RlvuTCeYcXKGDg8xG1X9jY2CBYZIPO9VHUGya3RLlh3w4
ALPeBb/HmbEcZ4n/mf+yt1LD4pabgC+NxAJ50LLsOjZJGBaz2zqc1/+IacoCz/gcPODlkk+5nJZm
i/5+06lpQ7talkV9KxP9+5gYymdxnKXIC6MQWiwwRFteMGfLTnhVilav7N59IfgRN4Zh5A9Fi81F
gKh4xFRER41Te+2c+yohgv29g8sy6dp7rKyuSAwzfhOZqtlzadtSzC1BdcaGM3kmBxWXHIzCk3OI
qYAuU6qE6JcN3GQir0dggz+FkIzD4EJd5o3u5VfeZIyKvKO1++cWvfjzK3B17msPEwE3T4O9euPa
IKsRDG1rK7Baf9IbizvvLQf9GuhWqUdnzICe9ZX34GZG67XaiJ8Z5hMFbgnWmnQgRwwqcbh8ZLX7
ZDeDKhU4MI1BuHFt9UFYUxpCE4Ihnoxh5gjCujtB82ghym5OV1f2qDLcln8rrQzBrESLJjhVVvmw
k4qM6SRn4ee0bFTZ7BSkBSo2UGEW0AQa++zuo8JnRyjGSWSXtPrI9oyPkxeDeFIlc+yguyTBN8tp
ErTGDMIaPatCUJHFC3Z5xb1lDVi9Rw8uwebc/dzOrVUuz2QJxfeWHCCQBJG907jcIlna7bY7P7ju
ZXGfLmoHFGnzeAzD76ocRglxlVYJk4AHon7plj2KwVkFDRwRzdS3/sHdGppDXn18ZKCxpihAb3L3
mfsQBUEz5+z9sy6G1O5rXR74E4UeQR77tOcWVYDhRWbSa2SNdEztFMmp8aYrboyf++ZaKO+dp+t6
Paj0cqAl2BMeuqm69iNCqTZ6HhCjxlF2w1VdCfyW82fmo9XehCF+zO6GRZBAG0z980rbe+YsPMSL
9Qk+hUdJWCGGidDWCgInPOTi1u0j4zGcLI0p8+Pr0WtEJcWC+aSX90fEfAEuwov/5w07rkk1kiom
xl/i07UN2Ef4zs0HOVo1j8sr/H0YjQ+KqXIASrCLqOKtRUefVbgVevD6279m6QRc5L973BbMzPmK
qc6YV1xUlohPXvuAGSoQvbvdAxeVLtDHGMu3aQqznn23s5sIasOKY+I9Hnp+INU6EAl8Edwf2wjk
HV34gg4rsstdlYtSOaaRkkjlvI+jWrorJymNkhY7YRQZATvrAqs310hpGSRqDFTFz7JN2iE18qV9
BeMGcpFdQLtIO1HLSVerV4VvPnVksQYX1dtpFwPuzDealEWS0ubR/MyiCDW87OZVXeZTGPezceCL
gS2ySVMN8V4RL3GD/L7Hy9GDWmK7Xy7/aFsbQP3gS2tZRmY99ev1KU8HxmsjdHaZFYOKQ7PL60pw
I7KF1gFTdYEfUuCaGHkY2ghMCJTAvhgN7cO6jD7xiLSJFRx+Tdu2JHgMCBPYbgLMJf1J1qRF7Vgd
GTzVTJp6/2d4zXoL4FtrZ4mfkajMuqEMP/nzzAPRgw4pYHIeYbKUFMI076fe9/O8g5O/7vFH5DDE
imzc6PIBq6dEj4MFW87i1Z58qW2POKWxpz8I7gbI7utgMOwHg0DXrU8Wa/iWj8dznpsJAZN6s+FU
RsCn/BGVm7lhy5ijR/qSkIw45YDVZxyJY+uPL1DavZ+LDUHUys2Ybh9wuNcM3P/88lrNZDFZtWj7
xVtUMwh50g95vXLMEYBSot+DW9LnTCgDZGfxAR07IAdPLOOletc/W2vV1B6hOdlFy2eeoJpD5foH
XIH+vqJEmugRMPMyk2B6VWxRj4Vq4rIDOrTeGABTbBYJPrYBG1mjFuMEZdRfPv/7tHT447NiLZEV
/qUdesz0rgqq4QBokBs74pzE3miQJLvX5Fw0lUiBw+kZUMktGFf4/QOYbEVzj8jSTG4swW1SQTx1
zqEqJkjQBpG9tgPJ3Frotn9RW3DuLUimGR1z41aq94ygHRzaMXSJpDlKUgTaY8hJ/zX6Vj6ycfZ1
0HZkHv46wvLgOYd+n+e3obTv1qlOLuEQbhS1Q4BrjQXFNDiZGMWFn6Iu1HSFRciMBN5DZBw47mD1
uaI32a7fMxakcPJK/nfaCNjaPnJT0bPGw/VHFVtMcEsHhARiRddFwri/FL1EDbBsAm6bIl7kqTMO
kNn5TsdbxyDupAYvZ2NOhTdY23apZWTKdnUvQSZ+P5KcKXombLRKaMniq8qBPwu8O6hghrHz5gvU
HjFEJGtQN8Lie6hnOMriKH2hWyf7m6RtxYqLc/7syiPK3ZI9fo0/JVP4Cq8ZKqjeKFdbf01OSXtM
0D66IRpdFxCYl7LJwBE+lam5dwaBuGJT6PEPgIZyv/kzlcizj/imbLQNzusG1zbpy7CMHHuj4BVG
HAiFRcOZqUO2Dc0YkbZJMeIgz5GxlxGl3VKSB1ENcgiUu1yhwa4I1WO1HD+8DUrl1xNIvPiKAxQp
2jZBWj7yYeJxpYN62P1NSoe6UbpzKvISzQOn5Fgo4Oj+aHwi+671TU58H3jaALi9E16VTmVaHpKu
1WBu/PuqmUjclZQ+e+EnJ7qVGiEzWwi+yfBVmmpK4njYxBIdUvGOLzjxkFcdqulyd+Vh2xoSW5Ey
vB1HUCF5NCoYu6Cjy+4/UgtXNRfjIaKPVwuEqAarLEb4w6MhlgTHfxgqq+VCmSzgzIAWTePvZnsJ
/1M9qsZBD5ubcwoHRQl5iaRrzccAfxgtZmiFO7uCIzDBOMaI4zQY2z/bpsSLwUza2Tl3yniQOEs4
qIg0cX08ayRSQ9LO14+6ToJjvpbjXZQc4tosCOnct7mXZuJMJmZI3ONGcC3Lj8Rr3zwoAjCCivDK
+JsxPlR3l7UQKN4HrcrREVbtPaWxEjDFYRurZyZoeEwIN3cz83sYd97vPGlIcjcAZ7zehUBLVqJe
pALxT073MHmNIz7ZitLffDmF1cj+Vqx4fsAMcT7QEVDWdYy4jMPY6jDhJ3qz7ul77ztI28Rpxhy6
DmYEMRzOeHE7W7qA+VOCrm6+0IVJD54pEVPgFs6g5piF75wMxU5+P7Xpn4wl5IEv6hdnGUoWsikx
ZI3ywBHaLF9CBpiWvcX0O0IUok374VX6y2/Eivl5iQZlQdflIrx4xKJvBSrS6/pQ+TJXx28RiE12
yGKCEhfV/i0ZmHGlesazIYt90UIZr5I1bL1Vl0iSlAIB97VAa5R+45FAZIGwJRXLXLjXOt0OZWD/
VresQwXfb5z2PjRmk2YrW3Q10RATxD4BGztMPh73OfermGgxnsGrIGnm/yKgXnthgh+4xFvRiGjq
dUrFLwIiA7AVD0kAG/KOgRHU5WecCRlm3/7PAZAzjUlKVEPVV33JUcFk+t6OgnsGvtqa/4PB+KFr
3HIeKFqjbWTOQpoleEw3KNj4is+CPnS9sYktobboDBE66QY/23U6qwcXyIf5BhljkmUcTgbLb+FA
RQef3WCojMdTHY+Bse68sWqRq2LLk9JA4veTF3r9ad6/113Ld/SUFYaNTTM7wMMfttr3bgLdVLrG
d3OYCtiODmkFCGzdVTE2D/RkKJ3I3HZoANdNYSbHEzXoBWf/cNu09TvB43we/wo+ykaAGWjs4MHl
LJGUKdiPiTCwB2MS/PFZ4f9H1Q6HO3vr/ppF0Y8QQrVGj07fQN25PPW7GYqjAYx9pfRjOEs/O9VH
fojAgEcaiqBt1EYmlV8W1fJafyvusZqzXAJk6aFoFOSk1v+ozQp3G6mJsJVu46Z7acFYANnKrsDW
4edf5a6IrFtKn552hjo6LoGcLUkGcNRO0KFOopJs0xyiNkX+iDoPWtbSxWYDSph4RtZ4Sr/fAtYO
FGdxBO8ywefVf9I+OmBkGRlQrBd/fw2H5HTESYAvLrjPSmkn5zbyEhazKoB7csEMzHKYphgWqGjm
XM57BWianuLmi24cii+K9rr3ao1TdCSl258Vs/OoGzIwOi0D43LysKyrrap+J8Iim+d5QqTOi1/E
I/TrhfXNtoG22K44AKRjX6UnnU+dppYj1hYLt5qHbEV6qSMsS36ow4bWuXjU6hg4m7HmyUK5Ly56
KGS6TuIydGS5Xm7sf/8kbWacMyJxnC1dSMzZrk5cMOhxfljwvirXAa8mvKxErjg2vZUbjCVJv9zn
ohC/Q/lUSmI/BqucoM6tzYi0bzC1Sd+ybQAer2NBhqek97SMRTCmUohARXTR7eA7wx9VCxaIPOYy
olvlbILpUAz3H4OnsS3KklfsTcsgCshxsQ+vrs3dwWr+kpx8jfQSR3/MUwpW1EomWNKj0Xms9N4k
8HI2pbz6iARm6wGaI3GxgThxTJdcfxV1iTDgXd1fGdbzNeND29F/8ZvJ7CmXDhIU55K3ses6vb9P
FWBEv1D2EsShzLzf8bacvGsjiIZjIZTEfXWgCGENoefxVBEmsamARathk7J5DDWN1jDl9IP/cflP
c6sRD6J4So5wYAvlha8+2hYK4WnTwJvpb5jSi1dNwBO7GHf/ARsne79GRHPblFFzKBJH35zEsvMa
mEBzoxdTsey5KY6w8UA6o+4y39t98LTVeIMsWEn9XMeufMa4UKyJzEkA2nbAeEr1QTlhfi57HHFz
VsrMg43aOtiw/3WkmkiX2S+4Hsbqy8FABrfmdW4Dn4bMy1DCzOQnsAG1Iu7MU3vwu73KHT36qDxf
1lgh3DjgCfLupqwmVFoV9WesAqCsI+sksJ/nBPXwgtos0OXuARM5wVIxFQ+vvSY/SJF9nwXPuQV3
cNHSCBe/9TrnV+8/0OyVdRTFUYrgMZ+dZbaNIYxazHjlSa3FXYwkpg65rRWt3cs/RoEGghCLpam2
VMvlX/a0JwUm/VTC3M6DlP+Lv34KnFdI8oRBBS92EJwTQEMuAiox1blxVuIK+Yh+xEvb6+6zviSi
LlmVfd3AS7jyAxiTorgCYMsLOoSWtLaqQTjux9FP0dVEg2uq784476IalQHQZuECRQTiHg2NJJJm
A+ghgWvJtkonVxJfs6AXRX2swQmJPlXbZjXBnwZ4cb8M9wLcrGFlhr6fFrfxkBcZIekVoi9uEkWP
oF0/66Pa+FR0y11H5DFSwNI2Nq47h+c3LgQXUAx5OkcJUDifWx2z++9v3O1Av3HCrh4p8jSzzo+R
tVE3eY1h7MUgTqk2nRJUCcpsZXNfcXhX6UrJdn3y70wt7EgjozNiBYeD1W7kglAx9JKaJ82t/bpr
c7OI67x8DN9im2GLQXazacPFVfT8w4GytVIb2CPOHHPhx0afgsF03HQCY3Cjk9v0t+rMi4LJGLhT
t5Mfu8BWdccjAJd3h5/mbvUmOjaFgo7rddsp5B9Mu5slqFa07+Nz6/Bu7u8j06+Z2LA6S8v27NLe
l3ieFKIHA9d7+3PKhaAejfySPw/h1k6eU7V7E+/DHnTl2iqh08V6V/wAaNh3F0NgihpQt8vX6hmx
qt7Ay/k+551Yt9Rcgmqu0ujYaeqCL5BeyUZUY5sb0HVLkJhsAKREGMzqeeEm1EwKNSsfGT6AbSZq
rjDrDUD7JFSOV8ErW9OVh9l4ARxQ+5LjsRZ5MfWUmBncJ5REjhSx8ZpFeiSjTOrW/5p/aEoFEFVv
YmkVfsg94b6InFywbLs/xAGJw3lk+J1FsDsEpeLG9HkerYhq9N3wDZKHPd52cIgnInwJBTd6idy9
91VZk+kcgG+afwGyYSB3VDBeDMUdW/YnN7Ypda0DhfQ0FHZhIBxwHrm8ll8qHc366aRw6AY1Gx3K
GGVERWIoP4iaqhwF2Pwj331tzn6hNkLR/nCm4BD7wUQ6nFwc6uXpNvT1P0x9kOzdUoepsVonEx2h
FcQAO3U/crm5649q3+FSuGCCFcjJjsrVNvS3KcX875bR3l+H2jouijMUNyjMA5bpZRxk80cwTNA/
Xabt0QcIUpEK8/ZZ9ZLTx3uPHdkb7Y1PLDes5ydAvvSSHFNG93nnqA3FqTOeCf5wqvjbbkFfIfD3
wMK5sz/2PcgC6nWP3l3WAPTB/nN7duBswjCV8FW/Jn9blDmmbMy9+EcrTy3xNxjOo+J1fFJ7kIOk
1UgLeALdq4WpRii9X5iqMfTSb7oeyqUkQdP+1kKKg/y1sspXeyn/LFjzvKFikoXsWkflapOZ1KvZ
M86ofgkKZa4Ut2DoAQxo4fz7q9PuqH8aftGDn9kpnxy6UdgSxOJ5q4gFEpMNK6H2lk7ccozYKFVj
qCPkkHHBs7b5VJZsa9VBsLPL17tAs8PfBb5pQJaTKBYEcmvbJQqI8WM19soJpsa6prIpWFKj9x7a
WvfcA4KW7zhYRL22NTxxGMJ9fcgCmKtcmRgXOb0bdcZe61FhU5HB3vdO9YI9n5OSmstb7X8axfjr
CUSERdmasrEhSEq4UAWGEJWsysAUcKqF9BUKKwVy4Xp7cVoPGnKC8D29xFcweHoRiVXGPGjmEdwg
PFcN0EVVjdVp5PyCsdWIzHDBoRCJPUfDbham9q24VK+XUW4/QfqlY6Q/WgjmeGLStLy8qo0yuyCk
gQVfP5t3CbT7q8u7VSC7P4LS5olVwzaAe+EQ25Tr5ePAON0E/DKrZPMQoCoPH0h+NyNxwU+Se3hJ
I31cgbNyG54/jDH28eGVdbHCrKuV8/q2cmXxt39Qgml1sEnRRQDp65lxWqnDTeRoChGmZyjt+lOY
qTnBkYlrKHvRy06TT0ccSlFHs8kUUxBO6969njkyAgXnCtJVK7VItGZwKgG7JOGjCw174kKu2ig9
x14FhaMKPXCMlZrjTnAgEpKByiLlwqdoOergEuukmw3zet2Qw8Y21cN2BXtE0SofmmpEjnzMXoCU
yW5xavpKcW/o0vE7wl1fCGwQ+MfV/o2Pz/qttwSaaaepq/fbuLrWk8zLKm8yIFZb3V0PR7kuRr1V
tADfndWYo9jXrVihs14fx7bG9g5g0t0HVBSNrY40m4e2hKPzmOg2nTkZPHAZrjekR8vYMSkKX+M2
JQLb58wRjoJAc7g8QOtQehQB9iq8mfj1Pv3d882oDLsGzfLLebx5+YWTIqE9loiD2CwQbLKkuHTR
1legjUyioyJ1bll5sYcvnEC0qE3Mk7oCmYquY0LpiSPPhZ92P5H4xZMSHWrHGa8Wp7iyQOi9ojtt
5Bd/oqrkT7ojjpFd9H90F055JeJxgsZr2N4I9s/M8D44KC2GMM1XgV9eCB/ftqqIm5lRV/rUZrxs
4Ndt5zn7TxtnRTC2UO4rZKR+vL5LRau4aXjjfSgPu8Qgphw7J07FIAr/N8GKuDfAwNv+3bb/oH3h
F+tstLGVsubIPNvTZzG10rMUIhetbT+yx1lyarycW1lxnX1UjAPIxPDxdpc5B3L72vHbECz1/yWv
FPRick390r4p/MiH9CQZVaOezos9H8XPdgj+78sT/MkCGMyQaVxsK8X0gQbVhEjlFOZVJ+Q0mnCN
w2VRi6kp8/Ldj19ckUIwV71io6++Mjyu+xKQnIZMB+u1zggaOi2vaFi1KGso5nMRybJrvmaiRpKN
98ADjHE/jO7KwyHrIOagaqHlSM2dsefNGiOWfUdkiqgy0H0hfcfdMiCsELdylHw9ZynrqTEY9ipa
B/NGOb85DQcT+ZCPd1g0Aw2ofPw9ok4oHWMUAFLwPYNvqaCfiBnTodkjW8jNPX9zuh8zuXBNl3Us
N/HY9sPBsywfxL9YYouQiMfKs9BgxPNGrUnATf/KcTme43brKEtc+wuiQnF/uQLQ+/mEpuOt1T5z
D+OPS5Ue/As7UUxiWT5oCYrYFkHpAfkM81CTorCiIjx2tIrR6UlIoAAsRSWU2QDofgvvF6zBO4Zf
7LA9dV9RP85Ij4RKnwqZZ2AfD2U3r24J0pRsmZAG7B/UXkcfDxGuNja5QV+U21GrtlzK2NXETYOP
iESaqxQ4I6+Xm+bEceI43bips2XBoWT3m1dxDECnmbHOshSOvxovok8WQ9JnVmtOemapZqHJxhEn
mGCC46eQ6fDfK82kqT1RNMKEuIs91+cqKGcremMZ9B+KwFT0ozImDvwlLFtKYj2+eguHHRrrBsGf
nd/q4HFUzehxKxavM6NcQlTnc+MCPNlyO3crT68B8tZYyOfXEq0ZCW+6vS5XxzJK8fqxFVQRwcsM
CiqqhNSaIDUeLqyNqH8I7jEzKo/k48T6Av5/0/AdhaYn3efajTf6CQUwE062kIr9INTjF4RauIVK
tIeSli+oZ1b0gjmoDMFdfeEdytMVBLLTzEAE+B5s+MXA+7usMYgfrKyXHU7d3DIo6tNFPXMcdDRZ
WF11A8DieWHbOOczybP5kDKfOaocpISYx77+kZxwPOX/ztrxFWK/GE0xvNC1g4NbHzFq5MZxyfp2
syh1dsMVeIVSb4Dme6H9GTI5ZCSqLqvjj/SIESw2rtZDvv2snuVySVCX6YZg35G18/UwnPUJrRF1
GW53eyGywve8KL7XZFMMdNvKdBrLrTAGqr8c2KMsHFe3Tl9k9ggPwW5kEWWKiyhZAxCruPAZ8LSq
l/Ml5PVKeXKznBdImUUo2urN2Plh452YWtCTaNGG/7ERcYvUyX/3LEAiLeD2q6X/phPFSHSGDPhA
mSunxXJO7LbL914AKcsR4QtyWdMsyegJosHslNawS48TItdTvh1p8RrAI7nRn6b7/NUpS24DHUgQ
p1gELbAFbOzBxxVDyam1OwnpXOBr8d6sCGrvwzHqGcUs8ugLc412Z6o80ofr70uOWV35rAKS5hM2
jjbCUftdDwbgtZRVE9l7vyrhgsGpS8qvX9i+E6V+Ohvku3XsQvZALt0ysuYpTgM9/tjXyeE2jdNT
j+55mc9P4Qk7VP5Ua4w/p8qr4TLRl9MGKXzonhWr5nZqiI0KWU50QsNL7ZcgeGsfW2fkKIvQzdqG
WCUmbRaDuTHYavH4VMrN9I6Yi1jFgWGeJmpxzgDipus2uZ2mpTQ6ZbPE2TYbJ1iQW3HGnM+EIcCj
s+bbfcGC+qK/446oAE7bTZVC9rU74u5M1uM7HoiiqWOnJshbb0fzQLJvV6gNhv9gs63jeQIFoBOQ
aJMODwgseyal+IW7/c3bY7dFj4lUwEV9FHR7EAwqSk1TDEaFj0/aQd90F2sfp1WNkkl9PxwPPOp5
uh6PoKTM2SwvKSGsIIlRI1BwDeHrW+iDh/Q7rESFosbxMaMgqtHGLbNlSW/NDAuRFeUsZDrZIjkl
WfQjwHd2elu/npw9t9FzUE6R6ikaXs9jHBz67w91N8x0apdwMan862ms65+ixNjzeWAc0LXqwvSm
eB1PwfQugNVAC5xkg8SQyXnRnLK6kY1wHeUaSmj19afRLLqIHBv2IfYmpf++WoyzcwTS4Z7ZgSyg
BChJ0wtVkd4z1NoapNgaSJmBb19WPfrXub8pgmIwJu0O143tRfh1xSR6R0Xs8zME2WyBqYW99W4u
aeJYQ3O5cNO7tveyMnDfxSskkp72h1Nk5OqrD/wweZQegiUwJHUtTAyq7psHNRitGBgCEM5Tugie
dlDBrycfzyFcSTIqCL1Z1bm/1cKytuoXxtuw+EAhDCXefR3j+ob+pENJURw+zqEuIuES2tpAw7Z2
nzLAQ67Wxez1YSnUhQVDgLNopmzNOqTO2Xavq0NBIlYjthSqHNv9qrcCzYHZ4q48SBbul3zBYSdF
iRGs8idvnEH/o/N/gtTmUCb8dnwLGvOQlvMCWsyLZWEfQ+11PirQnu8anR2NfHvtUAo9++Ws0SRJ
M2FFBU1O9ACEgbWhfaQe/ubrEUftfFVmIqxnyhsY1cB5Zl81Nq6t4jkh9wsvJCvs8/Ng1KRLxkPS
AoM3Ya9yVuJnO66JPtyEXylElAzLiDPzbJHbdULxawF85E9iD0qQ8/uIaxNkLX0Kp0y9+CsOp9le
h2jGL9wYzh5olJhSUd0e6yxW6dD36J2iKwCUVdKYWOyYRRbeCzE60eRtghu01Flg5cTCSLkLMUab
Exo6B7DOvNblkyOmrYefwdXg7fUq4K9XmRnDid6oca+wUWV1E7LAZKIHfs0+4TXFvRLjRrpxEqmu
di5dihhMdw7A6RI1VL+JmofYzcy3zQrvKlpQXOCmS/1mGRJkznH/x7LvZDGyOnIsuKilBKGJDFuS
ZLBQn2n7mdNz1Rg3DngoTKaCND0GpbVWmtdsW2GDadNa4ZvxWDsp3EEQ47Bx0VrlBtUzi0v3uWsL
AlND3V+LjMpRLtztl/WqeoN2OvElgXbYBtB20GqrcpEtjcmZ0cmBk7t+qVTyDflrKiiTpJF8BUUk
heBt/fe6iXqD04lFcjoA7yMWOsKxeg28vxOl5Vd9fAx2lABYJ0XpNDTxvuGsDOyORzRewBb+g92E
g4LXPkNbjHtny0B7/9EHMMXBXwjqaQdDx7nU+0k5FbSb1VxvVTq1dONbtwaPL5uy2ASUhC6Ja3id
wbOSFPUpWqbyA7DXFIjBi2Ihz+vNMrWOVizfi7OYPGvkZtuPJLQJ12N5PlHDVlqUOkfdRnAyn+eu
XVCfZX+uYx1seyhthMHTfn2Z0UuVRFrCsTWCbN7bNF0XgXPHDm/N25JqkXvlbDsPeSPwcqHZgKml
uesQKPxwdB9mu7xwbglNaM1HbcKs88Gj06NblwZtsREXLPcLxiBxLOcNWHZ9lzmq3cjIALShXKEb
dJ8FH9E6YX3dPaOYk8drRJqSP/ZBjk0fmeNNdME8A7a8VwD1SmVAoXh4fXbMTZw0/R1gZyh08lEx
phNi1nl3pWD5MVBe+vpVXilkwSXHwBpf/g/+ejcB7BFLX2RW2zRN6Vu29V6LD/9locxThE9fQXZs
xGcd/iUXp0Ici8MbF0mmUy+M0Gd2qexhyQMahSlAnIFRgI4LnMWOLS0ymkNGlAzYJgrIhpHpIteK
kqdwijupErzl+bPw9/5BtHijT490Ziat7Jk8IoN6FEz/aGMZhe8UIehlRvhlMJcjejmOzFjlvW3u
weX1s8HJZLaqnW92OhgpHNxF8bz7j9QsdwQupzgwt0wT1V2LUiIoExPzKW3aPI4CAWJhesjR65ro
jUxwcmq6GilgxQbSqBfSDUVxJVFmDiRNLXNYr+DMCavfprsL8Vq1MOzpnMvdNGHAc8Fiu0UpavlM
tL0vT8Ifz9zxsgCtgQdXGbzcYOI40wwXj+8fMlpSRDAM7VyWURnCLk0BmxkWDYXQdY8hyrl+LsbC
2kzFwXifFJHhZSW0kFpfqXdBU/h80ITRAOg2oeMdWgRvpymUs1kofTFFAgAyYgeQKLGbQLViDckn
C3o6Sr/PVKZ3sFjzWQ6YVmI4Q26K4YJAd+3IThqCNNfnBIprczG2tkcmGk399A8cUpLTvzmcgRld
uVnBp6HBxbZEqI7Zo9RnoM7vJIcD7cJhF4RQrABlJXJj926pj2S1I2yGcaLbNG04x8mRKMZwfAfM
oWzUMpPt0EXqJ6G14Tk/UK4G+5yI13AvSgFfsJPidGnfHHf8oKOCFTg7+3WZOyP8dLhduvgTqYjQ
cMzy7Wd68Vf23ZCnT3IvRqYwL15AOSpnkdF9e4KV2GDSdt1bJC6gBFdhmawyMRjh0FJXsfcoyoQw
NKZjW9wkZjntB4FamSbrvwvtbej8cGClL6p1z4C4VqlTQtEslSYoXqaIAZMuIEOh0rCUnazgE3bn
4Z9aO8RVCLuH12nX7kVyb7iOa5JwwqEiHezyZ7vthRfLGd7PQHltkuZ1fu/7p7CrBD5F9HQRGyeY
c86hjpvtr4Rf5OGm/l1UPwAoOz21fYABtMH3Mc2h48GULR14Nd8ctM2MBGKdz1ST3HBpmXZN4vnK
MYkcYT4vYIyTtUrfMsGsLzmllz/VhKIzReC2FRKFmcyhD9k2vB/QqbMQf7ot9EMXJ83IwTOLDk0T
VLtkMyLJaTVET1D1RVREH2GY7tw/ER214eWhcciFEgpcZTyx1z2EmgfcnGq7jMh3oCoty/7WrNUq
ZDfJRIQaPQ0HhDvIlQPjLQY3Z0HyKjDYG4HMxp1ixIV2dZywjdW9TbZPipWIMYPmY+JwEqRUx5r/
Z16V8x4pyFjT/o4meQNznVpkvQkZGDJ1qTuFzxRVCT00YvuVUCWoKeJL7GdASvu1UeQn14VTpjwz
Z5Vm4+aDspTX3dYmn7u9YkMKtSkAj6tKGy/hqeSjUwfH3EUzyHsaMpnm++h9vYzlfh7SAXPCJDq9
0qW7s35GTYfZkI5ZKeSV5ORwmvcSL3UDDOJ/VAVyyjVQwf0ZHmh71tTkm3Tg4ISG7CuiyyxVbuaR
o4pjjTXvz4BvtwgIE+RokZ5FtPeAscrGu5Z/y7qxxhK7gcOhuWOM6qHsgGYGV3x23WTKtCCslOer
lgE82qqMffZpjXqA+EtVt/plWxc9u+oZ7pfE7ZkPwBbAjpSIN70/MRaTqU1CeRwvDqvkUtyEzn+4
+j4N+4dPMcd3SDUZezUuNI3xTtJ8HSwRNjfth0dlmklYtlQgkdJl4kflk655hV7c+bFdi09S267g
x837HwwyKIpQHfh82hk0M/0l/vUtjihYI9JuyHdvOyc7Vka9RUBeQMI9v5KZCgjdxBmKwJPT1fll
MbmEqx0h35IMyCx8wqHyuiVRSMZg0uKWxtoV6kERiC1cXm9WXgYNclE2Rj6uUoF5pcPPwyi2tRj6
K3Y2P5xKfwyeHS0J9YXG+DTchKZKjZ66DT5uFdTMtzVN874C3ivPO2z71su+b7VvV4fTjacTyETW
6fI++ijeDLlOQ2RS2EAR5lxJHj0sSElVecxzYhkFrDN3RL+iR+xZV00WdHsePALXnoFT7g0PaW5P
J2vi1d+b7hh5UFO/WmUKqhb/iYkfItV0XRbjmr1Uaw9G3VaHvAq/EmgNSK/h7jABaEWILOQ/bfXU
A3iuFyVc9hzXETdJNSA00EeDtYTWylZbFUHfiIoKD0ooxW2NUuhziX99tFP/bvg/jVriTdU+eyuC
v7JCgJC125/KvoQGrkqC8+mqWJdkOVyTb4hLUovrtKIMohucaJuN+GOsD766GlLQvJOQNto78Ugd
163Nuyg08HRYq+oWF3J/qEJxkYq8WFNus/l9mXvKTe3hyfg4d3CCinFJ4BOf3g/7K3k3Mm6ArYBs
tXU8/GX7IzebvXi6LKw+64on9T2+zsm3zbNUs5EjiHpl3V5k4XzkOQsCK6W7nbg6nJftwH90pu4U
2J7JIkNa7/j1PYTcEJTkqNMNAHD4JEfqNT189B1uYXyH9GwL1gdD13OxKAmZzNo9/f9TYm4BwjM3
6rnKsjdXvN087fksfCR61EoCF0H62zqr8cgZTYMiB1v10vQSSTxGwWZ1PQT7qzn6aVQz7G0zMaRh
JmlMoipIiZVLntFgxeIr2iD6WTAfYNZqA7xqHII+q3Bg5p/V1zjSkvanhKCmPkLZ3SN2wYCF4Vax
DZg/ByUz1q/KI3jVuW65b5IkXJlFxO//WqSI2+G6zGTZPpKKURJC7jHpQYf3DkmdHj9MeE7+8hIc
iUJz6mATOOjzJmARD8X+tUX8AEA+1nl9rWsvA+f/MGXDu8cZ8KEE/YH2Wss/BnsfpKbJWg9f8AyS
Ril1Zx8TNngU0nyuuvhHK+ueoUR2Dz2evSMjYudXuuulKZQmzBF8FkONPBEaPq6Hih4Nm+XKckSV
u0r6RRcTucvzGRFjUmIeXk44wMLwddMsU81gwKC8zDS1iAiyu6Vukn905TdTpH6FOVmlbmg/zEYp
pAOGUbYiNpoGXLlIJ1hhVgNO2O3coWzxQ1i7aI0GjNrTr6ZAOWl1p2kIIBvL10aicz7CWvmMWLu6
drZHWBoKuwdS9uz7tAgzf/3uyzSXeCJq3IY5EvQDIWs0StBhScNgKDAxMEKIEbnt7z6/AHjcXDGn
5p8yBu0hisl9WlVQ0e42W10iq5XsLMmN0umFVKsA5vOHp+px1enI05m+FSBRa0/9SvxYfPcqZDWD
w8gsvITfPcIIsCBy0UygYFVu/XcNZ8gxZK2exX2vzKUASE2uxAWUNV+eQLTaL6wH+Wn0/GV7Apeo
V2pJqZ5fMhGmzzAHjn2x9tayFZ+6+54/fk5dqhk94MVVT0jb2++u5hNUZswuxuNaYZ7QA9V2UwVp
nzAQ+kdKx53RmftPy61IzPDuh/VLf6K4yieEqMT21/xD703DdzKr7l8ypsTZBuiQ9cJBbIR7U6/S
jNJRmAuyuvngd7ru9xxrmBJGh4yd8VcnPqY77OjouauTIDoBEsLXmO0Yq5ZAEPs3dQ4yS7DX4i94
xqp56N2tCCzzNnnvRPSsElAV2Y4n0BfvuMCxVoONaRW7zlSy6SI5AdWdA10YxA2VwSTD/jkcMU2p
pJX4PGl9J8n+0UFGfzpA2G8YHU+hJw+pGCrreuCQ5cMk7QNCaCgeKh8i6IKAM9iNWuP3e4Oz/ooo
rWwWj3vmHiV26UVA9HsGeRk31v4glsEIUjGt9/0KAI5oZm8UZ3PQQLLx3TEmYeRDHyvarJiH3/RG
PLo5IYqr/sl/J/qeihd2+IYpgRmEb1dD2hRSRbSvRBw4e23sObmZ1DEQtfAkUYdE5RGYQlB1pIex
W83ffF7DWZInrWWBHR6QCewA21nMbU+8Y7EHuTaVCzEI4ggoe0PhooUIvy3LCAIA6K465c88Cw3o
t2aGqJc2Ff1wTcwhposJ5WFS9N5jKXHMJx2Rlj7vjAqqabWODKaHFZdB6cepy5a1Ka90c/CNaFH/
ZThSkmOzwMkG3kVlxW9up68Pz7N2LgLk1K0SBc++BFW51rKaGUmJlKssJjNvA2OXwW1HRFlhRGNn
GQO0ayTU0GMBFu/ybtFIb5ferGxT2H+sZ9GfvusAqNJX99BYYhmrDDE16K/ATtxZfyywb/POyQKl
moiyCrYonScEyOs31KJ0WnSNS1C4XeOhERYGO7KQVm36RqlXQReHdogx/53srnwj7/rF6hb5bVRV
MVELZgTvTv6RvnLFvuCfyBRhyZo/92Dgq3BchmvlfMKfNruMAlLH1qNNeG92pNCLb/i1QvGecyz9
Erefw2rk1nd26vamETuFYHFVlqam8tpjSU1VNX7ApNdh3lzuLuTsovZpnIhjbzf+/y2OmdCvB2Mq
5DBClzS49FNuzUWZ3/p4AgaOIbQNnUZ6xv9bN1WRLYxbtFLSjLG4THBpfYnTOIOF+tHcXssp6yr1
vIPZJDc7SrFAJyyCNYDkJ0LYd19zArcEdCMLhAnaV3c2gy+rrmFG2PEgPUxeQAQGVCRmjrrSdVXi
ZH0PdYI1fJ/l25ULfE8ud6IK1m8RYkrAKes6S7DqQp5JpYDwazHa4YSPDMid6PME1Exfq1NhY8Vs
7GlzH5eZC3D8/5GnlCPe6Jhij648jBMA7TrRTjHxWGx8vPx1sNLDJVBhSuvjzjFbs8RIEembGPEM
1e+/131ZGKcZgc9K/UihXaIhZ7MWKhzGJoUXz30tBTh0JrxfVDqW+t8N1HzSKUXF5csXowCjeqn9
4c/FUElu9bE+QLuagMyufFilPi5SBxUrD8Oeq3tZwabxmeP9ol4LVzVHURN1nNz+sottpRVP9ePZ
0srRzIlKNwHUf/iKGKWq9uMS1A4TYW/DPXV4AR64Ka77SIjQZ6t95t1WspWqVk5b5IqmKHrzPaoM
tzCyQ1HuhT/1Xo2x9xYu3KhHLyGN3T7HHLMzEzBHut2SAwadn1vUM7fvFooVCts5WFezgB6aBpz9
RH83CmcFfhVC+60WxorhfVVMLL4WltM2hicb/8SsfpreCR0MwWLw602wANrMo94ENBacTzpSliLl
Qe0mF4YUHz28+tp6wKBhwuVT6fV+Rv/P+NudvqGC9TSV97jEIleJnJ1jDZKJqsAw0/+C8Xn+63Qg
NTdDbOpT1kGxoSk2/KonX6MMV61WXJyLgxARvmXVQPSQPLYsTwQMEZb+jJP6dmnI1Q+OWJ5pMfKV
PetTSN5Y4k7We8Q8WPF2yqrd+gjpCDvHwaFXsHxGxdsOzAZb3vO/R6VhDUiC4fiFk9BXd4BbGYCx
JTpAvOtoxfHyivZDxT0ZcqQh1wfslve2Pv0YZESBGLj8G6CER7V2esYR8olttqiqgdNBV3fxY9+V
97AP9m7tYb4kZuQ5khAWodG/z6mdn9ory73pu4VsaZyo5ImZ2CD//SAj3uf0OTTIlI/PHUg1BRB8
Pp5Rmw3MqYS1KOmznXCjXUVJ7gV528ixxsD+YzJL7cfzBYBzRbhWpJEXOTkuGDMalHjjaO584kE/
JezoeSSoUWP/PTpnqaECNrUNoWpPN8wP04F4HloJ1WSuRNBL4jiuuLsDb56QSPbaH+fMTRNWl9T0
4Nj4pv99YGLxAqWhSiVa2YrYOIX1ohKXm6lzBdS85jKLZfNwXqnxz9FgaQE95lYe+BsCl2da6YWP
PyagyJ7atcpSjVFcgAeToiEHHJK4UYrjsSg9QDQ4y7qmdycHH1ikHQ+qWeWPA6zI6GI8Z+q584gd
swACXWdyoejB2TcSDzme/ZaFf4wfE4bT8x572P/RUiknBlV3K6iZHQnB10ZofCwPzhvNZvKSIYSn
MBi+uZVpJaBgW8s+bYe8mt6jiOp33YZNup/ec1802u38O+0QZqtVZx9y/axT73FoaZKbjUKZ7gpg
hBuHQTk7zm//r+LaBng4xKX6Lobcm5b5T/5NUraNVmDsRMBC3qmJ+J7Ri3vlMx+KIRp9Ssg4MO8y
ndnbiiwrKTIHtt9PQJDQh7eqCNZB2ZfpZUB2Y+E9fcisWmyqR/h5hrDvJ30xnmmhbrw1G9VllipB
cCtXOC0YYAg24rVHnhMgfP7Y+HK+QabN75wevYnjMSQu3UoF5eZbl/f/7MhTIfJMezdASza90FUl
AIz+1fPMD4B7xA2h13pTX7ab66y3+WtTEteJ0LBjXbkjnO6a+gab7TS7kU/MAk9kX1a6xkrovmp+
ZmXCaSi8uYU4p0331MPQUEDafL9bUQxa6KcLNxhnsDBEm/eNF3QWmjcxwketf5guBiMs7j3tJcoW
RKbpANg+O+RQk/+yL6aASlAqSJ//LqzF63du1sPI06+EjeSubkjZmOGQzcJuU2rIEh+VzOC4DMKG
ToIWcHa+vc7dQ3p8oaoCC93nOKHVijDWZqiyrCz8U/WrGZeWISdjWRzobLTsn0/HLrStB83XKAbi
SPL3l/No1LycoAKubt4Li5BG9mFljhqy0/ZLHInS8adAmOabVRy0nTnrCU8iUPfOH4EG5/zTEQAE
yegpnaWpsTt4IUu9ror+Nqmq3xWT4gBOhjLMj0fFQDgUNC/vEehxlrcpHoRSfQyCw4OPKH00z9KD
4KsAAojVs1+0O3qtqb1x5v+723zoSpd2QFBt13LwgocOzLzHx55DVzLF7YxX5IP/3giBWowaVeaO
x0JiXAWh/IPjVMVx7XD7OeOYG9MdQYAfxkpQvyl1tdnRYkqHxHnNS3ByUVnKuGthRBSwXcSIWxS5
CnnLrVmvsGjHol85F/L6U+7OHzth5cxz3oYSYpdu2EN+Q4vwtRb5gwBu3td0wfPfTchymTnTvny+
Wd8dWxsdCuJ5C6c5K2JMDAjV4Z9SKzUr7KtOOPZzM0WqjDP7CyO9TSi3mu40HmKoOT6eUkMxKWDA
yvyWOO7oiGS+ym8TcTlwpIH7+DgXWqx3U3zqV1mrTuoa86HKp1ZJ0s3mxmDaYNXiIfg4KViJSpfa
5e2T+8dhqoHaSNtDjuWLn++xrC2aiOTE+PR0T2tsWFRKUUehRovR/3ldjzQeCJxdXEqXU56btXp+
gdsSZOrZWavS40Yv74RCL8ivjLfnkEgAvJo7wa0EDdHbfq6/vnK4/EEb/LI+Gp+KysK0VVx78ydf
JqbdvKPOL/i2Tae6K3LIE86Kvl8O9L7A/Ca7E47zBPGH509tmxkwfYhD1Fp14eNuJBu2Wgisn+I+
zYoPWdW87lWrNJ5F6DV1+HAyeIj1P17JOg1poxh7U3qjJqRrkBC4/yFR4lmNHa8xexqlihVNQTEv
FwmX/iUqCyfdMEIZmWDW1DZO2mGjoJx0UwoCIipTsBenEPVW+SsQjNM0LFQk7H6Igu33XDRKmk0u
ym4WfPXmwfjpdog3Vq+0sSHmeT5UFcHiv6uYsUxeXe+lTwNqHF6Rz3rgQpP1H843UIEDiidd3jbz
/iU2ztUKjqHG0HjHriJEbf3fHBG0KjXMO3P48LdA+4hw/SnuuAxSNI6rbXV9MdzHailun3NDH1td
T3OzT84GW4vAjIQeSMaeh22ZiKu4Bx2Wfy72eoyyDdFxPvqnhxN4goNTWWbBrq9ulq6VCbVg2xmt
DkzYNc/N3OwJxl1JZuckI4/S8MLrteHvTxDvEE5efukJURBYX27sXxNZARKeKnzzgD5BD1U2xznt
JHnVi2a4pBNLRcY8dbMdBvOW9AbcyqQUdy/nhde9FMUTIUFh58ulAghC/chnzxEvphB5eNPr7oV4
BYMCWiaCR+qeSKdbeXwnUonlIXLxMWoMZzh65aoT1wxCglPBNA5aVNG1ezwQtfHjKdeO9QOxrXX2
kVBtKIl7Xj/0BtU/z1d+y2VU3qBS1L9U34gUBJ1v+xk5XIBgcqezaqVh19nLvKsX1spGVfpZHhol
mZEGI9ayC/DF+kLTWKCl4P5U9IcCjKI7yrBPvAXpeqSz1mFQNdcfpu6dJqjTMJuPTmUnWOc+NdBM
q/73fCLSEE/LNjR4S8iBAyiGvsfYqGd4NNLEZikAv2MWokASF63LpIby3eguwe052/Fg/F3rnRMg
4aeyz8KdEVwxCzVL8Blf4DuJa6qTMIuP+fr/UuBsZEOAXzMOwza8Vb0WhnNFISeC34WEyfxNwuyW
JT2BocBjQSag75P4H0hINjlsFuPONXL96AwIzCtuS0bEoxVksdvih37aweeJE3nDX0FdOkZKvP4e
VA76NaiXRZvg7e5VIaK5h/fLr9qisY8wsG7+sUxtlkIR79PfJfHjCktD/PnbFRD9sFQYQ1ZFl6ej
mXit61s0Hoktg+dtQE4qsqy4CRzF/Pg351kHXxAGwVeyhP4RgQsXYy9ezRCH8+F//Odpn6RFBDrZ
+fRKAxUisz6VXoGHeaMfIulhgyb/25BlKljMi5F8NFEtTqqU9eUL1WOyVjI9R+pjyfqAN3L4miZQ
NfBzsGIK2+Xy100p3g1J/jxfjBzz456biUbt3Ixuhdgu0bgIUwyTqAyWWVfo7hD0xdVY/FsbAM1G
yxr1ruqXJM7g90AUCegOWm4gfyqpvf0ann0mjK0GSpTitHuXo04Y/wBdif+BqcyBRRxTNGB4LL2l
bfCvI+easeyYA6h1LlUTTArLzgBJk+XJhdfu2T4JUqhL+ramzXqmBGSc6vN7LiMDIvhbzHFlQVrz
ub/Q6XpvxRCZsac6ae56nVwzrY1cu4BrZdjFdjDN0vhP7Mq32VyMsyHtSlgZSpALJab4KZaqJ2B6
Kzou1pQIsbtmkiJRJUHhbXO7uROuaRHQSOdQpWSvb3jRwFGrbN4vdLXsNDIz8vHEzg1VD8Y6bjov
OVqYwwoceCaqvWxVVTE6Wdvy4qC3XYKijoCye3AAW41fqlmS5hxakrAIWN1CI9rggl9jmXX07UeU
uEi5fVzsMhdVVOsMzn/RzJG+kxrAd45r8hChmcAfwX03NsDVvXcgM15pQY/q3qD6VWVlWV98j+v6
+sEvdXmtdgUswEJuuPBT3Ci/Ga5CqgMuUeIEIC1wonyHZ1/0BlDWmGHDVn6G2px/0VHO3cS4ypM0
RyQt7IjtnKf4Vy3bJiDVezT8R56wkMUBCuZm4fvph2QezR69kb7RrNHvRwcsIqVsgP0QjL4bfTj7
QjbBaLX9GELBzt+4NUmggdGLHYV6g0fcqX4CHejtVVygu3W+qEyeW4k6nE/j2R2OzfpxijdHf3yM
LoQftUWVbyIcsOfugcOT9lZ2AWmGUD9ghjKHwH/TI2vNU15wW+gQ7w3aqdJAznrpvFx4wcuNiZBq
Ps2VMcqg8pOnb31ivqHmNZAM3yxvsWXOBI+BOmlGuNqhl7K80xPzDkrvxYnRS2ER1QcRzGTxCchy
ROEtX77hw83ZT3NZtq/xMARqPlhcWjOobNbCreYoJj58THMj+ltIaKNjhBUFjMJuMiAOAAz+HWBR
PTRI11OeHCvouFheRB2QhYj3ImnGfmbHzvwX3l8Y0ASH6I76ocyBCwhPpBOmETthFoNMc4ji41qt
WK2v2KY98DPojENquYnAMIPGkg7OIntoOBOgGKoPERPGhEvwYa8jYrOk38cmljAOtSyhNTv1BSuI
Uha+oaQASByITn4o1yocjnDRGZHrrtTtruusxrKBsUL+LvKAh+9DOXob6GjoHMpd6rLsNmLU8QYA
v1Ur6iE5xUcvmK9lO92aSPXR1HOv02hB9fqPBNMgJNdHqW+uOzfgX1XVN4Ce/Ru6VG6n5Q6JjBps
Sh5hEQdql7lamcBDdxMeglNofmeHasRU8cajs94It2JT2vMcOv8o5Hl3WJ3zYUZxoyuhMEQVor+b
mfDc2uQrNNyu9utxZYVXn1xCgMx1snAXYLiqGseN+MHrHEay9405BfFIXIDQXFMiz7aim876ViC8
QSOs007Il0lCr+kD0DWzVvU973Zy10ckT2daxodfowEsAA15jdPw4ee+49bfeFe3XEV/WitmTPwH
2KVvOaiaCcOB0vnhlLMM8oCSURxWlpuDIjx88hWoI4cVscggaL8kQj+bjwXcMnria7KMZpj2Vu9B
5wIHr66iXw6tyMgQNZyRyGd6havcc//4goF70e576F7OsioXMeEvdRd2e6s31QKfP+u9Dm6gm0VZ
kxr3ubjjHI8hWo3IuWRbIPDo+T9rQYV/f2T4Msweyt6ym0E6fXWvaW/yHw2cB+LuV1clIw8VWG1+
KE4lAmSgGX1q6Cu8P9o/V5y3YsgoOHRJHMtSL0iJqefLaXmLRcOdQTobYN6MCkS0AUQlR3hQ+QRf
pvrYFs36NW+nGBEOr4npPF30xzL22C2DKTAdiUP3ruFvUbulMCsJ8vA/ESS98jUu6CjojvVlKz0O
ACW/wpeMaa6u0Jx6OwAQ8kBJmmMGTQD6dfAT8GW/Lhs53MbaYXyrnZYKnGL5XrfB2ed9Y1gfIYhS
3UnMHhTD7OBaugFe8Bh5+R4kQpuUWYfmo9fxoqAhUmlAGmVvnALjDejoMhPLVkU2eaSPgAAC6R16
Y7pSg0J2pEpNfB15+7KQhp8d0dAK2E5IXKOT3+4Ho61vYOpBlAOmQFZAu4bKtm5ZIol24/IgRz3P
hCEMJ1vlZNTCek5txglYxuE8g7A9AgGMnfBi3sk0DoprGiWwiGUmiXe0iPFGIVahJEF2aIETUH6L
ffrowgLaX65fIJScw3aREo025SV45O+ikquFhtoQ4eq0HsWRxvk8lgQe4N0ZHerpv5px7adJdojr
5vtnBdtqOvdHKLx7d4AZApwxy9uu+ZmBbeHVwdVr+GtjtE3VIhp/VNu5g1SxG+HdC09vvHchaTOp
PhuA5IXg9+22zVt41H5L1VYKT6MM+PZX2jezN2zghZOULqmwNuL+fUqJZjg2Txafp4ULBh2QblZC
7pQq/z1u6UAcT/Rx6R1iPae12KFuqqnqLlD1NB5fqBEzdYtApEdq8rp6OXzDLsyc7yepkXe8MYNz
BMaRGPF3SE9JrT4xnIFqzeWZeEqwSDKZEaqPhp67T0HbPlyoMiyREGgZ5ZwOlvZRj+ZA5J1zVMg/
HUD+Gbll6q2U6RWmBcXe5+VkAUjfHe63syFE7cs7gIQiWAPytLGMw0rqYTrxAeIYVozl2YsmifVh
hr0sQc2Pv17i58hSwOQpG4MgVFAgHk6JU17Hnjwopbf3IbwDt1TAuyLE31pUxZKpueG/K2vfnFFn
jdiAhOgK3EVuCyObadv3nRwbgNbzjbhRDpKvfx4dZ93wyU+uqG/UMPaTXej59ouloM+0lg5r4ruV
1/cwFOYhFz9z1Kd7JjmxQgNxgxOEBukHMmc2ySrNma/WNzp7dhFa2dT0Z4XUuLwzZfbJZDFdK1rj
mqdcbrBGA3vTX1ipf8JF9MJwMYdAtl2Mi9PodPLmBdmHpcmRKcJjuPZ86NJsEEZUIuc2gPLQYSW3
7ssU0f+2Q4thz8bDKLljFSDJwb8+0MBBWCkRcU0uy7ijmxaQLkgnfwVGeN4gIF4L3YUJ+q/HJSSD
CO/YX8LcNW1+GeBYQO4fl7/RRNNOzLN65c+si2EdLxqnq4hzte3JfuVmEI8A1TcOQGHWUv5SjhVn
H0nw1wFbyAIvO234Fv0XWrAzz0iDmBMHPMqPz9ohnF5h+4cQYpvokayPoXPM5dXALNM8LOnmZg2J
+hAssAfGk8KwV56pUKuMqUTDjPYA4thnHPCoQgvlAEoCMAUGcY+YWm8rhwC5A6rEcN1TSVXxbab1
W0/4wBfgAyCLnitEyCItaoRurajScDpcJi6ZEAVkJCG5EgOEoEaV6IKiyFjT+IBl+Su284wUVDrv
jPG1UrcP3RqTlbNpADVrg132eUsJ2N+aUrM0UCGR53mgSjESmV7tBICjCSrGJXz8nWXBqWUIeJAT
qRZO7CKqt1SnBh8KiJBEIYCHij2y1G4D0piDQOKSND9XULBYf1wfhWUSHcorFWJ18bN+kDGUU+U4
jrKKj23RfLZj3PRVAJYK9VXgJhT7cQ8qWXJQwUdILhjoEOgjtEYaMtO7Qb0An7JGolZR7K3NSF57
JANAUGXyTBHI8d8QyZoL8qlvRIR/0idyIT3q2/kDQ29uPD/M8aAwwkRM0nj+8wbR+d25Rc6r4gf/
Cl1ZNeZ4wz1xOS5kbrzJQqR71FCg2DjyITsvj6rItFoZ3qlRGsJFj6cXSHfmTxf46vh8vAYofMZ5
zJgfzaWrRaMC30M+MndTYk+1sSe3EzkVmzEwJoOj3HhPYJY51RFZ8oZodYiHV8W4bin5eaihzguG
yeSWNicxxkhgbbi2xrNoncGVTXXjA2RWHGvanduP0bhV0PX+oYHWXe99Zc0AZ7m6ihmEcs92Eg+z
oK7XQ5MH6RgPf5nV/9iy2nj4HKsowshRp6YXS5+UIrXaDJKe6HsGwd5jBE4jo/xjSJNwmOJk/4X/
JMJASLzzjiek4d+98LUyErKbb2i649aBpGucBJz4az+TV7e9WjRC12jSIbHfiAY7EnxKsct9saiR
rhZvTG0cdoUe/epz8eN0lhdQ32eVZz3/g6e4Z2v0ewtWLmdnPnyjjXf0mp5lUZYTEqZEoq32P14h
5tgIzyn9CCM/8sn02PX+I9XT/vq0pOejSYjl/QZvb967GSFWHvsei0kjX5Z3Zkq8TQ1UcAiWLkQP
dhKgfzZx/ps8G9dChHy7i9sM0ZJ7IVye9hhM3hN0buzPo7DoYo/dDmZAGcpQs6vaXeZoWkT4IlQc
DIND86+GNN8C712Kg8Ru5nd9v629SFwxrGMloPoPluTjxOE6nQAEYJRYZCXKtWpFfF24Cb+m+CWk
/SW8xyeP+j61Z1g/31hs37m2qU3s4+Chce5rl/VgnxLCLMfQVOjSv52ZeegFZNMiOcFq8nrMhxV+
udgMymboflyd7aA0hkGtSf1tYJyCgWquk4+ETifbtQUVgGXMd2RefEDIqTCs7XYo/fu6VtNdbs/s
blIvW5fr+bOPLxBqS+9RwK5S6qFv8t6O0KivZJIkPlN5v9hJM1JGzyr/DCEnrvpbth5F60OGnlVM
Hf5biMt3PcQK2A1xuM01ehuFUPbryK+6Eepn8QqfSx8Z3YKgBtBZ9eiu/E5faYb5DgLa1c10y5E5
SVfu11UGgAaQoJAniN+8Eijk3V9uIMiYY3lf1or0aKqKoWet8IGuPi0eNUo8wwnic3h4T+pZK4ue
pZHqz6kQJ5oLkT8Pes8gWm/uYiEti8jbYnRymSN0xgeKyG1ew5+2fNeAvKL6AeLOFSGMUAVYZm3I
+Fo+aeumZDz40CWG+ko0Q2cjDSyNaiT4vzSjUnbDAi+1TlKaKsxxpcgwFUuVTBFEIIzbB/Cd8DAi
4nXU46b2CaxOMbIKBiRZy5Df3xS3CFDK7HWtjBTBPu1IuJhafu6EHyoh9SJ9UOXrI7ArflKCCBrh
n9nWsDz4TvvKKApbuDiFDwYHt5DO8V+2MVl56E8p4VFwoK/JcUVb9FIPZB+76ZHWCMzGXFlyl5vL
IAum4aUsd6ircWMddtZfOJflai/BWAN6lGb4tidQTQCq1ebmaaHKzAWGceBw2Al+XP1wk6olQJbA
p+v71JoqXekZbBCstV70LWwPcTP1lScAkGX7BE/Q36V5hxrKfEIizcCSPIFQVBCurrPlQGjsFEcH
P+y+TPn6xvwpEvFn48LvCP9zk9vwxTioQfE4dxbZZ835NOTI3CA9hR7aEGcw+dDVdthX8QynTsmJ
Eim0TSQcoOy1uDELZ+P7t282ArzIYBURasUi5k/sDGRCG4YIRy+Zahkw69gbS4N17PtNODEnOws8
i5Zs2+SMUKKZ7QVD8+MeC7YQ2z/PL7rSuaawErnKoVnsiXH+c4pnigiaMh9LhHN56DNSh9pYBDZf
iBG35M9zQuxiVbmztz8olg0GsYVvjToc1XOxSRFRHJs7u2XUaoimfTB3IjlTy9H+WVfi/k7+nzVR
V7bAFPz+agaHfkg8/dQqoxmtBo7UfiSvSD+cJw+rQYA6aeaZpcWAnLRwgb5IoP2Z/1HapVHzQAUW
1zYKj9kQyiSE22kDyjj6lq0ePdkd/zeY1Qs9Y8tH4DpkL6YyU5YiFk+BJIcPota+/3fchMvzJ9Es
Vl9h9nLCx66LjKsdhBBvF036cSz2F9Ug+P7xQgBq59Ar2hFkq5uxNI3UJJAh0pHnkob/XdqnE7A7
61aPD8pdMAfEFQ+lkSK3DOcjTk5ezXGrVg6nMqG9J3W5Pe17DbGywTXsX+QleVb5PDKa4PIGZWQi
54RSmFxUkPsANHZ+neIWcLgSuEtQnsQ6uMrD+l7/n13WimqFP1YtjpGPQYMO7AlISQhxKgUkpr/v
LGEnmN3CnfDu+6HvBGMhbhzYDamx/EpTJ+yeSc+nBxIcHdAvWeoScfn8xjTh/113m5TrkAw0JrsW
KnM8DJEy9iYBGwPU2QCxxxQVyCZ4YjF3jz7827P2wumqdcSjd9oJ/YtVd4q2YVRLl3rGd7kUZdCw
Iy49LfjLlFWGhG+SCksKK/HVpT9yo4YShtmjptqjv7OMpVH2bOH3rGgDEAATrNWu/gJataKlkib8
bpFxzb4qItWoh4JeO4sl4xXA1DIN/d/0GdzXa46CMbXNbHPKzxN3pDeDjyysE2z3IwcBbVg3M7Oh
RZb9iewMl9kDCeOrB6x0qB/3M5ectNgcN1tM7f6Y3zUG1ccQNM0YrXwGmtcBgYuvA1klZOgXxuzA
LDT3JkjIRu4nklZR7fkXxRVnIX+JsyDSgmv1Q0+XgN7dhZItkS1b4MCxY6+huC3/3ms5ap1b86gF
GS/kWiZaVIGyz0vBHV1GLqOLOiIfheOTS3SURmWlX1kzZVxSw2LTcv0tMMhO73b8zvi6VT1+/E9Q
b1nQ9WoPfdQTg4Ch9duSH1O8lWLQ2Cnp1tN4VvBQJ3HjNSS4Fyq6is53x7YlFGawoWw8RHArvgIP
CGzB8v3i1uX3uYybIdzlTtImGrq3YVUqdWJQo6PXT2i70Uf44d6HMd6Q/x5MBzoPO5g/42KUhDFE
MY6WFbmS+NKqEekR+w7ioN0Vreg/82YmVsDvRZP/wNouROaM3jHH1iGKpb4lIeFZ4a3yMi0z9xEK
M5QxdkXqtP5rwBQusKi8ssGc32QWPaUXxkJhNvz6BrkDFgBK/uc80a/tayx1Fa5KhsqtC4GdRFOE
Kt8zNSPo9EAmkTZjNbxLiq+FePD3RW66cnHdHCCKlzywOBlC4KyHIsMWaAwf7+JnVlzoBMfDqIwg
fsRAVIXEfjp6L1N2Qmu1znGgSF0iKm6kQRrXAKmBOURqeYXmGFswYnPjSdEBU94j09AfNC3v3HKh
gxpKU6ZOVa2MAX5TxLxbgjI54a1LFsdJLhBw1FaEzSrP1FTos61WHwdqSZgfzPzg4fNe7ZQndQkB
PF5ArZ2vq23/YkkRhb1EUAH8hx8Y3wTk0rTScRAhV31JBbXwq77FTNHQqitIEzCV/Brb671mqJW2
dFhOSSPX/tk8thOWJOCd26AtbMUXiondxOXDqJATzmjMsUUX61dEWTmTz1eqdqnfxZ7M8kTfVoNd
FgWiSaWd5pXUDFpbWQL8po2wVSCxCB5Nk25wS3foKhzwKF8jZRjbZ7V42vRE+67nqZvooATUjAph
BZ/P0b6ggel12CUO92KQF+FRaLNxtJwUpbg7XPknsHHZ7EPTAs0bMkt1O4VoyeU12BPLpPrvyQ/U
vP7MAkFTyL7MB94vkmQdp/FbzJ7rcFHcJOjt2/YUUAfeEbPRASANuqnEkKjI+cPBSgC7fVNfuAam
px0LtjksoGNv1z/7ZoTTiDzt/M27tlMPXMfnrSPxdNriPmd4TZ/oB+mIgXGcs796OwYkKfIi34QG
6KqrEz5uTMTX47IW6IZCTeG1ZrvjlovaJX3hHS6CA6U2UBHGWpmNZYcwPpHgtfdW5XbUwKfSmLGY
6q0vQ/SuTi5ZOFBN2X9bF1qPVx3qYHTp6ldZYrbhgCIYuPcMfcI+NJC+H3vfZOEGvtwSl5PfwQfu
t8OOshfxa/MI10m+BuQvIiyfugEFF774g6oQMOyTVGq6zaMQ7khGAQYPo+ydV4ElGQEeUK4wqE/s
m3QSu9FqlPHVPN8rU7Ncwq/s9GCOJhxkGI/ZRO1+/DcMNA+OH5DpXuD0IIEVijXBwo0TD83pWhfF
FwWcgeF9rfA+/cHXIGWL00L6McswVrCyD9ffdzYvGAQCUK0rqsKQZ66AyFLRVk8Xx1ofw8qd+pfz
D6Yry/obEMHkfwiiz6u4lktvfvmwh7eNKc3GUzK86oIWgNALJTupOeEnrm1ka5dWZvfhALW6fiHT
STT7ySHuL8BVJo468DKuhdWHXuySYOQLi0YQ/Pnc0hRySX2f7POCQR1MrZt8O5lamcDO+Q8m/Opk
RC693ncp5IZ9v0jzU6q2L6Pk249sqO/G57TU972OYDEsp8aojqDt27E+3NtmGx2AIb9dyS28cXgR
QHXyvrBLy3x6NUM9OVH6y5xdZeuLWdvfDj3LBuUlOJLITzs2DtbfaHyvWrdVISuzCAURH5QA5aZG
aUmmxyc5z6kecVx+Wir831MQ9dQZvmIneYjNsk3tvrj2mp+Cf2O+d0fKFO0/WsiCS+6ytIFfhuR9
Ca69kbj5QRj1eOsW95R+p01BQBB+yfEnwAvANqhDxvbLOfhCwdsWKXqiwCYefU31GYyKcERCaTt9
DLGqCWlYtIF/Bwbi0Cq40k1L3oL1S2t/C1ghud5ps2iRPvPbqWF814NkR3MdG1jvvooIBhItasi7
4zX7yUcZuNp8elRNDulWTSTXke/3fCIfP9OyaNS53JKRMJ3Bw06xI25prKl4P/fGxGZkMZz6RkH5
qQl39+6YdPk5+M6fvxSE3AFIK2d4pBwCZBdMUioB8qZqdahbvn98Vmb2ob5mIA+wQL+QyQkWXmvr
IS9BUR+CdzIsG1L54RdqBzBVw+E8Ywro/FnFBlaH/sOvMk3YOhAZysrnMvv5PZpPKBZ1VOHxOye1
9q8rOz/2r+5bQ2yYPUtB5spRbDFCkl6/tfwXMHRvVEVPIqicJ0NmeSQ/x/M4XCWSsPZCYOi+Nutg
mP8JeNmxZFea+uB1NOAWYYIEpWby9vj5kHJIFNjSCL59hHpCdOh6INI8B3AscLj+57RIQ9QAMK77
xXLDFpJiUcOQuKNmAc0X9SxD/GQgOPhtrqKERL7VUK0n2MLL0pY+teMAgSmH4WdXVnCbhlBH5ihq
635gq+UORIVHhBPV3IJvgks9U3+qiNSPqHR+GeEX0Jl6bJxy8IaoIe4tSm6SGO/Ir3dS7JWjhYPH
gBKC4UgQQFr93NWEF4L5Nv1ogwGvXFfbtgAo+/brmax8vQi0+YGQyzpEEQBBdhcW/u+Y7Qabaxg/
3VBBBB93hLtOBTaOMKyaJQ8pStDUJQRLJcV8m9wm569XQoWqlJXYtt+T10XtMu2zJMlJ3vdtGDI7
UQLYlY38q4FIuO+OVPTwaTOKG357uiljo/HU8RLnfKX0vYWeA5rnugMIhrSqV/XTZhI0DafVN1ND
lY8tPG2muWmIcia8smWDdin8PKz7LHdc9nuALd5m68mWG8BUTzTUDozBvtoM7Z0xjNWy8Xmr5z90
XTyGf9C7KGuFy8ABpMtHK+n6IYOk3GA/OzjMxDtTjwSO9RDGUGCcUTuggCQudH3e0x3f6XHQnDGK
7To9L/DmgIEi7u+Js50dN4O8/onPvYj5sSMr8critNDDIGJRsWWeqO8LtZuUfBirqqkgn9anaFF4
qz8z3RHu08L5OQw2bXKI3aUadz8AbIfyq9h/BzRUHP2fZU2a45ljxGGtehsEOS7QpklRm/qlpt9T
R0Wphx6JJHq3Ur9B0R/WBHVsR8MFcDSFNqNflFSfCB9wCeCnxMqbZmRUb4k8G51UtYz3zIKkeN0Z
90MGua835KwJ2pt+TQ9bHV6+OLDLP8tPrDpXqCXu66LdPOATncr0dxc3P4qEa5rgL51iuQTzORhM
msVDdwtI1rMSABcAbooIkPwVrzdeStTyXUlQy6WOb91scxqnpDBKs7cW+XL53GcMIhBrUOBSGoiO
NyCeJUU7xWCHG6qsZAoS7JAW0G2FxrT4V+5AcDmPTc799vv/A+u3ESZEM+gSfZsWKOJk6g9tKdvL
KUT+IIR7RrydOoAex3zPXCMpciqZiPwiootte5WAaT/Y3mb7SR63ONg8c3C8Zx5/gha29xLBkTKN
I10Cg9jl4epiF78q4EpxTYW2V1HWzzPpGJfFsZXWYk00Md0ECx0j9xqQlP2qIQL3pZMQVBV2Tgcn
5CVwJw7hNgegLSfHnXE4qdhoeTRQEcmXZHy3K4G8dh3kH/OmcX1lois0DJSaNK1wnC5b2Jq02wiN
4uwfsKaBWXwzx7ylOagRTOb8zJJAXBNx3TYmml4vBuM3Y1txSpszp8coC445GBITW9qQcFwl4/qB
dLlNr9eNlVfYTifydC7bVK0oMouVgRM6kwcksfdXu/+Uo4klLlOeC2OCCipVq6Askjjl1Mxjc8WJ
i+KSQ8EHIN5KQjPA1xq1ccUL8a+b03feXGEkXN/ULCXQc6JZqoTnPkYqYJZIJn+tVYZHJJshOd1f
3Da0Uo/bakjjCctfElXYF15IXUuqd0kGL8Y6o5iPL1xLIT/A43vGVkhAlt9mb+hX+FzkpFGJfEYe
7kwzu+OpfYRvoZ3dWxpsfFXZt7lASRe0dpT72sYSvPsKBbBRI9VN9LnForifD9wlbz6UwEs6li8p
UzC0rD4RTYfLXSPh7GPOiGJiJlKbbIBALpQ26zRuVK9xAQM9NfMPkLx55KgylHFb3X/WZI/YBeOt
vtFvPsQlcdUlJxNPP2Z5BZV3qJS2GoKLs+c2SkVG7EMjTl+tJtl61WM4mick8o9NnGHMrRL7iNYQ
vnlQHeJ+GuM36eHi0CBzcU0vYVOYTN6F45JZIn99dYqxiZDu5GyG3Ykdp5MDS4G72biDg1c1Y4WH
52ULpx98TsuQYUs3kFSnNqjpePjN9WqF3JJQ4T7R9qdMNk1zeMnQyyC/cgxIUJzxpW9Kq7AREDLn
uGr53p8O/TBHnFgJAa5052fDKkN7X1QcdtuC11Cs3O2dxRfZAevfpXHEO8JTFrXr1vWCVSDWl2lL
ObZ1mW4sjyjFeFYrcf2YSUMfL7G6T11yqpKwxAYPwmlD2iuUxT+wTWjRmFL82Hyi39ojl6on/N2y
0F3HBwiDheaeuIiJnm8Quka76D+gON9HqRdZ7EAx7ggIlNRHD/EX34xjFbDzxE+f6yu48V/lpGH0
bwg8FULoGvF5ooH8ZcQPM5tKFcYvFWOs36KlMu/1XhqDmQy8XD5e7+J5KTHo0ZIf/IZl+xdJc19P
A+/lnLyZ9DCbCQokvqpLZF/CMjWFnqFR+vyiWUTXiHEmsdk4LzikweONrnoL7wly+TCtuDYc3bfq
1mnk+TaWpo5HGYunVK5tAlxWpfms+koqoiJ+VLWpf3C/ao3mjLMa9Obbyu5vwX+ge595Fy8HzNCc
RyGh1HSBPyEtytCvL3bMtFUhkb3YCq5fleJVliknyKQUS9l/5kq1MNYzRNlbQPAzSxHKcuOhYSz5
SNcUSmx6t+co8t2Y+VLhFfhxSRHqJCpqIoBASUzS3ohcf04FTFgyhWGM+6cuumz6tQ/6O51DRjDc
dZfoz2Lw+h9pJRkMbmsCZgHlSyxR6TNkjYJsR3XFClZXvhN5E2Crybqn8ij4aOtXE+R8C/OdYV2B
NeJU2bjr/f0vozMPVDIlN6yLK0F10TszFOY/wuc3L+PBJWA9HlOL6OLXeUbkZPMD7eAoX+EftwOp
VXHFLw3VuyjCqOZkicmLVH2yf1WO7cjr5WSJnebKIQgST3b2/16o433/GhZyibiU7eWbbYMj7TSk
ura+ErcOVicW2xJQZ7/9A60NIiTi4xrvL+9G+B3X9gZnCI85i2/wHV5VrxmfqbdXQjOuP7PfJ1U/
//UX7cTX8iIhe8m0dI/wyUbHutWd/EZvR+4mYkLU3XIzu7V3DxPpGrsVYFG1UoTeNw+ITsq0iDF7
VAVp1XgiRt7Cv/kAb+g4QiTG452EYvRXsqOwAr609po8vpuvk4nqmTEfmtD9Q977m0m8Cxm/9R7C
7KvqeHAFlc1LTn2NLuyJq+Dzb7PUa6QeZxwk9kss4+kT7AIYNa/yVnSpCtrSeayfdAUFBc0eoknh
k4RCOdN0wTURscUug0Q/GmjOeZn7efLBHLK6AhGkN6IXldZ+Krgl225xRO7U7QrIWJvCJh69zskF
fxaoVj//bD6WynVmGA1xnXvJlJiLZUBejqIFNAP/SwE3u94WilfFX56kZNHmcjrC8run544rHZFA
+rOtJtt8cjW822fDsxBU51z3yqOM0/DXRTTflpc3vweEOt/6lcdje82yOfKk7GCW7x2IqqqPPD45
QYSy9Q6M3SvcpxHDh33DnQc+BBcdBWTlEaaJUBG+DDKrAFMKqLkmyjmThHTkRiaOSN3XltddmNTU
kvNiFg5KcmFvSW0iZd1OESbUpK2jIvZ0tka0Y8AN7n1ME5PRISgErK7Au21/WPCZyaGDbjORN6s4
B2ilVSKivDzJTyiivD0O9mhhHTmN6lmK2mizbtPBTklWuZQKEtBfkBWe6BVnO4vhqXjC/Zb1lCzq
6nLFb9khWuO2ArDzOpVDiZTHScPgjYJ8tOHIUOS4Tt/+h/764GgkPqqU0IHtF0VGxbM7jrhMmSsQ
fzoP//mkXNdUviSI1F9wpZXIqL/0leuSjEJEnIqXipb/Mld5eUW8QbYDiC45xERIBgxBk0Ii2hW4
JwLVKXQvu9F/afP+fwnDDQCXKQ+eGlPzJIaYCfAcX2VhY3fACOSW40eGB1TZLwF7Y7zi9s5rTqxo
Xn7S06kWiiXecH3Q7A/vwd+58FU/EpRkKy8EwG621WyrYrjVeaq4FkxeS2bE/V2AGnvMWJiDRmJR
THTEVdRblago0AhPZAe5h/Fv3FcK9R8b/RW4j8xS7QXAOjnV3o9wM/CErEvxhFVZqzItdm+oHjYi
LzLjBSVQEflsavciv5rpYpz9MmW5QeLhE356ei33zKHIW7gvmTwEjVGenWk4SCH5a5noWQLvwQRW
LDR1EsApTcUB1yJJ7gW9ej32MlCwb2E7laNYe5oFX3tIDkh4KeXdqRWleq+aoX5Od3yWtnvQgsaE
0qktsPuv1P3NWsIY71lw4h4H62xGRiBkWbhym5SQ7b1fb/Uob/OevDB3EGnLDyojm9aKWgTwV1y9
J+xvhC5j/eOOIknDVB5kEYZDMAgVnZRAxnIUeI8j/sgyTL+P8rVoJ0K5Lz9Pz/5MyIvdjnh7FPOD
D7N5X4TjY//U0elvvV9OQ5/a/IJ0FtDO9XSHKgUxYmGgg1b4MwKrEACP5QfNbA3PkFGZzKqCUWI6
i0pVpsmicH2l4oSTM4BSlIUu3Zpw0TAVGN0XfkbT5GAtheUgPLCuvkgLL51KJcTg5wGOol6ndymE
fvR9siUtYgG/wivFTJwFbNMMSfGWhwxg21Nd5cNUtAGjZr0u+ebKmby+WGf0oXcxPm+kNFLAzZsq
vMMLm9Q3+sBh8vhu4s1CTa1XPn2X6QmEqPxeKc1mkyqgFRnQCZLsVsVSic1roY+kXUluNBVgDAWa
ow4KsVve6lw53no8+KZsKshhZIouwFPaW+lvJS9k9zFdQGo49RVOtHLcIkMNxM+KvM8Qgl4dSvu6
HUw+LxDhea7V6wWFOpgX/ryQuDyGBdz4eE/YiUNKGhgaCejAt027dKKr+kRalfRtC3oeJvqIsumn
tI9oK52dVaUmyPf/GbaiMhGJeKdt6gr0vvLUd+VFmrYk0+6ouKIQ4hDc90hnFQ78MbntkmFpavk9
OdxvBeSyWmGJHBRINVifIn92bHa6hE8R2dNuo/05lnKjyiD7hlvcxkmxTlgJeMvUbhIzb4ZjlqVF
/gPTcCkQzC/xeDC5pABsvPJheyxC5CqRk9AabOp6WecULxjI8/o6Vu4rOtr2xylQcoTc9MeRz6Q6
ntrQhINdPqsgLFwHzeDxwmJPOf9xF91CvsabG0+2nR/71lQV0/nJ/E79VrkI3FTb6g9AbXIVZLr9
EeEDIo1SO86cBKWmuNrIkvNnrDxfcxl4oK/5ummEYTjM+/29DCzMo5E9Od+OfX8EIVo+KvniLA1O
quk8fdbmWZjEWY8lrewggR4HnrLoaJ/EcGpKkmm/QhvAMTzx86tgnUBavqsO8RkxYUHP/QPbGCxE
1RUs96X1PUAw5I0caCfEHm9G+6VANtJBOj+IV1Vz8ThH4H5Tm6xAwF4Ud327a+3Vz4QTvP7mOe0o
0KLnmdLw9b9AeDtn29MnJluE94IrGJr6Y74lkj8ls2/gWwb94IOso6vBzG2rbGXxcZ5KDyxrM+hn
k9nAz3PjFX1t340kdTTQ9PzS9EHz+UXMY2yMgd3FsUnk15FYjQY/V1sfTHhXXe6M/q6/psdDe0NW
MZrBkLHndANqLGmld1Su7oqEstoNCd3eoYp3pbqxo12X/Yf237LdNUanfioPZHKuVQ5V0s1f40wr
hxuX5ic/LbSbCd1gNkWSdnBkKEuxEuRDCyHFDuruEL7Rp/a3yV115ezmihjdrxEsppNxQK2Blblk
tUl/GOxRqLB6REyHiDp14BcuPrVuNylA20FS/yqn/0UotC7kSE2Ob9wwuD3R6jsfzRoJh1JEa3C9
gFbLvlTZjhwq+ISBHRDZJjBT6uTgdaIA0FXxGcmascmmKau/vbOpK70BU9qXnpJTAy074X4tCeJN
3OwnoBPdUDUKzuvnJmjN53hsU7u4eeSxPprkHDcLODkotWE2tRflNnm6D+PoHcqf/Omnr9B+B2xI
1zmVBlg1QzQyjGLU5VUBF+wJ4gNPAcJ2CMTSte7uqfjrdpeppzH3tmgDAusPJs7rjR157HJ2sAvK
xGXiwvYS8kBmKYCZSuQ/RS/J77sYlKidWLf969TjiYrI0H2L+gDkf/fHQ4XFvib85SyRaCAzWwXJ
eP+80lBsxhoPjSoEQFJsLHL0Nf8mJIup37zKaVeweWIosB9z7Bepg1SG+CeQrPh8/qg0SRsNVSwe
CKSD0Z3Tzs+9gj95po5JJwRtdxDgu4rdbIxX9Liu9aG8SyCde5FdHELMJdC18p3k43xaviGH4neX
9t8I2AvRUEJ2OZ6RRJpVJ+OJM2YcgLHgEjZjM3iHrtLwhBQ70ZyDDs6/wjzkIcPqI8FFQOW5lo0O
lbQrgbaR5UQ7Twa3lhKvIC5X6H67vfEOrYpt9OY85QjCDo8ajSm9R8KyLb1r1cHpvn/n/cqXWumg
mUVBrD99acMdcMcMJtmExiB6z/Uki/lMb7k2F0BdjPoq5X633J0Tk+8QQWVl6ckDtwOGETPJdjmu
Y9EdP2+1VlxTf7Cmlka6zEopkTh4XsLzDL9QVxvW/4si4pCtPgKlEMQxoFPlj3EKWc4Yf0T1R/w4
mFYDqCzgiiug0PaetQkxnT+j+LjpFXDW/qn9WGlznf9gY8xSFpaJdK0pA0QjTh/wMNGQ8BQPYAoB
BKcajHIS94W08FRNPigY/xJ+OOBHjpveZ1gNO5i3biCky3ukENbE8lL2jG50rmujyf1aGw73s/yz
N5RpekPBnfeyGGSAtyVn7c9xr2FcJ0ur2GM642Mf5ilttlKsGVyt/Qack4hCECQHz2tz0rNiaqyi
dS27pzb4eYymDq1QPGLKTAvKnh3IN0rUURhPGKw1yzUYsK+A+OzU2M3bXgXM8esSu8soWxK+neXs
x833sGJnrwtcPE/H26XyVW98ftb0+g62jvil+sb1twL7sMBEhsObPm9c1iMQGQl8wQXdvWe4e/8j
vSaWToJUo7uU7eeIsoLqgPhPHba5WPh4yW5Wq4HFRTxh5yMvT0VQZse4qQdrRfzm7reD6xUqHddD
2dd8zRWVkj9VS7G0tYp4yj0NjZzLnKGAZBXL1bNhU2S2N3IKBAB0vy8RyvGBpqojKoWVe6BPHTbF
Kn5dr6+wf+xbS+BRGGC1GW9z4UTrCiANY4k+9U6ziPTLq9JYzTw+1ulTMp5mbsiFDd9xieqoqxPG
5D/q4pgrHcc69akSt+HmE5z5FHdoB28C+TVQm2vusObI46WzTf6zIxoIMXL1GkmJB4fAdL66SsoD
2ZpuaY7WGlnB9cOH1HuMIGq70OnEA+PDfL0l3Y0MNCP0dDej/nXBLVHz6bftd3EAAc3cqB/hFGTV
d6fndBjaRRAt6kNmKBKFtD+aJxWSWKZ+KuY16X9iC/4uEx/APCjK5/HO3QowQLZ+qcW9fZoBI9yk
ZlNNLpNUuLVcVibwszUtkT7gYbC5LQ+dfoXZ74KKFscht3mEZpl0XoFHPPn61bkpsW51EqccItc+
Fz4R+KtUD8YHUcMcd/nTT6BL1H4WUL0DjhRlA3AXW+1PkUcWA8Ti1N6vGA1pSMJGfn6wPWrLBL8f
BlO3/b+DSF55I+ZEs6Q43vVKphbKr0uHBoa3P2Lp2AR8oDpBZyJUBtaZxqTOxz8izTpaSAmASWqI
nN0MD6m1ag5/nWgOSrwDdBRxm0dUyGoEUl6RhMDxLF7BpDYGJqpcDHn7DGOIg+wvnbt4gMmy2Exn
nBMbl8RySVHN8R6paKY8lhJ01kaerwyx/okjsMdyxEe2mn4jOjyolJ3fHkW8OikYN/WuGD6vGNno
wERn+c8dCkQ6g6uIvSXK4rrPQvXRKnZHpdctoHjgePkK7Bw8q3yHqGG3KLILGYTx8FWjQZH59Qm2
SNPTTc3zBpugr/wjFXnf3nmJ1M8msaRFK+s6bBet6N/XXxlFAwwVjmGELs49zVg6/VpiaYs6pdFx
5mVb/pVNQnl9v/9RIw0zpSI9xEhpngHZFhfAUe34jTeXMz04dZ8WPWq0hUSv3xWARAHM9sz9xYsQ
oFxF1TRzQckx8X9udEDR+j1qFHJKuUXu1ikAywyZ05eWHKRxRhXHXfabWg/SA3I1KudAE86FteQR
C3fzhUdgqHGfIMeWtTx05eLrbKs7bGECcHW5C/y5vDqD8PP5ov9NNOOTUyhk3/krXtiDYHmqzgZJ
H2fQ83Mm/FNwyKSy17SKZ4SQUQQgtvAzl5z0EYrc1PfGCiFmO92KXpIMs6r+Fh/8sYA6CMdrFXlQ
qKwiuw+Lvx4ACaYWRSdSRsgQ78i0wdeeDeeqlag8x0e5UNfhioIq7Vt0aNm+3AP8KoW38IkCz/wx
bjP4EVIejVB+XbP4eXXTZxidJT3oVIQ0DwxpIaEmHIRsxZF6j/QmXc6MOYCqDewdB4TGJJXDK3+F
5+YOLsvjRVWR5u6tmK5nQ3gTElUnDVkvgkx7qlPki7jJ7nUVlZf9lhsrEk3NPimHNiu12LOW5Xy6
c2PoGAqT7Kic1ryR/Qyc6OA7qJcOzTSWqdgZi0Qjj5TZj++Szz8ajsqqVGLwnh0PMTGn+u3+019E
IMwwUPycIfMVfncd6/sCJD+wVe6zOhuT+vit+7ZktCEXjyULQ3LjCLrFG1zO8PCCfWSdx2Nu/pHX
c4Hqoh+3x81IUdpHfAeiRlRcl1H7fAcqeK7pVaPa48XlLH5J5agie0bEXCbZ11j3ks38U2/qjgFk
Id8zsNA14pYU1zfrnD1DCuzje+aEJ2ZUHpr0M9CZ1WEUz9wuAm2wfZuKrMyt1DTqgS/1G/0OREuX
g6jZq4ZRzaI5e0DTJelRtrARDSlA+LgycoVIO5PyojafWVaYyHK608gx1EXdLW+k9Dw1Wm7zD8Kx
OfgYFBLymYTvWYS6kawD9sjzFj9nXk/q7nwUrfREoJmH8d13wi9jTcjLXchdANjtBy5UeZ9R41Du
jEbyibGgqPEqbsH8lcU4CD4CMdR/zUqFnwv9b1A4W9mJHfk2+27EFSt9FM8pvR5OCwbrJ22/bgkB
AZ4hiljFFhfMUdHnaNRYACG7ZOZidp72omkPn0wDdRLq0p1+fKLxoVFIeeeiTOW3ySAzoforJ3ON
N2t5DDTp5aLPUkPEBaEJQKMzSHKUoP68xCdgvPjImuPEld9mw4DgwuKWOlhZKWfUpBIVkh/Xvjod
O2Eu9v1OuJo2cqZFNeAgZrPbHvsIg3uzvIF4eU2B6HY3e/Gn/KxICqHlLMFl4hsvMDuREearsigt
QC/8x/pQYKhHz/mg9FbTicDNYyLjBWCn2lZFMgzrXkjPdrKcPBoChjjiiDnbaoaJK8LoLRONDAXj
FZbL8LWh6D4aFryAMLjQ5TZP9cyIF5jBIgABDganMDV2JVVsYGDvwpE+dRh96n1po1Xd2bfdGhyg
V+rwTKZQu9OE6kHxUgVBINatv75Ffl9Ebdte/0Ed7BhAW6/GzHs3BMjWtHFm36HJ1qQ46LNxlaoG
AnAxt31NmN8JfFsy/QYfVCGqRnAdzRj+lD6YGnZKO/jACo62Sd2Mwj6aXZWt+DT6M4m0FHXaV/42
f+O+WzU9+CwoGu1PU+NG0iO9TfNuwr1aViGSkLm+kFG6i9PVgMz1+Sfg9hfIGbNuMGR9/Gh+5eVg
jH7wpRq2eHiuh3GBLw9e9bWFa1EpR/ocuzo8h5HJP8w24PT+wMq8F1Jz69CnWkGX1lxAeIvBhOPq
5XZ/h4zVTzar6bi6ckk9kh9SPmE4+w3lKHhhxP2mRrN4JiquQ9q3x6Y4YbjqeTrlssIA5jh0wSEx
UzM39ZTs0H+F0qDx0JYg14JgBLfr1PXolXcqvkEWj2PTHvQ9mLooibNVNJrLsYj+2Ty27JZYLTzg
TxC9Vfb1AB9ZotpVTEYNKYB9owiscw3drJeG9tJmX3XcL/xJOfcZJZd7Ghllr0inbyQZPd3PW/GT
04pb3v6B/HACbCYn599TLBBob4ZGmezhKndj8zPwEJuqF+dO0qHa9237wKx3P1vL32SJWSqp5bPm
64UaS5t8290UOBGt3Vw3jGZ9FLIFh3bbY2PZwhaxaFdeQ39NKu5mRcjjO+i4k1i0DNgxTJ6su2jo
AhEX9y38mqO+4Q/QhH4piTyx697BqJ3SPsTQW/bvcPcts0w0Hgv7l8tu9FaIfD331PFR551hX8iR
z3cIrNjJT1DuaomvLyVnw+YTGeeSlcDFUAqc3a6j0E8nsqn6jK4p2TpYVW/wFY2hrzm4c2AWNhuG
38XZ+MhESqWazDN1KhAhqZW51NmdxBH2Pa6ip/iUb/+ofoTLGw9U/Ph7nSiNil4rwfEKb9Yqbybk
ZG2Q0zq7iIdRMq9z9K/bKOF+5wcMWvu/Swb0uNReNRW2mRJgludlH41ycg92TLqVTLHqI3vXxALC
eu38As42u2HT6IscQUFxoECxj0D2+4GcQ8hvloMdrS8B/GnmieG2rAB1OMUgkzwELVYvMzcUeZFm
051LUEy4/p09GaCIluZNI2FfUqKDyTF8FrlQ0Bk1T0CKdKVQ/WPti/9FFSV60IlNGqfx9SrlVTO/
mf+qs4FlQaRD9pZaqWCtvfhDpqPi0bMfZ7qKE49Ksba6IxLjviCtJ7pUwc5slPbauiT7CjT7B1kQ
lbJtaPFDo88X+HuqpyfTJQZASgQlL3pdpsvFd54BWqYeSfPSYYQ2kUAd/8jWn1jv/57vROp9/n/n
9CZxMTxaVPSlO8TzTzQcR+E/HLK1y9K/OSdVqaEtTP2cOdGvbNSR0u4IDPwI6nUu1ho6g3Kuvwap
Fp3lYJ6gfabyoNtfks/mzM3wJ4Ot1JPA8MDE2K0s6Bf3yiucKOBEMbcdkW08QF4IIFxl8mkSCHeZ
ix9M+6K1Tee+6kfY4Qc4/ZKII++BFZMsisGDdtTqLKoQzTXvamnz83B+k+jZa3m5egzNNMlovIuG
EbfMjqg8sZtJlmN1kO2C4WdW8Xppvz7+c5ew0rEyliteoM2SXRp8b87xDd9d+1Giukj9NuSI0mRO
XZtA1kMKKXHlkQLg1W7NhNV7IIe5ZykNcSP1YItiq9hlK7VJwtza5QrhZ+Six7ggOjn0dbxDMxTe
1/70apX8IRIrfx88I3YWRqYBYpI1eAwaFrCIz9lrOm8+w56o2LyBSqQCzpzAZrP9246f72eHxdxc
DX1g4Wr+dZOY29bcR2ldwqZinAX5rsLGfnbDd6lGvCDfL9slbaBt48Gg6TC5cgIW9W9O8vEJljYU
ZgAF8WB7CQeoZ81bDsamplppJYZI8zWrI3pQYcwp3QwURNJE3YcKTlPEGWvBaPTbDvRM/b+osynp
H77GTBhFfsWQa3NT6Lsqv/6NySldzlH8rw/O6qvvpl7qwp+FzwreIy1PXFpWPfsJFQ5rd8J8bnzT
H0C0HX2ozFKBqQB+sxLgizyanYhvSK7E24FfaEvA7tpBcSclUyUzmR7GzdmCj3FdohrUm/XPGv4V
xSgihpKNk3PA27u6TKxPbVspu0AQhRgXYb33zONlAxlF8HDVPrc7EEZQ/bkHdTcmM4FM2gEUwx90
SAImsfzASF6VxTmc0zBzk9jQFnt5mURGQB7Y7MmbFtHVAx8hfHlrWgi7pqeEU0bPzo6fDsOWuV5F
6U/pZfwBOiLVFfOdwI8RgZNMKF+aQ71xTru5s+G5byJlG9WtKCRRq8jjsNXGmfJMuVYt8FPn/buT
95R9FsRW4RurCyFfAaLjbtIHJQ/OPZ8FoldeebEytOSXZnOm4T5PhAgfExUanGX6V9v1xRPNJdFy
I4bMC6CUbw7O/E+5y8VBvP7wvoY31OOxv3v69RPAjWQRqPNxOvsjF+MZuIwTfh3pedJP4teZSb1i
tMsbWmANQoHL0lVPl2RzMpb9+kYAhRZOdvaLQLeT0JhVcEpg9ajYeEQ45AL7QPoWvwHmh2QyCjST
BjXLIoJ3j5AIAo2JLzZduprrkgCpYhZzDE4i3eRcLfkmVYUlWZlItSRDLzVrIJwFXsX36VP9Wib/
EmN2mS4zSu/S2BaTEH1rCPVMdDKC8v+7+q9JhzLEiNNI3Beg3tX5GjKR9dQVJjrKh4bBLFyVIQWg
9udMM4v+oFDHABtPmBlQe9ai7UERoYzb97QRp3LoSXFfGGo7dnlxezi+TolxcTe55UL6kJ3jGUQQ
iwsmoVR5F2zqPTnLXGGkRzkld14hcHP1zZFIyIvzbMstYP2+m4JUqaoTD2WGTqTRsjH2M8N5YG9o
EfI8vmkQe+agodrInQQDxA8Z+qONjUsbpp68gHfnYeO4ZhgTzzcMtCUBnvcwU5vQnbUTufW+TZVo
Q/W/LFEKWSWNlv4mbap0SMkSYyVmH6VWF9gE3rQZ1U6vkyI6OxDO7COBhqAGY2efgX30eFlI7fbW
aAnHIR/eaoVXooBkdvZ0TFpcnrqk1IPmtBC7Nrc6Xo/NHml+vX/xO9DVFWlNTJ1nbWWIGKBmNZkg
jB5jlZKaqT80aAlk9ajsU6AHAFO8lIaOQPBWZYqJvZAc3FmzO/cuPVi7M95aGF8wDdTSVryAsJlH
2mJ8JzGjuHYXECo+A0IIQx92OjP/3EF93Q3ElcoT5ER958/yKxX+9jfnCX8JhFsWQEvE5rHTgZDO
vQowO37cNEsB2Q3ZU0dMr/dPwMG5cOwJ7VjDfZeEMAAol59EgwaigQ8/Wwe8Rh3eLecALZf3wRoU
BmVwfkxXsSI7gbvgEkWWfOmq+/qfjw5rlBlbruMfgiAWC83JBDxclKBLToGkdsx07BGOI1PNqNnJ
HjuT9LTYwlH7Mp/9e7nXBgpEjfpAkY0vs5zx9rylaCDPsW2P+qItkvHQh8u5pNfAfV3mi0rzRjjp
qoTqeGaV4in9R232bn5pfn5H9UDBIcwtLFjhYLdp2j/DBeVb00kLOLx8OeSwVxOTMwW2dSziycrZ
+jDR7bdRaYA09vlPQra2O3hczWia+wuKVKTTu7jtVpotSeaapmrt0TXSXKQptzipwMHn2pe6GgWF
Ofp5V9isBOc9VZ6bvUxGkJV2jHIXCShv8RGfh6GV86jElQPPT9qAnFCdT+S1i1tbSuMu7U7LYpjt
fq7KmQOjd9aQvPdFMdw5ibkvo5FR7biaQIKLSpwyDmXp0JyPRdOpecrdMiL0fDhl4hiEUaANWORJ
dG5uyIdHSpRO1qpS/czeWxbvP1AtCRCIuv+fYY4imcse0riPWXY7fbd3YejzktZnCZv2geo3CtkI
ecYdI1EEoWIDVhHbP8ocp21I+t9Dvpf3F4NZXmIf0wxjDbu26JKVx2z+zHa5fKgN0qBnbHk3DcBi
dWixQ+rfBYieY5myT7E3MfuFAquYU8JjzfPXKtopavicvzuJupqKwZqdVCeISTeRGus6bT7gMTJs
6wsxmeqEIgTZTiGZslHm8Zbb9V+mykx1/zRNK+T4X9/7B/HIZY0vhTUzVq1LoMVPXalalI1LDCJ2
wRFL+2tX7DkEypjPLFbW9rDrM6HhgcWPy+KHxhI6Fmdn1qGsTz+KLtC3dPEDzAbppVHqbYZ53zRt
98CAJ6lpoxGVvFWUJltchJ/PI+fWcjWuMonWboXNLEj7lCRltzAJLHVsbVrTH1QV/BbMMH29QR6v
WlBylgf+aLSji+zNXyoi3BZoPvVEar1oVN1mn9jt6ImgFi7UkuRLPtWWnwXvm6+oNEmWj5NgOrmF
uD2U9yxGoCSfWmq0vZraSGoQp3HPWckZB7gIWCTmyMCxh2ggRepQmvd0eTQVDZjB83+/dGUDY7px
O0/zGpjWPGbAyCtmIO5EskU4ArA/w/pnVaFYonymrAsigWSTcFMUkYQ8TzFXdnMdi+AXhTa7hui7
na6U4Rx+X0iGQ4dYTVENbBU0WPuIQ4ZUzG6psV16vp44h5H8NjfYntF5LYJN3jX3+CZVr1yL8cKl
UicPHGBKbgPTmLjIpy2Ue7DqCdTnVuEBl7gfcwV6ZcW8HYJq4aAT4OBxQY1f7UkFzQTnVTTo5Y2a
jN0V/+f34/fW2pEghUPPzMa8pMKQ0RdxOpla9uZK+9/wvvvKBYpIOVJP1nFKhBbPoWiyBRWW0ve/
g9XEMOxRUHDsnWVuq5roCwhATErNgIIDaD0R528QVsooEJAlyU3x1mZ7/hvnDsUv+0tMI3aZEhOD
7648Xu/0jfrNR1Y1vPlgaPDcrjTVXAHw2OGuLBDcBKDe/PJHv71/zl8clbS5zbnSqrnTSnhi4/ce
bxVD9h93i1LEnY+Iv6kI92ABu0qfg4pRTZEko0IBwwgJcgUQsy4zpzay9rg+kz+BSxdFiuMhDvbp
P7/TCJqu63MiG1IlRtIRfuygVSe804O4H/XrCAZ3x1YVwu+IRBunBJmM3cEm2xQ4thkQeM5w3jy/
gmmCHnfW+z1q6x+W1Ok6dOxDEzpVC6cGFrejvru1znsaGWQk1YiWdlTnlkOeUxsoc8YDdtNKlDJr
lwIPeA6n7+nypIavG7zNYyR2YAbAgOYyBahPaB+hN+3DpUrlXeTmLaLdRKIY/8Tb0bbPc43XLsht
rkPGb8ZWwAwRZQVdtdoAGovkYNyTuEXuTsffVmKAeKeqgJhO8fR9fPuU3TGZCvmV1nFU21QPNe/5
bWHhKgxoSp32vV07ayYFRS+A1IIiCEk5u4DAJgnhw3ZWomvDz5TGunlgHpjcCIHA3SytpZpbcX1n
BRYxRF38ts4EKsbiNs2tecE+xDQf2HX0nw6pNm+2ns0ACuNaVFsHaAtCXUJBNAEitI3BMUR+nwsU
Q2yxK6R5jJ6vEZ8aLyw9KLXgydfoL03UDT9HDTEfX/VtI4isziUuJrIViztxAqqjLuqxytVif2BJ
+2vphgAnPyAcrk94Pbb4iL3nzoVz5FfKKWvG6UfouAIwG/KRLsM9kGGbUJUNQBPotKb7q3WpEE8v
KjGvKVJqHoBJPwxCgNFAItg5w18zcMAuQ+JYmEx7179ByW+2Ylm7mkBmLhM3w0Ztmxm/kcGJLfZx
Ll4ICfSWCKiTZ8V9aeea3Pk1yDAezNV2rTsyiaHrMY6u1bYcx+68lnK4E6qif0g6/1elLMVUh0fR
6dShv7w7z9nHedzcU3So9FyNWc4vFOU1MNoqacWF+sY7Ex9OvBpnhhyQZgEL6XEEzjgX6pOtmbmW
aMi8gsYbd7vljT7E3Vp7t6WLnaVxrlNeffu6ILWFGy4LZ2+0ak32t2yAqQ8DMBbaKrkn9N0tMMwC
DbhtgoynSHkAJl5Bq0RQtqzRwhTMkFvUM/5qHshghByAsU57BswiWpX+jCe8jzXozsEiRuCX2wiB
3dT3Tb9Gb86U57QCGbjn/O9mM79V0KiBe8/B7PQhqTI7SvW80gCXYSlqhjG84HVg+fS7HzYz/mHm
tOGaLOBuGF+W9gpeTNUSAvA4M7WWz9AMS+GfjQdLR42R2QcGX9nITBXIIUl3s287qWjO/1tU2W4G
jQYOBWBZY4iAj/xusqJSSQ5MeVMS9EoZTZBbMlGbVgKcDQspJOoVwUJnYSAb5cgHwOj2PIM8iAMK
TCNy5C4jBvYA387vKGfAMheBbAxGLnG61piYo54C++7+rOxstpCmDQA5DqnnTLSeF3q0joylqugB
RwJOxsWurvIMHd9mK4jhyeDEpM0k0innRQmy+VY6KXa0r1QndRB1pMQY8z6RzmKzjjeyztkeY+Jx
yLSXSq04Abw6dxceQAYETTpDVT6VuCiGXRdlYNF1a9LJyuWVK8GuunM6YIusmiV+iI6OoW8eBs10
O1M0HrhD42gFWvB5VVZAx1YN+4WaK9w/HhJKiLpMdrJn9ugW8kt2RwKt/j/Mk5OZEQYXRVtztPwt
DBH/gIr/U1pbPEebbr4iNqpMoylghj02z5Hb87FagqTbJMeJGSx3cuT33RrwgieWFV4TmYcXDFNu
eeTTPNgLpy50Ea++rTQ8q/XXy4yhilEz1YabJD4qG04riSzqU3V4ViSztNV/gJTdfHUP1tB/hRT9
Lrn/+rdT7aO0dN59251rxpefHcg/mzKGD2j+W/ufUwzhaG7u5jwKdyc71sMX03rVejdvX9Zae96y
y1Cw2W/fVn3pf50+rUx0vWiFIp2vQcDINkSWDYvjWcP7o4CJ4VwnZPI70n2yJT6KkZnaeG4yImPC
6QNAE2R1ZiZLbXliARoI0FGwoAxoTLI+5GPvLFIUHlrLk+50TddF6X+Y2BHvaSKmfFCs49ufRxAc
iMx53QFDFFiRTfVzCO55ePMmXpSAIrKbuqYZZ1sDNL/P5cJWPkF3T5UQE8nV7Q+hvwp4TeQtIxn5
O0B5ylW2EDGzcdF0eJzdjp8HbsOjND6R9gAUJGPJUNQ0e8x6z8ENZvdHM/1hJMwWyobT2lAF4xzz
tezb7ZdiaGtf9PzkbsznZG5nQH8j3cM5P6BTh0I+VBVGbCFM+FP+tLlZ0bE9Xz5oF8WUMgbFl6zy
0T8QkolkfeTdzzYJgfsEnBVOi3OmggzhwLRhGvJpN6J8MsoYqPDJR7gDr7ZVxrMbR+jnmNZszTZN
7K550izKhBg5O8mUT0AQha0G1On3zVohEMt0pDw8wWcnWtAoh2Wuz2+F6hSMktSQUo0akg1N1MgV
/Ed+v66a6Giju+8FNEvWh1s90vLEFR28Mn5kS/MNgRXtmQeC+Yu0/Tsph1i5nAZfb6ZCS8QBqK0t
EQT2RVbJ1DkRFNNmZUhstktWyDjRewVxufUqu8QDNboqNSBCrDMlP1BNu5SDNxO05OjqmqpIdD5I
MJGoL1AJidxXKzoZStL21ejxVJJZJQZHPRW/faTb8gNRCzwI0R8jCvadNs9UtUQVGeE1etoVjTbT
JRiMcVZNXdi5VQ/elO+SVpwCdcj9GXhJ1dhxX4mgnYHGvfeoH0syLoe5+WXDkdXcRrrVW5OhMuZI
lyTk15AVA+rNYwTJXbCAYweSQI2/A8m9tIZKNnbbKC7IyCVDTSUNY4C41/yG4KXrb+0x6Mq8/Bld
4nwayTryiqB1XKc5n3dJr4TT43LkfGof0I+eOnGdT25tALIXsiIhTg75Xq1Th7M5rOO5KIGrAeUL
DezCbmRyHXaJum9vcKSdaVarTVF3Z00x/A9xGL5IvuldsFk0c8Bt4Kudb2edeoKlAghc0rau+Nmd
0LMTJk2WpTDNI5NB1Rqra+HYTH4tJmXScCaT9Mkx7bpUd51/FmN1vnvsnEy8MTeGk6w9FvAswx1D
s0521yGOZZh4iONZcEVtAm5Es4Y0aj4QF4/sKY2YQ4FpqnqIampPc2quBTXAxZrC46sN3anbHdch
ITrKhF76d6k5e01DOTsnBVlchyih+u23RFfyw/tRz9lRBO9hiZVwa/rSnKRhwlic/kGheCUxp6oD
cO85O22WSbqC1IpqKuxEdSdrxaIGiONDQms42yrr02CG5dRF6WOz7QlOEFh9JTAyEK7SW9Qzj5+0
Heuod81eT2r74mFNjxGtvFx6zdZw/PW/KRCwEapji6nEiJIlv8XMs+KXolHhnpCGYayGQhvdsuQa
WO/wjRcFcVOAZDqkOe95FuYlDJniLiv9L/RcLpmqq99h9hdUXLZOWf7Z2WogNGKUz5f7rP5Y2Ump
h8BGo9XYQb+KFTxeW9UOn+hO23RF1SFNSaEDHAfkaMWyQE4QND04rflDobGrE9oaw8InELA2eo7T
c76yqYhRHI+X4cwAuBEcHq+V0YkXEztAXBn2tVJs3jvt792tAo2jAFIRnTS5rZKCsIBEQFFtSUs6
ZvLYYpplDLvoaS8dw2laEELvo2HHtU7eLjaN0sxUYWzbD9QvLmCkaeGdVjQY3Roj8KvRg7TrOOrQ
I1ToClwvssJcnuBZfVT1K25081oEfiJUk/tBFm7BvBUs7fGPG0pbPBmribm0lPRfr1RCn0k4lLFi
bZLnVVzR0StOl8N6u9DP+rwDE3HqKAGxPjf892rPWZFLZ9uFdWW4ksv2bXnZruqfg7uKapuR+ofM
HU5Gr5DR25qtEchwlRa5G55dpn77kiUQCyAf/76aHvGKlmRCH5UiCg6jOmdgX8DU7zsxfYKdCpuY
NkXOnZq/AVXHGHp2fmclb3OO0inLBDSBQZ21xDI48DiydON6yAlWlqNszZZeDf8Bl9P7/2sAhqg5
GmyfOTytj6Q5NG382wXgK99tqJUV5eV/LS0IPrQmE1MT4AlnXuM7xRlexSVUO2dmNDIl+wMIaAPT
Hcpsu05knK5xV6Kh1KZA9a0EOXfMsLYHVAHmxAdeZguRG6CoKuqAoznogvJGJYXZhMdjbQ5M9BgZ
BDyxblDyCPUCN+CGu4RfjBYKHcvJaSg2mJhPe3QWqAI/vGVnatsTGtlJeWHXl2ZbjllBjJZMHX/a
VTXKUOuaAtP48WtOgriCH/fXQkM0fztYTB4uJdKXx2UjV3bvdoju5YgbaxC3DCnXrRkEp4yAzW2R
bjCyW+yNddXr9T/ol85+qYtpRHhkCtUgnw6MFTHgodpdOQHkjs9g+eNZHvWeYy/FgOu/ECvBeD+c
k8ys7fUKpO9ab6K34H6ccKur4bLiC/olcTmL/ozIaDr8x0Mj2iMd9fVve1q+c2ivFGfY+yoaun5Y
IIyZWYo4zdpyBH32C8kZfZHPyYCcdAbD2AJwRxcGyhlgUD5B6PRlCS5FT/j+9ZYREx+LEMHYPfU9
FoD4VZi0WNH5PibulxACYlPiuTQfiRJeqjoGgw6t/v/ZKd92yKbIhatRvHgTc9R29vUx62ZNlAQs
bdwAmezTdEev541L4oMcr9RLJGzG8xceu82WFSWaN5uWhdvAhztZEHQOpFiO6w21hCwKHiyZUQDm
WvKpqeF/vzyYuh3Qc+t6K+Dc8SEJxhHd4JPQL/tXLYFEX/UTFiypxZU3sJE+jquAgLjNWaN1Gzll
mjYalwsMFEEXiHHCU8VMPIPJzzIhh4Sq6JtK46aqR8rEERSZpS+z/lckU6dhzR0Bd7UzTn9/WUJS
alhrdjiXq/U4qj3V8+XQ1gxHAMsXjKcMSbGml5/XiOBHOhmZpCl38z3I//ChiBfYai45E1sJm71t
YYaZfLY3/5XRBnG//vLtlRn0/44WdFCQuiVjvqhWH0rskFpkdzyX108+OKmDUU+81CCzhg1llxey
lZ11VCOMqrUAXF2JkmVvIxStooT4MPoAUSdsXfjPB4dKrRmgVm/lSn2U8ghvgVMCEFWEt1bl36gW
gDFMSc4hSAepFz7o4Bgjy8s+gCj7bAhkiWT16ZRk6ConqRo3EQliAjNqU/yt1St8IF0lmfwIC5hL
HOW0ZUHi/DBgF+vINKw/ZGMgiOSRjn6X5sWu9cua2OaRzH9kk8mMkAHT+d9fAuSOxCgACRs/8+it
5F3htrEsBCXxwCK+xg7j0P/VBT7bcXeMiIaD2GjqZU5lj/VOL1BCDJHcLM+yp6/75c+NFlSgB+yD
DZokpu4wg/nQQ45+tBzYo5qQjFR3pIrYDQrYviFxc+uNFl35txk57O2+H41DR7R/JAbjmwgw6emA
q0IdbBHQs6jS0GeNCEmVZbYprqEbEPMqVJJXX35coTMS8z/IPmBzet27iXJXlHNA/S8JxV3WbcSy
vyllZzUhX+U2zUHoqkf34vdU05tgXEsfuDjiOZwCb1ICym6RhNwyDQfnl+BTvivLcGVcMzsXFrJL
YvWciCoG+lYCbUMg5I84QMwssRZOpAWCBjk3C/2niDtOngv+52ZT4MdOhYDXtZMkdXwrFP4YF9Zv
Fjx06Z1t3rOoXzu3ULl6SETanZnA84Yo/nwZ50JJuytVgJwHvI+PKhp4WS8ftoaUoBOsSGMpAfqK
D3gIWZZuaUP9IJpTxkJRN7WkDYqiFhmsykXE/RtH6h4f0Fr2hFyIscyIXbhMD1+9c1KA4cT8aLyb
FM0kEKjgPAf7UFmuUwl9zFtK6pGenDarlBMnR5KHNHKfNySoinkVzu7oX3itQ64P8X8IKFQsqwb3
1koG1AZbvFKhZJQA46crzz0sAod/bLy4lrSB0IxSqtsiH4150VUnuiBP+NTe9ON5+OqJJvO0x8ek
WwuZ9jW7trHhETPPabJ0kzJbfTsRLjaeuJpuVyEMKMiX0c5IIOxm3pWR39+yOhhjnaPTlgfr4oUM
yhIU5+KXuzFeFNFH0NmlKjubVmAxz51bUS6VYSUW/PPBwxz6qQ9cZqhyyIumbL01eUzTc0cUHUyY
dh5tdwAaW0KA63wRrjPu/JiIyxfIObBeYcY/8azIF9thTgxqOZcvhcblCxaSK9z9rlHn4hTHVvwI
cYD0Fcaa22T4cnv9HaDSRsiAZAmc9ZkEchq3ozHhn9WuEC80YyVH03X5cyDEGW57AJVG2Sl5MRwV
IoeFlBJ3qlYQqu4gj2MUYe8jh81mbRI7Ai8SKREpkBWq36yB5n/u/Zc8MrIkhPPNzoLuJAbT/NvS
AVXNHl1niGX1MZXDzd9g1ErcXHExbjc2z+R3KlgSae0X//2oCCl4uwK6GezA6Lmp3RO7jt9EPW4y
sPeS5KeuoYgNA3KElJ0JFATaWWDkP03vxBJmoN0mEXVdzaICVK/fNZj4yGOn9XrAEQ5tijwYCfmH
2ES2NZQ3KDbmO5kGXPqiQVmpHJpwDNo6TczKq5Kutzo361BoKix4rxA9kaJOqL9pcqqAjdjQCjNM
oA0T5/ntBoyIy1o0xHUK3JyzGVSvCYz4vtXVXodvvT+3Ktf+bk/7YAZMfJuYj1R3rHfkGIlMEAgL
RzXjNKOk64MtX6mQ8/cl/45CSOV154v6G1Dn9TJO2AUzCobU1z8V5tz372UajFj+BLvYx+Zd8RrO
5bWpJ/t7QXs65REGmgvxY1vlCZp9DIu7ABKJzo3DKSwCba0i3mUET0ClP4mLr/Ir6cJyMRvkLCbN
Z4HuY04EKtKaUyBScLPY6MKjiciTGk7c4Ky8sP9bUutHp8u3ukmUIxIam+CXSUPytvjAuaW1TQO7
rVn6NO06ROt4QT45bWK7JOb0CRDmbVSoGa2k98T16V/S4w0FymVE8NjWZZy6s9EczFSVU7uGZyRy
NZvwiiyiqDR+x/i0IgRCipgRV3OuCPhOoqmaFNsyZJPxnD+AX/M9l36MSR61PmnkwBc43eu9K5im
+zde78u653gB9c5AlIMvhIamoJLehPzZbuGIIPYkzEs9pFZfiq9v4I8uGjRYoxwvEujigmomgCxF
t/UPNPb+M91+6/gdQtfmccbvqyqukLSJfjQ8Ni4QGDlqiHqOplCCkSR6Oh/mAS+Vw5LPaYOAJB5r
PSCNKbEIu4r5LLMZNI8qNlYPpbrfdeKZAlpzUKKHoi469+8P0bBrJ1cEBUGsHQ033DMmOAvbyh6q
FKppeOS3DgukQ6t1IVFXyfp9SJaFHGM/Vq3qPp6ieKUOU7tz7A97zaonZz2KmQQz1fpe7Hx+b0oT
7NgURr4NN7hmqpe6hCgfO2LiFdfuIUU/XN97QaWB/bmKNXG4RpEryuS5Yb6BbDPttR2pZSMtlyFm
3BFGYlz2Tf30eDrftZbFTrMLKeLn8eWhlyujPnqzcJnqtG8KvhzXBRcLU1SY65jAr4gDi9k/Vnsf
lDnurSPt4aYXi5AXMg61d9+6JKm/ymYa117BFEGmGzAA0qyBeSIq/jRmlaBYOzlst3Pvg0Tl8Sl3
SkyfqZl9O2nL1W19KwHcvbjSAB2qVhw7a8Zl4TNolIncaq6cUX2yJdvvCHHErr/GqBEdYf9nufMX
cqf/Wa5rZkANMYnePuj04nTIafwRT1Fiq9jKUnTuXycP1DuKF6nATRjf9BSCrxZZc/24EAPyjOm2
BGA6d2tKDoBLux6eszotkuS6Ahs46vVuGnE7yUl7ASS7ZOWtZmiZMuB4zkXsXzVklcous/Tc9FGU
AFTIcPBVQROv7CAwqHEfntrwqn76uk8zqP/3NdqUR5LUTKh5gvwaScpalkFq9xvhwiNOpA3t7ot6
04ZMGHT22coImg3aaSiDOcaJksFM869CuTU6gEuNUosMZ9NH4U9iP+mUyELOT0FVQWeR2iHBgBuJ
tHA1rPfgoKohCYGCfQyfQMssgwSS/3KOlhPG+0UPsCiGVFgxaXB2cCcjqhpr39fGBVSoShcF3dN+
gwxybjYId6TmttkYB8SgwabYvS5Zhy8hBLy/VICTR/nGnSe6JLGJFnfwOyCwQGbY0EPrWxaFfooX
17vlJKzFfH6OIGcZUT0lyBlZl98x1U6GbEQfO//DWMBuOf+LfAhB2NVZMItmP9bWbGbOSLANzTqP
wBUGgxu6m/G5Fhcsh614q5HwX3OTVudwhUrdU3ua3a5N5nm4VPd57NE0FEMstwygQaBwJN1sYbNv
KIJ3p2ELG55d8eZlkd6bd7awANHJyxYXyE0VuPaSWsKJT6Qt/E793ZGrrIsHmaR64Lf1gqXW69KJ
x52ftDHiuyVIykLJ0hGPkuP2uN73wjF6NwvEX1c2lkQEo2liPqyUJV47R0RRy5N0l/+0BB7uZUEg
xBJX4XaM614aOkSy5Vy0RA2mbcDa+QzEaXBSils6KE7LnzbNssFvZeTpy1sBgVMTa4R8RGUNVl2Y
irXpseeHBbDvLh43TFi1qcqtG+8GcIu4X466S3a46eXneD2uvbogdxj1oAL+89kAUD9LTK1biysD
zd/Re8fg8fjIt7Z4VR2gRKhmAVCANvy9YbqihYhOMTSdUIU/ijawAg46Bk8y5OitUCrnZeuMN3FO
1JbPtO1G4Cl0M4eQFL6ZcM7QGelOyClq1T1e93iqIvR4/PpRHQHNOPmz+jxZ9AN9J5PAPlNy929Y
fa2wYpyP5jSbXln8WFuZY5qzAz5LdAs2RCD9vsL8nzCfY/P+psPu9Qs9XU9heUbs+zBQINuSefk3
A4XKPCDk9BUsrYf4378g4jSehcui8n9Hjliajc0jRKvGtIWqg6IgukipuIJuodVnDkdXkDyblOps
4IdnhoxbBum1xFUK0U+s0KiPEdkX1VlMCvz2+EIcGy8+f0b2fyFnkEO540Q+UWVz9avEPjchGNh0
pOeI5L+mD3O9muKsjrKrIH1EZ7aKvm/ZPeptxT1wHuuFv4ZAm/8yjQ+8gQ6koX18D/VyghCC7Dly
8qGY+vlfBjOrngkqzNjzJ5HIzsOZwq/ziYzMvem82xe2u1CpBHb7iXWtHZtqN6MozY4LrpMd/RUM
Dg9TVYmglMFML2PmMQue+6jJtwqQI0KKrZ7xE7OEW0Gsp6TfKuYk2Eq+odryWdt1uSsenJOTs5Kd
ktwwbZZNgnCHZ37EPPnPSVMJegh3Z+FrZDxMPWm3/x7oSgfhHIY9gwJ7/sz3rxPq93URJtrCIt9K
Et5JQWZ3rb6ihQQ2kabwerl5gC2ZwHb65k2hEsrPNfaDsPMBaFPgtYygX7W4yAp6kyvc/H7tT1mH
I1NGKvrcQylbCmVlbzXyxlb6ySLlU01kvuF++anzeIcN+f8/FQHMsTbInSCX4MVfNDgenJk8qi5Y
k3jtrGriiTxpFh4N/nRDvK2syqoWY++GnNjbgT2kfm0mFjcGianoAzSyanUCKdm+BST1+kwJmjTg
QEkn58vGkibf6+mftttLSSJmpqc/55za4QS7y2UENixq6fcYKHr+CNSQ7FXkm5ZmEImOe6DihVqv
9h9Aw/hwlafIj3Kt3NC3cuyCSzXnoxVmt65AumSM9Z91VEtvz3GjDAJ3NpI7HgLPqsYEQP5nZdXX
sRs5YoalziEvJ98AXCH+zmCMz5zUK2pokPQKgtY78QeRWS2Y5T1a8trVW4Vdn0ZvIYHbuEI72Nze
Kve8A8sjKbLKqc3EeqtsDrRI/D67pd89ZDYWriGCDW5wpX5txhni3woQLObY91WAQZ3MLVXMv90O
PPxRDOvSYpqQKpQB4rr/AnYVLqu600ZXzMOKe5rI6hU8FX1zNAxweNve/fKtf4aqwka8CZ9cqZAS
jWFZFEnkCHs+G8H8bwDD2MblVCWhJEnaYKGxZcAhhFCWnULcsoPugR5RdjNu4ymG1tF4NEF0pacQ
+kv9AyiaF2gCFIuQgWzWwPYmnAMxtU9XBfyqCTSRvvbR00YyAlgRdXSCM/LA8hKrVhHp7vd5c/1L
zGe0JBqY+Np8Q/lji1kQbRTDX29NdMiMgHnetoLfmYZXwfpR0MwIWi+EgKSqb4C52msDskhS4CKU
UasUuZkcEBj+BId5kSEUyaOzFZOos33NqcBaYHuA+Ll8msR3NBdb6IIlFzG0gKwZr5HvzsheZ6lW
6zyG+5ZyH9gg4Ca5Rw01uFSHBlE4ZdgDbkx4wW0mp+U7tWdi7oLhMRT8M+wIxZC2YJ9KVq2A/tnc
yo199K/oY9SqWtZpO/Hk6oA/5XBEM7jnKPt4WwDFyhjJU1Ps1H/wgxOAmsTrQksmK9hzSF0kGYFY
YqYzTXrTLh08Z0ZpTztD1d5EMhKsxq4kA7oXhdhrtI+dRyj3H0cH+v6N6bBXW04VR2hZTJ4MTp9/
aiW8/QHtyRo5VzwESrp9D6+vHCbZczB8/lh3ehRoi26sT7wshF62gyPSp+xAGa6pcg+PSZNFhJhf
+YHLk9oM/LojUj0PjgF9s54WsM9GHoCDHIr7d0BkODXTGrCijHlp/3/i7ijA6E8VRcPJi2aa1irb
gwsrP/R4NCdcbVn5VbIy/Vr5rkqbPGdXLPoPbIBRF95pLPo74onmxv7hC8PgFakSPM1/jEIT7fRI
RVXcyk6gUPGkSzodceUPNc0HislEOMOKV56csb8XRFch38oo4V0euKH7gFeEtDXwYhO/+cw+ngrj
rj7gKgj7WhqGTEtBukg5GEVI0ZPWghaQtBdfRrZg5358WXxGhOA71CJXbqdHhkQ/jYYAU0DrybUp
PPPfd1c+kCL5NnZZ6UGQcUWfuAzeAt0htoyBngnNgx6bL4fJCQOMjbEJgOmSNQ8TqrBAwvxlrQ5g
k+MrR5zXrEEjhK/Jpuy0iXneoC7meSD313FuPKYRCIBJn1OQcuSz75UUb8rs3a6Se1OYm+pNDi1+
NqfhbT6GN3FUjmoo5XVvMEe7Qj9tENsBZoe6AX3/CyBqfMB9qLl5DT+ZmrCfYDoFMwcQE8ixxWrQ
RENH+sSG7EeeoHlf6PY5r4qqY4vfvTc966mi8DtmgJyflprEfG29lQUYDANGybH5zfr0ycD9CI+u
o3TooO4Y6GJuZXKvizr9RS9mWhk0qCYNAbFdYXyExQym/T6vhpTFBl/c3//N/NXLgcOduE3tYMA5
aE9mzwXyR461VYgHIdDG32VCg15u1SRuX/U2171SSSZPhU0jJx4yn0mKJybYmJ1/wdwgoBVQF8RH
UgaTqH1sl8g+UlA825Nj506+xNAN3tbLIy1uoCNQ4tlZFLWR/Qfx2TCAbJ53U8eWNZtYi5Sx9vem
ST1sXJilSk29tDXzaIk3LRE0VXizQ4OX9z5wciK6uAJ/GZwRmZtyEzYRpgoDuppIC59CqkuUmgh/
JjWUNtYDixpygAV8cKpHsMMoFmiWG7a/ZXLOWFk9QQnKF1k3lvI9pxA3AgnKnfIYmeGMsBklQ1Sb
SOCVwY/tiSm8cXYpX/pNPEXYTejS+BJ4yYgZyfeEDeBMWFeuG77fgSExwQwsidvYTN+vWHA8dC45
DS6Lzg9sIPXdTSBlITqPFb7lyEsfrUCszamEeO3QNcfeUTkeGQ5Rlt2CVodVBoYMRKgKSauO+Erb
f9l5OIP+qg/PLycmdecBHIpjEdNizVEepFWgTiDELrDsBBPYFwFcX1/4r+k1tzOqG0kvXH496Kyy
HoVw7fFG7g1m7wsPvqBYRGhUiKcQo3RMqoqSGwdW/kM/lnzdF/TMrRTCyycAOoV8+VBJoikovv4E
ziLx69ePehS+CxHiwzoR6YWQp5bilqCtA1+X5zwTmFICKV9lgCQG/0n8eDucOZcCYAuTBgwZybZ3
CPuXRvUls1kOKpSVfoo3BIRPWyVuUbYCTVOrzxn/oe/pUkKepeE2foSrSmrheKqIesNIflM6xr+W
hMZ4N59q27qCwd0DopQ5iDg0mZnrjuJG0bHGLyMkYrJ9ko/gcSJp6zMgij4qTvr15sTqbYQ7cCkU
sMKoVEmTvJpPhlio0W0CX5QvasAo+YleX2kKZNql2Oueb5M8cQsJ7thHHXo3qQV83zOIk1A+ZIVk
b9d1kfoPSxYzHznkQJW3xhFV5sRPhYMCobC+n+ZOSTjxU3MWmKUXq0GK846fp6xgQmybBpsugoTZ
3N9AQk0t0TTnEUpr4bsBtwKFUHfuxh6LOLL6ik+NT1jw4HlWu/pGdr5/SEyM+Vmhvbs7NX6SsMgc
PUHHKUp1LXHgAC1wc+9JHGbhOJwwiGjOSrSo/TNEc/n06duLhz6Ms06R1Gy3DOxt4twGPbsp/3dD
48/RDjXkPlLJAQMx990C36o4lcotIaDWuu+DTppnJ7Opa8jNZAdFqbGMPVjSH2/mk483IMkCLpjH
I7MhU9NQlL3bsUXWBFt3x19A5oAbwoo0YagN9NWKhDuqx3BIRBFy51k/lJJanIouk4MK5ZTG6aWB
nxcQ+lWE3mjhcdGzcvVIuRgqAZjwDPLeRhmZkP568zVG1y/CuKYFZAdzmXwxlgUrpk8AjUle3ma4
dpbcz1UZF3VgDjQGTBvGzNPzqXjew1vGAhIb48b2t3qM625CJhdsQ0L/YxZ24c/1Yi1+nLD92YuC
sVo54pnloHshPGKOTlwYWsmwx+CoTE8n1HHqNTpZ9tx0lERqPSvSkdWOK6hMQ0zZ+k+UPCnt+vvl
zdfuHMHGld1qET/A9QuzB5ErSyHrwz0Mjthp4YQPvCNO47XP7FWhrZeiN0KxupzvUa6GQ8Iz7GwT
iHKkafOQUpGcPxTZ7DncU762vdgvDCYlEZrPXq2qb2uCe16DTaABmGTr0CtIWTJTHpGjCkp73OYs
kwQTTlNRnbDfebKnCt9np+KhhKYg8JgUQoKUzvLaxkr4ebBz4t75o08OEuLqbosErvOttA0lCoPR
e5iBJmdKHvcwHd/jKkLw4bT0KrIG+EgsqcmM5J/d+uZrSwowdv6LzvrGFz824/t7PTwOf4aHYNiO
YW3qdl9kDHMV1cYLUR2gh4BzSNr5ufJ00f+xqu63fBpewWPxz27KrmsP3XSSTslAhC0TtdNK16Ux
bZESFJTtmJG5xBlYMeRb12bnnyDp7I2m2fJCmo7t8/fBH6RfAcjS9AxR9ATtR6Sqk3NaPbK/gZA6
c6Tio8m4KVsKwc7O0kUHpPgJ7Bib3Q6a4dK7uMQrkeOMtaBls2fwgDfVfzyWDbPkty9HLm+RLK5T
7EZF5oRr5YfFV+9hgUPuqNyR5lzXm/J7/0qlSdn5w5AF1zj6tbFuhFihPxI1giMUvc15Mj4TFJq9
fiOVhwRLe1EqihTlCIk+PRh4yJtYBZy1DWJnLpNr19b1DzG3rcBDa+eFsuMN0Fm9qsPBOR66BiMC
xdGzrfXzQ10xivaJKnJTZetNQbZNDXMup6AOSHM9PSfY+YpH+AMUjB+BOMnQ4LdqK87e+APKaJv7
d4lka1vE99UcgPN/I2AQ7P6VSuvkk5afEV9WJHiH20Yq/Tg3FlMPXY8gTfjFgFHoiwxNY8OJNVTd
n8HCalRCOvYpXhD9KbWVuHcpyg3qxSShlMw0vw59uz9MiLA8pP3ZxMXgLhMB5gsS6TMwu8x9o15E
GpIKGdXz5dSnAjMMWytJ3AUKF43dU2iSU+6v31o27PgGoxHMTi8WJk4Y8aELa3Y8jRQCizucsXPv
RDJ44BrDsFZmKn3OPlAs+8eJUclrvgbJq4wPdDlPhwE8hcFj7ZlVxqaYwzlO6SFvX18vJQfjMsB6
xjvvtbWcj0IJxTmqUXCIkKzTM2GAs5Sfi3HTSeR5eSkSmWZSBMVI9gBqCG+sQJ198pSK3lHV6Vtc
aZpOHXhtjAJKN0ARpsHBRAWJ5snmme3hhs6quWBjcKBV1Rb2WAhla0Y2EJfPJZNPl/hax8aZ7zEV
15PasJWMujeMySXfpR27dqwm1Lt55zyF8eYjjA2bo6j41P16oD/AtvUVGEFnehbrEwEoGIwDvtxJ
dMTYivEyiNHPys+JZrYXtT1STcYGR1RLDrPsWIGmHLdaq15kr8mVcoVXcaeavNWwvb8MFXWfWvrR
Wn9TULouCp/jSiqBiWPumVacssytVFEih59OFdakTjgnnp1p3N/vX9/my4XWG3alCifbUmtsxg4M
Z14pBlcyJY5KljsB/40AlxVgGpP+swe+JO+ypNYbL/WQCHYTjDRX+wbcZC/azO7h0HMqzbp/n8nk
zTPysixUkul7Vp28E9ZDqswoQMRPbEmbo05TBOc8Ctnv3Yvvp7lC6DAr5DguxT4Yya2q1iM6cK8w
leGazzWp3KggpxERMZq6IPzJ93OayJBrOv6LFIvZpd23DN3VWtH2p8kWSKuvdAQqjiFhij92miQr
UoRFbvTmKsz0rSSLIIyO9kvO2OniXyWQLm1wOU5RiC8vdN5Goja94EuRTTfj0QGkuDq/LR97BNL4
X56Sm37OwsJ+IMnl5OiyZo/rDj1KIWGYwr7Y23DQIFnMjUtmsU6ou7YQ97IVFlsZzVVwaeUs+jyJ
jexD8M3yTgdsGKY36FUyTToe6VWGKtYPDOu6K7I3wFIRhzoK1I+8BCwl9cAOkPjlg8O5regWDCFR
HRB/51ac+JjFLrY4UnyyUl8QcwZcG5tBidbxiUAmlMJ8+tmRQrpLvlvKdJ8vBnH1bx7maRE//sxS
6qxiUfdkrbZGho19btTGScahqEA9QINlOQpyr9/4rLrwh5z31hG2f1GEX774ZyJ/JbbZdEte5Qfn
xdehgkaVj4NpEsSLY7FgC/SK7MWaWHFgV3IudF7VkYplJIKTNN4D21d3KICVp6z4dGYMr1HXKhM8
ovyh2/CjHpnEKlwYl58o278PaQUcvcnmhO43UIfFaZiG1Hrx6UTaeUep3fiFswKOSS9xyka1AdrY
sBSpct+BCUvVdB8qBcqh/MYCqmu7mzIF5rOaxc6zY03KQ8hdvMVOCwT7hDgmn0w+ZqNJ3u9HQaXW
YvL9izGUGZr7n7nNO+jGCf+xwRvIGrtBJbDM6iotRaFNW/dIPoKJZBYPSnfXrHBHbWLdZpgDAsJg
Owqe7MPGDEjZF4bmGKGTIz76vjBzo0POpwb4CJPtyQgsaEsD7OqMDMUNMqB8kaIZ9RNXdhqAAolP
ujNqjOwgB14EjFpzrGwubyOVaGb/AHZjAbcYTPSQvLByjNumTqlI1F+WjSFN7YWle++vo0aoxZv5
kX0s/hueORIWKJQVQue8+suMhNEzJr2YUy7To3JYYY9S/XwyFootHCxFwHoR8uK/Pwfa6h9h1Wia
sf398eAMJzeao5h4QS2IzrGy2bVVMVRqEDIqbzMmvpekTfsbhkFucaxKap5bVxAWw+ojPgSP++uY
pLwnSF8mg6MsJb8DC9Wi10OyqoO9fw0T1TjYo8Li8PHTGapSrdshirDfgHaECgvOm1uN5P/2TBAu
TT7c14UHohG0dUMXwcibe3OaRfPFxYSK8GRZ/B4nO0bu85d0lfYtRXpgqJ2eNBu2kpPR1nRt9Y/L
h9Ibtzq18cmBcfo7Lkr3JTd4LXnVKHWmd/fyxcnkEPYiiBUG86ONM14r56FfG/KCrlTyXEC2NTDA
vEuTNuxW4F4gXz9M72G6zlu/APKfcoRehcx7jZWafc4JdgayP8DOXNTTAkIaIy4G+qYW3XybjKv/
nixXYWmfoi/FGv3nsgwUrerb70parMWxtOolktWGCDBuuAn/vSFlynGRfivcqYyCX4f31pUJCiY+
CaC5h9nTFn1tDCLj/xqJexrCEC2lX/zMrLlzUaYy1kYKpgVqCSYDL2cG3VH2Qq3sFNj55P+v3zfS
E61I0m9bbRC1S5bxjxB9CSQowd0l9mI8KTgUEbbWzEeccbja4EY4+ahRAyz93d8gCC06RneJk9W3
WeKRzeX9jdSFr6r/g+rTlH3iikUpsNGtBj2Mnw38o11Q9Hwi0azbzj0kVivVftn9uJeZcVIzjJPt
Tt33wqjLKQLIFNKx4Z+nljpHjdpwga5EViEWXCe233pfx/+t85f1XMlJigqO7tSLiMqLZFnUVJlP
VBhwEDytobL2t/dnLaUhkwq+U4L55p07MiQPHlhGY2MFNpfsaQr6+lBaEvKyZ+OSrBLZno7mOswr
8XyqGHp6GZnR1u7bbSnRp3YNOLnjN1PH+aozDbxD1bOUbOJaa2KMpSjcCsUL/6q9V+maIz4/032v
mawk3i/Ky2Tdfwv5qZzNoZBBCkm6nNcBZ0EJWd9YAGw1kHhE6b4rpHE5X9H5CLwSgzyKbQfhmJQp
htIHviiaBRk18zdAwvNTkOyIMzxcYh+/XeI2Un20nTyKNE9c+2e866Ht86FIBoyJE5PPZxoF+vcK
qC7OQyTcyIxyKYUuNfI0ImqQl2Bpek4IfAAADN+7pMHGExyZnWlm/lLS4d3u+YBKD0Ir8e2TrPiZ
d/pWkmcqxm+8uzEqWSR4kFVRx5xAhrDSYURMjf/u3KcYWJdnzZFrITmZVc/xRO0VCNoMztrLYin1
1E00c4ZCdUVu7lNKGZnBrVbWEqoa8pkaAgh52sR9G47yugsr8TFSBYnNAIlBN/hvLrAhN3tWoxmb
F6dD6vjmi8X2R1Z+BhLaj/V4PZibTfMq0Rt/Od1J5+fUFDQrJ/3n4AOT+BN7PNYPBjJDEUF6PhFN
LsT0efd/tjZ/W/dOjACRgw4GJ+FQonxBOVyt7NfnAcIGCIakTEN/QJ02SaNQcsfl1YsqBUmncMiP
zAIHLD0Ap85jS4D7flXQwa3hhLkTQHN8uOeIiKB+4CJLJfunH8XfHQJLC1XSJ+wtUDn0U7bfw2zE
taBcoJZo6fW6ql/AHL8nVv/d5Qn/60I/+ArIUK0yk2bag6BRvF6456wJVHMQLOAutkNUT1CIjst3
m9+9TNz7wZ+gvlskb0a8BGO0PB4HUoaij6zKPF+PGi17kjWGpNtIyfhWzQ7jsgYxp9SP6QSGv+Q9
8dDYVZmYaOdXRkD78uwk80KZfnRv3JKRCmksXtoWrmT8QcdsnBqY1azAS0qk7ZlMeAUSh4J8WVQz
9ljsUhO3JYdfTSSXd2hvt/9E37OctsVmJmD3mDjRPQMbobNUJGsP8Hx64eRv4KRtVbbPsKcR4KmY
fzCY4eU6mWDIhfCBOQMb+iz7RFZPQDEe75h5/JkZm/T9DUL5I1hYnAWw/SaIhd0MoFXg5FTLOpSX
m7JeoJU2b+0HE2iMoMjcZPkWANn76r/6VCk7ZTAHMJt2SUJpfAzBeRShAlHM/rIUwrrVjqiBx6VX
cneullQVMRtsCOPfIGKcFq8D8NosOJpon2ebf3KvTq+dk+O9gm2Hllhsf5uCiFDX4MpjAiGgH0Yk
KtI/gEcOk1Ybf2gYMJTEZnCuKAj0nbt1G3JnR+svfz/4E0h/R0/6QiCv7So4R+JJCbotXaqUKFKY
kRy7DFVU1KCYXfwsc2TGEc/NSKuTIhBGeCNku5f3l7JdIFyyi3HkvQjHhrIcwRI1OiBXsbFVpQPL
Q2uN8QTd8FfPz5RXVGOfcpmQvucIu4bOKH+c4TenrR9uRU3crK/kxGKl2Hgqo4M6YtpCjrNBdt+i
Vos3Zu1PKqB74KkMcIOFrnnH3qdCauZS0Iy71erUKdkBjCQDlSCRQ+Vn8t1QX4pZwTWDAvDUQB+N
wxzlT96zRTLp/8ZM1xTRry5l/Njp7fUx8fw68yJljViywjc40Sxf1uiCSOUfmUb7ieRmnFPatJJ0
vk3VGZPPKZq6QLXV6c4WhV7KXmtR6EE1Yyybbg4UBLGa9jEzqAviufYsZSn6tBurKFKvohyGbFnU
z0xqpi9cHlPcnz6rtzA0R3xT2DGjKd2zwwjGlG1erOlM+N3/Zg1h6XPm4nVvEEsvkzO+XudhD+xh
OrdB+aN8nZKPbNtet2/RwNU22yFL4ndpU94bS7xOQ8NHoLznABtTioJnqX2KICk+tjdURfYjJHTo
5CTcNrSsFNHtdmeqCGqG4ZaKuL7X2ygWBgHcz40DhMWMiZap3ACQEDgppszDARzbLRVqB4qw+EDY
883ITEMts0DjYIasgrmL0pzRKA01jOUmpRcE8hMKP7h2bpCfVuocQ9APAODkEjNDEUOATWiawJdF
Ae9vUgFQAcEjg53Waiya9HIkFS73ikGwhCuHJpDD/9WxBFA4UYaeTeX1gVUNL9eTyrTFiBUV+8FK
aApn4pRr1cd4+0bUbMOIUuB/1xwTSN+0omUyz5WtrOV3u4S5wQWpVA6Mw/ROOwF8C0ZSEh4ucF8m
px6MK6X/qVsYgrZedRKvpqFer8bhaTkeNDV8G+0QwDVDpoRosr9+iQqsEXXoHf8ioZMYu2fcT4iW
QIpO3HHzVoDul+EXUgf0GZlMN4MVq9e1VMTtMGYuPMLSv960I/Rw2O+G/m0qqUUXS3jakD+Ctn5y
LdrPLidPirXjeoHtyHEh3ACBJBA91fWdAW11ch2CuKejrTdVDMZKYTeRZa6Ep1V3uFBmkfDUgVlc
u5NB4QMoFh1JkAHXEoMkEWk5pbBW6fprmTM6TawWQk/6UUXNSCAjk6VY9LtPhNSMJhX+flVDzg+B
IUzUAGrNgD38io8H/uvh2x1TJ3x3P9rlGlsW2yAMaae0gox16PJg3y9oROiSb9u5djygndAHPAhz
2xApO6iwucjpBLcySCqJ1bzjQLUrE8IB9HLz24U0dD6p0KJoYYdlpOIOyNZ8KNmTVb/Ez2sb9AL3
B1pVTyFL29RCB9wlP0eL3ktDf2/78LcZk2aZpWtmlZpBOCdS2LVyhV87/aZoEyXr7CxhcyrcDNBx
WR9mI0i7WW5pEshhfoq0jV6Ie3VaCenYpJ8g8sMEo3NWhYXQhWwOwbBLWj8liWWNGX05z2Cea7UK
7tDlvLnel/y0Y5i+kEtGqrO3y2mi7ltFqL2hG1VXOoNZHGpj52QkdPOyusmvJ0iqveOEx64360Q9
9uSpI0ChSI1NGNxMBB0UySqI3FlAk0D7FGVijqdhWBb2LZpd1z5WvxJgYHJkybIlnHTh0J0dPWH8
vVJvt1ZH6Q8OOXRcBhoPZkOcLxj/Y4yRY8jAdZTz15JuZ+CcM87iojQFmNS1UF+YcpAKsruA9Sd0
ks1z9aVRoeTE63yojINaLUiWyZ9hqUUrRbgdLcT6YOxfHm+WeLqbX2ssziuccRJqijCasQGbD5kA
u9gBw9nhYzECcmT/Y1RLvCajQvQbW18p+5NlMUT/RI9za0lkUMI2Epy8zGhzcnDldhxX4lnMgpIZ
MQIWaQCKT3L5dXvKEEJ8LUliIx83TYKeFGWSt90PxdsY3Bn3l0XOK2DT68UybIJv/FYGEzMzwhtp
aBJGkVwOod87sLPHorNr6zdIbLMN3ARMScoJFkkag/Id2jagQnpI8B/fI4J9lJ6dWQlKPZTrdilw
iBuMXk+hxSpXiu4ZcegIrlee9CzZfyAk8VxII7HrfJWIwpBDttKjdOuga8ngKwYKTeCRDKuG919X
JvpDCmxkqmQJZXFGFz8K3LteK8wpEEsnQGKNGpTWa1NcunZ3CmJkP5kBk+sGYzAaC6Me1gZgkIou
WaRjbEqyGpSHIkOL33bmSAONdbYKJhgg5c2flYi79KyuEy+8Xxw9EBl7BNWgUGjt/Li3c89qbgo4
NoqVj5mzKSngcXjgi2+Sqd9xtTnZ81/hNbuKAQJaAkKeh875Ps1aqm9QIiqB/J5mA67yry9XiawK
DjnwGRlM5PWbascc4ni14BP4DY8Rg2KNE+kvmkvobftdlvgLs+kv5y7kvJglRMve5fIrrYte8w2E
rBKc/CW1JI4swlY0cOmf6JfxAdQP6Kkc5anAQUzdjMtd9Om7aYBikGCamBDdvY7amT0l8IV3FQ9a
m9S4nOkt/l9diUn9LX6jUjdywIDX3fAMcYmSsbPoWRL6ZhEzNnx09xJp2CIDQ8JvsRgOKAc3CE/x
wkpgPK3ETZ4BAI+lXDelmjAf8ZoJr4JE/T/CSguiQ2BnwIJex+LnBDcnjx9MWIPvZirKfADnt1F2
VyV1D/+E7Bfg71Lpqy4N2bWbuynf+cu+HFf/E8xNd4Ci5tD2tJZ6Sr/xEvFEzHXvP8qeKe2ASYvS
swryk+GeD7o0zQFwDpb9BmuxG1xUPM89keO/XeLtzr+LCvh5+Mv4jr1/HfUXpJNXzjyx4v4TmLz0
wQbSP4iw49wB0NlmTLNMX1kmmYkc9FkvZgOnYYy2SOulisM4cKX+FwtGdwGUmBUNPQ2ePHtzgUW6
I4hGrKDqCaiRF5coSnvz9I1HAy0zm6MeOGedfBYDBoP9vagLQ3PGwVaaiFbDChl1rGXx0PCpuG1t
BRnLtHfoAVad1vVqrrnGOKdpHYaf/1b7GiHzKoq5oW5oyeiw9cEwDJoNVZirAaq8YzKp74fSvx7t
YJYcPGdkv+g3CVASErZruYPHr61QHDmY2JtY1kF7GycbjMfjw00m/OlWKh69GawdX6NgX1J9ggBU
L6MhV9mLclVtpuup3S0r85xdajUZiZhzD6YU4AGrU4YB8VMMpoCK6KYntvi5q+5sIFlbb6NpESoA
KCrTpknO9NHNKAhMbDj2JVE0Hry7gKf/wS0vpVGQiOSMMeRxFUmQ6fCcfCqymBD/2H1cM+KdgPJn
xBIQw40RO+rMGO1pZKbkItqmAKrdNQ90xvRDFL/RL8rTmmUVivWqYxWay6QeJ0sOw8xjkbIkInxl
oTTUGe66bQYaNPanP5MTbaxColesWptE2yjlqdECiHcyIjeDbrFeEkk2qUeyLAzU0pQQ5rPWO67I
EdAsbeAnFTwO0qXY5CQcWtRYlKoI5iAHuVqrOK0jSGi233WwZ5mG+FO0Qe4FeRYXzTdgmqkkFHDH
a8UsZN8VLDsMtWzQasVK5bvrOrxzgA3dKie05hpdn7H/W4xU8GkTe5z8od6npRPNisAi1zJPjNYq
cpm3AX2lhfy9gIBrcRUtpHHjkMMOxHlzNZge5+Qtfwesr6Dkqff9Koj/AIfg2MG7mbGavALF99E/
tYDpIeAhEm0U0LalBPYF00DREgYD7A8CtHwwyq2mUbiy4n20eLCoyP5gc927ZpvKY4hI5fVEcYNh
6o6V3N5K3zS0MRqUOXr80iDQMKX3NfGtViekz5oKqBR6ZVDTwCLEHu8DVsWOx/E67tyiTj0oFxvd
Oldt+BO/R4HyHdvJlnGZyNFy6cv3BGyZQ+rwleSzHEbPv8LkrrX8jmeWAIXsz0Q3vzBz8WwiTOdM
NcOtLhlBtyXT3dLdyn85UD/Df0UU6iOP6q6fplSNTzWCXivfLuhmMto9RwLYEHZG2Fu+Kw0KgnT6
ftmMkFbjmtsg9EtI+MTgZrQJXnBgDSl2ita5ctwrS7XrJdi/gAtZgNTz3j5xoxtRl98GhiU31igj
Wy+tU9ludo2P7Esy2sO98jYVOx6NlVVKo+TopkxgH2pbNLLJ78EvkWxEcN12v6wmDEOBxgeREWYk
yr71/qyEwBesEqWrwfipzQu5H8p65FKvhV3AhQ3JjqxpUHQgpMaHc0W5O3TvNRjKExAYyGwvuJyH
9PzSEIUDek0eAMBrf7A/5GTOPhsS60YNabnlHu0yuS/sNejQoOJYzoinmPa9l/CtaqevJa/7ch97
yUJd0/oo7zTO0LwTLdOLYgm6OGzrbx4jRMJhDqpBWeXemQi4NpqK0shd5m7SzOQH7jsgXVedBEYd
5ObxjziTqv8bbl2yxVoUivduE/VDufRFKCMyBm17az5Z524YaQkcg3emlbAKxi1DkAY4gmZqz3VF
gDg7JWKVrLddpNBy30Sp25tuwoY4JGSIHz84mHoOll4S15W2ReL7spB/Qf0tN9ZU4YuzFs2Cjs16
Rl9XVvjKt7mawHD9p7wNEUE5v/Z6YnOxnDRiWa4/2v0qGoKuwbJdT6AAvcXu2NeZbcs6xqU6eIhp
4GvHYRJVoflnS9KEJVkB9/pSpx3CqOdWjElbJZtbTWqUdtRq1CBm+VwqB6NducmRfvTfVtFS9/76
BEkUU5JKZD7tUvhaBZ/wy3j/wXvq055eoL45LqtHziZqd1aFeGmcpTTbzXzWRKytLJ3gMmq38v0o
6qjT0KZW1OmY1l6Kp4C3fsGN3Dz1XRspypxIIQturSk8B7GmMKpb9H5OAXj8Ae1bAD8fA5P5OIkl
ZUrT7uxq9jEGE0QTwPREmXvlfAzXHSZKvAvvwDNvLZIceFzFNU4UDqiIvhu4g2t17913yEuppJ00
rzriVZTxjmDK40H1ARBfZB3Z+BkdqrczY0UJjKRIG7h325qE4STwP6gKBRQZW7m/8Ulq1hDfkqtF
PoBVfdS6EdPIjOYTpTWAMYF1XJ+NqFPCtxJiAcOHN2mTb59uR9a4Sz6NGPR9/5C3DAsMcpIFiTH8
n77aFIIvmhOYfxTeayxKjefmgFhQHMiOPRp8pXAwJGdhsGBxXhjMK4K+OAghVLgcb0iNQD+TK4j8
VnA3lEfPm9+RSJycIj25um2IXIagujyBMT1e+pkGLTuMGuhpeXcJkSuwn6zVU0OMoUR3K0m2QjY4
GFf0szz7NxvJSmkskBZ18YB5z6SB/FDzhCyEhGhbw/2e33ijEOQ8tR/b0HCtbX1WQzPId1wDInXS
bfOb8TGYoCozbEE8GQIEfM3izKMb5ZzwN4prfSG3gItHfjL6EC0PUUOopVCCZVw7+yQS49gVXbcR
8WniJTtnMrezSfbrpgsKkxnArM7a5ND/xf2WUjBpTI52gOBF8ipSUuZnLlED/fwrbEAQXKsDH43V
Z15GeEKssbqo9bA1+Be4ULaEmuqAIyZFVo6g+vGpW74o/fLhQvHulwPyVioB73NBihN/yDvQVQ94
cf56YwpJh35O00BdlP8unYVHp2zA7NKWDxIpDOpn2emC6ZwBh92KtQhyV1GCWfcBJnkCi2bUpERd
RA2YLhI4fkr8LngjMhnOyeA1L2OIUuF0fvMoSFLbJEfthnMo7k+s83RobMRg7wW4Tse7vG4TdqjY
7NnnM46eCmkJYOxUIb8WOhrg3YpsjEEW2Buy6wclbZPKVmMZTd4ZesTPRmPS6M0ahIwaPz1H+utD
Qnn7lHI5+6YoFetnW4mC/2+7UQtqlMxc1+9qtjvzkVRd8q87J++bnoudx/FwoOWfhqpROc8cRDPl
FWUvOw8qHl4f0P9FgR603CpLQg3S+oEGZNHxTC7IVYgHWRKUPXzR8LsmuabXvLrTRtwCZ5jyzGsl
rcCvTKbcA3vcuXXGqcW6BcjXeMfczf7XPSXI3X2Jgqyt/Jp7UX+DxS2gBv9EAmE5FuRk7zXJCL/q
BGv6Blab/kckpVn4apANh1BdMNe5mEzwPPcjbDNm43EmO9deIOMYjHE9UDgnj8DiKvY7qcR2DuOo
dhpMJJurKtZm+cK80BykZlEQH9ymeIUOMgAqo9bkQSSZYnS7x49QLH8vuSJQKQN+4CQAvdb0UlBc
wfk8DsygWSsmzJLDYeLNOKqlE81yQokD6GGdZ/Fnlm/Pi+jBzlUQ6rIltw26bkOmpbjVSUmZRrsk
8DBd6EaBKDlwYOcy6dszcc7FEi4SveEDApjmOolJ23mWysj2JUdlYQL/3ZEJFuokhvqEj7jWtF3y
QfwYKo54+Fp7gbfowX11zHyBliiCQVK9DsBc1RuBiFgvB3ighq6R4yYZJ3ZjJNhA8UQW1C0zkOBi
2Tsc8hA68aKHIJk7GlYlecIc3yj0qUqxg3eKPxiHJ653EfGjHirUrhrdtwI5eHHG2a+Z7COn9mL1
K/sREMdNn2UhV+XMgf28YT49ayjs4xXtu382qY6d7Y/XqqodjJEz9UhXpcJ1asOM7Lo0vu/nyTto
LVFiOVzzOG9miZsZ16L9svjtlLy0zB9cpPCfFY9iljF9fXbNEjbB8DqDWTzpFczE5zzIZu+ANs0s
cV5x7zVd/S711xczMdUJku+40DpxTFGJkJ/p2nRAhNt/sHfVpD4IL8yv8PKRFLJapXlAb4nPzJPE
Su9YqPFunNsLV5jBQcw2tTniqcc5VWapmKy36wbeQnrLwh/ILVOhfCSj96mXd0vxPzjzLJxxjejg
6erd9PVnHUXnV+bv0xDaTvgObOq3OsPq+IL0HWRo/P2Ya0wxbfQPxDLXMONyxwdoRhAOPWovB40Q
rLzic9v6nvp/Y9awbgzQ2Lbxfz4Ps1+ZNAMo8IajtWDub4GF8dSL6DCzWroiXstW+Hrf+rzAeEfD
qyf9WCi8dIxLtXlnpiAs4pXtC+JzbQh7Q2vHcVOqiBpuBCMqJ2xdWCXjW0aIHNRIZwt9UUz2f4ay
RkxTgh1+LsTdWyrRvOvAsOSn3MSfEkjvIofAXOUB38CwMPXFEjEC4LKI5SpZhW6PXOrzuG+b+ikr
tK8YMBE/vvxxMCcy2rI4+MUsO2R8+8Kav47iiKLbspxpFQQpLhU8wKYjnkGtbkiG2BOzhWHbmehK
H0GZEX+yVIZZwTCcHN1eu2XjxeSTPfoUJFl0KS59lSeMHoJQ8qJbt6C9a9oqhTFBT6vx8HL4bac9
JNNhff0YdgJt50amkZxZ4pXJuJ8b5Nbpu1PDrtGb5TBUliI8jGoEJxv3roM8hHsjcEqNAnFQDKEz
S8MMJK+2wmGTpEz3n5tQkpkH9053eJUXo1u1CaflZkQ/7FmGLgVDPzvkSMTlHKtXLQWT8G4Bs1dn
LMgzTlYFUjQ0IBsLBErd8KwTwwXMOKrGww7PUjhc4G8y3egR/YaVDsLnOt9Mv27qu8GwuNbUFZy/
JfxxYDp0hqSMOMjo/QNwJ+IVHLe+3oIqS3eIEKkJQJgR3wI4vMZlYNsNIa1xTIvn7zeM3K7R5M1y
Bc43YnpBhb2d+oV72cHfyw3SXUoQ/joBJyHwCxEM2iVXE2C8jKklN2XrjJh3LyZiU+4wlgozTu4H
o7+cPpKWuhWPg+OV+vCZGw65T9pwV2f2zbOPXn2N52LLBOAsQLgbJrtO7osGa+G/SQT6CyF4UE6W
2u7noZKDfbXkzcPKsK+IhTU6m7hPGgMiSbvzYzZ/H7p1xgsiEIbseZozDfKXFXcGHKcmnDACdXDm
BKqvnQckjetKWCS042YHYc5gaeT1/T37xf4g4aVkUoLJh0g9zTg8JcTWnh0bwFR/yAUeVdGPCH3E
ZnOu3s7TIRrjRl+4j5AoS1VIasYfLRczWs9q5RPMHPC/URkFgxHBEZ34pNVmayJJqsyECaVMXZyr
ecQnxH/KCep5O1NcCSJwzK0zRSG4MiV0P0YmVflLy1ZNPVK7E/7OOMCeitSuogLpcjlHufreq3fT
T8AvFr4byHQu8PtnhUj2vx++UiBY62a96yj07eNSvv9VZc2cQlQLUv67isbg0rSspvKLMEHJ+rWq
rv6Bm8nXRiBreZZ4JgQ77dxEoCscVQdTFnNDGuB0xFdrJqIiV9apFO3eZ39Z3d8a5TxPKd9Gl2EO
c84N/ipTeWQcQqYOxO3pvPtCJZZKmwWXWOTA59+AKAKZJhOL36GIpYtEJ145BBrFwH00F5B7nRPW
KCBUAsLR7Q//sFHSr2kwgrmpdjPseSUcW0yyTaDVLSsBVjUlK+Xghb8M5cfsQwgatXMvBZeDUqs7
3LXdQzu7epPI937ZQncERNZ+oLv3wiJYBQOCHBuACxuJ+GBMpmDtRp01nCByiIRVhPJb1WXC63/k
ZHHmuAZFrSFVxfLcMJXkw1EPgPPgKweQmOF1iBRx707R5ZVU7nJ/vbe0XvU6GMWwEUyofJGHdZcS
mkjTo/KGUK23UMC2Id3+ID4yXBbXzGcjUmrDq8yiYtB00lEEl1U/R+NxBK+vjuSkLXJEOom+BPaz
7SAFVzIBzWu+kYzFXiXpRNbIndKJNZ03p401MPFyHPZ94TPyQFkkkYS8662FLPZh+AaJ4BwIGJoY
OFJEAK7HF5dp6q1a97W+vc71dDfkJ7KxRPGmPfx0NM6S7k8t36jhx9KolC1bPpNGmk3s4eDqD/5G
Kk/UPeqkRrzvlHjUhwVcD1z7GYH/YI4YTE+tfXZQkZlu5OeJbu4wZwr5v2j84kxxGiRLqydkyiFd
jFI9HsHKVoytQpB/k/4bXybOZXNmwsoIoBUtRK38OBNRle/30k70uLYOez82spQosdihZkvQLQKI
M87SCxOE8QaI4/dyXFJLNeO/o9cLeOJDXHv3sLU1YrrZCkJEJRnD2b/MxLwJ6RFIC2Vrbixcqua7
rQAGRItXJROEvEkpKmqP8eAtsFyjgsmwXnrKc5z1Vw1VryFGl5l5jxWNb++Qr3vNBN+PyddJx9B8
ad8F7kQ7jyL/qfTh9x1CicBXgZbKZcZfRGSq3Jf6A53dortEMg/y7OTquK/maL78E7ODRh6X+Xkd
0fO4ymZZV2ErSL5efmfKyza2KYB69jQnPcBl/VrEn1oYqvdquuvq0v5whlHnSv5gtAsNipjL2InQ
3XEGQeLpB/v/M9NAt/WmDoUMQoX7pCS4N/291tl0cgWbZXzrS0zZ9Y4kKs/IxQr+JoOzm0EZMTkp
mpEz/w35MvzR6FeCx+KMg7SFjObxDYibidcEVbGDeBxefUhC5/hiEVeEjz4fq/Ewp1h/OKuQ//03
O0XNXWCxcpFMGeAHxXBhtiBElts75FDOnaDlCi8xSGl36/wZeSGaJYpRS8vZriHeKFGSQAXC+Juf
cho77aUJpti2/jbPCY8bcvz3mA8i2e6/eZf4C39Ijr7D8ye1sRfsV5/qY0se7fNzHoZEEtse6gkM
TFHNlb81QPxYB5IDU4bJJ/b4luqVLaFv+o0mGPDhmkT4emvGNjOhchEmNMwbD6H1InrGHXSY1sP7
UI1+EarA+Bbn2oogLFcr89wq2t6D+EPzIcC42QPpEGaZCo+NmNYKT16aby5bnO5H9Y5RcOQq1hDa
moizdu/fbIFEPPgxOtQz+toajt1KPwxOjb8aBG42GGRJVh55SvlIN4VK+5H+0j+HfyRwmHoXN4oz
batHxPDmAAmoGlhgrLxWaAe+PV0HEM5wycrbm/vb7Whvk1V9o35FzYUeCcJ399cuN9n9FVAy7APm
GRAKDugsO/XE0v9lyTx5eK7m4foBfMrPSspYq7ZkKlCATQ40+KsmMB01vtdFaDZbFvvNv8YtCSlj
iP5I+fXIHh7xUQiqlCqkS2sFupUzljHeFMzOGGBpC+eJAouXwROiNEjFCCHOLSXvAhLy05xw/PWG
lPc4oZZMBLUvGdGedhec1wWlNcxe5YS2B1GlDP+p/ZU7S6ZJ4RjswRjTGVgccfpnIcpDE4EMlpE+
rT4O5qlDScAemkKlDy4DPsZ+x4Nbrc6TTiCepURbcyjhb9G1L4e5uaA/TgQu4L3fkkxr7noGMRwi
iPQ3e99G5d7onuOwb7mGPprsrIimYnqaHJImyhoTVAqojfc3nT78esoCDH2ioEGguZtrK7K9HF93
vmxy39+lN329GPAyBKJkE7J6Fen8He4ej8wB4T+TMYcVnLGXBCGOCctpaKUqmDbd8Kv0FudeqHxV
pHn2eVX4dKkPeEDh/opA3jdasQyUJ44NOpLoEwAYsex9MNI0zzMZgk6WGne+00QqxbbtIyAc1Bl8
ptgFD8ldUKvhBdTrZH67HFygk2yEtUt9TXMZv8Me98YhCySjMrHkeva7zzW3yHDUhX6QycIjGMby
l+z/lE9rbwyGpylXrxFOs/5lk/dY1ByBPT8JDmt1LvyZkkE8QUjoEpLmdRWvdCf5pFTrYYo2b0kq
OWwdwCZsB8GhYwWaznwLpx9vZWoRPaxeD8zK1CgcK3GpINe+Iyc6TZqSBmlQ6puvRbRehREof5iK
/mAP0XN+mR/Lv6Ne9vk0KBwUxrv+lTQicvqfEWd+l/VWfvc88rEe3sHd0r47qesjFjRU+Yw0W5Pw
JCHFclgjCbhRj7biHdNEFxt6mn5jxsgOPlAsmTUiF3wyyTim7Z+zSREj9atGiXUbCPT5VsWOInIz
A46UW8mjR/23a5Z/ySCGj5ivOzNv5IlQcXHL4Tj88NviQVoDcvovuiWSp1crMDyWVqu+kUbBL8zq
FI7b2bGeR92T4Slr+t0vIV0y5lqgTu71ezW/3e5ggXb3N2YOm9vRXCcH1I3OTtbTO2UTJAKSIPta
KJXIop+YK9XebsNkF+EBijsXPlR6LjsQn4N/W1ISmVhAQL/LwHuwMLz5M3pffhefwDIVWn/ackI7
47yc0h78NxIHiZ/YeGx2VcePkXFa+AITmQcpX6XkvcsACrH+Wlj7gVmlwXc1g7TJTDwlydlpjDzg
iHJ84GJmwVUrF3hiNyLKbO80fWGNwHEgMra/ZXWGxmLdmF+isEA3pj/lyfaeOGlOWvSX1hB9bDWn
dSfPK36Oqez9/YRIGogvhnjZZZ1hHwkT0+Dz4G6fTzVjWGG1hbT7Eo+xoq/ztp/SJYCWmyYqNioD
/l74BTZgqP1NWkzVZmmOlFNOXVO8EhbhD7X9fO/d11KRmuLBMztwiZvXoUjcfEZ325o9G1/4QRMM
EYNg8rgTi2m9DlOkchvNd0rEJc+ZIY13Oe4HIIRuEuntIPG0ODNiTEQD7tTAqor+wY/ylsc5jmC0
8BN1tQ27Pu/jlQa7aOG4zv7UT4dtwqPaz900qLwo+S01CgOvSdvVeCHrXCdgvdi6Mg+3SvMS64w7
n6gmpMYpw30YvUWC3M7e0wLQhfxxHQFPz5zaNgc08qccaKW3jzbHYJfSImbPJfc5XWKuMeD1o0ru
N3Bi846hHOdumO0MCRP8A6kj1Os51InwEbHE9fcucr/FOFSwiidmgX8OmQa4UHrhrC46ldp5NmtJ
Fub1R7//UBcyy3xQrtDpwEC7fVwPt+1MynsRU/vrK/1d5CtdAiDIw2JCOa+F6QF8/Ormf7+DPVzB
rahQNSoNb9A8P219pl6tvfu4dGOXM5lW+VUN+iOvlPnMsnaQDSp9drFkZUnC3XN/sJ4XwE3ZvUxy
Nj8yz02dMOmJf71ZYHtLG+p44U7Kw+aG7IS/EKrjVT2w236GJU5ZI8zgjuLcnyTy6FzC47ujGYEy
e6CC8IbTiMLQGP9LjHVh9kHL3OnXC7LAOJDjpUp+V0vzro8cQrwxM5abfcDt1d5UXsuH0NogMMAK
+pldUA1JcAan3maGUBc2zch1OeqGuVlfMkDM3u09QPBie9kQRtEOw+y/2uivtIMW4nWoW8fi7vGn
aGhzjZVcQYR9Vuzf0cxaScHuFtevey8P6E05Bswln4+vm1TpF9NjuuK7pfy9vMR1JKKg3L6RV8Rt
XUNVekEmhu5mI4AIHUGjSPLsTNWibsMvK/a/aJXhdh6Ool6Lsa95Xs5KgWQa0ckGKPxEXKyb0J7Y
Mn0gZxvxtYy9gVqYBkq6F5iUYaVhdp4XDtvUXHo/NVBHzbo/gOJpSgZLTAUE3SiPLn2FAnvNFufI
LL5LyQpTUFN9QrINtjPXZP+wsXIjIrh+8hDmeCFT0wDlHKy6RKr0jSAgNh/jMN/YykVTHzGQv42K
f+ollgOEK/gMy8FmmgombPbcyOYD3FlQS6u7f9hKnZXxIpxNmvMPQNaJy4sSeBt/XI9pvDeqaX1n
33ONTiZoFzOmu5iUDOSI8nlAzOQ+z4blOuhVq8rxPKwF9mEVZ8OzxE3kkof4vZMqrpb1YopGLWQ1
lXuGmRROrmICJvHITXenNVd/J0AIxZeAc1lQ4ZPZQDOldXEUMwsxwOXCoNdDsTt8h1oujB9KArCe
RxqMkbVlF89DY1gDvXI3UU0+cfxu3/tkYxZ1MHLGL6pQ9lNrle4HoUXJ9UT05TBWNPNBIiorfToe
aYiHuxBPc/W8yR2v3AKAA0zFMrDRKku0u40liIyqRi3u4p7syq4nrPwPH9DWocfNLlJKBZiQoHSM
3fkfczbR+6SLzdkzwU+snNASGNl30o0RjpB7jmLYKaQvwcbSNUtaJeBs8fqH00L+oaZK3ATicxf8
+S04L+qPGVRyRGRSyjnVesbKV2CoZxeUuVSRVeS8jSDJ2ezeenQimyGDNSp9v8jZL5ihXY0c+USJ
5ceAutZHetENJlT4TQnMOXxBr2/AWVR2jVUYBcja4TNw6LqZbb2eXauiEY8L/+IzT+XE9PE2SXVx
lWKblDyNRKU+k3dp9WPqdgtai2or/W7C+RCxVI8AoJN6AL4a3TQ/pB0b+FFNhKFyX854NWRYeiuw
bLQhDHW9W/DXNkfRptTtFg3z4RlyO5z5ssu0Slw/7ihq2P83PiZc0qQ5WSLA3CkFw+1yme1LJ50D
n0NJC/6S8lOcQqRBcjpiWxe9tjPaa/EeMSnaaxAx/QT1+wsnHuyP9I2EX8hHUwpNkyxxuwaNsETG
bk825Z/cVGbUHBQQvhlexAaqlw0dJZeFzIzH33IH4Nv1Scs2C5bKAOrvNgj118aWSLWOzay2/pz0
uL4UkVDX7qWaad3gmEz8B4TnvN0vWntKHFD/Qtk1C5Fg8n9ay2A6twscU3KQ6mOxZWK9kZNb/uU2
0zsKSdnjUhUAA3+VhxKk7UwyUSt04Ct49A7fjfT70bU+K2Rgd6EIvgwdsRdCs2kmAx+g9Qz5NP1j
bUtxEIsPFeZYN4q9B409maWbIp2BTmzLnHQdvv88sY3dZrBRDqXWNrKaAzHhdgvm9h45fBnLTML5
dtEhqJSWHcrojCq3dSX+JPhWXsuEAi9yhvLCK27nQ8gV5GbHt8AVHa24HdqZ5Bhd1exdQ+Wt9llv
MpllP+U/AraiQZSQ29r+3gSNAm1KQNkGyZvOsQVcrTYUyAG6obmXkeaVISeEgIo7u4h5cih2V40d
o89mVpaAhGJ8rzGcYhbqc1nsyTUDSEpJDj3ceikFIYGW6MdbZ+TsrHJ/TuVzd1/zwEYf7bmEBTZA
up96fIUES9vTQQn/kCajSQFmSMjyYyj+N3ZDACHoHYzSewHGsT+2Roor91s9Fknp/pGtniYf/kk2
iWqWZmgPnjHif+GVL+pv8XiueOYhCgU3BC6gLP2i61nx+JSoNtvEAKc1VuzqAibhr2nx7AQGKpYA
/5Npyb923jKyALJ0vlG797/T8xPAMV2Z2Wt++Z1dMOmwWRT/u/GsPrypuLySGEiuPL2VE0LXcYHc
sk6RauYSIz05RgyYsTvEY4tYg6KzOS9fHaADX/lmi3MIBNQWlhJBGKM4E/mByPzfXtkhKvycT1yg
mFAmjLrU2kjwF5Fud4z2+prBM8MzbTxp3nNcC5k88azQxkqldmO13dmhT8qrMNpe8wTlE25yFa21
rzaZOmIqvfDABMijJw/Z3JsoSiDoknCPfNejOCusXZI1s5K9Z/FYWlDO24kQpx+HzYoubpttYdr/
x80up39hCoOZBgulpJ5OJgrKOeyAG/GZogTW4nbLAj1B1t9FsT91yYcdTKMxZwFHd6XzD56VLC+0
4lxcBHy777G316/kmBuVbiaq7+awHkLDRaNrBk0gFjbuYaFFoQpamSm4nyuDKWWSidYp2BH8x3DK
BaGuksVVEUMKhcsHaYUAWeFWtdxlmYEAZ7bdraPEew2p6PdN8oD9OsMmCkJs7z6RgokKi7qmOHxz
zyk5mrjTsGbHPZuFt0YWvEfePBh+TSBYDeQJ84dAY+4X253HvfxMY3wIIk/dX8J7SZWwORHBtwlZ
QE2CL9dudk1/PQ3LUDQ4V9TA+pF4CIIz1W9wWULUnnBRk3XnLkapTPVyI3CFiE/k4igL72EYooaF
/NvIhpoV7IYak6KimtguUu9qv5MCUJhtPS/evaoGYK2WmKlqQ6O4EDsQIldRzrdpbK8wzMLllOrY
CBWF2pnds6eImntrAPtDloCBRkUwsRGRu8FUh9OqwMP+hEJb2mtqdxUOPFItnpe/eKETLCc3GCr0
lAWjCjiiexfNusBAJJ0wEFndk64/esrwWWoouB8PLi+cxMK4CVp3lGu0SXHHJ/f4f47lOYzVL89G
Y4GmscwbaFQtZjR/EoGJ8z/f/xJcbCEYeeSoONwCaJ++TpQQwpGVs6502XLCg3EkvaiWXfqi7s8G
LaN97M+VLrVL3BYgiEqOPv3oYa35Hn7ARFFO/oM72UqfPDimcs7EeJC1PUzSism2oAatiPtkYrTY
7svRVuW+Bmn2L/FRGLU8kWLoJSQcc6FJbDv5yJV+o+UaxLuJGlMUYMsCmuYaZRY0p0uKeSbsSvIy
uLYgmZ9LfNSpy7u7mppzDDMxsJyQyXz/CnYI5jxMIWyM8lL6K/FK5ZBApdLWJg/BICe6RYcX4Vup
glnsaHAxV01s0QAwELCInc9YZRqfsIGM7vlH/bJP1CfgYim+nLU8hScaben4AashuGvu6WTkEaXi
bDxWq2PVm+ACJTKCuupST1eofICnSy++Ydh1CcnUeGtInMt61iIP4Xins6giqroMae1WrOY8jDBC
tsUkWMrfqc/1nngG7DEx4I8Me5aVH4d34zkk7SG3oPi5sotVmUS+Msw08qmWk2bBMa4LABZUjVBX
dDYK1wuIgpUKcMSfFe4iujCiD+EocdBZ3GHYUcINNpDkoawHKWRUG4MDp5v6jPAvNCZyxNOD8JeC
NPsWoWA7hlmzFxQgdNJ//N25WvGXEoV2qelUPrswNXaDDmsp9ROksKXglUUG5zKSQXfnn4Fk8QRG
hXoVxwZI1Tp0f2ZwntblaqK4LPNZrYUEim1LfAiBG31OlcOX1K1LfwsCTDtVHMe5YhfBgWxptsDh
SzpqpscV7w/+VGynk/GsfKkuikmkmO1ejIHMYZ1TyP6UbiN1fGZTCJ4TpQSUgknXfEIqB1BWkIxq
HsNX07akRP3I4H08CltJlUtYcL18Ua+0ggWH2ueUubapK33ZAXN6WaEyDbCRVCo6sNQuvXIpRqBs
d239IuekUzrF9A4+iSlikjH3PoxdCDWGBZ+lCrIR72ccx4cg5jN1+o4y2HilJxQQz3QQZg7G2lU1
MzCWK8fV1toJfAoiPdA9mdkp6BEXsPK0Yk9Pvj4Eef2Qkkp7MG9qCES8nlXW1VWEddAAArbAqKGL
e1JiUg4m17p1zxPeqTaZf22VAZOBKMzvvcZyGIH9DEpy0hytIDjhXNR4IDSY92uwzmODziCyljXE
DK5gxxx/YscvyxQIYxNeqVdKI623XRi9/eQhaYoOhwSDJyi7WSW8sNnex4rNNVV8SlyrMFRwCIkd
wI3B7ITIy0ov/3i8T4WjaNyTzITu3A6FKK/Lqwh9wmuYcFbQpJk/cvnJmRl8kJ2ff7fURmcLs14b
gC4d7Wxij6HxoednMPolTwCoJiGnsU6+bX9WBkhwDWCkn7Ue3TT0JJHCJjCtfCXcgWn8bVORwG+P
cp8pD0f6e68UcT1dBnZqp4opw9d1hy+i/w6FrDQ+v+iIwj5U9+zDisQhCGpC7GxwpftSNCEvPtNO
OxPRcE5BFSWVqO//Tp5L+N2VpjlsiMkWyyjzGMFUwjbvjjj1W12cvbHl2WTFbaAjDHQHDwwmKT/3
TY71PHg6RS3A+yfEbG4FTk1lO2iOQ09CRfs/kQb7SRwVo0Jz2SyBHnrY/s9tp/UpMaRXEtEt9xSy
qS5eS5+YcTkN2MRyogGydQqvz9Y1waHJCvQ0R/XXr3P4HtpIRD2dhQO99t6MWhnB2Cv/U7gNFKry
50OYvXko+tp6LJE9YhTVKJYRz3Vv1/2P1TbY6/Mdi9gg7PBSizqHc+0qL+WNxHoRF58NZmQ6EJvd
7XI1CSDR7l1YLB+lO0eYAyvBBA70zZCp4prmadGwXZGUNh/08paMBkCnhwbPMRZJyjwq15FJct48
mzON8ca9efsLdlT2bP6BFC53NmyOVIkyMzm5sivOY5rnv5+yvgD05w95uJiyMhDfHMOcZHp7P4Do
QyOu8e4gESxwo8QJwWcwSB///L6H3WdbHTRXq+CcJOu8jB2H/4yj/nueS1GzXF9ZnHUX5mxo+iF2
aDBysmse1ei0TWA4UYNGsnqPG3o7hj4h/JG5P14RRomYCYQef02AieAiuKwixTeauwfaToJV+FcD
yYWef++ZWgY8jmV0UVIm2CI81Jc99c3MEOjUBHZKB+o+fSbG6f+EL8t24s4crmLMlYA8dHANDcrh
6IqZjAkAj0IpeYww1E1l01Fqfoj8ONJUMoZprssLhAfXmwRqDNK/rVVCfP9g4yEX92/EMAelQae5
p2ysfw9JkMXZlZmarwq9t/M5QsRKq3CDPf5NXrtKVFJJATXYBRExZ/Fnc48hrKs8QnwZm6qmQLRg
l7rI+4RXD2cLXby9CpMLUEZHwR0fgSKs3f6W1ij/QrVSiVqGakd7FFeUYYzXhzdq5F/jUSm85One
Wkhc3VPja7wHEWQPaFo7xtnmhL3ZX8/9+QiBpUn9bGkBD+xMYtKg8iPMQYbwcJo0Nxt4S9YYNUcH
RvIU2e3m9ANuMmOOmcYS2+W3Q/XGDg+uFDiAzseeirkywIvdLvUD/5Zy6aQguGtu3DaC2XJP3yzD
BtiSVEHsYEctBjm84bfDJncLlXAr2uCdRQmHz4sT1XZljEW8crj+BndyDoGZysCfzYjE7g9bVkq/
ddn8aOiAQe/zikkBQPIqM/5y1Z52UCJCHDKeA9GKTP1wtddNmr1tQWmeFNnsYfytxLo9Izg9YfET
eOWd2s3c32/dN8YCt8ZlP7XuzGV6+Za/MebYCPCIDaxUDYJ01i1vcCLKPz0YsA93sfa9XLSxpyxL
3F5eeiSE/+rkDY59XjPnPBYTUJ2aFCtKvTqXRtI2V94LYINDX4VudgUTDAnmMOvzZj03fuMwwekN
6BRVuazLXkjwaEUofLEEiUBUQOzOt1UE+MPHHeQztp7SOIkSpObB8KJPqiN3KEPFtk7kitZM4GFz
IKsSQWObzlxaIqKqKfWXU4rKegMUmfBAvZTBs9ZID1+hmjd+J466wd0vPuJVaW+Zt8Aii5+mUblJ
BVkfz+4JoJistrX8ge80qXxBm2SRwzsMeXyLbunLvUCthbi12cpznvZD6LZn/ZcrDSM+TCKuaCUV
DotqTFPOQYmPoPKzWkA9j4xPPP+xNNvxbv3uL1O8isi/FMlO/l84rhvWO3JbsqJt6tU1jFlNY2SS
yXdmISLUfTibkXl+8XGpbB75KIdaZRvagKM2DBCIAIpShaF/i+cBR/viOpY4b/qmjys7mivyEn6Y
+Vhj0J36wIvWC3MIWj4jMsZSC76k5DLIRz1j3OLNuxxE28DUMXiVhWzWWDRlop6JLODNqn8u0+PW
sNfxbsxJb18ILXNYvu5lMWSQdQ2c0exWOSMK1ZTlYTPIEF293ouGgegzmV7jFB3l3gHMpqtCLQfp
mnX4F0WwJuRZ8V1wj6Ejz/yMkIonu+5Op1LS4CeoExyqIhgkqhjBxRspb188d2CopOH5fbYespKE
PndXEQWTyqLFqu2RTaaq1rwLM6mL3/nq1uFo16/j4nCJJhyg7IquBHTkwgpkaqqJaLKYMmkRe4sg
wIevHMtTad6Ot8bamJ1pmCtlLNYgq75CroleTm9XvQTpldneInwOVk4jK93jhzh+SGjUVUkrHOAr
gmc8ioKTU42Sk2H54g03f829LVt2hVCAYuMHjh9mIlgmCzxkUtHyGiVMPiE+dVF+2YjPCsKci00Q
0v8OxvuYQTqw2x9rOHYuJaQFpT7AzqwOeUsQE+f+kaj/qg7TmpGt+wb1T0WVpyCQLtfF5Pa1WFlE
cT1twwSdd5y2kecLBKGZQdW9b00jJZO5NAFJ8xsKVJHNfTC8lcQr8IMn+F0IGypx1k0JK5qcHOKM
02DhR1/FgtuQ6xy+vS+UTgXwMcwnOnMoHAQhYC4FYTuHwyqgzPluqk5VxHMAf7va4xRMqDVHcPde
hQprx0jSYvHdHRYAvzPUWQM7aCcqptBYQViO7fgU2xJ+O4GhYz/hxsDpHf5SFCmpor2ACPhBryoJ
LxkflEc5z7Ta/jJggM7hPQKz8Y36nUTm4ur4bMTpSNnX55gXC8Vduztd3GU/ih7oX3KABARTA/4e
bFTgCrXvq+KvYXW2TDc82LqsTlvaepRvStWQN20sYDadoTgmJqDzzBAys0vmtcTixSaDW4eHBdG5
TtqCgy0RS5q6bvnRqDrCyKxh2+6k/fDROdFRdKO1U6omkzWwh2l5ahuLRCNevFGVIdDHbHq+IaRj
aT/w/8AyBFtN65mrqfRjoXahQT8FcE9eASQ8MVVw4ZVyQ5z3fCPtb18JdWoCf9osR9JuSlWmcNQC
uGZPrHgSrDA2QUTRK7yXgQP4YmGGY4+1850ccCEY+aMr9s7rr8uvcnFHmL2RSXuivD38jQ1LY9Nr
l4sstICcuHQRP1vS6x8T5DLyi7wEjwM6oqYP1zTdRB/WaE+pI8vXvHLEpVOemLRQbUkkGKC5vttF
sFV3V8XB9WQpZqhlIm6RHJBa3uDQ27jy1hwDL3WWIkq/QSyF91Q0ZM1iibCQ/m2q1+0/qJSk2Kjx
xtdUT7deUwDCxpdvtj6OhABAce3SqxY7Yd/cASwp0GK01eYN2Vc+upuOVtQacTl+EE7+yg73d2n5
nTDGnbUkjhsMb9+nqRhP1MzjsrtJMeJZoVNhx7dvEi/JhyXnm7eZdTWkMezUJf4zOlG1Sp1Ht4ri
IYn26yoSXB4FoKogSleIDsjd+hzl/DRKbUXNdP5w4ymOgVZdo3JCFCbDmeFXAshtkRgwey0SniI+
S9oekY5KFEQGwjfLbyFLFvo1Orrh1s2N6NLQ/yzwxI8hvyPcvdy884tyybJ6UfWSxzC4l/Non2Gc
0K7oFvTw1Od6EtffM5npQ421EhfvZF5pQs+sDHHv67DRDEBd8y3pwaV+zYBwGAnU3zszwu6IuNo2
pMMhTo+TrRvbte3RnF9RsVmUTIxuTdmJTa3m2ZSAnI/bz1VnXnHP5SXcFY9ItD/u9n1t7812xNFH
55VqPUl7sCazhVGEYrSds13QV36lXbaSCe5IJU7k0zvemlJlF8SGYznIW/ULM0zSY1T4lbDBY9Mw
SMqjYiEdW8XCyzuPx5hFuMzD+XkCC/EbrDI8e6Cdd68PtqCUm4ON//Z0mF+L+0xr7ddHExNvizIT
WrEZoGkylrBiyYtGe7RRo5LT92Rdh/6GtTJpxhp1MJCuDUyG+3M1tAf7nLIQ/BloLFsP5CP74b+U
Jez9F2Q1CtyeUsDUlwyf1RpJSa2c3GwS6PtjNc4T+5LPtAA2t8KrcikOmG/vdJKfvsTahNyzgK+O
F1n/7kxshqsygeSki801V3LhtSE2PhdRQvOtvAtu7SN4YSh/IZyaZhxBZIlpoEphb7gHo4Bunh5r
OGraMh7bIAgVHr6bJ45ToecmFKi3spQh9YYDGdlbCn8FPfj6bTUoWh0R3j9C61DR34jFLD8belnz
jlmdMvnqmbIn6yoDAKETlFqEimiCU1T42+aln9gtWt8mQxV6uCPV/QOzyh/tGiei7jcfcOBCKfAy
Dqdo0DtcWvtE0nckQqRC/FZOU2vduHnTaFDbYd7eU2SKnkAPC2kGMaBTVNlH8A4m3LVJbl9WJLib
fbrDvVKylPDq3JU2lBE4lsZMoKG3RQZ/G5SlBHSZv7hoCe6Fg4GyE/lRD8iSPaneWHAZGDwgEGpl
OEh1dHHHjXoMgjYch8CDudrKot2s0cFiT5Wwk7CJ1pd307Mt+7pk0izrWs0ViMhi6A9Ci8vz1D5v
hqNBg1pkMgDubNn41Q3e4F/qXo7CQa3pw/Q+gH6s4HZ7lUY85HrKdX5TKKbmsUKWRk1Clx4UeK5V
Ih4Fh6hKp1hm1Fe337Yx/WzRAxlxFeHwqSn5jgzoJfeo3iAVbF6S5LCaTHe88yW3Voy6eDOTH71s
FWhdqWKDby1fyt2e9A/6kh5xW+AjQNu3zfm8ouVFxIAJliw5jz5sxGK9W/o4vqsZ7wPi68aWvx5K
ZXKqy4/slDfi3BOqh46110LgLi9mwtOK0bcXi6VHsmvQ5VhcR8pPMGgFu80X5TAkZ4pE/c4IVDNP
mdsobywj8YsONkMHXjnaYaaWEoZHS3WsGbT3+1bpHw66WEnrwcilyVZ9b/a6sPPU6LlpOecR13uN
lEg8Yd1VAZX4rFMBnsuGsesxKl6RMRZyRoZErqS+syf4pHLurv/W96ZVVMGrcnJEov8tnoz1sKnM
s5DSmQvBufCFVXdu4wxwhO3UlB+bNTvrIGZb1YMi9gdayGpp5oniFT9rmjW2YbKgpRF5oGZ8fKiu
ArsmPu0XxcWpDy5fJjEDfvRNhfgnNYBz/wTNmQsfM6giwFO64PNZzC4kiNPOP081Qjc5BeGzATBZ
xTSoUPbPC+JGcc8hzKKn+Jn1USwyqa/6Z1+aJTlwPhfHCmJTe4vlRJRViRnrP4rpjsMSFOTkFpK/
kVBIkcgD8BHflpRvqKGHiUR/BX+SMAut7mCqGnB5D67hBKjUJucI7p3mxsM0oxXC5gCKsWCDIzk+
eSS0/YaCW4lJFvC/9l0MHb/nrn9bE5TTuIjUkrIopaiN3uw0WCpYghQjKn2480uQy+P8ceSlf0B4
tXgDxDpFPfmQiHeGi2yroBvi/jxWTaK/6uYL57m52X7US6keZtsF2LimNwOFtyEAzHmM/1WDnrMl
jG/018rLxMuf1pZz+LLmwjAgo4/oVI2l88uPphh+pxYaLslYAhYJK3XXQp4YDRvbVqF7ThlibPpZ
o09KCIdSPNp8CSd2hFo4HlMq5DRBjw011IiRHROi8fK0BED81oEtXx1qFbVPqcqO+7+9hXa8XRW8
YhSlmNW0dG849oMw2dKkUAHPDjOdx9b5bR9A+cCRNBUR0TVRJrTwf9ZkbfBA7g8R/U+V4VCBCnda
AdkXfLPbjIJK10NnPnfbGbR82w0GRQyBxUQYjjSvZQN+ESaIw8WNaAGy8uIz8wXiNW4sIOcd9E33
Vk7oPAQt0GKN37r7UdWYP7znO7U2vmzEXhojDtdz6SsdikHb/6x8+T99B2TKg2Ju/T8k6qjsWIlm
Fj7LCsY8SRxPWASp2y5oKVEpf3SOFF3e9rZDoyTpK9Wf/JNcO8xlw0Eef4s5lI0S1Vcb2kf2Ms6a
o6uFy0zsQAFe8xvJ//FPd0WydnLP52sJou2S3EK7SEFAb/MbmBrbMHJ2hjuc2PGKFhbdYT6ZVe5C
4XotlAnHY4/5KmAK6P0vlpaPAlxj6ODq03Ve4P3XUnCA6TqSZW3vTU8j/5nFiE1ViIcTOlc0Ktmn
RDR4am7XKgY5isjbojt7dYBFvasDciip9QmNzoo45ugAewNlrsfIBJ+fdxhJrth4f4kXdUipR7aT
70kJLsampC+7tZuJqaGWKap1KCigfsvTR/92cF92RcaTqCLZ/KfNx9988MNjA2SK9/0E4ReD8q1N
3sX2OMmfNU8KRBB5L9Mbd394QPesb1DUX/IsgY8s2i9g+xL56xDJx4mtbULP10Xmyx6oSbukfTaT
/u1ntitva7hkS5mF5br2xHmevqgWjTxscD+kt4xMGmh5/FzRd+9EyGgf27MAvscluxeiqREiSYgN
TcpqDm9QZShVw/5Ze4wD6QuzQHH/1bLbHuXMcQWYMUFTCEt3TwmOetEA24fWua3h9A7m8aubsgJq
doMnya63aZeir9YHoutxtljPS9EswzrOvb7f71EzIbUGrTu4vPWE5UmlFt/cti/mVZsOZx23mhTV
R3sthvVU4tCC9zZav6z6aoIKTbNXGn2ky+QdczizkbwsjYX08YFbkjFmEj+BK+1hNtYg+ww6wMBd
bf9UqQFZsyR1mGsaW2UyVyVn9wo7oxJ8BSgA1cps6o5sLO73yrNiPxIxYFl48Tjo43QYJp2vLcOG
D15klxGxUBzjcAeCoUD/TcKguTqIiYZX+4wb40sOD9U1IPtPhQy5n3zUMhqax0wcrFTpvtDclPkz
nEG6nBPf643+w3/7qF18tG32eyn8AXPcwQSr6ZQvuhKw/oGVahxs0qMZltZ6jL7NuaUy1EatHydJ
8tXJki9FehsJ3CZ/jWr5A3oa6SbtQn/fqbzyRcOuezvv36k/Gw74k1cJVPSfuOHei0nmIH0TQhXv
GoI3AkR9nH+sui+nVnjb+bjmX3Bljp07KrMcYHoQCtRufSg0JavYZm6n4mgYPmQ8FyIHJerUaNj+
ayShyfxEilj7jJnVVhX7uxtc5WqP3i9d9DCUSm33sXTEZz6D4qUmS/dyTFmOHgtFrUNqpQTpSE+T
6Hh2KmwcYzlsfuhmYMdU0AifAkvyBY3yEFydM4qetMIPMAb5GNX/Kzk481iYl4ScgrLJq9lnJOyp
1Sf7cVmhkhQ/UFKw2iAGFL/KnNV0hYJi+Wp5WUXwxvJDxulAk3MIldkvGWj+L5j1U01SGDAhXNCH
dP4I4Tp27/JsDpJp/ZRMh4L50w2/ks5Mgao2eRoiNABUrlRDpfweaZgqB26tZIHY4iVGgNNNseE3
heSJrHyiR1GXIRHswy25UZqBnlpeeyCG1fQ1moTUcu2c3lENRsPT9AupxZbkuK5OtpRg9RUV/Ag8
NHvvzppsAWIILF1hGQaobWok2ey6CEWotefrCBIstrcNEY4OKpqidOZiqDYelq/5LHe2Z8kAnPTp
scTAJ7JqS5Y02zmlyU/YMK627VEyqsOIaPdkf90pIbFngu7l9AAfy3c3QRfXhMWI8qPk2DoZAwG6
y3NAVw924FfUFMpqySc49ajK6oP7a46THi9TsNxaenQVJMdJ1ClbNARwZUOGkrU8m8tP6FhCOHo4
ozGJ1UirAFJKRpCjPaTQkiWG8yn4XKuLxyTl1JvDr/163yQhChtJW2+nhwnkq4dJ2+ulDOWCm85R
WWix1ma0bkt8BnMQebaYfRR7eTIWNLe9fJaSCTPg7CDbNHijjptmLvEIIetqbQwsCCqKiuMF5mAX
EvfaeizdxCayrUgDpupCPx4ILWMXVZfrFzNyVk4jL3yKePLT6fAMfOGMatbn3DsF0DHiMRomv/I+
0+h67h/E4p+65OIVhv7hM09bY+7ZAHtruUs1OLbOfo+2E0HQuVJlK8awnLT4EKh4mlZTweLLFLx6
XPbFhORUKbvks0kWtHp46Mz4d3RiEZd6ve6+Jl41pGfAyB7HNIE3E+QqMMkPuTMbU/aodj29ro3l
usb0WOBxViYsuqptXWUhSky9IRBVwDw2KZiV7P9H+qGGZXQAke4Ln8z4ABTk9jAo4Fs9vKQf9Kof
M4ivM0rO9EX7h8QNyuh8FxVhltav4IUveUF7sJCvGUPX5BVVoRU//TBd7L9vCwRQWgfwVr7LtY8F
uJmStXbiyb27OQ+H4qWS0OqASYceE3mNTFsH9X6cSyFbrDB+CfqHJ8N+nwM7lobAv2xMmG68VYcc
7x37p85FOhYOQ2VplMRJvexRTZeZaNAsF5JK4i+pJSoFo+tBMgWjIplhnUdLNz76yfKOBVoanOSO
k5bJXlFbda8bctlBnDYCjjVO6NcJTgPLPJZqsnW6Aneo3lAVMX39E6c1Vt8nP023KZVpQ2Ouz0Pg
l4yqNsqZhgXmBuh5nvvcQGP0P+N/3B06Uob4VyxAvK1yvi37QWtD5Tufwpx7g3pIFjY2LUNgcluK
sFryyUfZqkXWiWPBtMEwdCsR7ACAXQUrvsvUstTx0xGAafhN1cYvtr0uZ0uHWXIldCVKCMhScVD1
0iSrwSN25fBfLRgOWNPyB707XFJduDIwAGZ3dwf+a9adOgfJJTz/+xFvJhZQTbQ6lOknFDEupOg4
0FxxSoGGeJ3/a2vI2vbrtHlTbK7u6GqtKdFWETBcyDcO+7dpMFWUDECuCtF/hvC0kIhLRfd+Ics4
6PwJIMqfqFGLjPJCfFdWFeKRqlDGij+p98pUUPe2iD1gVWcTzbMR6HRaFjOZ7biP6xWiVpeepf3g
jT2gDnB6N1W9KH5SZouCkFKSSYiz6xi3sGyOasl8syevgt1nSMK1NPkubKNbUbnYMEPYx1gT1fPS
cVnWN1+/IpZPv3GiVl++4iTSWQtkWp9HdNcKAoEVrD3qyEe7xZAUiJdPxue9mJycD/5S5lu0+H1L
FKgXwynI1fJQUMP0oanREQDH1W7AHIhUXfMiHxD3PLKOnm6jwn4NLw7bb8uvMT1QEQpZ7/W38IM6
vpdBIyeJ5eQHfS1DL8IQAvZdzzH6Q7JaY7tVyV5LiSlSSNSzDrIIwvzXFmDgg0W1JixIRkbxJJ49
5d617OZigMwRDUDMKYIU9wtIIiTE6jUTdprA+2zbZJVexvOS8zVai8ZkSDt736OUY4drMHYeSqDv
EG0lMz/hCTK1iZrZ3JSJSIfToH3HjBdyVu74LsMVnP6sDy7Ya6Y8eeXuDGOA9ZzTD7nQikM+sYPv
No8pCng0xbaISwkKNMXnlKin8VspyloRrZIEqFGOIqZjUR/GfmO6aQ9+pAEjYvTNhJsWGnncwTup
QkKaniJJWV0wKvXIb9bjzA+JBRIIcVCxr/Veqrrw7U40Cmhi7D8u2z17yE7lf5L8Ki9J+xSM1aVT
EkUmP7Iyr3mRFqLrYtgbc5ICYomsiwzZJNfSYoo29PlsLGPbuJe2ObRG0AbggBT7x53agY6MyDP7
KsgcxwG4I70SLYNa7kf6KvkUlHTYnspumLmLDKYIf/AoQHbkaHQx9mVZOACH2xkiDEr1gIOprrAj
ZZXQJ6UztK1N4QLvjvUF1PaunGdYvhrnYjVdsngG47xV7MI0KFevPofBc42tkcRfOhpY1NjLOLRh
EAQ8Q0uCSIEdkdSXv79GgmjWnwbeyzwenEA9aMEFWX/o9s2P5NqtB5por5gCp+VfEdxoZeLcnlA+
HdI9l5w0tWSrvLbzQhu1dIE0OZlhYfDSNxs92wloJlyQ9YAFlZLWeQMGCndXiQgwArY0w/Pyf/Jl
Ct9oTqEt/j6CmiDh44OXvLin/s4hkP2A5W136rVKPGVu9ynN+ijMvlR8hD3uU8pY4yMirfv+jZxw
jDi3CKLT4O7eN/Qo9qQmnprIZOyzMsLzq+pQ8qwJ931uPDSmmiAQaBkKce/8sZKO4zVIdWDc1dEZ
rFojVtmQqIOGPQU6DLjo64ZmCLDvxhJvZebUhbafs5Ms/bZBX9IqV5h6AT71tS2+a+OyOfOLcqT0
AFWf611CjXp8PKPj5wmvfIK/NIrdRE5nfCYAENQQN5EQPVkdQ5OmwRTGbfBR7SSjiKakIfU42Z9q
nVFoAeYgl/GMy9FhqBwAdGTQQjfAndR9tFooFfLd5UAcihlHQGo+x4V5JoPpfiLZ/l4aRl3+x8z4
NfcEUTfP5T2m6uOHm/A2riyZ0+Iq/RosObIEB5xudU/ZWMgjFG3yRf95pvqPqb9bwD5Qi3OVfaC1
V5MeCqUwpLmC72Glzk0aMQ4kLnYPjP2x3nluGygcSrheSweesT0+MtoTTQRGBPhB7YFGOBfT+r+g
YnwUn6EQzze3XZOdOaon7TwTD1BM8rDSzQFyYIltof8aU9Fxj/juuVlKdtjCvSVcunrqwWSjfPVZ
xPZ3Qj+D7/POxcCBc1/mKR4aESxZuTXHFhFvE5XCsxwBK8GrZTASukvRNw8KbNOOa1ADx8P6WF3F
lCOUuUek24QZDa3kpu3RneTmky8yABqVwTKhLBZEW+TBGNIzlmmDw4DIMw+/qU12SB++TTvzL3rV
QE3HEl3eE+sUqxi6Dj+U0y8i2aHOzvxy08HI7YHuV81VlX3m3Nm2iGefzfICLiSDydRRl+Q/3cvy
nnVvqRhyGKTzrcLydEHUP+PS/+7KyWl+zOTa9Y74rdyj7U0KJXO8+57bRiunyWoJ3MBtj9VqBb2p
NX3R+N5xwu0NH9boK9kzJKxl6DDoDT+HEzbylHbrIcoqGy7ci95lk9mWLq8WyB+pK6hTfKcRnQSF
w+MBN9EnS+RcbjTrd/pjKmICWyl0d8drQY/iY/D3qeFKw/XR5pO7MZgyIthA4jdXHQN60xmfyfuf
9Ll1tOH+mEnU27MWmLhmg+g75Lil7Kr4H0jh/vFYOYhlEWCZMaN0aERm74XFGg9NxP9K9diZVGQM
8UX8yqCQFN15lITzEHkt/E747X14CxPfSTiiCIxDGa2a7iHWz7tuwe8O6/7yy6JOmRTo9EJt+zc+
NokCRJQx8lVKoMxAp9NFn7M/gGUr+Y6djrbVAmV+9mCGj1GXRfhyE0NHF1nOTEuCGYJ6e6aPhY8H
cxITpYTQeo73409F9+eNr1v5jxODWHRT3KWS30ZHFCbVQBYf/nBvdAp440ONmNpGudStHXH+QLRo
xhepl4xXxN094M5DbSZ7pLrNL49pVwoVY7MV8sGUaPhIFxlMTN0owWpTJiomZt+OKZ0M4pTT/lXU
2JgpSpR7JfNx5nXCW+/0XZQfH8BOqQPRgN/0QCVim2yr+OGZFyvzvktl43SQDW0mgcLqenxLfM0/
Yqj0RH0IPsL19yuJK/VtJ+wawaqtZaM8BNAeO1xTtFWDtwDROoowwOksfbOoF+eGEdCbcvyXPfGF
Lw4l+m6dShLbBzy5CI6Os4bCq52lvsXor/vB9k7g3Ci71gxVlrXdJKr7bYUaSS9lOyVWxpv2aeGm
GEJvWY8viKKWQtdNGKz0e1zGS1lTrBkWU2jkzX2FBBjZqxvvnN9e2sIJCyGLyalpCFir+boUgis/
Foxx3+GdHrm/ahfhcDoyOVwl0f4i/Wg02yDBxS5hQz06oHKREDeYL0zmxYDN/M03XC3QN6UHZ3eZ
qr7GJbqs27JcI+GSOZ/NAZEEfbWZttwipr82tajqRzPEJ6CxaW2TpnZ0DBKLgmzWFzwEK55E/7GR
90PIYFTQsNRbS+bFt4puUKiKwqqJJwIVTo8FtM/8/TFivpzPczX+rzy1eLN76N5CsbeKjMbrM5cC
akxSBbLChkiSpi8OMDYSXAVSbssJmQmBB14IQpTsr+Mt6mMIcjoHUXlPFEUiEla6RTVG+hX4Ah1w
Eh7aFKRLXBMUUg5NvdkKurTsOhCLroR5tSo6pWmlBTfEveE1UKxil8X4+cLMU1Hh12Q5vmzlV/eK
DjrScfkoAX5RPAtx+eYVkEzvnqf4evkstHm2FzygGv7zdBB3DDTSLHa8eKglVzZN0XuLl49nYx6O
Rqb9p6DFm0A4/fKrX250TNWhSI7W9TCJc2Y6IVrhX5oK/MCsyUiWSymZToqA8GnOpVF2QJsvENGM
PmPNKpsM7OUdKq/rRiR9Qz1Ap3D8pJggEThSH+irjzgf0ZhPt+4oxwtV5mB/kKro3vPfvZfBcYKm
4C0vFlozFHBci/rNs8yxWQAWY8nb0oEtgiKVJIkGpHiA44sOSEuODcMEifuILezmJS/izMsXrGhv
QbO9At7fB+XhcSb9W45ARxZUmBJOBSyD2u1mf0yk5Oy269TRGlJizvH9eio6R08dFiVb1JItSyRw
zsGZ140MouhDwMgz5VHvRI1PVS/RsGwEo8HkQ7uID6kgUOaIl37gYHUR2n6weB9e5smoAzGxUBwv
BV7YfdANYhydQbR5/Vm9KNFp28GHrqcKqWQaXMq7Az0Xta7PDKQ22ywI1sQgn5ijOkE2apAEiQ0/
7D6DUQFtVyj07CGMEg8gv+xNlZ+ztZYoplZZy+ROi7ClvsV+T1cfJrqsdOO8/sbANZl8s95FIR9Z
s10L+yy9AbHrGOPhLqF//ntspzXKB/symVMai/hzfbOrQibKM2fIBAm1Xo2RRLZak4GfzUanST8Z
yA1JO5PzZipzawHK06HTKed1PIyEVE8gY5DrYfw31741vayV08ONa+1b+WMHod9eHBOfAVWMilGa
9XUt/Uf5p/1/aE+V9Hm1pnHy4kCdsW9gLRm3iOuHBXAgMHX3ik3hxRu5CRXSY69/HWuq5CMdpudc
d1bVmSi9RfqoXEDs8ugjRmwBMiaTYMXf3CWWvVnEMczs9t4NmVv813gFXCYY1Lsgive9yLc+23zN
ngkhqSV1G5hSe/+qp8Of5jRiLuCzHyqK70XdDqmYfNOUaUXhtQL4qe9E6rao7gtBVYqg8EyCQvKv
FV4nfljhvmDowqQICW6R35aejJN3XiRO449PkuXYvvyXhcddOGnZzbFhwuzOsE2I6yUQd+RkjCTx
7h0t699ir8wgsn1Ah9e9IDyGZf0vvS0+sBO46Tjo2LXqYWOkKK8zkhJ2DIbAcurmYwkXDqEpjX9q
3F025UHTdZfMy3Bza1Wbt68IZTIZD73Js+J+ZaXNY3VKXZyXiogC2ATwnE9c5y+W677E7FTNf5Zu
Ph1V8m8ELzl9QHv3cezn0nUN8hYnM8aqp1SuxgieNCyEg0U9Lp11D+kYOE9Ws3VxLkEI5zOALAmY
zTZdmgTJOPU56LdH6BOHxq/6xIwS3P45XSydq4flLmW9UNbW2yvzFIRxk9wGRXe3LPzAH6b2m1aE
JI1JMbEPwENnAx+vMRnToMIXrnrjSmTkLJTSoQgxlku5UQGQHBZ1/GHDI35lk6TPwNJnkCYvqdIF
qOkZLw2EGmW86MoTaf0w1+JgRpeuAOaJlHH9MJV5K+0tytrUCnym7A/fT9VINSWyduxRB3TYL0xL
SZKZ5NGhwDxOZPTmBQNNm3qD3bxl5euQMUbFG1ayhXHeHTYSpt3sZeVuQrJucKb2N9AxfB+39zUI
JXr8anNF85ilSBiWkxJPl3UPRhXIpx4QPH5u3pgNUJobAgLF6AJ/6vrKw+1qzgvMHD67K5U7EyZc
oGwRyQrvEr6ckmU052JSdzwwKYK15O04rTs52yPktP1MKC9dbxC30+YJxhY2AmeFCnVBnZoDDWGz
SZqVMAVEqGLboYxtq8LGD19w+jT9Odc73/OgrQKz2kmPBqVoPFRlHlDew7aWli2DAoyoWriWFZT/
IxrAouPCA2WrS1KKv1ZKBw6RxWhvd9KNk/S6h6UiYlKkHpaMIyzJQYT0T8SL6Qs6fBdsvda1uzRm
7K4xEkzXLZia/IMTvq68mx+d2j0a4HG4FRNSd0o7KenQWxuz5/W5iJeBsq7QZcJTTfA0+1Wr5XGU
ON1tP29EKf7w1nHMx9EXvFuD2NqxdJgCrG9ylDYAQJwQdCjmgZPDLoJpUko0742o/qUgWpa+8age
KUg0ZynNoZ8Q6zB8ZYQGP9OwkFwR64Iajq9tnO8Jdsymd6l2VK/5YEuTGdDkO5g0fug2acRiOHR8
zgydhqBPLn9iHGHtnljTj7dTVKmQ8caziptXp0zabQcvszSYHZ6CAyt2s+0k3UKKIUJTtic5BRyC
8xWovyYsgPik2AamNwxSNof7xlP7C/gfux4b2nmWMWaHRIYpsmqccY39RvmJzi03pzxu3DuJ1gtV
e5SjoB25PjuM6iLGT4vnrYHmiIIAxuRt7szks8TqXycJQmvy/2mtZZI6YX13BuXeVvNcjXseCnbq
ZSGp4g+8TNbN/CTTCOgJzUqE/la7Y0fw+vo8f3qz9HcL/+lTwwZ7lK/C+6ScACuSUX9wI/F/vhgL
LP5cPvPQjZkL2wPjK8o/VYR4ouAQy9wToR+ajVmNX+OAGRUyH3wA6/J64iQxwnkzMXzSa1sgylPJ
gfWfgGpgc3BzjJ3PS9Z0uvRl6EADvGPbhOc458hxLefPp5mUCWWJS/XDjEC3PL+rHPgj0YTVZyek
vBzg8+VhjkwaMksQgeXH84LBSZdZaIxh+e9dKu+ZVboMWwnS8FQmmqIcjcrpBszc/VDXHeVMt2gW
N6+RLw5nXNIXBpd7o083zT2K+t7usJP/q/51W49RJq6Eip3zGIFODRkwLzxiXF0IwU/135SfeSQO
DBzQxxsWQPfF/7DIrYZIEGX+QTAKwR2Fp3kzZnWSacSksPvSKRZgEpwvyPYi8D4ZmTnqFt/5D7ar
dERtYFtFOcbTL9z4FagiIU3wtlKkGkNAlWgETgU49bs1FOBHaAOuNDFQkqJsDOmVZzmuYCFN6hk/
0CBAniSvYHPZAsXhndBUtnAveTsQ6rZRzUEIZ7S8FQhC5pBHOveF7id/qp+S7WzHCDILDnITniKc
5MlBbhy1jbD7Xed1npvJ5k5t6SLp9ycDfD9ZekaT0AfSsYVjQdrsvYcD7XxxyVrqheCaHKOslnF7
OMdn8wUiynIcbpe0bNwwk8oJ/9fdGEpswL8YcTQnQz6tz7eBx4dYpLZ/aGTSCA3a8eDiBh1fvXgt
X8om2ZKwi4kYFPHcXicogPzG9hSTZqPp0RomJV34QOsRtZrRM5Nob7wiuiPbjZzds5rxp7pHvgQ8
ckWjO2h1Otu1O5aooyGkm940uzv6orV2LXMlse2+JxnM1NumbkZGcqiwF6Eb5QvjjjJx72urnJcv
ndhZjd1Qi0a3bK5egGN2eulFAqn+UqVhmAvBKwu7BNQHGVdzAebZeQepuXVehzpWEkOjfGNmgKdG
yNQn7D+P79r6Kdw1K3CCIh4kklOQ8ZPR79cd4BgZU7M/8JHjG25XuTc3h0uSGPYVKcik65BetS6p
8xYd9mRitirYp3zBG7Q/ihr5vbzZfDConqBWvfam9ePz5lD29eBwHUgNRscWYi+Bd6BlL5vr+vX8
FT4rhLn3luEvqaIFrHtjLuEDNNerGGIpUOCW2SL8X3Nah44sxqtgW385w3tlLPqQSw3Xl3vnhGos
kAmDIg4uL8guT2uONYjVPLblcEJHPRxFezoaqLlqA7z90qTJrG0kf2EFY4fVHRGZMChHoqTeQTEl
2AlP/m1xBdq4HrUSieHIGpubUas8btwvftvxhRZVyKauV6I2P59fg4cFVvEeuqH1o3vvgNlekA/D
MvrDS5kl3YawJTBtS5SNIXJoyTiUQWwysKElhoC+LbE2w/cW/L7SRHOMwl5A88h0NWC97jEE0CTA
Lr1foGTudp+x6VaqOiBr/XzDZIpKz+ogwzbYk930dmIkVus32/aDRy2w9dBSgC4dUT9GFYP6bdZB
z6S8ASjWbTQ7sGaYwx5ZMI+PISRD8CYWl3pCD3WxJ+Mi5YwuV8mbsfJZ/5yfSywSY8YEPUlDTJWP
eTrVq3NhlIzSCiAjFod2yY59A7xbhmb57uv3uxNdhRyVDNgwKcP+QSvH5j5OCUj0OywR/he/LHvm
dp6IF5whBtbIl8SnNJe1EFyvkt8SvhDgyg/rbnvcLZ5BA4KL+zHgDRZXK5uTAGrR620Mw4oy06WN
f9VR0eNKnXjHCh03n6DFqUNxOTuANAAkdHDYRSwUtwx9TDDU3s/X8/VYPLZLVe22GCnS+9fHjFgz
oaa0o5Uw4xbHJytB+YWM0bC7oJFyFDj8/c0ujyUmLeRjFvSkdguBjhLWspNUs8Ndyuir0FE9Zb6I
5nGXMDa1YHY4JXK5S8YdzAVVbvtQ7wH4bTpYdsXPqmhEypXELiRM4qUphzYdTSbXB2hHIRo117Ca
5Vjlvl0CMFBT7IPLAWSYJmMK+yqEtUStio1eTDhQNSj3mGE+54O36wfBxZhGvACVyQomZ1TI4J6O
Np5bUTBIru5WhNccfi50Muf+35czlnbmUTRTVmyI4Wa1OtUFXlaZOAi0Y81LuVTlmvdw0Gu9V2V6
U5L3pE++v8nc8TKuz8jbTQI+GQTxFaX48J89pJiRsYc37FNw12EmfvK9DG7wrjtERMJVYUqunjLJ
rEvhcOgBwOiNwj0h4p9G5SxjcytcwnrW60cTvZhnVu7W5V1htzzCJ4coN46TbPbyAUswIau1rMEv
0eMgVD2/m4ER8i9HzKriDdC2815EM+1L7aKmWD0H8OEgAVthPvF5GcxspQ3cc+pLEty+wcUFfhW2
APi1xkoRYh3gQyaDE0aw0iT+YrvikfYFV1Z5tVF/dAFLmmaySsUE3mQwOovYuDMM853323P2peNN
S1pnvGbEb3iWb4qMGFIoy4PD8td+k4+H0i5KVPSscUHVpte+W2IewXyqf72RVWKGQOM9wVurOnjX
05vtVQBfVempMK0Ro2gcW0g9ot3ygms2NroXpmvYO87iMOPdEIYYroSjUouJN9nHWdTXR2TyyKKr
7VChosDLMJFzrOxPvSc1zZ6N9OTtQkdsDnTvUe5g0usd8Dqx/3K8DmxgEEHVyovyt0G/G5VdPiHx
COQpVIDOj9p0OoBXqhDOz815KyG7Rauzj9OAVTHXdVD8pnGR+/QYCXQPWJfwPg8T4PFx3MRQwOQc
y1hy2VxDXU80e139wTBEWBi69pvxOCOG6rCU27HjKIcro0w9/R/cpmS0LhcOGb6hP9fAQQMtiPMP
YrjIfjSxcy7jLbDAREEjpBoMbuKxHHGlW5t5wjQDy45aREQUQHAjJijuabYOeqLKhF9Hft4CcNf7
VzINyRcbkBRaTQLX/PMdE/JIKQqMu8fgn+Y1EI0PV5+oyl9pZz8jxbfTfbSeb9C1RniJsood8acp
g95GG3Q+5Dux9nBwTXS6I5ZCVkZuyKFh8TAmMu+Iz59vChO9PfQ8aYHZuGC3GQPid+w1DLSN/eGX
iHddnyxsLw3PWeZ0Ds3YeCxIXYuGxUhCSX4IEuRI2+K+78Rk8AlnBBQdiyz+2I2PRYbmst8MZm1j
V1tfCbgHdRtv9LbMdwAWHOltayWlk/7pZfy75Tdkb3fDc55chtalG/jvbeKxmkFTAGrzvzvAh/wD
w+ZJX6WMA9bTlPvHbRh2nKvSPqE32iIvhyaaYJHbCbt/kXjq+/XXfAQ8svI0ZWvQOEbA9IU9aal/
jXg+XxZFM4HpZWvCeqJd4Dx7IRBR/xT1LXXlmcqitPccC3KQ0WC14zJ3LwB7dfI9lFOYLHLo3U28
aFO7s9Eg1PaGxtX4EHV1M1E22JdDulMpfhk40ROyAFWY/FNRl1iOL2+Eaumey81Pj3XDXE4Ihqon
jNSt3K8CTKi9grYYv2jTWQnSe58LNT+rq3/qnZqsdFXzoLleBoY/ZvCAO+YO8MOhInegbi150b6r
qtQPXVszaU+YiSVuuyXwRsRT3YbNXhk9gLdNG37us3MmXfWOLART/39Rwun2uchYN0pHM2Qdo8jv
B7MrDpiQd1fazjmetD8mIFhIAcGsepouE/w5kNPWnucVe1d2AOy66StHv27rIWFdUeFNCdGJUKEX
FtN9UgSmym5dDIvc/wTmhqucroUUyWtNuBwZbIc+YSnGFByIVVk4roH+n2qkUHQ0NHivkSsgTfCC
GBpXPVQuEGUpL0VkEaujZxYs2ktNsqmcvGkp4NgRdjahABHRWKSnBEscJwtQyRK6xcH0NJj2Xa74
/fSZFF7KZ/g94siUNboiTI8229WdVmq17m41Aoa13vGp23hEnMg0TgvjzbPX+sKQoF2WVj+fInIS
buvzz3fxDM4Tzg0JaV2FUj1glGKvLglxwiWtIJUEHKavnZaiKYBMIVWs9A1xrDSzURxQ00fhTY7E
XsT53fJGVipJqHiZ69husA+rUSG+w+OH1SC5gQlQULJ0PCKJlZsyAInuYVnGFkIXs2ZeHR4V71B7
+nVY/9T3QkrTHOX+tIf90on+2EjtOtwr5JAiuG7aTo1qqKsZQVDqiLmcI6EZLWlE+UhCHrMXxeVu
Nz+itoQc/p7rbr+lIIS1bPu4jwy0nfPmQ75PH8v4MLg8qgvHn8FwsJVHB7Ywcg+/JIRJu6Bu+UyS
IkjHhENPDiC9K1LKHsLrtkgXvmiok57CXuy21ZFjzQQJCb3kp9OkGs61Rjqwx3fwC0OGLIl7oI6W
6WJBc1BiPZENsgZw6TxxaCKSTqC+Sin8EiZ+nAOwgaZAYqfnVcmc5YwTc4j3vFpWPE54COXoLI3k
gYWzS+x8ZsyetnctrPs+RWUnGpnca2AgMrvD98t4pPfVpmE88q/roDC9D0GWPIvxknsULExwsl9y
je0knmxy/SUkTz2FDRPPB24+7oVjarWxS1vaaqQnci8eooMPtM3WL/OQ88USrMRZNijrMxFSpz6p
QL9yzJKXEydIdsvfb9hI8F9KDKVsJeIqmzPzW90ng198JUOnPQh9jr5NqxvPjuWKewC/wo0ZhXTj
ChuSgRCVvi9+kUwhUkvUOhUr+jsig10MqoFn37q410EYa5avVJT2dSu0wHYDJsGOcQ4NiKPejycD
uLLS5/iRU6TQN0uHgxK2i44KBe+EPBJvgtxvcZk5ayeXmiBVsxI4u03TN5e6Ke0cGweOo52TILHv
DGBPyo5P69NR4S9FEImVtQnf6t+XbB3YzQZVrrxUpmzzrzT81SkgvJJrgaiUYrDfOA15kZnEm69e
NM744xNl5fPRNNNt0hCQKb54kxyf4BV2nsAwqsKwJ3yTzIoQuh9ZAoPwZlsYgyNwzW23kjBdY/HT
z8YsQXAhC7Gjw3vHjYNoiOv/qfYHj8wXQLB4ZcwLyQOF4d67xDuMm1jbUgqJsjV8/sZ70eCoFApp
/7nzhiPwPOFoTzyPwzha+7ZnqT0Y9y2Y4q0tETp0cuB7I73bhL3/pDYQeWiTN0XOEdb4rKHoRqav
3IqU/Scuj46uXhT7d2p3bhS2RX2H+QvHsuFBLinqquQqw0XOw28RSbpQmnTf/mU6y/BjJtn8sV9K
fR2e/1Z0ckwYi0pwYE2Uqt+SbfFNsCa4y8/br25L+rbB86m6eH/kHe+8/PIaF5qz5YHMLbjwdl5+
IXhClbSF41PNd4zoGMudmSp9KhWPYI03F55oz2eJm2IheidjzJO5chd5Fj0exg75oTq0y1rAfHUm
07imI8/ihQQiqK80V9vcOvYZe+xZp8EJxTw4ewug13TVtoGCynDtmaZ5C8i0CbU5jk97PVXgtmyv
myeFp2HIP1z9oi4z2jOsBTISMaCs5zBRAQZRNKGK7i/v9mP0g08AOuHbcMEInCtGgDM6vsoHcdrp
Y8tzb0kS/Rz4l4F46hOOn1KZIFrYuLkvmPNWvIMtlJwTOIXKX8vwN9Q22pn/LoYhTMhAvjw5AFV5
0cZwY4gpRGRP6FbwLWpSRbGLiEsEQ/tvr2Vlo0oDEcyaKIfje1WHHkqaTQW953yOriMbgxVyrHqb
IJwAdX5EIc926YGJe7NP9rIu8Q5h2hx1NN2dYSPfuWXaIEwv2bcNrnX6u7pSMS6DZcPtBsoqkWHn
pVc2kkLsjPKR63AH65rU7ODtl/jRZ/Fgqq7wdl5XwHXwyKJpvTip8+jWsH8y4zZCdzQTGr0PiyYR
WR+DbGmF6RNDmOBXHVseGBH8/4C8wh5iwRlmg+Gbai3rfi7/N0Jxequ3T7fUB1W13/eWlsjrWSuB
bKCC9ya/eEf9/txfTYyie77Y9KtBq1j6bsq7LwtPSz1eLTJu1P4sLzJy7mJxE0qdMJUCS4ScEO+E
niUHl5dU4mZVAZEBrcTfH/CqOM8XVI+H9ATgG2vkcPcuMpnROtMLnxSmmzdIudR5HNQrivDzo825
2J9LdK0lCFYa6kWf7CyRjgJQsnSxXWbr92yKLiaSGh3MnrjBz43X6FHJktOd5ouGMUjZWy67wiiJ
9PCV3/Jsewd3cwvldUfkUsufq95BSo8nkPgnyQijhxjWMS0qAC2cEDMLlcE372HiYgJT3/JPCkTf
73jbbEeOUsJOCEcn1kywvjdhsXdRrvOzYlVBVCZN7VdWgsA3+a1ggPKl8D4QV8gzQWC4BJYNhMp4
cW/F2kLORjVt2c3vH8dCkdvgSRYZGjTV5OvyoBCcJcv4QvZ2hmbDxeEFA64ZgZ6K5OKJmnyIfb2m
snfWSulmrTE9/MetPKW0dVbqH/qZhURva5mWemj9C33E+yWBvRWXj3Wn+G+necrCy456dFyqKIkI
vqeKy29bGuclluZ0aIG5E4YXiHaEv1XbNn3OUQgNtjWwJMbeQiWHMfVqKQiTXt7O13eo3kJXSECb
OdNkK5cKK6oITcW0dGeSVQ7eBh0O81hUVXamVGu9CumU9wGnxBdkkXtl3Bv/YLYsY669gTQ4MuOz
6uynv55FmCn51ex3rRnpwd7F+Ty4wJQMNSnGuEwPdKUx77WGeqDKKDVgOkgAwi8K7f+oOGs4OtkR
60yAIEUf78N/H+CqNju3M0HGEJFlRubrzujEBXAZpcIQ5MhvwqwcRT78Wef/H3IDyI3kt0chqWJt
l4omPvAdG6mxHc93nJLZ4Ycmxccg5T6opwrTAb40KEKwOFDtvBMb38S08T7g8OLuZFJbZUCmkocD
dD/HEHj2kXp1bazLSJ4g/M3xcILiMYW63yht8CpVTaxIuvPeIK4vjC+v204ltkS5NsFl88Rz0EHB
k/UQNmoynxliLIybi1spDAjbaZ8B/YB1oJUAGRQ5EdEKLgDiS1ApaP2HNrmpF9zMfilPnV083feZ
ST2ISVatVHanLHksHWaRzEFfrsx0CINOIFqrjINW8Rsj4ejYwpWX8O8EQ19a6CoFf28ynW9l6egR
XLb67PCu0lS0Kwy+Y3ndSy0MoPZBBOhs+asToH7x82u8J58cbyx7tnQlp5CHs1W7U5TK912u9Ofp
gVQY+SR3+Tucu2wVworSXXyotOy8dQd1gsj1K+pxovCf0ANrvegxl3HrGnNFQ8wpfqhovaGy9Jmb
Fi9+YH7vOHajCvinG9Hf+4fQnCoSiZvJaur4+sqd9tTb3ual2+9H9igrCzKYx/73MUmjbfWVAQDJ
hJ0vy2y7MBVy2LCtEHlLtu8xp2DVvrw8etHbKEmjUmJFTB4lOyZ3dQFARVsHcs3Hv57bs4g794Yr
kRkjLHu1WLCJI49hIF5P+ScisHC67JAvg17DTCNHmIhT5y27wi1eYEKFiZYMM02hZ9ybqtsvfV5S
uFcgXw60mdHkX7Qainz6+cUhvZpdqOfvIW5tfYZKPgEC/Zp4bBHC1wnNGUjpEr/BPUtVfbXW0fKz
N7apyx8QQy4NlzhvN6PfL7gPhPqychVi9tP5XIMT3VBWOa/uqf5Gk/FPdNWN3G/bUt9ElVeuMoVd
k7Qh2rZxf/ypufBUvjsG7BjYCrMg0Kaar+d8urLpGJ8xhpl9LJMVu5oHUMxrKzvDbGwdJH2RpSBR
w4yxewHd8RPTKd0LrndaN+idLlfbe6tqBb8Oo7YUZixUu26ZshG3hBp2//OlViiwX1czGLqpRUqJ
WddJ6SLeYdXhNM4JLwq9b247pJ3dYUfp0hbxmsA1lJPiuXGz2xH65czu8JwiMkoFyjtFZEVIpsq0
faB3zR4kPlwy9h+mA3YOsBKrMylmtv7w7g5wwnk64uq0+d5nv/NKNFYnfhpZf3lErXkvbzcdI7l9
SUwU2S73hFrdjdg1aSvlXADvldiBz6GbVWw/CTYijyt0MvUPQJjHY/OHzJozuIR4U48UdpmxJCdA
v01LbuyzYXVy4OfDLoJn+yhudQ1BXu9x9K33Omh988ZwRT89ln46Y47K4KoR8gQ3Sc9Y7S0eHTtR
Y3+2Cg+JFtD8PyFeDcxiY+H+EJBDtlO//rcRCDKiAdsBMDUxVB5v52KwOXKDL9MWKqfdveb80WrJ
FYCf0pMFerCIVNilo59hIw1sKQ/NoFBp+VgGUMh5KWNyL+ylNjk6G/ikAcQM+hDSnDhFDWOlnQ7o
ilXs1EKEbsOxm4/dsFUO2CfX8S/datwCoTQNS0vHUpsRWnh7qHD83wU7IvanPqsk88h0AI50cnBz
P6Gf9twa2qC+QeVDcQEzUrvaDeYMuIt5ABTNT6DcJIh6nltNJulcSjICX+3HWuqdjX37EHXfssF1
hDnPrxPD4M8WP/njwzfzZSVka+eZpttZu8k97TYW5uGsIBvRnN6uuNQuODx+fJ678wquQaPumHh7
jOyD+xzRAjKej9/g0KCJXveXK8ZyGT8+4/BvIgyTcujtuFmlN2Rpakx3YkAPgUg6Gp/iiUaqtRik
Bxrnyu7zAnjpc8oZ7cX+v00pJLF1AKlTdbG1KN4C3no8y7b6kR60TPDLJZsdUhx7+cU6+kELWD39
AOITjoUcUirUZCftasIKCC0pePVafm7qiMKcfDI6VkeP9mk3fVseeqdQU+GB8ArfJ72v9ZuASsXP
Wmquh19tdfvjaruIdbk5UQP3nGHI6BwhwHoEZDD+47DuHRGywbLRKgpHM2Q+lOdYCT1htEUrPCUx
IE0wCjGxHfc0l6HB6Z/IbpI/PrTZbOeWCdeCZI7YuNqR7Uxo3yUegfwMhUKiQgL7MgYiH9hKA7RU
KiOydV9/07PH1PYotf+UNq2wDY5+XkePmTntvjDMmm4rw9UooUsJvyDdgx3mECRbv9BW4Zkgthei
7SsQKi1TtYWlqik6FhLFMKEGFwlbD6cppoDn3tA5C2+OaDRIaKLAwpOfg+gnyORwkoY3PMoevMHA
04s46f7gahpP+Rl9Vy84JCavchihadWNQjlzrj+cDNhTCoNB2UZ6oPzHN0GNjcVcM8Mp8FGoTD8S
Ad9whC7id3WQ0NlydofS6FxkSzdcvVFaa++BJtH/iYWMVXrEUjpSsUl297cLDk9+Ngxv9qottQQb
Tozd+GCRPhgvkzJQimjDpmZ18mBHUUrrW67dRTZcsBkdeCdz4Xy3BvkohdzkXyooDsSUQTylisF5
7GOU/rc99z3K3jvfRhzwUlZ9vSA7mC23keXanimM864AzeTciAJJXs5w3LFpHCMnFxL0z1JzvmNK
XmqvQu0FrMFT+vVOLiI59olWB83WUkxag2/svb3JZTfBPtAuBwF2ZxXiGBcK0mmOljtBczb6B/rT
40U3QYToUpmYwyrVCSutE0s+tlawHIfslF8IxI/7l8j8NMAQnZV+RqY4gBVvdWgnpjNbpZPd/mpK
uAn/ksKDJZIY05pTLSpuDbdlELAKSH5YMNJ5zB6FA4RS77TUfDpnsVO6tY+e0KX2QPOScwDmCi3R
BTGRqR9P/C3uF4qVJrTf+UKi6WNpladeBWSBHzhMUd0XI7Gkl1C7oa34afYPJZB2xPGhsIWlf42P
aA8PTRZR1+9eXuagfH+zVlB9+TO0DXuK3VeQO3BbFAa5JyM/+twxIgYTiWv/5Eyg1aWia41PiXHI
gGljGQSsRKXMcBJbW5DzQNxMc1po0kz7qJvX/aQKZdm78V0RAI0KzDd+O6ps7DUu+fCjAjThA+27
PVmu21QDv1rFvSXmasKo9e9A4aOYFsNe31ioJW3TsmrIMoI4p+qRlDbJaHmtjnRoD/qAWYZdidpN
MM5QX6m76SeIaxTUcBh2/5TuaRiMOqbU+XsE3XKqu2OSj+sVImcT2w8NYLJ+e9xg3H9bRmzjjFy4
QJlvQ1kybTnuiLVtCtDAaVxSbiZvXzmKP9CLAe5YOJ2bzCM1dEE+5396/VxNTomNHT2OK2wyOJzY
xh1jkieF9c4FAVgUS59NhVj/rvN9BJDJTY8g5jlalRIvbiDEk4lqhfMU4YZjASYMNw+I+YXVJ4U1
NoC0LE/WKffp2+DcQzTinBNkUUyRDGRDN8CBoLPd9pf/ikDBsjByHqr4mzDzFbecPXLtblzCslnj
NVTckACpjmKUeSQJ6i7Nm0EVYkcZyTOglav7OeuYGkVdpIwpAVlydt0IzMmq1NRaqOrZbanDCMXx
hWtiK/TekT8kV9bHdB8Z0Wc9J7pXjat/7H094JuiXWNuYnaxMHHoRot8mFooM9+y9gXduQAAkrRp
nbmIxmXhKT1nPr7/cVJXtqChfO2ZRO2EjCEn9vQxIKn5q+qzZRnTAFnuuHQJch8APFOYMdfIoMGd
QjwVEbcKl1wx8KpSxEH870IDVsd7/ZQBi9uQFpkQyJxgk6tdLHhTIRlB0csd6gaTn3oyQMEP3SgH
IBbnP0G0yIzCWjehgkFRl5KyieLBvnY4kic6xzePvUXWzoAEQxwqRADGLGJ23oVRVtICVxjz3iZ+
9zU0vJtZQrVwyoMb7Zwt0W52k1kaz/boID2wK5JWvM6TL6Vf9PG8q8pLNnOCr6PAVu3kOWalMCuh
puZrIQ5h3xpUvJuIzTg3woE07D2RdyrAQKfcY1r1o1WM7/Fwa9gyesIpzHawok/q5MeZmFmuy7J5
015bMqpw+MAhFMohvetCSWHvqnnvWc4H2Z1KkI+9XJhmOYEW5dqxIjEkfSDJWjG5qz5eAI8GPINY
T7fpTl/i3ODGcy2n9epQ83aHBpvJfVeYWDmTsa59xuIhVi/iFdqXUPtYVie72tSFrMTNw9P7L0yQ
h4FZ6avoxDUdyOzxjcIdSAXVxcIa1WmkC6RGdUyyNPSwi804rJfl4WVZBruIhwteQDQduS0836rk
gjlKrqL9cW7mzJYbZ/r9KHAra9uWBmpUoQXwbRT2Vz1TiALAlZhwkJ2RrVXz/uHCgyD9SWcp0MfN
pGXVdYOGiY+mNPlDhchJbXLgmiQFJpvFe98mjRqSxgfEKK9bnBTrnD4ImTPGfsaF8hD34RxK+sqc
CuNDRR488D5Yt8VlHQooDmKsl8YI90VmhXdJFHDeIf8lIdP+xyOWzN2E3ItfJkGGGvzfxlRWZ3mG
rsvMKhbDigRICweHNiNkvxpuv3QWUOiT7R9kaIw+pdcmPbRoqjwdQYDQC8echqCVJPsL98vSgR8g
67KgSMfb9EGo7XjX1Z52WVdH3DTnQUCSUiIo7iaina4fmipoe4vaRGxDwAhtl+8vzsSjbq6atS4k
njqgqgmgHMIVJCMjRFuxV7k/zpTcRUBRWxzjPZvAJvuzuHdSuHmch99yJkBVuQ==
`pragma protect end_protected
