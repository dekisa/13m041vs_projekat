// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
sM959vEvMV+z+qaLA4AKPv6BifgpavZQsUC7xZQ0NI0gcLvXGl7WDAZPBZCsrIXb+KT4cDggHw3X
mnbVaQxDkSGySU9P0NI54eIXDj6x4S0P7+5rcEOQP+cIrpvuhgCr/MxMxwoXpUqB818z6wAr5LY9
h/JbeWYRBnNfuanDWcfK33UooN+X5yUNteFj2l+5syAq8kf4OeNzdX/8uklT5WGPVcPoiLTfTIZc
+ETi3YonjO9FwlQia2lNS4KCoCxTi0ULFBkA1ggaDrOK3Ey4CZrk4Mq9bzaGBQ5hY8cHYZSBzRuf
GZDJoFZY82dBfhoFdJaUaYyp1UfVQIP7SyH0NQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 34048)
VV0XGr3QJPMgfPp5nnyZgZye6B5RfkMbQAHIQEHgUP9SsMdwm2hVFp0LGA2j/DVfs93bQdk0y0wD
8ln4q2moIbSuGdyognVuHHDl4vL2FCLzy323aJQP5/hWeCmlvIKyDOguN5jTBJlwqJ4cg6VrRHIh
8DtFZpFigINvMh+JxfsUl22gR03HBRlTspG9ucDA1y2bA69NgJDi/hoizuFvozsBLwpAnF39Yit3
KheTeKCIR0XHluVW86kFx2or+avsCC4OJWwDJD3rS0zBmtS7/XtwbWFH9OG2eNU7FmY9b6rqhRg6
Qk1nEoeqnuYsv+NvzfQ4mFAtbvBlzMNxRqw1M//xj9jMCZnwHjWgIFBO0iBVrA9DI1PTOt7Q9yU2
b2qGcDupay8IypgDEzgjJIzNshpfOSnhsF1a819oVzCeACYUTdnA6nCSv/CXCuxrEgKxZktUSpP9
eaDthGxVHalsItU7OBFFXNbRxS8D+aFViNW3ueZNsgewDcA+FosCaf+xcwGiOzB+w5TtthGAKqXB
+YDeq+l+ZcmoEoaF87f70vjsuEcHp41Z5+CmyhUDfR3XGlfTzQKX2VicXLEiXc8EB5AbcgtHLSVf
wMGnfKYVT9lkpw2gViZK3C738n3Ba8+RuXBJgS6Nud0iVJWZ+F4t44ABj9L6yI1E+lVc8J7h5IJq
0OWXaunwdMkGarAJ5k7Dr4RrDwmbO6HWiSrJ8Hh31yqXQkbTaEfoEDhrq5D94Rv+Q5usul/rxgq8
DhNrRdQt0FHjRhQMe+ujuZWyLM227W0bZi5EFzyQu3qnocWOCpMce6qYOr9dxfrOy7DEEiOzmsFR
o6t1fSB/Lb5PKUMOpRCEB25JcVpeVlaGv+S7mUCGNRsLQiaeoGt4/PmEhvJy+ZIs2XgeslCY+tzp
kmMg4Jbl6VzySPggHKowehBHOXfQvWhJ5aIH5VXDdHvZST0zEgFUVb6P5a/zXplwuN4Nj3bTm9aE
yuwHpz/q8Ty3fEiEjIJOv2dRXaWpuwIyhyUStpCMmlEsPQ75ujGWriM4FKWghy+1h0sCPY5uVF/p
V+30pb41tgmv7fSBG7w46u9oNy1SYPC/o+lscxjJhruu+Q21yqeyWa4UZ5xdVWEwGg2zYPs2fSDF
xedR8ixLdXUGXPWHbBawiKVQI38LjMifT+hqS1WIexKM1N73wi/aTcjkr17PtIWpFVpgf4bjiY89
MAtoHZCyBzKuXcorePE/Wh02yGW9swiyriU8yoY+skYsfJHGHRt7NiIxqfD9QaMUb7jkmE+mDWbP
cATePAzKxHGJT880NQI2Avnl+LqDV0oMp5y3jzWQdSvoY9CogImn70yfyujHL5Y9DmU8AiJw1kvp
Wod2mvEphuchsARD0nfjnkWpnhcZ+A8GKRvpOPNPfFUcIHFqr4JuCvV7PZV5D7idHqMnaL5yOwO+
lPQfBBSJZ8iLgbiRXZfgmDoClMbirnxZHdfPQ1TEPdjPDO7G5gm5/ovVRA8U0ib6CXbFqy6qMmNp
tILGwWmSwYwFeaGMJM+t2klbRu6o0IbXotmSh0CguK+NSN5s3o0pEhld8KXhEkg6ZHdIHjlDbDrU
djgmfnTvAyv9wkFPATMz9EAK2EwTLDS5F6PdKwGr2nPuQBebR9uQWcadPyCeqoJwkYsjDHaWhMBx
h55bV9xwZKfwCgxpSJmO8xms3GHYAP9PmhdAWg2YWE67AUKPYLFgEtNoP9LRGX2RNfpjKE9e9Bvh
98FNB+EY+3UHC47uMn0/+2nqGDh8O2Q3LAuXfCD4LKMyrgUeQ/7k9B7vFGAclxlm5ysRv3mFaqsy
3v+txOfM+Qpl6tZANGqYrVOmtRit8DIIrUo+hlToIxIJn6RnCQefmZzvK6zEY51BuA5oZ2pVFHFS
OxXxSjQc7nW+S1Yyfext272U90PYflDb/3XA2+PTSnyYbxRRH+ZIef15PcpPqPrq6MCrIcbFA/rf
DGFQG/cxyziLL01KOJgj8mA0VPqUfSPS++lMYmIRFVf+6slg/N5IrL+wwmJm7MfrELte7cov5DDv
ubVkwElYIIDoIG+CrPplJAHdeaUtdwstcylHYJxPhdda8oZjTsg8NBeMIHJF7KIqHd41zFErhvAc
rROydjKdpvXYhdx/EzjZy2rdlhx6i3rCmAMiXxck45Ti+L/Qvyg4w9mMU8Xg4uOwTlpQPFLm6+WJ
M1uD0aj/K0FkK8RO3gI+empOGnQOjPesrPbSX3yXtpZ5BAjGxzetSEh8w6Pq4OWtxBGo2LbhAuKs
lC6kKkxY73WrmS5Jm9OwBrnMyURZQWq70qxnhsJnbGtUKZUB9rF26N/TNXsJTx2VFfmtb4vP+1+y
07a1oOCKJioxEwVuzMKF+Nj651R/se2jgW1YmbXBJsWf+6AKSMLLe1YmamycRvrR53KwSRf2MCy/
0L3Z5P+ejtxTwAbwtnmZJDghOovA84p/yi2Js4D7SfAwaBJqx8G6uQuFXqRZxfRRiNtfk5+Y6LRS
dT2ecKq7rZuLkQfOBdT4YVN4uieqJcF40vzKyXS8fFTmhGUu32hIoQ5RakqZH8RsOVv76QumPweD
p8MhIP9QkjaVKaK5BTIozN0ztctS4n++862sPz8Y0YJ4+IV7TYKp/+R6m+O6PD5jUZQuPvWdWxp4
/GpUnLy+yMOTtBM2MUkwpSUhYVf6V87op/e6yUSMZgz51SnzaySIYCFbnMwmd5jgB1Dce7MmDAGQ
8Fbmw/ntAslY3Qyuiaa5HvqUOq3tPvyBTY0ZRR5Zm0kQF5ZIUdV07voxJtjgeA4YMVYXYm/08JaS
s0JdcU2SCzu5vplnfSSeYe92+y0OUSR7W0mgu6sjgLcuEMGgIeokZXlm9tjhx6ElwYMWsLJSF7Mv
72RyBM+vuw/HhuTIg4r6PQMveS49Rla3EDqtPb9Cu0kt3XmJ2B9uGtDGfoiV0uQilza/A8qy+z0F
MY25jj27cWlRd7fZ125tyymgvq9Ea6n7NFwShPPz5HPDu72bnFunUnV9A0kv4rnDH64uA2T/kcoh
4pbip08POjFkmAtaygeb3G+q9qaGk/AGg9khxCS6JHItn8VlN2oPKK4lUb9LRmNxgaR4D9HI9SRo
xLZ2F7WdyA9K/b3OTpEuXfbRatImPAlgt9lGn6c7twWFaGYYmdPTeLVraOp9cLof9I6oS9O5c+XU
p3FMPxVHZ5UncTDuYC6z9UcMjmQH43Q0RvYIWRy6aQexawCMNLDEZIPhsfuhX+K7BA5F1A2l41na
lO7E28f6B/rl86/eF4UAsxFHQssljlw1i9ummU7a4tPi+VX7yZPAiUxzUh4wHRF4Eh9BSXLSBIRp
MHqlbE4Hgm3iNTPSJOwOqcSK741idaW+y7M9RBroNJfw+szeEmdfK3hLLbcXiL3xbedwgCyGm0Ow
0Tj6jkEw6GZkSSebhhSc/f5XAye8j4+Qfm8wyPJkpi/9FYkbTNR54LASDDgvfrC3iwLpDTRgAwBQ
g9RmZh598jIJ7CgS+HFsKevafIlh5bOCEOTuLMQpYo/LPogjLCGklLb8zgkF5bf+/Btn57RXpRoj
/Mna/8Xo1exOxpuJqHvGEdbRjCS9miCeQN4qxEV5HOCZGylnuOFaOJFTll6MDL29WBDAo1Si1R3m
HFw8qmzCpNgEV6I70tT4su/6hmc0PjUWWxxHMUMfLhB1SjQc9nCJWVEMuZD9Z+/pFo/h7ZAtkKpg
WXDi9Uh22rE7pOxykfBGgdBRIGk5zuGZ2zKpPEttU9M46Ei10pPjCUYLNYPT2JubowgePJcfM53W
3flHPx9FS3kdgvEquSRDkw67it+hBATYPlua+AMW/R9xKg/D0eVDOxZ3hEHcXcrXIEpCTBRFQBIN
zUY/pHVZ0MMKqy667NKycoK18qu3URIcWlkRboPrUmpkOL8y4pGC/aX9VWDG3SeTJuJGfsnskyDR
liR0q4KxUjHjtL9NOJmZ5JHKDhwIzIXdr2y2576lzjXSNEhkGC6eOUQaLs2kavjfT4Qc+Qm0uBrP
TCdkKF3CIPcVE9TUQF5h1MCOGZGlv02glXTuGOA/TokHNv/N4iC/oY5m1jlNmEzvUfHq0JC+NlcE
diUxpnj6rYx9n/fF8DOhFp9zLTbxSKj7fxvT9Hb/Qgon6k2Gcw+pFO/pVcvhhMR29JQhn8SXeFCX
emTZ/r0uqbJLBOgJ9NaTrgMD+aqX4qAWvI/C7uNpSeaYrY5ZJommTGFNffThEW3LipUmvKSiW5nR
GuYa1dztEgW3LMIQ4wcrst3YrSxb2+yYhBZjR7RyJnjpxULqfuFtopJZLPfoYOb21CnnW1q+vL6q
BKhZUub6o172WW+w4+Q3V1iEki+sZgF8KYG6NKWU85Fec+zQa4izB+IPe783j+MUIrkegB5B6Pjx
5zn6ra6AknhBUYQJjYRjwZZZE1bdse8esteagDlDSA4ib6MWPlJpk8jsG3J6CxEPR2eZf3blXaSj
nJVQzw6Tr/suMd5byTO09nqgNVpXiAkaIBHVJ4Uoe1yxJ+6TgooWTryB85E6f3prr9dyQd/mSHhs
nEYnmWC/ZyIor8Pkpmb8VxWVkz0sbwkK/03HJ3yznJTBl8Y5NC3eSB9AkGqLEedljBiynUUnT1vf
wAs5cFwBIapLeVM5pv6cIRKb254ogQrEEDemxB4zPT5xGDKUYtrn/eyks1b+m/rZc0GmP2fuZr/F
x2fgcttFN0RYS1+z1tYMDmptr0QgiTlc3yiTBAf48uAFFTDzaT8DBi5/6VlNWVwrB3Lhda7hP5Kc
/tdcbUNu63DHms7SUZ4Eefn/SdSMvHFfORCGuWuiNdqxv9WlxtM1MQFopLO0P6Fb5/IDf885JGlC
y+UFU2qasI9YBGOdRSyvNRVATD7z859/q+8qBSYxNxLGqpdSaVBe33Jx/LxcSTSVVFfn0hxOPoPu
UgJ0fasrdXpUs+rZDvCoRYkNVbat4Cz7VOzCsPJIiSvHhD3rVT4LLZzBW+J5X87m6pffA00ey2YA
o5mI7mK12kPJB/AMQCxU9F2GzRy/04pQBPTnczdt87Vc05mFa0Avkap4IrxPBMO3sqxXmALsN0WY
eajGueIQ54QXlcje2/MuCZbcyXe0mhU/GRB/cR27vzqFkOTucseDqbi70d7CU0Acg28t7BBvqDNe
V6Is8hA5Cz9BYiUakrLBCUKcERZv4jniyWCb/L1jYmScrw1SQaplS+BqILkuKjDaWCb4TzkSk481
VvRdze0Gu3cjEKrN66f6OCtkV1F08jFakF05sEeCewd0vhH8TISZtULMR4nwdSMGAkM930TbwqDO
zqjxwwfZSzxP9Zzo+0ETrfQGpGacFRiiOO2/F6Lyh43tqrgZFQGpqHwBuYc5nRLZHZwa6aSBaH0u
LGMBTsdvXG0ECTQy620IcgZH8PsDp9ynznhx8vKHAjdEjcOVBUVanxUcaXDeFrtgz2pEOop2JxKZ
D+aYnKQ1VtAh+jEuV6GWfkH8TkqVnU7Y/YxBy3+ncYUY3FOjJdhFTyWVtaLgmoK7ZEpNdEaymedC
pW5IXwuymhHF74c4I1KuWliznL5jTyxlB/MgpYkv5uARXtlgI+JBhCVxDY8cmzMhG/kI/8DkNDDv
ZhEJvdGnIPyjH/4PT05u48vocGiV6hlyRg8fy5TlQQuw/iQK4pljisw707qvHgne2vulYsSmW7UD
CvdE887glGDb9HsovrKgZwauogoC5jPJSbKMRQ2yBJxai21SQ+1fr2CRs5APEVtD6Ts1VpxYd3GR
mmlL81xRlxqZbGSiNICgSXN6shB9AyaXiBre/bFwBJlPqqPNp4tkI5YFGyUdgb4/glZiRu8t26iK
d4JC5km8q9dTnnloDimk0jRftqLd6XcHJC7+mUktiYAfT2XUfAKyazQQoHIiOmyDCyCI2nQxa85A
Tc0SUvdxzGnaXtjV/7rOkW7Jscc+/7ljtnQg1Gop6GEiys1rb/IXkSE7DxTfYM2t+YhHD8BKGAtv
KEv+U9o3oAkWM588uKaILDxIsC/C0+kj1xim4rWtFSigIik7EbumGw4/9npV8VtU0Up40ajPnAq3
fyqmAA21AxV7nS4EHusX8ijI4hNBEgghkMuPHfvYca6o0c3bgvHwwvEh+Wwr4voVQHdKqLHZ8gze
b/BYRH2dW3iypUyHSUM4JdhXmAa6O6lzWEPMsd/kTU2Il/Y+aCIMIO4bPv2sqaYTUautILftUkN2
9inWYdiwDj+BPY6PmYRZmsWlnaQCPPMo14GwWWjpeZqGYMuhfHTGS0u1RPiJcdNb9jXrWqoesAPI
VXCs/514ji2cJfKfpEDTUWUz3SLMm3hBWx6DYH/XVJTj0J9F66KOgPvfGv87ctb8Xo61M3YOprW/
b9fGfmfa4pitLc7dWwUvyApKGsnF+0Z+zfXQZQ6LsZ0q7YNpXyZwOxldOoSrn6pizVFBWFifElUz
oXbCu92eZlrQP4sSDp88HyspY3neKiuPKu7Fq20sbnLfAOHRfWRoP97quHOboiPHCOo9tbRvv8IH
QoffO7Oy18pJMFAlq+9egq1gI2NAx7/dNQ+uiC0103vDbpwjC9ma00ZR0qwYwxqD/hbnX32C7BdC
IbOP4ymt1WxvFsde0Tnbfe56oBVjoDrBCxF7XbrwixNr0+J4D2U7qy//PIL33wBAy0OzHturB6FU
sfFz22xqzTKjPcNxPRNsQjQi8BtX04W3YfQV1TbxCsMstTMcfHXS3qQqDu6nhl3YdZb7o2uKtHmI
ZOtSmrZEbIUpPFNHofwuPf3pR3wbkCw0HwSM8fvkqHjggmhTAlq+e4+7nH1gRGp6Ro21/Rx5tc+M
POuj3v9RHHu/FPtVhjwoQQ5t0zT/fvyy3wcEHOWPIxA6O8R4BZJv94yQlaNAqLwcZDkDgiisHxY1
3oGlE1ATYrWv5mq31N6e6tspMIRLIcYBGT2WQEad7BEAdnKCsCMSG+rhvaGV1nxztI6YO9aG3npa
5mpqSeO2NmJkqqoqWnmvUBcJ2unCdR6iyaY4/ZFckzT+R7ddvSQJSTvzBim/yJy6N/aZgmwp11Yd
zs4q0sxoYkXon15VENhX5q4Ew1qRFjnO5U3aUo6zX5EnySjIj/TgALPqIHIjD+taw6kMWno/zqU0
X3JY+WQ9w19pzhL98ICT7ZHUIuaBL1dzYnSjHavJFeopsuf5jpHyn3VhjmW+maVbD5XvK0VyAGAu
FFquLMEyJFhub+kk6nnnoqE+R3lS+Ga2SfaH9kHQsJWIfloENafmtJsG4sWPYSNbL0ipUWDMprgC
4T81xLSg6GCs6OW747CmN+/BjAKYsEXij7UbLI9LSNVGj6piD+E7LJDBqnfjjbXvU4L9VkyRCyt1
xwmataL3LKzaY2dOpn+LynseS4rKHJSETavwkogTzRad6Z6HjaKNyUdERz54cwOJnmwbpxTN8FRk
nGDXd2380AXiWhxc01vO+5R3pIMT1ou1YBb1ZoybHfEpjOCuJmmbrTDLrPNZRLm44jSnLC3aKRQ2
rx22o/WBkCvNoFqWNNPMYooV5YRw3WnfTOYR6ZPq8qH6P5jZjv+2oK4aSvFqXjwWPnyfgxltCpc0
O3wAy6nMfgNYM1r4Per47xFMMan7XPHOXFhIJ3cvIbJJQ5XKVFBnEELrGvMzVyQerErRd2kwzE2I
WhDVNbPFbx1NjSYFZLNBRcCgWbJABojh62jV0RJ71+dssaKdBqdnhhsVQ25lhgtRnDv2g1m3hxZO
7BhYWMUmc/xqLxQ3/JcFqlpSFhfjKDSu7RiKflJ98Cm03hYDoUzhIhfpkYy4EnlH6e4bhGFgv1ox
/USug9wTVc1q+T2EgzRPx+smi+fY25K0JQ3GeWivMNpFN3gGj5hJ0TcD7ShUYxAq4SGLtlEIV4rZ
535ddgHGLFC43HfpIVA3tMOgkAlVya+Yado4n20IdEIseCSLUBcvrfRdMZUqeqWi7x8CXkeQu9AL
hXutZYYtX888Xf90fCapYOsRi3+v0EaDAjzFulMzmFNALL8mEGb3vKATBm2sbXcMTRycdlGZN5VL
ktXlKPjRtWWu7ih+HM4ZwfyIUMkv907ZiF3AfHQDTNn/OYltUBHqoBGdi2urk+HU6ZZ9ZKK7FPgx
uqsJtgwxSR6F07VKvpHIQiLKCyXBiDXJtg8vnaHbdnbOjXxD1u2zt7PEI1DFKbJgat/Ieh7+LL3d
0tRvpVnuOKCvh7cUrXSr2IX9z0bI3tX3r72PShHEsrl2FePzPNxcGwzIMLxHWv3om2KuCk5jZOlY
lXeJE6YBGFVIb3NFUkwMM3sQh0xOb1R6Yf4rzG2BlA6+SdLb04HdYrdfmWQ9zorOdZGzwyRgFOy6
8irLXuY5h7f+ZBu9vwlHHp6hQc4qfZtopKJ8lSA3gcCTQQL0bKVL8yhyXI3vOKd6DkNqy6YnpH15
RiiOqovG4knFgTbEIQBmEKHLXXXiYG3TmiDVe4biJtMjge6Fm+Va+8coOcTmtYhx2dgJSSynj4rz
sXxKDCpFdGibGGjKPM5n/1VXacdBk5IxT9QhN1Gkbsu3gPZ2Ft2l1dU4titY/To6hqp7sGaTfYwo
qhliq7RTqyz8ITXfTqq/RwzMMo5pdsE0vwYjS7ZdbQck/8JL35Iqtk2JWYRXdxfCX+MN1+hcUQvb
+3DgahbuGTAA3mYT1jgUHG/AEC41NBOmNj7YT4d0BHXr4Mzn8ZqxUtvAX2SYOeEGig4VMzpYNT7s
P2VnHx2+0wQgYIatu8VZl8YxWfUAwiNnEdyJMTbWmDMBcjuiVFcQmlqWKA3vQyKGjqWuDMVQBaax
VvJBDEPD0zZZDGawwJYUbiHjh2g2OSrAvAu8ApgMbW9oRLCASaRlZc8vLZgx57nAS8osGsdFiPsj
6W02K5N7Oojhdx8WRFPL7ye/r4pkHjcBS7GF0lJfxeig+iVjrbZN5pq+GRYvL4AzpU2Q9Zs1gGYW
tGm37e1mu1kriH+QvjWWKfXJ6x2Tg7MmntfJQvylsNrXVwz8aHJX4aZGi5OyP6b2f4h5ruZNgkDn
XqYeBb4+n40TujOcNPA9h2CqlU1dcFvidbsPPyXGh2Dgh8ws6as3NSS83bLuWSO2XrEgJMepo/RB
TC+Es30cbzE8a3g2uCJHeM4/FP8lQojEg3tuQslLOXi1KWgo6NB0+nW3CCDY+gWlkuu9x/Q45CYh
Oo7KiNrCuHX5KYLoXM6rU7D1QH2gcWYogZ6AXu+lGhhJlAIE2TiLh0T1REStovGmQysAEmUeW5eC
1eYGjCby8FFGwJCxgM4D9q6a27Dx8vsXGUThHZ4xxZFbID6NXoxRvG5zeG+/nIJ7gC7ClGxtG7af
rx73AhQNcbVuHEDsVZmtYxalNsy5lWTS9OoC2NMGgkDgsah1nwAJXiOgcDUfz5B5I8vtbsO7hqr4
n6v74Uu4hhKGwcJdBH1gIAUTKB9E9dC0D4g4OYVgzeEvhW0IR3/Sbb1KWYevjzSCffvCUxGpCcj2
zApJMibzTZoVc9ujlgQ3hC76o7mIjxnflZdaEiMuvEuhPy41oHMiooXvtok0OyNyO5UvzuZrrmfH
acMzTgoVvWPFHNRUoEgK1no36M0Fvsdgcvo42hLRxSHJ6kBjQg5LJrnxuvoGvifAGCuzHC9O7yOX
S3UoMzXh2rDTuXUpzpN2D+IjdNBcB4diUC7jf1ZajIJJk265av+2/AnWBeTwjWm9GqzkR/khGoqk
EljbnOI7nG62AE4wG7vqSMQJTTQZY3E0vN86qrkGOVz9mkAtDVMtgle1cLeEKqzFOIywrel6mBUq
Sp+GD4KlueiMdCyugDjpDIYiH420V6vKtRWePMYAFfroGQXGTNSQRnzNtsWb52JsXcpwq0C/PlRH
sGgkS3LkA/5DXMTmjL8L5Ptj2aFef40RLZdz0RsvswE1GI50mnl8oBiA/dkhwOufCDTDERUMtF0v
ORGhrtJgm6w+yTGm2t14KfNQtL3e9KPCuuHAtoj7u24nAPL5lS9A23yAUybOMcJm0Qd4lYIkBZZ7
GdqRTDB5SBtW9CA6VG110Liw+vf+vD1arvD4Q9n+RsVZdDnZCfb7iWID+e0xF361cRA3NtO0Q6xD
Co/3T+Spj6Q2GT+XX1be2d/aNREVBfo8/dax1k1F0kY0/u8QgX4NuR920HkEAp0ac9Eu8XYmxaR9
rtxwI2aCthwPRFUUTo7c94J0bqGhIU40uIqrEU2OX/piaXcmbKBbDGjYUpi1iwTKOt71E98O/HF5
2xb34nR1vhaTKo1oKf3seD66nkiMWy5CiG4IuUnRUxrZW/4wjOsiNFs9rSYYIAz2WFGFGe1uvL/l
YKzLolw9iP1a2KsuQ29+gbxME9mfxWPi8TdLHtEgv4d+1pUwEIfQxLp+lv/8B3CTH2P6F2AUj3f9
MhVtsyNeZxvfWmpFPdy2TUWDzmyDXKmXWF/g/x1fOZXBTyQfFIw2TE01vk61bV8Bjbt2OHt4L2XK
HkMZvFapfaow+GTbCkxcWg8iCTOnamsf72tNlbTEnnWq8Ej69lhb/G86YoFmNjxrapNKn3hiXXFO
ZDVo4THUXTUPfiijLexmpqftaFFSyNclYQlEs6l4wmAyNMoRVNNYaeqVOTOhRmpjBh+kwGMLIFqh
Ar/uET3Qx/h7qq2Oid4jsm2wigqhen/dyqTHbu5lzvyoC0qKYGfQHDkhkVP5U+6gatp5s9C3x+i4
zAYqFHzY5MNOizEB41akBFz7gYEGhFvx+byehAMMlEoBQg8voLGn5pPGWyYO2l6+Vic/3QhKGAFF
dEezU5Mh+Mmxxc/9D6gs+ERCwz73wnkOTRbbEswlwHJ7ZACgzK0YuFkmKu0o6M9MmypTKdCwzgUQ
H0zvkrfHX0Ju8+t+YiRcDiNy5+SRNNAkf08Bx2+eRPC6Ra2G4WHS0a+Mo2Q1rtkF9ycz9rhV9/JL
kzYWdCtRNo/rl4Up//NslhGPF3zPwXSZEGvcajO4cEExXhHAtuKux/g3nnMQvtATqs/SwTCSb7oP
9IQnqTocm+AYfswb+4Pjlf5ZwdJhfD0FelIls49kPXEs9e+0ysjr8cbPdA7zGaz+32OB9tnHDV+a
XAuJH2Y2kqV0PHl6b5wQQmUY07zcnD53Fo6Hnif9JLz3DDd3ofk7hb2Gk3RRDxVeWm87zdaoqjAu
AK6KRUn4HJnFPRUjmElUS7DQqdoX4WY6vlZEHYVUzcDwOnO7BZDPH+C8KRypTuSJ9tL4TG5LTEy1
jxCmCSqFntxr5hLfO6Z9xKmyKcf/j9NvZsPIiMVn1gfrzZHP/DQfWhdxcpuOsy7w70Ncaf8MT5Ul
5nI4VGxEtmdfvjQgQRv59n47yjMctzQyFBKnuaHLii9vXgH1nL0iBxnAZOszUs/B3jFuWKtu3KZ/
SfgRNC2+J9VoTXUqqke/jgKHhn4tU5+sJNAfbDVf/HmVW8LFFu5Bah5x1fgRBHjxmocfK7AqeIrZ
BS3GyDBFA0ogGqvGYln7un6LMT5qFxRfhwR7sEJ9b1QQCF4zj4MUJdCiOJuOPwTYKYwLYywA+Dpo
0jWMRUk5+m07pZQf+U8tucydwe/39pXgs9wIc85I0W0B/EO43S4fOkgg479aYoUCrpekHBVeJ05O
s+bM4JaimUcUc7RusfUH+bir8xvgjg1K4PMzX4HHDHKMI0MxqttCHyR5wkAfNHN7fKSS9eYL0oFe
IZ/1xpm2iw8xVdvuGSV4FeyxDJkcDBxakRu+yvFTwiiW7hE78fJoTHUbhZrZwbC4ips5rMtGphds
J+5vs69DyuirTPGs2EUb+ZicKjsFAXeB7QCsuknjtNCRTMLgnzhTaB3yTVBkb2bV3XhH0ZeE1KpN
x+tu9IiaO15VtLvtpH76QTtwIcfFMsiVVddZAtOFdfynIZZHHC+/BhPT0ylJRBGU0Zomrqp8JtFf
rz3xWOrZNnK3osOHg3L+nyuofbGVm+Hl5CxgoS34ZNCNGR7vz2DNR76od9Zbh/ahOmgAwKnOCF0l
TZA2So/ghGvzMsG758L2xt6OhqQ/8e3kdIBTNMNckC8pwQcGTxObJxdOGIHGuwxweFe03BOMVOz8
+zi+IHCh42CqwUoakIZ2s6FIjN2iWtiF5s/QcHHZdk4VKn52LZXnzJdh3tx9wfjzd5fSoR+1HSCe
as2iWgvOW52MWbZ+XoBrNEV2OKg4XqTM9x12PWHyWWzelnJtWC2DdbiB04HyI+nJQxkhaF3izlvY
8l7gZHs9N/OeP7C3bzUEihFDyl84DrJtoyefzGQSEr2Yl4o9yuo0q73bGQJu2lkryDl3BDPjOONl
OHZ9+OloQgN/xUMOoIQ3aGsnTXbblrr06g1IMEOz+EylO2tXIZTLYYJH97AZjB+LbMuQ08sepJ4O
5JYFodK8UgoE54QEmZhnIFNMeHsqP6wnHRypuLjotBgn3hsRPWQ0R7Ra0IqSDNMNikyoRIdlDabe
49cikUGQRDTlGr6lACZAS8VWwv1ycQQLx1IEgdQm+RFE+bjEeAcrvaF8bg1PPP3L7i0b7mfa8zHw
w/K29fOIiTBDkJ+nPNh9aVMSxCn6Aj865tKufIE8KETMU7pXPWqU5EwUSJmZlU09QesKQuSGjMGW
27Q+6vC6KP+jWcv/rJjD9vLxdITl2opelt+D31Nr8SzRLVp2pJlki7hlz/dPHVNlWrJ+pouymENE
wETkE3IxufszZPS7lUv4EcIOw0eBbnC50o4MrsbCjYqTKKpplz5IxuOpZEpz9puvh/UkAtSoyEGp
qFF6n58+5yenvWJsksuNT6yRFgQQjerEBtaWYViusI0hrIoBZh6a0k02VZxl0F8ykZ5QbRN+0LyH
YpNF2J0RSLSnBVL+XMrY6aSFn7j3yHpHDm4tTEjniihYD1WOPluuyAx8y/ZCEfyaO/ufRlwDUPBw
ZlWppSUAii3rHuI73HuCpRJBkprNZek7mZF3r1IzGSW8Hhkh+K+miFnL+uWwktYgaXIusIQRYT7Q
b5hyJbytFhQ6/F5iUMHlOBpo4wwRUT3DlrOu3OfBZZjqlm82Rg1mCV0tBH+vVGOwjFbWn/Hioxen
Dd5PvoKm+3Ra7hapLcS/ByzJ5agwWPfdMsB+vpba8G38/HIcvt8/uC3Sw2PP3LDt6eB9GSXl5zXI
QxnSNvXZvJxpZ3O+x+yJFsVZKbTlXtu8sFsKR+hNsQgKfzFeZQBUVHzkCDcqAtDQpj+BjG1vVqok
+TWMf2+Sc9gZMkCMX4iqRu/UtP4RNtg+fMki2Vu39m0ktk8PKetdQGz0+08I8SGyoaifPdxAp43m
Xm6ZDp3ZoXikwSsUXfSS6ed1yX+cAoeS531ZOb5cS4Lok5BIVtIjRwUHwTFzgl22P4c4ASmy+32G
CsA5kwUsrJNVqt8A6tE+Sqh2JQ8ElQyLaXey8C8V7dnt3ZG6RIIVEf7t1PrZFaBXc2x5x/zSrrhy
UBki/Gn1HHX9FXgp16lANELr8Al6W2B+g4ArGvQAcxKsv+nTdPXb5nwPCRtrGEDI2i8FfaUPS93u
BIfk5+g5g+i+iJ0yhp7D5e5WBHzl+74puRmoS/PkcIw/dr4OYAg4XfDcGYvZbq3dG07dMHyBncAq
AZk7S20YujkFUWNK8EAPEArit8d5ra3ozGcnfjIwyZVFUb/1NfWNjxaH6pVUN0wX5r5dDdZutNto
NQNZr1rmt24f302Wp0FGf4u9Na8CjxrGLxD/Gns1OvS2b6gZBK5NiRAr8o3uKxSWGl98NjXBjyS9
M2Sml3wvD0rlj17iIyZP/fJDuVg+Jd2XGI3DsNXtju961aaU2RhqUpaJTDxlA1I7tDY2guZZULw8
kSA4bi+ccC83pNzJo+35Rj4j6geXdWFhy8TEg/EAzQ7tyl4rq9WYBYD23DnncTQYMLIF2k8HnGt8
2AROo9ls/ur24hDpNuo9ecuOpP+nXc/S1JAJN+F/OhDwyF50p1hKmTw7mYXcwierJ6iqFBF87CGt
PvBsd6gmHZFNxwsQoYtLayLh51DJDJuuuy0l+c1tZTLUyMI2Y9WWa+U7zLsUGX8oUq09DPOeIYao
4NywHdRiZtMtCs/UzCWiz4FCKhjXmJ94ejOhf8tpSHZogTGoHztOb11HiSy6AXUBqhi5eMdBUJY4
iNlEdYjcWdfeC3XjhYHkCD0QJGuJyD5nVEI7KDiLVkvZnYSK+gH/U2EqNRfsfav/KX8i50EqiTCB
A6P05JXXl2sfPiRMBoqtJkqDSxqJiWq39udJ7VSpQOmXDEbeONvuiPW9Ws1xTf1VSlJqRG8+9F1e
eUSQ/+6jHP9yHgrw2k/1H6DWdhoNQUufeWXSu/Hj5Kbvg8Q0qYvd1/5wUpGbc1eQgy65dWrOGJgI
egfBPzzSklilgngXczHYFLmRJ1mzGQNkB6HwFHNJhxtIc4qwYN6nR1fUCvi6cgku48w0/mCTgnBF
ilnQCMiIjj4QTCFEKRz2xS2hJOIiiZyKU96fP/eNJ1eWxaTDamGEIf3qsYJ9QVQRpOHdr0Jl1kDo
6cW7LmPg+MabDijAkpSh/Zr+VIsOim6dEm/4cRc9F6wjRVkU9I8Zu462e0z7i0HGVOv/qjC+JylL
vgdYu9yYqHQFijSZPb2c8fBoQHKL+x5DhEdhXgSwV4A6jA8BytXW5IchYAZIVcRRnzBrRvTBnvIW
6ydtpC0nUGA5ufxoeDKQh79ARCBOQkEeaDNQJROm3XCawZFwA0sKA7X8uFAByBhAIiDBDjHhnnTZ
akPhcxc3DKBXUz4V51TpXR04lwyw6VDMJXpEjAHJz2CZT7NVRiPMduZyBnWKHgSE1CMMbHB3FSCk
y5wyqz/gErt7+ZnjGUpPLW517TWcgcwo4q+olwMZj5xcbUVVG+wxgupdwHiNjA6OEbEa5fU0o85T
s5slHiedBDLckDqvz1olwAWqI4DRVyD88b9uYr91gygE4fjjPsncxO5gg/u09xT4ulwj6T6tLo1g
4Z5nLTiXNg4bP5gqYEdIXPSGGmCwo8bI7isBAEKl6O6lRzoAZ9P+43HzGd1SQ95luFpOn1/oSmmJ
pe4lw08JryDrZ9J45/1CzdCSYfVan/HTJIR+XHpCXzDB8o0c6MwxCiIvRXKuM8f8Ic61QQAc/CtG
lxoGM0m8FHegeF3483iZa1elabJycCfwKGxK3bT3MCoGzSO759SECpdh78MDk3zvoSvc4nAz9yf0
wB4BcAAmIdPSC9lCU54eYA+ho+ccBCTmPWGpSzA9hFr3BEz6S6Kc0boEEHZVVifFh/py4QvT63Hu
ra15SKJ0M7pDbd8OFeHiKdw7+htAoprUS+8XUUcps1EovJ4UrWsYqH3AzcQQ7hOBImuVo8xiGhds
ZMygLMV9u52sC4049Z3jHdA9JAMWJxVR+Cu06CH8GjbK18jFS/Xt101nLa7c/aX7bBhbSK2AK3nO
6Ms3IyQFNrEnkwAzqxVXdYejj5hYC3K2KgyS4jDJ6geQJj19jMlk2vw5GL/IcthDPey1+TxDCNLU
VU7F37w9xCLPnRmfA9a6rGOIpWzOPiJPoKJbU+xL7YMTVAJpV0oZPMo8Fp9odzKEKvtA3V3C7HwE
zWPk/7gnIXip7dgf8ZAruK+S/HE4XdqoVIXQzonnkSy/BJzGneiGZAWNKukgMPolDmsch8EKgQA/
/ZnJsCNwt9RJIlzby/q+DaaKL6Uz0G+agdNetKyhWE6r2F7PCbdd0utOSGI0hAwVm2tJfavgMCm4
ww7jRscer9Zdu8p6DxQMU0egRBs/Xkjx6sY69fu3DGjZRjWj7PumOLfKDVS3cb5mhXvlHeHBt9vh
+U43e4s9VI8yvY0GHJDp5fm+XS0lkqZR48CsaxPHVsq7vqpIFY+BGF143UyGNTiCmRa8xmZ9ixP1
rc0Tv1WnA++uZCCEmNOgyq0RO+wLSzBJIbxmCXt0z8rXTSjS8ejy5Y4LA+ENR2Pzmj6cC9hn9Xpw
H2tj6V+KlIZh0A9/yf0pxjuZhz8wqXR+uh6yxCoqvJrquXnDoR/hykUYq5sOJyP3YjPwChTk9hIm
Cq22vFLlYyScZwlscRsUdByUcgt1NhuVzKyAePoYrbCkQM8mcbBV695WhFUaymM3PtfB2WOyOID8
NbI3LTSIPMlMA9TwYVOSSp9ys86ZpamiBSI3WzUnA2a0OG1d27anVjJlrjWnomm7ke34uhs8dvqS
ID3sMI+GOdjMYifC8Xkr4oFecz4TB59TYfw/1T0nUjgdcBJYJjRibypXz6IKcpNroKiSP768V6mH
4AkzXsqp9oXoMrJj9fThQ/GqU8j2fXDZBvjNiFRiY9BF4/VR6owzB/zM/yZZ6EIu/jCv3d8eR1xB
WWigtbiUIIi7aPtsHGxOQmBZuoEyYoOtdlqIFSCXm6Zr5ymQWJr/O8XJhHwHEvcR74P4BUEcpCUX
1YSzhk6qa35ovXYMKhdB9mO8sQ9RrqXbbzdklylbV8dq0vlGXwltqFRnDcXr6lZCqdVVhXBzeQTJ
MUq4k7AyLTK39GNFjH2M3PRz/xaQOJQuIgidriZ2+22CS192UudZH9WlyCY2GOZOS0qGVFpn80/z
ZphcjwIdW0C27DAmVLMp3MC0tdCtGEEtjQSIScTNN2GXnxAOe16pUnH6GIRdpan74i/XtvbDcr+k
wEgeR1dtxVzWD6zAqdKUg1WOeLZcxgLupzXIgqLeHF0GT67Ewx5UXI6dEW3qH8t7jbmTabT3emmi
LTTz/lrbEQM7u3L76qwwg+hS2zi0XqI82r6QSDI1pzQf/syefc2oSD3Z1FC0780mDCzoUL5I09UD
5xUmh/3TX0HUYFCHlXdW3Jbf6pt2qYex+m24gaXDwPYOpepQAIMj4CopS8SJfpUOi3XBClsJ9GL8
B3CGMDrTWstqX1PSlj6OOZMLDYMMt1e7Sy5keLOct/GMuP6X0Ec4mNMjalC2x/cwKkFe3n48ZdJC
vm+irQGJVCckMeGnumjhJh8Z3z2Ahlns4Xl9Zyck+G55x5Tk+V4h/hBPf77bs3JvmphqiFQU3EAz
zqgYfO7o/lwK4t2LU884vgV+cu4ebq0bHisTi9puthjNBC7qUACkeIxZmj521w5/FGohCfQzCjp9
qUZhr+Dc8HjwK95bT4xlgHJzDlRWu3UWRUi+C+Kcygub72xSwscV8ZX5s+V+P+g2g7T0qr1CtXYg
fh5T2ebypfSGoEvn57q+Ou6DjusaouOwbrTqbt7kGoUM7Y0kxyPi6AbLB071c5K0ZgRnFtcLmOqE
3G5htYdHYRh06MfIvCnrk2iBkeK2EskA7LT2BhkJoUNRuDId7US5RIVff6WDB35uEdHoSi9rDdGb
6i34afMVO/+s+ne5SDwh0YiZ6TQArsuNcnymrawy7l9dJa/62Y7z6maN4RwXXjbN5KZLwk0Lgukp
U9wnpjRIQ5fP0rTN3YGWz6ZOff6WU2XKLPYGROBJ2sxwTqM9le8sKdvuGcUeAO1+rPTHkCtVnIep
WbmJ7bcQUcl5PRtDFUeIKkWjvDg4xpFqS7hazvw+f/9HxZu77GU5gvUibjLU34xdysnIHGe85y9x
1vVxYKj4HWhAEDntgWh6X2MYX2uIoAooHHduCDd+cgjisr1vKnIFrRv/r2PUbfySkLMA9BBQAOD3
vuuxqg6z3S9Fxpx2TZyjoQKZmVb2dG/xtI+WxDMulaFBp2+JG18UPdtM/hhWwZ12GFWnOhXkHuJs
RPZfqawDwlgxHlyrUEWASd5bHqAiTnPifMIYLLcLYm2NC5AUu0effp5iU4ahKFK15bJv2JbSaAvl
xyGDm31y2SqkvvoyQJ3yX3f9AXt+UwbKS/dD+47LL4SWnNYnA4VCi1Tnl64MISge9iiSQn5YHWsv
HFv/3/7VyRgvACCGu/taCAeRThK/gbw5+DTrGWPF1m6bRe91c3J4QdtgT9EDlCRSs7J1PlYMToLE
A25+QBTgCWnH7zrLpaQlHZXQKssLeS15a8VhSDEKyDr/Xp1huFH7szWkWv5GZjmfSDZpxBRYSMdZ
pwjHvmjBoZ2ZGwdvMe/41oT+s4KQK6G+TD56mPQMlyPnr0bigyB8aD6/sG+SVP376Gfo+a5JTb1Z
uXVv8EqiliZgFMSF/1fP4E9fv7REIwzHlomJvY8kyMwOCWuUF5XTtm/TYZKn+7cW+fGMBErZgB5Y
mY/zu7FMWxhKV5ANgPOVkPuBi+yHiN9HtjOBEjHNKW0aztashiKBmoDSU6zldQ67cqwie3XckmwF
mDggvbcHb2op14W15AKVJGiR3G8erKE2obRmIT693IQz9qwd+l8NV9jUSWkfY/Kq3TLUslkp9pmL
Olbi9nsiVnssjfiwQqoAJyDqrazW8CXkV44JqgKweLvBfGJwAGb5rIqY8W4o4eouo+EIKRgVQtV9
TvbVYx2AVvKYDKPsqMoHvbLeXut9r6lJp8yk6c2/UUCUTv9QRsIb83mco1peJ97KflpQGgJXcoE9
WW9tmrTpV0GdgWJcjVr3Do+Hg9u2UiplXupKPhCL1U5YgEE5FLx3EHJHyfTBLbuorG4CyK1VdyTR
AhnLYpFW6EL4T2YAao2Ex2yQurElebbdMccxAkzwHRfShq8nZm9BYqm2cS+CVCbO3yVC9wqdOyNg
NFfmc0povg1cSkZdE1iFF4U3QoaoeEs1Y7Yo6iF9TbUkYq6gqN9z8ylyvCZSuXXg8AlskzlbyuV7
ZuI0zXnK3aVMrVgiDqsGnozZIwJmVv0iWVUgQtQWot//5JDnVbMlTnf88JOhFepoxXyV9H3iAZ8q
of2G2X59MRWdpmgzFUHiRlZ+fQp3kENmxIuFIXsqPGqeHPHiiMLIvM5Kvyz/4djIZaZcTJrCuGEQ
joxis9BhdOvDjzj3udJ0DLBKogLWTHH0mCb1NP5Wi5MdLSuAJOFoSFwJD5OPQvIjp5Y+UR086/J2
zmklMpFdOrlMQyyXl7w7BN9J9ZWlai4b1nQzBGLTwwDJ9m0dGhuqG+RcjWzEBgEIemsqG9DLmywo
SJ1OcZLSKY753oDrYsGUHNwvJUQ1jZbkCMrON/CcgoIPx1y9cnB+jQBHg4jiAN7dG8E4GPMTlPve
3lbsXpWjqNau4K2cmcYX6bV67I+pX4Ao6ibG5MKzQDtboW+ESg1AOsUSjSvD0MhX5bldoyOwgsPl
WRErMTvPMMri73OQ1b8OclhbXkkHqG35Y2L+eeyzIHwVUBKR0XtJo+DMH0OyoVta81pETrSpU3c8
Fn60vgXS63iXOBgzOEB/LMEX4HsJRPbIotxEjpl7F6ePHg4GmK0EDtYsxnXOQ5UP8rAFfhzsMpz0
GnYyMJFt8xqhabYtCI6lgjemFQrla5GiU/VXOLTo0wqa5WL69OpKQcJ/dgeg2CN7c4Bll1AZQHWQ
9nqpmB01GYjrrC51h3tuYbq8QPrNXo8zmZ4IDOPXmzrAQ4rU4RoZHg4v4ygWJy31Eu2Ro4qI7+WM
qJewseWnAqrcgjcJPVbudJN+yR3m2j0cYQwyiJYTi016gvXwU+XkEcfeUxkYpZ2M855WQsvIF83c
JnBM35d6FjDrVBTtLxrvUJi18Y0S39UxsncVRu26ejIiLiP9qzmbN6Uq8OV8804q2fu6vlfWziCB
xKsFJOITwERYUjoUo5fb5aRE2ciSoAV/RiHQxABw4BQiBUEUMBKfF+X9ghl0EzJoE3bLvpaJL6Iv
ZTkLleUVtS09a8T2ExIz5bFVchsg5X5D7OgKmawst2aEx3xTI/Rz/2QY2o6JnvPPpqNvJvHD8+fh
dk8TOnGA81H/tnHSLUjDZIzfyXARudL2AHoLCFqriu+Uxmo7tjQ3FVc5Ul0HbMpQqypv58YfdLYJ
yna/HJuHhytvTvCYg+qUNl1WfyJskCZ+XdADD/jVTyzg1moF1KyodQEtWaRqrfg+sHibdGw+Q27D
3uuA5NULPbTWxVW46ABv+Iewnbp95mm1bPPpEaNAdcl7Tbp166g8VY+k+/ygDOdym0BDC2vUEgh/
2FEgH+Q+g1PBTm08dBNo50OxSpChCq+LW09HBdNP2dwLx7nJLr9Lgr4GjpBm/XDkic+EBnXxGifY
oh/ToilFxHjloY4a6gTevLEqa9b/cD9sWC6aypoLTK/7729IRGlEFAdgMOWLtrSBzFH/fcCdr6J4
bqFzlbgtsyLZHzi+C2DduTUCGSlBBC+/7CAt1O7ykp6r3BhXHoD0MCr/XAMY97jaRfOvtK5a71cU
2MNOhwkOB9CWm2vd+5F0mBjTI+gHojiQ8GQaq/OzkN4/9E8ePdYC6M6iS0HyCLngz93vYQ0/ocpy
UNzp1XZPRNwweCK+RsZ3MF5k9YZD5VpEuhOxdXbVpnam6REzSfUSB7VcEf0zXRx8w6QM/B0uXr0y
QbyY2lkT9SoyyPT8plh8x1Gw8X0lOjxNR3fj9yHUVlecMJw668+dOHqM504vKAp8FKvP9UiDZQYO
2gLlfbnXdcSXg+Zz9cZM/gFh2r48TFxKyFoCszpwSEuL8IWicJgmKGXx+/Z7YV9rosKmh+LYSWuk
IsLWugf8exo51I7rCdRxBdPE/c5poEgqXHtuaGmWPpsWl5MIkmaD586P0V2SA4YcoZCLVlQLykoL
4WKXtKaLyywV8PhHDXOTgu8rwfiyUkaeTuZiNvFguzIbxzYa6zukkccGXh+cWP1JrXxTQOvaVbow
Txw86svqDxxM4gDzxh2eL8YzAU9z5gn2ljRlwslVml05ZgB1y3hzVFAChnM6o5oqnPzxF0cN0zML
yrVeMcNfz/KfvkQSd8PnPLpzbMutBj03UACokDcfnjJvwWfq/un0jZ+bULbRF04POV2WjcPNRZHd
dFHOvEEuE51/+6ImHox+qNpdSk0Rjrfr36jNemALvD3mML8gRhH/dKyoJ+hAjd8y+s7GmQm9RFcx
aJmIb4enltPOAvr+g3GtVGoBIdJ/EsdsKZa1T+FbpXrKqhse0H+Hd4xUm476QOl+d2rrLqQ3puyE
IThcz7dltYVXP6JJVvn7e7PsW01zy4ix8b44lAAxynTMU7kyn/dh0t8Bt9tneP1/rW0PYqXK545Q
EUUbBruxt3bia6fjgdGFe92oDG2q1UbD5lDI9cXM8wCkDenGXXs1G/WCGa6TcUfZpNcr/2A9gyMC
7YaNRSJjJyH7cdd50zz5TiyvtpQyYXb4pbjrVAzuVxSU6hJtSYd7L7zCvbBj8VnFpOqu15lBCcr4
7QBmCQO1voHsxDZ+TYwmlyEgr5wKVSBymGxpjCgJbSBCOW7vouFYeZV8OiMlG0XEOcXnQWqs2K1P
tkgmxzp58DqXJTIf+/ODEwmQ1UMgBY/pUOymbXKOY1gY5fLcfQOL0ry46ObxExFeSH7LR45dSDTn
cE+cwSzBLKO58RJYJZgX817qOzKvKEX/k9gmyoj6hh241CjVctk8bo+T6h2dX/Qy3vR7mONnTkJy
yE7VPQ5kLkju1nDcfCcp4urg12bFEOTkI5Xoq7nbeT/8Fxzu5k8r9BdBKVP6W+lydp4E1SK9ZC1o
UsFzGK2i0FkOI0d/s2iSTukcgdEXqBaX6u/FStjkaaOyUoLAwNi1u6qIibSMuCisKEP7+K8MSQmR
qDg/yVVZ2MF7BTkC3vtOPHDfbkgyD9b/Xbmz81QQQM5q5diX0Wtmkn4mALKPstiVY4T5LOnDmKI4
2IcmIrYqQWAOoyVqOpKF2rlBsWzBMmps3u+RBTA5cIvFvv/bB4QztDCwetvPnQFu68HlME5RWCqf
xpzMGW0VtaKF43Za4zQHwi9NmrS1lFsraFwLXJ2JbbTbNTKLdGYpEg0PwPbqckB7EZiVoANf9gAj
7lQXsuM9fNRGZC5FW1ouBt9KbK4LoDQCD65nP39o+OvRIIFeUF2dnMrUxmCVbXatyRGOWd/5MrcJ
gLNEVnIxUuRX7D4oxLrmNyahsxYiKYlsBVtNVGb5qul+wTdKLQ0jBy0S/rZ4H8fNTWN6oAUcq/LP
VK7XE70B5DK+pyicUsboqxz4ireBwQ0A8xS4QM8a+od3TPnn/vBIvyb12gqatolEa0IuYi7fUwqw
psKEKIjpgHuolfOTlU0ySlfN0LCip0VlB8lKauH7+vjGtqdMFjh2yHy+jQPv0H9D8vjz2O1pMDNy
bcMAsEBWH1hdPjFY8pgYyLNt5ZL6icuO8a5zHN3RieoyyySId90zdv9yw1/C3H6JXod4jULHDqxU
TLzLztVmeX+ZU+dtSgCKB+MWcoVYRto4inNZSPsqwbG8lh/xVdEgCcvKfNBxi+QPRAQeyDxxrwn2
kdMMBR5koLA1WU7BQrf3VsST1sAKD6ompUmu4kKhxaKC8foc5hdq225KqUx2BIxicOsMRVSXbs4n
SN4PLyc8Tl0ToXSw+ZF96gXIuDZBHYxtDUFxZredH6sXr1mXdtms3IF+mMn3cxB3o33HM2f3F/Z0
7bcHEHqi9ntJ1n2bPvynqU4r71J0SkEr+0Scd/r1D7PaRVyW5VV0Rbv/XF1n6qr9LYu9rV8aWXY2
AlSOFqNIW1u68/UCX7aeBzsZFbVEInW+9F1C4h5Y46+Kfan+ObMYZhTZu0mNoX6zIKCjLX76jUUA
s6avqlDbDCoR2R0+1EFE+tWcpP7qNh3ls9YwvYnZwPZywoKPG6RIUjDe5eoK+JQ4mlCuWAbAeaDb
9Cth0iUre0IPIY08LRGnrR0/YxE40N+5zS3EuWB8ToJfNelyBPqEEgn6XRrZlDxQR0lPNkwXPiJA
7s0sEXEuVAqRx/Y5uN1Krlw5h6YldYzELbJXpg9Cot8apTF0qoHhRb4/55by1qVmFSlFcPf8k6wR
Ymb/dK5Wmp6dHWrH0geBzfK4Y+0EDhPw/PuWN4iaK6WtZhPuWWcDD8Wup2YB6e2D9f6nD3n080Al
jyXyfzQ41slHnyOBcVln4aTYF4bN/Y0CjZTvPSEJx7F1Uvy2rG66EBWWs0d+0XbRA3I+zgZu6H0T
bfEusSv0GSim/9oyr193S9FRVlDPk/b/V9+0oMFDqmR783+1ldc0u8lbCGUf2J6Hp0s/NN/MvANZ
EEIw7xks2fCDJIS1WDowbHL+rKjkwo/EUnubzb871Ish0d45GoXA/kkWRFLfc0Y9sQ0uIi6c/j29
aVvQuOtkAl+IiR68oLKeszVaJRHkkS+1xEo+ylNoA1cfIcf1IXeP9XO0kif3qficxKK2yOHRcIA9
TJmE55D3UrgdXCbPktdQeiIR5ShIP36W1WQjvMJ1xHOYkkLQqMX5Zc2Is2044Zpcji1xzSu8Qv4B
7FpwQu2lbb82ILxY+J++nL8voBZnnVKm8nA4s6+r2svZszEOZ6opzUnnh01IoTuxDmz7qUbF1IWo
nfoaegCu0TJC3eSNYVoPOm7KidEmsBnLm+zFN7JUOx22oc3uGXUAtaW3mnKpWWJxDLs2GScPKDCU
CRkyW8xo6VDzr5//SWZeo3V9CduhHT5Ow8Pa3kevudPWzanDJZrE5WFkJomFfgTqIRYgMPN9j4d0
sS+d+rMXLVJ5gnKEahPtLgUI4uGeue7py3F+qGaCxAtgQNNTwBMfuZaUCECMrMrCuZaFrXKfxeIo
LTBbp/yacC8kEgO1fQfCwZSR0YSyxEUHOZ/U9pHXsbSfX5ZYDjFo8LNSMYfDTFNW9FLJdI6fjy4w
CfzbQlvWEtSIdEVuxdfUXXV6VtNbyGbLxdrnvC1lgFgBoqKespPxrzHLI5Gn2OsUaaEzDDcM+BG2
JkslqAqPHNyEXq6uDpTj3mTvUskvGbTmMIyBDwcAIgd4lKUwsVPZsWRxajM6mXZosEPnVBO8totG
xect/LRncOD92V02ICRcjzNOB7P8F94ucQns9vrITtKn9obcF+3muO5oiX+kilAxHefOve4yXd5N
lzwHnL5ZRDAU4sHzp9tlu8hphFrkwX3LwIeFrooedRMnqp42q5RZpogkGRcrbo2W2zvAyV4gAtg9
my8ZEFtjO009LeJSBkH8dnZrK6nwOf/T29eCatM8U7wrsydHh8wsfbcFscwF5PAs/pN2M7Qg+ZQr
7QVe636J9KAlPnYrkOEJh55bSNpmBrB7QWkYhbu0gC0DnJuQcoePUnseXc/3D12i/ypNZ53d7Jhf
rkiS4DyuHtGe3Hun+fsxDC2LwqqkdymZIKh1mRearcL5DuOAoYTx4XT+OJdcV94MwFnUzSt7f9ZN
05RH8LrQYleBx0nLm6ZzZlF0dEk8xtvFg6OnMI87JeBMcg4ze7+sQFN1wBC8hCEnk9vyxikCsttQ
ZPGmYsI38gU0gRQ6WFPk8JJD7l0Ak0HBNDg4yIxe0eOned1F/9+WVyRjKm/K+Ink9Jb4D2zeUcfw
V0MsT/JUd95hwzrmuj/SqBkqcIvJm726X2+we1kWh016IHJ9VnVh11T+xBh8wpDu7O4lgdK8eeQk
RWZ4MIXeJoFx8kC0j2P60uRlPhSDEYlHgHUwLud96LDtIIBigZAesmyOUscnKmzEiDBD9n2iQV56
KMRwY9CDT+eHfEl8p8ijrYRX8dyz7YVFr+mMTyvwu/oBUBXN/WE3ZIhBV5qHfELjqHLWGqTASGDo
ccrwC8nbILpSBfkq9OpgDDphxNFQTYa1purLJYVOXAS5CevigK4EgmyEQsaZqdJmaeok+2UVFDD/
XuYqFZa7Y0fOpQq/P3JvGxeAIKiu8GCIUqyFisz6/VvPkslEGuBtTBbzcP2TSfcPQrxf2YHe8RtB
9PDqreiuI9WmLB+Gv8vqc267x+CGPKII0oxyWTPEB9PsOuaV5oZTgITGxodE7ghCFXz06aCLKdiT
yqEMUgb8JPSOyfWjFZ4Vq+U9PeeaIA1RFaU4Z0qy2IDqwNu7Sw39iSHHPl66i93VDdgUDmG73cad
jHyn19Nj/e1xE+cYUultoaAGWYPa1OwjzgsrUpRqIjRulwuSP160JE3mvtYYJbrfx7F/aDFVWlwe
U5D58U4+Y6tKy5x5vafGcF4zWuhDnb3t96c8oFjZtVr6OnNZuDUcfFOxUzzxqi/sNACX0RGnq1LJ
PijwqbB1yr3SHZL05LpePgeqciHfRaYtKmr7o7x3UShcxTHro7wAjBom1yYFP8oZmYrtY1g6/X+H
5S2GJQe3sZDh1THA6RMaaC24rUsnNPS8IDRnYyxTDFprpX0ompdxA1fdcwQFZxybDEeFa6z6uBqe
6FM8Ozeo8M54RFrPfW+FmdunqhUhzi3LanGFnqJAiDDNQX/sNB+23Ifpez3/1HQh4h2Vl5uJz3xf
R/vUj+bEaE93ALEwh9gSNhwvgJnrudcRqIMC+VNqD6C5BON3tzsAo/aHW88wWQmztLiphPgzFDSQ
XMNWyKdKEqhNPtvTw9AesCVvVbEgfv8Z2zQlul2u6EMoTDmUNzPmEMPETvBCiDqGP8epFMMGYYfI
bRXPkTj0qJ+AZ4gr/FGgmpKdO05+8CR1wS88RNUKIdSTIJfg5kpBZQG1KavWyglRhweNogmS5yNd
ZmOXTX8YgEuIrTgD73316m6M3W71RC9oukKmcLhv5/6w4lWBDuIuJD0ABbhuDs63Mkt6HcoR98p8
cZdBCaz6Xi1q11mWR+ynt+ZBsRYXYR2fRXuW/j2mhO1u1+tm2Rl6ZDWjjWQwkNkBKs19gNYrMQ0f
RIXtKOv0Jiq0kCCrQIEWZxYOs366MYRv0H9W8hQeSXj237P7egEWvMrclOF4zMw4hiFxJCPWKdac
VnzSBb5/oVoyFtoHIgsH3JRByILcgetr8MxDJVrZ+P0D+2OFMT6/kdjx1hEWPfgOyEQ3oQstb3Il
vKgq6m4Rh46KI3Ov84jV4C1eWk/MfRcwJPbqcEtb1ImGvhwVz1lPmoSbmcAcWl9dnEs9oSdChLpb
xuWvi9X731RHgDiE2Y7eHxWJpBg+xV31oQJq9heOHqM0Rrr/MhLJPQ4v4s8Sr4R2gp7srO3LUmIx
ZDT2bLqfGdSrf4Zu16CjMIOasrMlgSNvySzxJIi17l1i5TgibVlGCRfUKcLLssnAcBZ4JPDIyExZ
U+1gmZ/eiIvzakvuQ+DYL09/3AQ0NRRmNKzI7FoYXf019qb5RQw+zQAt/96J3/S6KP5IkPwpGsGN
wGo7oQMmAkVWfPcGRMERBX1eSBW4ZIpRBGi0/k+8cccvSYDBN9r1rVIMhlf0/ie0POhWY0KOQGAN
abR5CHk8F+65oELVZXdOSVvQUz3J0mfcdWNHVFDGkjAb+q6hZqyh532jgDlUFd5J10b1qEw6gXGm
FfvE66CoI5KEMiT0R0zs7S/LU68hRW71QwgQz+RE7F2GH9OVJIBrl2wwnmDDNUs0APJ/80AUbKtL
ksCi7crKreEFh41OLcT4tnWWELXsquPONhGtJGe5MXtFGmF883U68m3rjocSSo5bNpieUgLwoXaW
661FfqVcYVL6rlmqU48Tt8nBqHoWdtf3Ew4sEYvKN4uytK2m84MFjN93/foi1yLkw5bjZT6GyRYp
2+8+elqcVaIu3kTw3V64FC5EPVKOt1usQYoFKA/H6XYTN9VXBKeX+Ez30iOuJmLJki369Jv71QZA
UFrBwQJQUmYC/FeWHKYbtyqfZVdPwGzFwGUG0QdZEfy0Qe6hAcL15EhhiJ4fgHuMKpQ9YrZxJCfP
C8ww7OaTQY1o0lj+85M7AtmmWocUMBtY8ePaaV6U+EpReIfzjACfs84A1LBR8MvZJ7q6VygUUxMG
dKKcqVUrX4+sW5Voay7xk5OdZFIqQVbBlzWaIpHmM5QPls9/m+MhQES96yOT8C2u90MFakL+HRcg
h3ui9FY1kSwZKuYdnLs7XWNYHG41BquQMjqm+0pzeVjJ5saWuT4DAcGP9ai/we0E3PszSrY0OvSH
vEalMzV0VBsvb5IIQdLCk+sQw/dyN5D9OdH4ziOopIzmeV5YOiAIJsPtNEMXH+vUuh+4tacP8ICk
wDlqpwMwmix+hVs1R4VHVpH7Zr1Pxju+USMm7ZS4qb7pNLRGti85rZ+/He4PH8BpAlQfPApOz2oO
bxvAwsEp7/KqY+p/+AxjwcIshAtF6UEkgMQMnwQkC0McJdhSzSnaR+YmrcyToWtghePJO1kGPZbX
M3MuiA2Pc6ucEPHAhdIvY/00OrbYR+atbxaJw4ItQI4NBiUHuoyhWgFVq6rHomnU1VBULnTBEle2
2o0Ir6tOVmjD6w4PteiIfa6zVmnYDvfz7RaO/tfX3/wScI4U1FwAjiMT6dycwDhssWKG2SahweOY
P/mwtzR2VLdCbA0AJP0r3XlAJLZ3ZtE+bdfa0wqbb5T2WV3vlk1AAdZoVECaugZJzomm8MxWzOhF
XkB64MhI3KVJ9TZ766mxhpqBnW/Batn1HkZLJDzFZyigsVCqhrVIxZ/u4JGxAImyVPbHzkfudiEi
ybaZlLIQwCt0STKtP8FzbahiHcztgwLXzSObLBpwg+n9u2Wx3Fcvcux7IH4/0QKzQ7lcf38pFO92
8qlVU0g99BIjrh16MO8a8EgRgAHAFPtF2lfEyM9La6c49bq9tDT9j1ZgntCBr1fpZJ3KCfXKyflO
zM4hGN9FqCH0DFrSb5MgBgcqiMysui4sBfFlNaYVqaxNuChN6z/LfRQ8SHlOj0d48B8FNHJhMos3
TvCjRLah8CE8TjwQeo+iHOgNgaxeL5JbGLscIctRcMrPJzbOQoMqj3T/6JBhFoyNiXzbOoyV4pW5
TMmHYVlnCYjQCpiI5rzGHwM3RevFH+l3Aqdnk/6RBEym2+T1v7/D1SeQYVVUJvlAZRSaVsJlU0cc
no/bIA4e3nkIKVKnoejqB3BGbYA1x5ojfH/wMx5jlQPib7WKyj0ndhYPjHOkPtumOhx5GjRkCr4x
Wb4V9L3OhuhN3z/6kW+PExVuUbpzhd5w0LqUbf7+dxOzN3iR5Pz3rGnEI2cTwdAcpk3P3d1OgsoK
l0xCdW2JWWU0ijIDSDzfx9MgEPiXkvqyBd0m2hRV4b+KaFmRBBHv20+z79J/V+HvkohM1WvOrgmj
djew1YhNp9VZB/FTS+KF5RUntrG2Om2O1PLySpre4bg7uq3JD2E6tDv7UeLH4HXG5ifp+IJTpdQ2
G70N7SZJPfoGANZOfZODQLcg4vIcIdFkmKn8R9Ljzc76Cl7TQg9d7KHZQbvUINQ+nklTHiQPUV8E
k8Z+/KBg5dA1IYHdbOB6ggiQ4wZkpVqtUiXJFUX5agNSYk/Ae+J7rF6zaBzQhl/rLVretw62hLTO
d74zJlSvztQ3b4lFis0YgMXcAFnT+OOP2ZvYbG1EY5GRmBoaSonYfR57SluUgkGsZzQROOyQbMEJ
EFF2C2Z+Ci4vJEgx0ISIXpMe10UzAqwIPKFA5y0+81mDLEa1rvtHT8A9EezO52q3dZ761rVtfMOe
oTXj1SHyIHDPIjNOGXXY1xDOTq35BPEnytz8tqx6TPKxZKV36IpcKOwcR9wy4Y/tFond9e5OLFnV
L06scv6KaBWggvOcJhawVnbJf1Ivu7cKCq/PTpEqyd4fNBO1I46pVakyW+yhe456tPHKMbAAkCwo
vUXpb/q6CfmaSgq5DVGKRBfo4F5j605iRElgDERoeeGjWS7CgCyrHdhbnn+IOA1i2ylw1dmMlLDe
U+wJgpCJ63hPF9ODZZgZHQMy5rwt9sWtxtFLK6pa4M0syIYhpg7mb41Ica7GQswxZ/7qjkmKxprh
jNH+OI3iOMInmGG4PqCfh1e78sOkPCiWnS/ksuIyDLNvuxBc6CxVT8I34rfmz9scO8SaKSU+5+LB
mOGUxMyQESWs3ts6rR4xBina4Nal34peDUYfDWXGyHINthnIBps7D81q33KWV68qWDtFOTkWN04e
OwTW4T7WoFTj4rSYhgj7ZqhOl+XBB064ilXMSs7kxxWI0TXi9Qwf/SlUh8wy20GbfK5BKNElr8Mj
LVoEkiEHUAO61X4AlB81lV9H5u5/7QRYCky9eGk8P29pad5IedQQrWKXCdQsVEdXTeH/MxpCgMBR
j8dCF+9uFC+HCOd5qdXP3ufjDrjYrWqcBPsXAAeZLedMQ8/a3W+vmaLInl1tebUVxhTZFNm7cHnQ
MLTEONvAv1xzNIAFJl5f/LqQ8Mgiypjo/F/9gmjkatLYm3l4Bmg7sB9PB9aDdh1tnWucjgrDaccA
GErqMLu50+5YnO6Vl03gpaxSc2QPHM10qBfbmKT2agqIZgVc9pETqQheylRkXLt0Ckas98ZIhRMA
8hFDN+e4oW5Y6NBc0aaZNSEIF0ptBSjnD3C/6PJLAgWxJPLh65nOOFUW9t3FMAHQg2VQ9+6kVjTX
9W+fBYtBazk44cW3B3I+o9x3AMNn/joEGQr3e+alXjSJ6kUGokjSDeVNTXtunAvXqIruZHLfapB+
otv/u5QWkSnff+qveWv3ABamYqgTmpny87oa9I3M5oOrceiUmnT8Aaez8/HI64MyVk7BPrrOhf9s
1dqk1ScbFh+4jNKhexk7Hks9DD9AZzH4COAICthmEy8HPxijOOxRka6xAc+uPi4iYJUEMZArCk1O
eDJnSMbTN20RcH/9nOg1OrQXwndNv03FDu/0xVIqUgsLeRlRLURXHPAJDE9q7v0pNV72HkHfK07U
3hTqbD9Slocw+/IKXjGKZbnOn2n1XUnVB2qBxQzvxdT+g38fxEbnr2eFB6I09Am3XmGlUJTo3R0e
oe6juzsYZ0LehepTFNsWaPZdZUTj6Qj84SqpGxtDDlsaJGqToK/qq8RqBgA5351hKIRdbWKnLmol
uywWPv1d617juINDFavezfLsoQyCIj5TTDliy8+EU0tkVNvGha4T1Lo0UAsZXxO1ECPJBqpJZuy9
1vgGPSNuwqSIqkTSVd8mPn4h8NxzwMGBaoKGfQHJqTArSxstZxoD2MfNG3E6B66V8RFLxn80Mcx5
D0sLly5+Z/WsA3OtfzBPsqu6SgCXBbNnHN9im12YJKZr/URvM4cAZgrfhOgaf2T36Aqt1ojzdArd
7recga5PNr8nsx9TQfkMsoNxjyCZGURy7II96N+J7/O6NQNTGq6i3Y0gdliTF1EzoXPbh78aFwXz
WK9q2X4siBK8xKPXDUPz9ZITGi351Fst3grwZIgaUF8FwJ/ZdRP3Ds+xKfrWYyo8P8lHy/pVDe6R
cmsSqdNKXi29mIKB3KxHqXhBuCT3xY4+QiAsUqKkY9IT7U03SL9NyYb+y+EJL1EwEnNdpvfCfSsH
vH/BcuhtLV05D6w4GQbq3mAt/vjxIc1J064vmwzRBo8mrEuuFWFm5E2+l96gRusau4U7mBaozJ4m
vNg5jEaP7C3Y2p/PXUmL+LZLWqbXR2kRozDtFiOH08+Cyv0o0LSe6SwrNyGQBbuuffd/pfAHjSrN
vWWwPdIhosV3/BsINbpzY86e0I1bEfOjlbQj6Yy8tI/1qJIFT2sZGVcNk6PMfLrKA6zktJf3gV10
zJdPubLnY1zyj4Ge+erAZH8R/k7pcsOXGgRe/Vcic+gplwN9YIZVi4VD7vflOLODWXneeV8raNMa
50b+GazlAS23n4WC/yEruwpKVzPhWTd+GPgJzbk1XYT7RZjDS71tXYG+p2QgReOWQlC4pSliI7xH
vMTYxtC1Z6eT78E8YuTjr/MVJPPdvha4CcQmZeTyLiVVjTsJwK5EbUsW59LDqLOAVBFw8OmnFrUZ
rimp4WvWaE/kQuAHQ0TYqQYe67elnOXtdP2joLrCEa6Kx3APBSBlPqReR+7NUcI2xA8FIJkisLLQ
SOh0KkpN0cNZgMmXhDn22yUNrDtWBGkrCTnMuuHiAwefRkCf5wbffwgfGjJEkSByxYBG1PHYaBub
ac4TnreI+oUzWW2h3//qp65/GuRQHCL4MWRGduT/vdyqKnV/7mSMIMdh9ZYvFzlC3pio6B+Q/up2
bZPTfQInyB43r/Y5puo0R8z80IwQG5X7aGrTP+ruN4lWiCyqDf7yRp/XmaqIvZNK2k5+tDzgPUAf
1VQjwe9QYCTwvCILpi3gy5NqpkvuruoRPqbZMj54O20TheDXNo/TQ5K00aUF8MxpcbVs4CGsFQNq
bpC2cGqwnozxVKOEWHx/DizHLUkrzg1Ac9rDWu58F9BB9Vs+oQbFe1i+PPFn6QICzDHPQJVeQh49
90OppsLPDmj+ZNgfRbfhfhDNQNVqkVTpFcjTJSELwqFEIor9J7WkdYYPpLyUYvN6CE+DsqemO5vn
en3YVAMw3BBIuSBMR7acP8yvbkROxrylXyBCa94v8Julhd6Dx2fF23GXfLgnpGvSySspTRigzRAs
5hZSh+BvtqoD6gPKUdTfk4gBCadzHzhbRG6xrvTUwX8l+zG1PkFi3JqR2+yD3fckP4Rk5yrAxK+d
/W/0s6aN08+6hamOSaLwLgK3tZRhVa9iG4ocQ2ebaj6ojYTCcUazqZis3UTQFZJn4sM2AFGV3gTX
HRE8t5F8QfV+QGkqLA5k0y1TsEaV09+heNFkeXBVK/aI+yLCGweatVqbGMsFtmaZEUBbwGVL+9H2
er+j0KesA7OxwvUoouUIdDzPPpmpAqIz/3N2k6VxGu7rLc7Z4vUnKuZCJxJh5j3grFbknKydJSbi
3JyFyqQALXK82tccWYKnC7fxezn7iVsP0iyjYGyCOkQkjPBJMpdj+hytUANEPUl7C0fDBRcRIPLl
hwOE/gtSobmy/i/DwvPek+II5IdCZeILnRstQH2/+9N4+yvsIud7ZayPd6dVeWWYh0mq8G9h1nnn
GIgF5jAjbc4VbgbmnBmPeGIQLnzO178OIY9hpmKptu6qwgTZLKSTOPonkD9gwpndpYYnAeUBVEMv
GAaMBV7DrLd+sQJ9fK3QNYFWIyyI2HqnfxnS29nQaMg8N8LN9aNnmxVaMqGokHrhT3Pu0ixcEPbh
rPjWO2DRZ074/Mx8HWoLoYTHVjUbW6CL7z1E1yQQ5QYEXTsBa7/4fNxEea2sDyiVlxZ7mGL3F8yW
/Vm8THMRsIHXIdejKPOFNOi+KK0xYhvlM3QwpsMvLFuGuQlQpGNQvxg/yLnjMCM8QgUAekRr2FTF
P311WHcZmzBqeZrUa3xLVRB+EC/LdYnv1F02Wm6NBa9kwoYx+V5XLq95+2s/1FwpuFAzvxUy8W2e
gSLq0nOoTQvL6q/IgBnrXwPDIROkayrdvBohT/KrY9jCzcgwD/0VObdH0IF5OY7Zyk54YurnGXbu
faTdXbsUky/bDJvbxx2F+3mYjJNu+dXlUgQj4lb+X0ZKPJP44VSgtMh8Tw/5nXmDadu36B/M9Xuj
LY+X2mpwl60GyGvHtCtXqFzsMONxJikL+tIFKax4EcTGWkuJbNRGekGJIUh94Je3nNkhA5Q/zykf
9+zlK1Fj2/X6lmf6hkv1Pr/SNTrhdYhaqo9oOvivzPVdNwJbGr/kFiEm/BEZaiueBsSPK0wMJ98t
BU9nxwUnao4Q8RxxmtL55XUjujv+dx35KxGG2HXfFMyiXm8zk+iqWXfwIaXX6cGHGF1Qw5hIfvME
fUwXrIwVZrw6y5Tdt4OrG2ZLci9Yraj9UW0ZM1DpkYci9e7EvP6JKtR/1Mb+RcLewybD8+wmgbCQ
xz60mYfuZ/KDb4ExAMlMgCGkBORJBZS3VdjaeVCvpqIAaTOvmB1B+ANi2ILiIErQc75bAV2v9k4x
WjgJIpUuhUJOUIy9qH27AXnl0O7qbzFNYhwmzqEuKa4v7A9DDEJljVSfnGMsGblV2Ptf4iW3OekL
98CtNMNpdU/a5Yk+pwJYUUMOrBEMuJyUKtRTNtEtWVOxTHVXT2ToIiBwsBNOthKUaJFofeXSitnJ
9PX16zvzYMJv9Y1FFtK+wYBaag35WOfANMPdb5S2uLNW4Anb7nf3/4Or51OkhNqi4Qo8TAfrG0CQ
cGIV9U4Y3O686K2SDJGHs9C8cu2AHtgVagmG9FfM44TxM5O40meQB2UCT2sqjttNjpwv1EA+Kolb
k+rdeQ9olvSzZhKNPzllgSBMbI3V7Q1HtsI8oV2CTx3FEOy2b1ExWcEn6j97X7DmcKI9VvT++wcJ
/f5sbGUipjOHUOuNGSP/6kdHZ7m9ACaKmE9m7BjINphv11DL+JZyXJRRqcmphCArSl62d2TaPLYY
l7iF0WUA2Yv6LwbLrz60mYVXZJddvPHwL+ccg0WO6iMC03xmi2rwUT0nAdj3RZ1jP70EDwEVndZ8
eLBRdialojChXjINBRfR2O2Gnx+J05cQiDLEl+4/R2Ae8aK3DWpaeUAsCmVWjLYdRbHdmGi2B7jy
hz6IyL9omEtKkPqK4SKCtYTMkezyc7uXsr7oA2yEGEliUqLtb4x3Q8r6Y7iUyvWuAROa8vI+iLxj
n6H/15MQFH5EfLgdjTuz/dpbClFLxx1WTC6lFYiL5aXGOUZcbxumgXEmM+nG1NUvc7B1081rCFWt
j6+JODChzENfnLJT4izyYltWC4pMucYh2iQXhECC59KZF6GcyyjCs2bZuriEG+dB+eL75NXbcJUF
FogyY6YoQF63YA4o6273JJMzCMVxUOVYgbTZnH4YoMSdTOxdaTulAyvBydODSAYMZyfUTYRj2f8E
OMQvGKa9upz9/tRvweshXIFmtMrQgxw8DGDJlIIhY1F75cYmXxRts8IjlB0++8p7Fd53CiUYsV+W
vGO0s4madiiij11+vXDg8GwDE271UI7IfvlyOMq4/vofNfkqmhk69i1eUArsNyS9U/EY4tzBTmTQ
xZ4LaXyIQKARAgV15BJl+e9hdfh46N05iaj7NZg/YblUDDElVJvfgXftCzw8spkIIjXpsoLLMeyp
CUoxUk1HxnL4XWRlSv5xoy2kVRB55s0LFjmH0qecZ1rVXSNOAl3MiW01j/Vb53NnKLCfZsTKDbWW
OFxYjEGmFkfg5SQOLUUdQ1hGGS9pjYkAaIUeKkY4bMod4P0IgrKCBfyI1LuHH46L3nDhS+H4nD7k
/hkga/5Hsu4zQ7AsAQ+ZYB+0Y4TAC2Y5w9+bLl+nm4J9DJWJEd7gcC9U9MCnOrB7GPV6VJ2VGHW8
n7tf0HJuqPR4yO54G2zFR2izzy34P6rf1h7xAdXu+0+IFS6iVd5u+08ph2TotmppouiKdat6mW1x
q1vtUig2VwwZWYTZsVcf8YTDJxX7JlW6H6YoCY+eUz6EaNMY37HJRoWhYlsgrl42pqxF+Lji8rzX
oiyN6zswAFcUlclLFgbQNnDbDOEDmPp4TsIPNRAdHrgpZtMFJRFBfmR3R6lRx5K45EsT1Lh6Stb/
16jhdjfchZLJwnCyA9EHS0hxRGXY9o1PsomPVYkDVIO4aO6zpYy4jfEHlp/eofCIVLBZnyUHm0qc
/b/gWus1+zOXi1oOIqsFNPveJ7MXmrrCyFgZGgdUJbUIv7zn2gDOo4PWA/l+s9Q47SM7bvHVP8RP
vjmLrDWETf5ojGJ3geTAVUBBaXkcCaB1LdX6Mr2U68VVkcnf6DbPvoDLO9quIamQF+gZ+0mDmZl2
R+dS2wLU82SZ+3kwJOO66hM28qnf4g6yxJHM6819Z7+DSdZNg81gmlUf4ncgEn685H9Sdpngll33
Ljw1C4AJ465Zkn2Uck054BV44gdsoITc1nXg8XT0jSYMVTB40DLBK8h86AlQ+ircDlx34VRIr5Ts
VGfmXUae3CwZBs4zlmkhqVqNXzZ6VkucGq7fGxIkSbHuZ8Ff/Aoc2FKh6Cavb3DuthaaqkE/E0TP
gkpA7MtfpsWmY3yvGcJH73VEx+8K66/Vp8amvWyG4gTyJpnAUFeOG/5tghG6xJdal4f9BauGXyOc
fyzY1p7+hK8SywZIzfeSnr36pZ/ZNsdF1tNHdCG5B9l5FLHGkYpjzbdYoBtJKCWaA5tRQsUU57S0
ftWhoFnY2XSVVOA7Di42lkl8h/WCqG5tqM53TNGUr2a6tUYPb3scGha2XcCMyV9sBnuHIg/g9g9b
KnYIJTBWP8eEVZf9fpW3f1LTH7wA24HDMK77gbzqNOfuoat7Y56BjVlB46Us6FvX+hwRY7pWAXln
4GV+DAQtuCf9mGly5mkuOa1X7l6/lZ/U/npUxPPS/8IXw8ZgyuKq3XxT1/U6pgunLXnVWa86e5oq
ECg1HeGvo4I//DNWa4wNz6n48TrMy+vyJoIvfb6qu3BcWHONZtiNo2IKIruaPmcZ9FwEAXUdZRhi
nr4eN0cfkKjlk0DX3ShMQDcxJNU97t/QoBSwFHseCzdwKyvc3DY5S9UngbHV0ashucDQwtJhMye8
yoB7UiFDb1nuFGshEBpzO+QcJsX1Ohw8PMFJ9MKQymaB3lQ6Kaf+6jl29Osy0Lfo2orjl+TRUNky
mTKda5AdCPbQTNhWaL7fExAYeUFSOGk8z1Bf5cbWHAFnvag8pNy1Zbpi61TS9wFLoO7WSX/qx/6r
AEAwU0rOt83UMFEiY5Ve0zB2qAkBAAFUmAUNnT0DC1wpsSaDQEDFjJFAQEFmdAdSmlvyOVbc4MDv
Qf1PxqoFkw4XcWoznezx42Zy7GLPhRxCfqId5HS2I9wl0RiIeaW+T+G4cmR1QNKXb7aO6Uijbisr
4cYuN6WNoYf97nsr1JYDPJzwsEd4gnCUe5RYVcBcMLiY7rGg5e1Pkrc9h/uHYQQjZbRvlzaBjZll
uwj+8fesl5PSFM3t2BNhYfeKPwEmAXlCc2l6sG2BZv8r2aQ/32MTkiArs7kYpgtz5ZioEDcVCsIq
/A/wKy+tIgHubD/w10AEKfep5nMZVJHtvBVMAB1jMEs73Wgrqt1xW5sXpde8KynjJyy9AibRMtcH
oMaOt3zCeZWHvwaR0cQTipjMXIZFIhtKtPWpPSZpbWQDiV131xHnljDUyG5P/b6OUlyU2Z8Ea0YS
V75sAjK+Z8gPoDn/SlUesgoqG+gL9ruFVkd3hAA9RdX41XL0TJjiLRCZ7Gdi+mPGvj+MJtP+LUkN
UvwbN+hEEKpmK0T7hW5KhmtTz74miiaEM/12tluiT0Bjr6AXgyVnvM3TbWnMRNHQ3UB0aMueNPfZ
mrM0TPrvrPIV0f/EwDMBt3Q+iHJJkjsODJQQLbNwcUG07HBAxenM6smPUYsekbWDSwU6M/IFSF1D
HCjpgqx1Va4WbhrRNLvAJ8F6XdgArTBFB5bnZSnW6GOEAtF954S5uz/RflwxRfgw9uSRJ7FTbv0v
c++TFkToytWQNgA9r53E8F7KzYIC3ii6/WJHe2d+ObmYnP4ro6LWY5bJK/XxUGf7muPxgXJ3B0iv
fwd3z0gxKm/NqeVfDYzxqx2DH2qQxfB7EwOlm06+kTGZbpnjiWCdLOOppFQfLA1i/0t6w8KMnPXE
Y9op8iaUGlUT6ReyrmWNsY0Z3qXcJ9VpyJ9fPWZydIU8pYI7Rh0iOxeZv1TUjREpkFmj4mc+KG0p
s69/C7qhTNde49xsD88npkVMsKhA/ZLH530shepTNxMAHwawoZ3fM6HzCvc6kRGv7/sqRyjOV39z
toJUDxLFWM/slxIx672ge37EtNWjWIqq85gsnx5EJSL17UfSdbYQFQfUlx3mrButFojWYBGVlk2/
/Kqp2CvW1DwCaKw6inVOkxyvrLWVrV5nJ9q605rUml/oGJ410j5rQ7jbf12jy2Q0+Cz+6CI5KREi
xH/2vO+mkFoVUxXlwW549rl6Ljgg4GboXYECY3oPqk0wK+WW9Hj6mLOe3ZktcnHt1iW2+J3Fyh+G
FDLSdDwwBHe3QRAJwiOCA4YdqSRqF8EbsCdjukLv6/D8Rs0diMn+ThcM63BwB5zg9Pu4Lm0tOctG
8/8FKXu5oCmMuC/OGU2gkgdJRnz+XyxxIyCPVmx/Yz4XGdOosAHi+H/PPkY4MPBHcg/eQe2gT4Uw
8Wo3GPWhhSmwMr+2PhYZyFq5xBbDIRfENOPzfBzWT7DzAVgwiVQfBShvyUolPkuGDX92bZhCpFvk
7G7XiFVsUrWZS4nV+bf+bz2G4zixOI9vMAywgAgh1XqlNTsQpec4i/oIh9C2X0iGe3M9mzeRXqYR
vItUIU/cN4siwTKQ3DAfw4PiFSwqCa1QzARToUpUKjPUfjLPa+UG73uNkv7OCNJp/8F5+Y1K9TSn
9rW1RKo/m6OhDLB+fXacic9AiS07c6u8+X4XerM904vzox2y55xn4t3CsxjyeFYhAPk90y0085LA
FmzlkB8r6UVtNVyH8wtvYnrAMdrh8ONLMcpvfc71ZJ20hmayg7nfxV5hGnRfaZclHVy8QSAu5qCL
0uWaH4redSA9ReTKfvvUL6K5ST6W4awMd+sFyAgaEh15g9HuzXbWTkuW+FcCNZyPWgF3jRlazUnd
0XCUkTeZ/TZWOWXjRF7enk++IQ4f05mpsjuod9Py1ympcNlxQm0+y9ARMy162Ote7WO3GpLyoSqL
pmPQg5wGmHmNgZDeh/SLF33BzR7SqorJIaWus8euQpbbUTqMz7DRzaYIqZ9x1w8lZ/nSobD2fwaD
9lWgIcp5baWnHpLw6evZQjJpH5aFLvbv9tNVJd5CdY+kwpu0/KUoMmrCunlyE+EDqMPVYb62/mYi
faf8irCByAHUBYQ6DLJgxt6L5Ttc+4A9dPvCvXHzSvJZz7mXepJXhra5kPMHBI4BIQ+42V/nGoiG
x/vlSLAFNkFAFevJAdWBBM595BERXL7RsyuiYDx83PggAH9akMsuWXCdTKyBRpsDRF6iq8VKgSJT
R/DHPs8Dm+vCGJUfFxe4KdHyBXxfooyolBPvh9w+DfxwkOJqQoywhPan2zDhRaSP39M4a2K4huvs
X2gUBnzRq4YU7DDFIn2/ypZgGn3H+CvUqFNHHo+XCWoNsJY89KLk/9Y2mp20XXpL2UybI68+W4as
D1DnOvmoWVWQgE8J2pWJcwkGI0wwUQsjRB/s48+kaHTQLJcBDCQLLr1eVe83ArWcu3xFjvWCshJG
14qiCtntoTi6Gt/o2GCqg9ye4t6kIjhcpu3deWf+R/exF3YtwsQzf2oTTe4ZcBD7gvad8PRhVPUa
Fh1pc+21Gp/rRdzxZYV4Jxm5pPf7TBk4L+rGYCRVCZdUIpvBtyjrBi7iPhhKIKu5VU0FGC1lWm4M
fN3RKumFw1kDyjfsPlyBaJKg4Ix2fs2xtieq8W5QoRzoM+tRb0pXNtledYVrZ0jgp89i6YPLJR9r
hWalF3JZkMXhF1ao6z45IcC00pnXZrQzB95/NQaSijwm98yyTG5/TowPEy3W8Zw53SEpABUvQywW
pqgE3zMW3jjMi73ikLKeC9UgDz921pHXU1B9ppmn6DUPfS9eGbTxhfHrML6W4bBlEXsETzLPhhe9
Sey7GwsBP0ABabY8DnLpRDoz6aWPII4/Or8Sq7JGuSJLB9YWUtep39c/GeC8bt2sucxt6mgtwqVb
Q12Ipmt6chwaIBlDo7C3CmHXOPAmROPc8T39xNvp6/kcOLiTrW91Ni/LkJiTTum6dsM5tbmVEupb
f4HOzeDmLhVBs7l71W1+2agBepisJZD4Miz0I5BP8D8Nq4PTqrU782MqUSI7sYRmd4+X69LMPbqk
IqJf3Jder5hwSax4qKV5OG5Zz8zE+QRRct614lJ0DqzIoO/ueijJ0GMyesOjoW3nCyMCvA5WpdXs
2uE1Ui+/3JjJLekzyZ55KlDVw1y05LmjnMChOJ28lCOvJMTbHTeQind6acNnRmvWjVYukGcvAxHx
unbw8Dq+ieKgS2MDlGxO5iFXvluQdhEm1Cm5MW2bv2pyZn1LFA1g2UryB+pwQOPETIYpFL27Kj+s
buqX6lDItn72RrKQLdfVYStQ32E12HJRhiszSTqAM8ZpNcrP6Afn2/pNOqPmT+QFzmCa6bf3PvsE
rdsMHRX9GXGdOgriTPlg3hixESGwRzNzTHbWOTkH9RTeSham7JoZXxrddSUYSfdPpJFe00TGMNRP
RbNWnwFd9R5mtC1D8DTIOY1FiXGVrGESQ4CxUzlXe3aJbO0/zcVkKcHwW674VJVWJZc0sIRt4Vig
0xYXQ3Pw5Mpua9iEMlIGo7JrnZMHg8UdHKBcj/C2YimEwVdel4CeJxRWsZTjRKbSqdZch8nPE+wC
pVAnykqjCZdxmWxEpG+ijW9vIgbFodHWj3P/N5wKtvwErpVE2lOQaB7V+sgQ53H477FcGDbNY4WR
FOi/YORJ0GiYnW7+CnH6JKbj45t5qH+w/ZfOCLjL6pxApFpOdqjKSzb1iJ9592XpRLlTKz19pWu/
iukz0M8rKhnQ2QzGr+nW/dDWEThH8qejV7H4IATwsp5eUonRiNNqu1SUS48zH3+pQw3MnsGs68Gm
gSn2BXFXp2LC2tNQmQOU0bu1IGWGueFKlHUs//UB1GYnIjP+9tekZ/4Z/uStRFlkxIAvP5RUieg1
TUozL/t2lixhrt8OHBKsoac1nhfBCAwBsK3NXOZsnDL624s3pVMZRdmGMIb4yIMM7i4J/tusOU97
XA75SqSUWTSMgNyk+3355FXh1E0HH4TDa2ivCnvXsxIENFfDjn77B5XamYG1XBRLYAXZLBBODj+/
om5jH+ak1X4modu/Fdqb8N/TYvuFSZlgpXkrL8CyRuH/BgcuBPNbFKeTv8MGA7S9yDV00ACvip1k
QMAuiCMa95qFAeR5gfI7dmC5dB7724XHkTyfTY7CpU/uvDQB8Zo/Ue2jRPhm/+x2lbA4ZVAWiS2Z
MArzU/ynblz/ecwc2Y/G6xMt5pIrlTtjduHb2rh3odU7g2Z0pMHxxrj3mYOD7PgzNoWX/0ZMWyyh
CIzAXiFXlBAQf8U/ugRCkmpHrpABvo20BjWoif1UauUj/3utLiIz/LV7qexNoqUTLAZcJx3ohiku
0n+oicTbDHBdmTlVVa4iekQwA5uNr+yLNyUucr3Kn4HUZpqhD3yjGku1rGJeuplDCy/G8mACiyHK
YRCkSTSVwIcyx4hVNcuEtzwiRaQ7eCnkKc8JULDdomdDwYhxxGgVO+iOFKXssagVsZoMpr7JNLh1
a8g9ix3UBgkuqSSJmVc2nf7atFUTrTXSrye7S+EMtaDmeKx7ZjVdv++RFZ2d81R+/kWQ65RqzhfL
h5kIr0rzRHAehwmX4ddWDMKqNuMh7xVxoP1X/6jiOeHm/CQzrgwgDzURxVESTXJgBhMRMWz47bTG
hqqiuOnyPt5eoaoNnYlIgsneLB0nORiDkYf2MOyrHytn08+14a8QXI4cUHW7ElFOMIorbDxMmbi2
yalf/9/GyCNswHzODe3VK8sLEAVeoJTkgBXjKFq/CTcn7Szz5LMSzXGos/qMa00F4KDBJOXMW+xe
lSDYKQq6dCef1QM/8ayBQGdgpUJ95gYbZyUwoMuMeKN4ITwzBYvdwPTR/+kNCYc1E8MBMgkmiYG5
Xzthe99nVLDUv3RsIqloHsJlbCMHxb8bTYgOpg2Fu63OoY1ZWiYmGoUbr8CnfUrBM6PmkFxpu+OY
2NdxKGA5umrdOBX4JJ7/fMJe/I2v/n1Z9tRpqA5iuNcnchSggUxM/g0k4OjS9QGRBIceZ88pCDfD
BHiIIl2snOGn+XM917BCVv32Mxhp+fh5Ibptsfg15hi+OtbrWwnBZOwkOKuV/IP1WWjoruiUhUqr
uAIFz5OS1vAG3572JCOsTRwOVV/pfAQy5uj4WY6sJTs3qgJmclA1XzG/VuCiN4tRclq+LnMcJx2b
XKYcDtFkbWr2NRg3gyVtee7lOAaMRST90F7eJyOgDWzdDiIK4ir5B2PIkkckL+TpqkEECfoDhtDW
uAL0arOPpz/ex29CBSmPgcBxPY4cLzvTv4nQz7o0I00gZpHlOpbbdsGug8gK3F3iFxVq45EXKnar
WzWvvDS35YrFguzdbW3I1zaUfBMhxW5dT/KmN0k+rU9k99anW3THYVu1QnnfQbDeTmsimWbNUJvk
etRszmYyF1B4Uk77lEGggeKcSYwBiV8rH9SdORbdEKbklMIH5EibRuVOzkkpFnHKf6OduM7Zr1Kr
gVNjpXrJqHlaXEli9QztGZ/dkWiBsHjMu86DxvIUi8Ep/c+ULfpQp+RYe60dHw8W0eEV7RXTwMO6
o0KqPbCCHpGeCICYePcEzH18/M+TV82rwKz3gfbaLdzZN6X53XfbezILcIy0Qt8gjLFZw7kuFTIO
Fa0PrsnZ+WwP8SLxBuQrJsHl7DA5ViGalYKz/6N5Z+iMvfkiVvJ5VWS481ILAXBoWoscgbmRGRfi
stjR98cIUC73itiZdDkdGe5MgSuaay2LaGB/3SgzjMRAKqj1NrhfO4mEdU8Bgq1hznCNmemGRZMK
oMsIUx+DqzwJr670thurE0RhRGX++YXnHmrPl6HB7ixjWb2ZHynRf4ho+ISRWP9UKXPmwxeyer4p
tIumPi8JsChjE5wDDBUQp+2nS8e12BY5swYp67k8RUNgY0UuSdAHyq1Htb0ZNuJceh8aiEa7naJK
53KTwc+Dwo+ZxAYFabugF3pB1WE84Kz2rG395XvXUO0+A+55Ps6Qb8THLjFjRTPLW397giH4pk00
jFnKkgxnH04pjT+lT+c1hKKrNH+fjnZJS119SkTxcikCJaaEF5rUoI7LRROZRdvgNGxE7VytRStl
FyIkBKn5yosJSyj/t/A24oubFbbcR95xjqlaBqWw/HAkrHl6I/qeZZ7urMm9S26Mp5n1Ak6SQbhy
r5S4MVVldb6DnsUQ2H5V8HCYpllhgcds3VxNjYNPsJN3R1mRAi1yuGmKx2sc8b22tel1BpchdeEQ
mieAx8iWee9vdYxtugTf+PHks9qmpiZN3yuYZ84QI1r5tfh7O/22/SPlIyIHPIMrCuVR467y4oEA
HzHpTCQL6CitTD+oGzzI2rmaDUcI2Nyoy7FH9Typcek4RwtukXE8DZn673relKKE99IQoCOD0Opi
QdfwyJEOQ1WsLmH/va4lZqMV4Q+PPWU4XPmasn9doCPxhUAI/pATHjO5i2Gi+EQmZWKX41cgjqEp
X5QrdXdHfpB++kr+1O/iJrOpSG4tMo6exDsVAwOHdPrw29U3xxSrrcWbKz2Bb2/QVmq15sYjSUVt
J3dHL08P/qCFFdswoI98+gxWewjhl3rfKC4XUJlLcSxdBTVLaMmFnSIJcUvOjziYvyGdVioJvwEf
ib+TH7xECRq4JLA+GxoUungjrL8FQfk4Tl5kK/dM4PG+obFm07k9GseN6JDWSxfCiZQcJjjR7ZhW
w81fWTcXQyiqvLWgy16LiT04cTsflj0In1lySUB/0tEYOh9VfNDWkSAalFX4kGuhHH+R2M1Aobuy
ukZHveYES/st324AkKbrE97iXG8LTFro93WR5BDyh5jYN4TxN6ryAd4I2vFdhhMsaufCUglLHJUa
9TBthIb4zcDwkmnf9g0ntVDB4SPTvK5ROtXOWQlJbTK/Zrfpual4mDjsPV6M4x3VhpSVgG1eXAwN
5vrLruQptqUYxAq7zWPDEq+IKSMPs73u9sp+uojvjKJBN5GJqM23nHoD4OHG4KsiD0nMXoDxk6re
tBnpKOenCr02VaExBa7dWlsN4Gn6HpXJZ/QoKwAa+TIFxQZKfx9COmwvGjypFN5Vje5ww64IDE4G
3mkfh1VQDgXXcLPy4PxjKnrB+fTJMlks6sDPGxQRK2NNarQU94aChlOmtgE9OJeK7U45IYByreUQ
I8h9erZ5+kEt1zg3bKPMwfUAKDW5LsqhhE6WV73zao5ySxY76R27256Mf4JJnIHb/iTt9JOAJO/y
MGLiR0NArKv4cvBpKa72KMSY4BnemQOIfUorwvADJ1qMbJgiMaHu9u85eJLM++0cI9w1DY/tVpFE
f9Ipy3lVpfwTZjSza/R/g6SQD/ZcR8gLKpo3Jmpkd62efCe6ll46JzSp3ZZBIxVOQdZxMY2sFhWo
jWvBhq9vJt0L24EjduJXRzEBB7ps3jK7sA8P8A9RxPsHqBR3bMLLIdxuH8We4TJr+YSwkS+54eNg
bh1FJczrVBp1O3umnARMIpGvVUYDS3J500xXZotzFzsCRG3DeLUhsmrC038nmdh2bsIE7aqImayN
kIAix/Z4lXNZWNA0rG7bccbSTZQZKTi3LPDrF9mlo2MUYL8++NoZZhUxIERvU7r/wHKUtqO6qsvG
4nbidA2QuYnqe99zJ2xn+gog1fUGZE+g+fqRleyfNMdFZu39VLw7nTs0zJx3B5Dy3KxeJkSmcZD2
mA1M+K7vvOHEh2rZkmczHax/jzHPlLnM2qKMKG9MIrFPJ4SumSrDC89PKtreWtxHEBUwLlGso+Wt
4H9OtaX9x571eFdbg+0p1k9e2ZGg9pmtHGtx9/Rlchz7hcFmu3zhNPyV+pOIxTHpeq9uC8a7JsKP
nGEUGIWqhjdWyNIM8AO0pOLoJ4ztzCAdXkfdimzD5jT0FwqjXCMp8+cywHYozJvdXvg26NxlYFQq
8VnOsdnGyfI8r7ST/rDFCxOdflasAtXx2eLGOS6maqwO6nC8minIBKDOgYAE1m1DDkgslMFEtFIC
ksnjwYUEultYAgJ/qaBcijZgPYnITqvJz9qoPj8CPWGN+48zjiYOCQVgwvw2EhooHf8kmalgFkkN
VVNCT3vn0dFdxa4/SbeFRjv3oRDCQsJHhMGoQjzY2j68pPhrj5Ux8TASWOc4x4PPhWUGlG1BMCmY
2rMqS/dPOhNyqU4oehrPtdApnKGwu2qRiJ+v/KozlGYaxpIzC2ZripAi09AsQZUKXRJl/DkJeBay
G5sCgIkusD53geb29pjF3BGN76g3ApefmvvWQkUqWZ8qKJ915gymQxkcN4EsOs6l11ALL2K5eI+9
CWE0Lb3qvawkUsFjXcEYlicctEqtnb11EBI439G+sX7bFrh5cv3gQsgFGfgZkg7ymsInb0lbd1x6
j7zAgT2hcHTGQ3cPWdzPhUe4NO/Xszzp06CjVYedGDIBtnH58r7wTMQKFH19RrT/15wxUaBoMd6X
1auUxAeHHXGszCjj2oOx0CboOSSRqAi6yecc4M8FlcfUiGqUT9RLUPzp3PXlrHUDb4PYFd5rUh2D
wxVF1q1V/K+UIfeDePuc2HF7GRmOxZgAnNV5ynMwlT5NMbv3Ra/rLDRAobabubquOCOu0sirwEnF
oEKLm4TWLo7png0gPpS63nUW1ZYp4zbK3TDNGSXcwNnJ09mIRlHh3S7+GYYJ9TrY7jQxZ0dfWxty
GwYrXng0YaJ5IP/LgMsHJPtq0EfsvvnHzRnVw9tTIMeoDT4Ullpl34lxUPGE15m2pIzN4OSD+AF9
ExRB5tTUeNEKfq7RYJJSxmGVluR4o1Yfr+AotaUjvKUP2kXufYnH1q+eCvORWit9u+I6k9nyElZx
Ky7qx3iO/qOkAYYoHWU/sEW3eiWFqFnRRwCsjCtVU2M61bW2xOnfn1qt+bOxmeY/fXL90e3f1JRY
41glH3L8z/QWb94zbTuEursyYOHsXKiZWWadrlJ7CEP1oxfmZ45ZT+VklZqoTwxRyo+IYHpBYDKp
QccRg1Kh14n6eWJ04aGxaLctYt7Z+Q5RtBnJyEcehm/q95kXXtK0k+Uphi62DZerl1sEYnj+Bzu9
SOeY8Tix9mRVGgIJ5UTOV73yvloILo1dsEwxcXUCk8pMqO3oXoXCmldgyaHXFDk/BpdjXDcliMyj
mzrVWHQ2RfLusGG/QUHMkjm16slGeF/nPOX/98q0iSPu7TjuKC+/zHXqOVBKempRlCbR5m5/4r+7
vKWPjmNm4JJY656gpd7KK0Z9mYbkZcNmjy1EN/VEyb+s8eW4EnDBa1kI4d7TcCuXihfbF0X/81Uj
qdIoD24H1tDtwziWhX0FOcuqNCCMtiW7McYtngHLm2aVfuGKpHGtFCDKm5VgUTO/7HcU3A0ta57e
BoP2fueqfcYCMeFm4I7ye3ucW29wV5mHq/S7rkjfr5scYa7qyILyQ16/3eyGwBvVXvlwkzh/s/uD
nFEX2UU2SI6mcynGkhEvHnY8C+JN80ZfR0Y0NtHyW7TTNCr+xDX96TzT6Cuabrrgyvg85j68kt3f
gZ5Q1BCcwtNnHK2B4VZ1a/pmVOl2deS+yDSxVHpLDNgF6r9A/eTGgkWB6MX938mBQNwbVZsJSSEl
pO+p93WtRo9KRA5+fbS7aJkozszyVi+GYhhEgqwX5CKT1IN0UAvX+sObDDuE7n82p18M7KaN5lYm
eaxwP+8iEA/3vF1lQikuz4DOqidYSv7JvvJeJOnbj9QxjNIitEuTY8RZtbWPUrK5oAoDQ/HOe/z7
qGNItHo9zeOSh4jj9frSWDZPlE+sk5x6Vqg/JSaZAWhSN8ZW32MdIL1UBMNtPQp85pJFNAhIwPIo
UaVSyid4z7VhRn2Z3s0NOsOICvC25fltRByEMKfNTYl2kGTTDmiFzpKXdm2cE4n15fsnnjYszIAg
Op9Qa6cbPNfVR3i+eLHTqZ1IwSGQ71F12/VpyZR/r49kc2ZOb3FW2XNa1sbZCqLjRFL6HBHOJ/xC
RlSneWHLnVzaNQBkwWAM34K3Gw==
`pragma protect end_protected
