// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:17 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GoudJyi7TKFKwOEb8XOVKyxoCk0BjpoJopxZqQH1iWro2KhnJ8NOgReyC+mBU9Mg
fMJ6sZIlRkm6tO8i8JSYeV/FmQC/zTYlWztNUzQ6L2q37L7TQoDZfXtUIDRfBA7R
oW5bWCE6Ms7jxiCpAorRKQNiQGEPhX09gSw8tQL3VVY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24912)
tGBIIOfGW3rfgX7s9/1ChOcTHFJ4qIbUm0AHJDdOHTBryRHvEyvLzNaiKrV51HOX
4pLRIM1WzX1GX58R47trYdDh8Cbi/cyLcL8FB/qksoVui4ABIrFzZnJvf4a9JhRT
m+3Q7Lli5LsRq9XlQPQwri7Xxu7mjuGAcgrokwZpAR6B0FBGazEu24wBsZMtoeGh
1TEz+cwpcL58vQfLfxKWHudlFYlP086eOqqchhJdfGHCuNytA+A49XXHK5BoMAlj
WB75+yRlhE0KpPZfB/d/+Ms3uUBLjssmud5jYwT7jgT6rOLMYIPFX3knNsHgsdO8
57u/5mX+FlyAAB42uSV3qc7ekgLBgpJt2fmWl8OlyzWnnP5V5727LN9nXHriZgxZ
XY/Z6ILTPMUHDEJBURLn+Ppc3DAf+swUmHFz1fT0zs8JgysDQpNU4fXxNgvxYcDC
/MJqiMtJesIyQC31pn5A5DT3Vzo/jJ8rDbHJgROg13zTG+LuA3CfdtePNj6Z59vk
tU83MC8qObM97mGY7q3TtkdsOIIgkacqGU1VP3DpP291x+Vzb1610J5c2+KkBLfI
f6VnLh0J/hcVVs75UP1jLBRU9UKnCvdk4AvSpFsuPMRqdueLuNroDC0KwWroalE9
MP24ds7tUhAIM87bJUtPsHV0AkjQKDbtqEIsjmZNLu03QHFSlBCMxAZb54qQIdvK
oW/I8+d9GxQ6lCl/hZaHGUHtYS9PLRkcU+9Vs7KQTWcs2EI2yt/ZrvYRf6Wl8qBn
TpmI7zDYwRUewTH1k59W6W7GDORV3vTE3fE32NPnpKxL8RMXqyXFE+z+i6ptPNHe
U1p8VyGSHu11J+WamlI8aeJqF+gFpKBHC4DvAjb457eBs+iaIl6kKdcGxej1KG1e
3N6dNRQORlYx7JPP/5UoSGtWN97eAP/7u55LMydAwxEPZSB3oi2j/x5jVmXz1v9e
78cBoiWamoI2SwK+oGynkbLz9Rnv42iDzYKH7e5/ogAlKpX9kG86nJdoVEVNBxr8
OYQdA8dHrNK2e2bW2rsHtuU46ir01Jhz3CA2K8rxvtqc8w0YkhrZsjBEWGhX4YsT
ALC0Kmo6siq2C141s82cxFz8EP3J7PEwyPZn29uRfVlVhbZgmy+CYxh8ZrNGVg49
WFe3eNhBf2ZVfquDxotFy/Oq8Izu1dv2dM6RDVWqxvi6t6eOW4f5dYiMC6I3skpk
vdQPA5zZ/wFPI5ZRdNcw555Trybr8pU0nc6MMgrV5mTJsavDsySh/M+9uKVJwTkr
CSSnBTCBL+RAoxZ4ja6+6Zov8IdmQbsP/CAvkREhAv1m8sAdsuHhRjmsrzGEngvh
l9e1tUukWAgsg0pxqwZQzJOFBwm3PLfFxHX1K649pNPA6+4+ZLBnHNThzVnxCD/Y
ug6/edS3RnTCmKlkH9B6T/qmw6Uu4yMpjoeTLaRhdd9zchnasqTbutZjwBBD92G0
L72U/brf91wSArj6HSBylGbCbxxZfPGSV937w0euZeThbVMuh5O2Ll04ztoe4yM6
7XZlz3j3VDMqI1X/tXUoaaEDph5Ie6l22hO+mlIE7v3TqqqFVMIPNkMB7o3Y++I+
m04dDjO04caUSe+Gf67Vvd/iPHZ3YvFEVefvcPHCLEZoVNKywMXgS23I2dr9HY0x
2/QZ+aQeAlLjWvKQYEa46yKsYLJZVn24YL8fkkPRJjnzRW9X2QFp7sSl3gX8agyi
rKiLe9lMQDycgQ9l7Kv7AhA6GflFNASFt401PJ2VQ1LsoyxLGtrq95RFG2IZlj+Y
qaSwaY6l9suX2z7smPKEZ8uvUfMZvJ6mRJY5IeZaieo2WuCABk60J4j51yuoysAc
ExuXXvgP5FsII7GeIqpSGPBf9kMcv3TURibJ3rzokefxVofPEJivG6LBIBaFxBmW
MKQzSzDhpbxgZ32MGj51BldPlp4Q0cE0AcFSRXXFwB3LuzTgH6/xwLuaA1+SKLr8
QXoVHlvKIDREG6Wqv2OTATDDFYVw5+uj7nG03oya2UoNWQ8VNpNHqsbYMdJucR3+
iA8uNOqkKb7ZiFeAuNuaXawrmTMGRtkT9nwleDNXXLE0yVlE8/7rTaKmn4up1qzL
tzLs1iojL7Ujqp5bHg2Aoxvs+szS8Fy+cXNkXXhL0M3u2A7LyLe879DBxYsdsp1e
QghpOCXmP5tKoM5HcAe83RJhazKEPxDZ373NHECICLzkkPGtdVlqdZwtciBUCQTa
/Za2hETh/xxbE1Z7W5Faq9p+mV9c6lGpb8MvzByfn1UFIaqUXeLjR5Li77+kR7Ex
Mov8KKCsilKRV+pp2FAghnm1v6a52XTZqJwcJxv4sMk5kqaOR2we65gk7HtURmFR
3bwGARBopkp4QnMjnfb4XzwTgeG63LfTVWzrK3UFnZ8iNaolxw6i4UqxQaUdABm0
phuDeZ5TmwuPlwGnk63TmtgV/RSZ7lJaEsZ8YCmZtsSmAp6wuSPptpUw7t4SnbAl
oyiuss8st4430/FjtiFMqjHMIWxk+D7ECKtrdIziFYEGE2VI/v2Kawef0Yula1T6
YdsVhA4vleNrdURRvZhDI3u7qaQnEeF9SFld13m2paYTnLaIAOMGiL5EhG3jjTrZ
xQDXuu1nOerNV5v+VPZ8XyqjMEwt9heQJ382Myo0OiffGlzHTnoCXxQ3Eb4yAMI4
w43p09xntBkJSxnTMMt2stjpH0bprWuy+ZnsFc6Mzsh/fbg4U2yHN5tm10R8fI3B
2BqyN4jwe0qbzqHHG0aCV94ZJEVQR6uiaTDGrVJTjJ7tUfvPmKtwYkFKcfmesFeT
wsis/TeLwSh2bJdTl64lv64m0oZlbI8amE/iZ9Pi65v6zam3UrKMkR/T8ZFRgD20
AsH2pkSuveZxdJ7vyQ1IodjY+I640oiwbXQimmX2hjDBLL8lrs/XF0kBTIV4oGRT
mxHknJ13C1Xe4t9quiaZQbvWNe5PDp2gYaRKgQO6Qqr4xyrI7GertJSy4lXWQz2c
7lTjXgZQanZqKat2gZ0vKQDPjLQR/QQPWJEZ4eNPtOob+KPVeGfhgrChPd43LidM
4Pu8/9o5lhBcRVkI6kJSoQfyu+rlYs/gbky2dgWwIBazbfhgG8Iu0vD5icW0vu08
0SKCfV1bopmEjv2aH8m7j+6nk7jWOhuSGHTueYN399xnr/F5Apy9Pm65qHCMewwK
8+/Bn2zt24PdBcAy0A9uBs7TWFoObdHCjAcIfUGM4TrswwP3+UpvEYy65+12euOE
q7ouIHPob+ztbByo+9X1VlzXMjk53SCNVoKT/cSyfYGv4bXpJyQ95qplioTGORfD
SgR9kHS0gaSJB22kVHKa7hsJDolXZHMILvG/dPyG+UH6ICmcuumdetkSluIKIsoM
sfp4q6NpCkzy/qV4jH7/7oDQvQQNTLjHnv9w5T5RZkije/kp+Rii0pcvZlH6DTMG
yEcn0xDgo1jFUAWsdDil37EIau+ZGnI+WPBaDYLtNL55aQq/L3Veth4r5Ec9PLJv
pmFIZJZVw5eK+EXagMNxbN3PT/qiCu1WDl8B1gzA0K/jEW4HetCfNylGi2iQCnsC
Rg7m4bbYvxDD/WFn4QnwO56E6lwsAH5jvwKHvnIGT52yTobyoVZlb2whqZxtlm0L
xmbIMgKhsGi17OZu2066Y4eH7mLE0p4isE8VCEWOTNvcdTQPdRgoSNJhwTpyf2Nj
Ks5zEpk53zY4kmqT1HmOTwBhgvpj5ZHEp6mJsH8yxnE8MYrDuATRAubJm102nJJ5
FaXONFxc5Evt6xkglqiLM239x3krUnjCo4e4aGZLfhERW6ofMpuk+VARNJw8zf2E
ybBPc3VqVbBbNEsuJI9Ry0HG1KiEEc/rEiKGTHNSb+QiOnRpb3wm53W/nTtfDjfv
d4tFncZ84cRu9hAfszf42z5qSw0j1FBTSWEtIp6uz7mbpGOVOHz4/29tUu4megOR
8jOd+9kuwmJo+fYztNuG0eQk8pDAu8TGdDtm2XQboQtDsPs7xL2P8MdlM2WqYYi4
b6JrUuhT/9DOosE3iJuSAQe4Vgm09EpLJtixjs4psrJL3dqx4+FMzSEhi/+8plTH
U9TakEK1XBYWEm6y2rq6yzZgnFQtR3jpb+5dY6+E9QE5gAImfxFoczBVi3jRyk0S
p5nxBh1xkMIrtLYbMR0eybkymiA13InFj3X2Na24ErdJ2ofLdqZSJDnTJfUk5YyF
+bp2BhGXPogSNmefYsMsc5EMmzhbSJ/qhK9nA3WnPDEFQxGT0sac40i7U0rkyJ2H
yvb882udYZI1dggypncJ0L6hQY3+WtV/owSKC3MWJVEGW2W8XMWYFX0jmBuIghqW
JOPGJ3wUe5Uv0HbA8uk/FYlzI9JijcDbYY6oVAn0YcsVDSgNHOmsTh0jQ25G9/5V
VkkXz/KcJP3ovqxX3Ymh0IzA/YwKfDWm/auHouIUIZE6K7bvi9Z2UwMkxauKFfxi
ddUitLcDHvxfUiLSFTyVsTKndnNKaL4/xQdBn2CWkeAt63RX9ert1DhyFmAGvPnA
c2DoJw9U3fRkYo6fvMZd5ckuL31nS3od/O5UtjM3d5EgLY9lk8/Pg4Hk1b75JIqQ
yrogBTJgBR10Rtzs475Ps4ePFAE15zFCotwwBEht5fVhx0aGDeGC7HQFpLuq0I0h
+C06SDwxT11pxXrGP0AL3wmPYu8fLzbLvNUmVdNCLSGEaQLlIodI4Lh3FwVQhmxd
FATwdi6rvTqPAuxHS1K4WzVyRS5co2Z2yMtOHMgNEeAU63HjEvgdCIXiJ2b4Ylns
yBtVUVKcK3Jg47WuRgdHtl+tXeuSAY25Rq8eLy/uI/XQ5ckHZplYBgycGxtuhbFz
Ildr5DQaOzwEZeOJnHD8W+Q7YhgFeNLsdbdChNh9SacwU56cnFASmjluBAkZO7+r
yuNHmdBWSQJn0kG1e6iRQ6abA4SeTRHP1NiVUaY1SNLXnEuUiheYYEc1jiFeW+hZ
+gw70oNomEFsYHZi0hDi4cWZ8H7HPd2DQJxg0TRfXyscgyS7+3QYAf40Dh9eRbp/
NZm4u7oFN2pYrbqt23EWi5rtIWU2IlbPUNZK+5rVINa9aL14TghePbO8wxEb67Z/
KVlT5IGNjKOwfiHZlc/TO2OiVWwOEq16rHInV9qptigUa0cYnosvUpunUm6iM5hO
uHx4vVQm3xgeKgwCb05PstA0IwjpTChkdfTj9U5Gdha6LXgTN9WKV8cgZl3buJ/z
nlHaJaSAJpRg8egwNQm2Dg1+s8SMsZ5DqQ+0TBpuNfO0dQpEbtcQOcVR+dNOXXjr
Gc4UQQhaebuebSBmSuZOkeuUiOM4cxpQmpdC9TUQbAJTwoFfBVSvD3beYc9bUOXe
/0J3R83Yz8+t9ku88JAyXGSsGxc7jOCMsp3FwbIwC/yG4xtoRJWqezBvlgtCI+I8
nMsptScFwuXaQJxLcs6XpEDlOyiN9AltpnzR2iN1T138DPZMZRJRysPzHBBHsNda
Zv0+6yyDXYA+0j5xTXws1j50fy9c7AQ+aZH+vKW0mcSWkfWLlnpA1b0i8twfo46a
Pg4oeUUXMlR0QO3/874FSYhmhYcVrSXP4gNCHvf9xK7wpILfGpYzPQI/UGbaITAj
UuLHw4H+5qu8mnHr6K41/ppxjQYgCMNMlVJB8xZWgTxT8YMyfp0KJ9VoDri+smgc
LDtisVIkr6KRL3CKjMSnTzuqLqtIMIRr10hc93/w/QcnRiUtKKBlCCjCnF92/Gke
5u43zn0GPJXyE1fisAMjBOO+HyS+X477XHSlth94jrqFYDyEo7MOIDDbDE/3SrUy
Yc7EWB4mPvEh8egWGpHWy0cSYIPVZvHQhKOqbEHxl2oGin7lcql4CcPqaxMm9Ksn
cNqjCfcv6LRzaV8+4JQd8RPfaBkHf/MXYA3Er1GxB4ahehBLtoomgOiMT8qCazh5
BDoqnT4geoWU94y5Ifg+wMO2RV7NRNeyff0wrQIkQGvmzlhAGtZxo/VvgewIFV7T
L+r1uD+1S12tVRYPCx4iriKqeqVpZnKf+XCqJ9ZO5AdkGmqUSwjM8ulSBQRfqgDb
f/4XWRhc/49m4pFNE2ZC+/z3lyTV+TKr/sdBke3qstPhrpU+vWEzuqGS6ChF1h4/
071ILsQ7OTQwHdNE//L51Z+T8KEz79gjh7l7CHNnDeIeqDRMAmEkFAEu4RdR+QS7
B8zWNXcMorfXpOZKwrkXhfnJce8nctz6louWq6iTeRsi5eRf7NiDf4Nxk7KuAKet
rLDoXT266DMp6qfCHxdSd4OlINwbIE3T/c88uoNt7iWoDcvwNq1GECFeEc1tYSrA
CEBZ7wna+x6rXxlnaoXWWRThNDsVUiffJw7A1gHiSuqwbBSwTg92u1KKBGgXl8C3
JAzcnUxRvd/1ZheVksF2BSVEZH3M3HDCB8xwZXZxlPc57/HtS41gzqIJuQa5u4X/
qLFfG1tjM0ApXthp8aJiwe15Kax8fxCeByzDC/ak7GzlPn1To2isp24/NPE+FYZ+
N8n0IP0+G+8YFRCupiFpdzdEHUAY7DrGhMigNwvGAlKv0rhiqujwqEA2UTIwJEXR
BwcMV8wYHm2zPv0MI05vHuWsS/Z8YnSctsPDYJl/CS4Y+ZLZMFGR0Gmk1CKRKWNW
qfCQfbFxJtB9VvcXWJn8j73MZ8RY8DwnjpW95nCBmqiMZf81W1sfEcKdZ40oSdpb
qMF0Tj/7zAI37ir9kfs/3rulxTcNF3s+Ra97xw0bS2P+ooir7kGv8vZlDTGcFEOg
lQbjqpwO6ZYeyiK3OehNh/G6+115bdPyBNQJWxpaPyqiTKYX/+BUJgAdUMrcZgwo
peCq9YpcL8+LtX8McsORWFcKu6gpUpFZy4yYqIDkMbqlkdAFs95geMHcvC0cEWJQ
EIyfXvojvfuy7HkvHMF6dcSmHgg86id6E9rVGmeBnNDlxBW87o7cfodXDuZJSLSG
iicwuNFxOmHLw+s5stpCO9gzxFgHIBTjn9HbUNJIR09OR9wfxSVkgfAA0EzTuMAp
7j9SpFYdxK6OwNOOkZQkpXxHExMzxJ+zRvfMFhHChS861GMWtiuGPZXnGBB7DBav
i0HWOcvaKla++TmD1Szgj/Se5lfSwpwcjtiHHBwyZrfS1vkoyAT7cW/xqukKlRcz
+EVKCMT3CZLY0mjrjoObcXh7pUvT05ynwt4Nrdh2gqtKVtHqOrMt6/YPgV4J8C6N
lpBCssFfADH2BRxG6KdmqOFSbnA2l2tVI3bbUoPgrBcc2FVNpbrSJ4QsNQSNgLVT
j9lkagCXCcG1V0NFYIsL6i+CoYmCxEeA/DisN0UVJX9NgLa4RQ4yjKlXdUAQKcXI
Q8lxKNwJ2K+tBP9IMrtDyY5jYCbHQY1PtNm5qF5Q2QWWG+Cvq86ag9vTfsFvVZuz
lIXqvGLldWriyG/GdeXhDEPDZzEw6acyzQqc/K/GRYPN6GKJ4Vqra8ZurCAz3/vJ
6Nz66Qwn5RYjTfD6tBmfu/yjuyimIH6xkrPC0ITjK4HmuADdRzVMY9eQx6keKCgZ
5AWfK4nUq0e+ItfO498SYMOcVMH2gfjjMXVCnwxLT+cSnStE1xGaBHjgvgu2G6Rw
gXFjMSvDptsGtZ2nKLyPZuFe5eg75JV9AvqCj7SSNeS/dTPJxo+MOuK9miVqs+jW
VFWHENsqusYm/pMECilH6C8EZiOSD/Y2QrzIrjDL4nuI/HTyR3MYeaE5A4M5d5Hc
c6exsjTB/Tu4FHk/kZJMsY0a/j+UVYeA8OlG+wF85vWSYg5rQZ2HmDKfXhJwGeFO
F2MqBhFtyTi7zQr4ExlY+VUY/8iCppahkJ07Ls7PQeTea9WjjPrArVlb3UW0qnsJ
ABq13KsC8RLYYtlA57CXmOZuPJ7fq2GJcaeCmL96bEWc4YYVwZNCTCLlumiwADc9
9f4hPu7c1w+7skgmfaXrvBGUkl9dAAyNReSqaWdZxpPX8EYlEWBrjJHdsdpC50Gc
Bp6xNGkFrs5p2MnaQK85BECRJCdDFQwWDa1luGpopZU0fQx5mLMg7cDeluDS0NRF
xOs5XNysYDdCl4c4M/q6CYqWlHZcVSS6JoOEUhVGueVF0w/OsGRllJgKEk3FcQ/S
QGH4OGOUHpoOLA9SYmPzypM8QQydCT/EESBa7dS5wJUjZvKMKufOF3UUdolkTDGd
VPEn3oqAxTYotlBYucQuEh+r0vZXJ2YY0UI3E9RIKHku9GaxlJUo6q+ifEFBgPNX
3bAhNqVf0pBXgigo07PT+yqvn4ucJn9rq2YPA+juINZH8Uw6WwW1yH+od+sLRrkG
wTnrdB9JZPakKcKcjLxN5Y56dTJSMgM2q1Pl6/ynHJ7z/wTA7ceYJl7A08RmEOCC
qoydgu6LFM7qdogAu5rjb98114ETYH/g8VdtlIzdPWnOxaQyJOWkpFyW3bnPW+TO
XNjKi76xqTCAgcqRCBT23c6CRMCGFqXXuN+BgCZdtBt2GLv9zC6T1YL2cRCRd+x7
M0nCQO/Vpx7REckG0EHffda2Wx/tLPMbaHw4fqMZN3aWECj+mxMOgDJf+CrMg69d
wpTC2/aVXCOKppUNg4YAE3gDMZCUK/tt1zBvCZMdVIaKHAC/5I5ZTldI3g18c7eG
yS02Y0zr2JQ3Fb5PAp+m7XYOy9erCFVq1L7Y2JugFLweEuOd0hVsp9ZL0jaFaUTM
tbN2nmiemsfb5labFwoYyqxVflU4+pdY4Ylqxg+DlIsW+RhlH7M+QqKA8jNRZaD9
0xJRAnP84T6hz1Gi/c+MXvcnRAoqTnon3eYfVTus0OAiWQhBAq+E+V/IJIVn1nLM
XIOJUiK8XLek5ro5GkxWTLCS25+e437PYhGtf0uDIE3+FZjpjYGpzon0taP2jwZr
A/F1ddqiqemFmMPFe88R0kbh7FFIi0JLlpWOkI/eF7Wjg1j2vypEzEJy2F/XISd/
68EcYZ0uo5QHuaNtHDSFzF0zm2WwjpMd/HNxe9AVQGCyQMHZbQJIq9uXhSJYZFkc
fHqWH6KyPoH90f2s1XSFgoehBYVgyTcSJJwK4RNarMbcKX3JawxUkTSL31tEwIPT
WcWy4lKDh8FyLKbR9a6boQKYObJhaDXCEnJXRGy8VXioV/yDXwV7B43LfihgXhzu
eMN17PMDELwRYtM8aMe68LqS6oaZ+eGL+cLNwFJRXoSfc9JVMUWZAfxmBdueHcYC
dX3K/b4bd6vldYnHSTTg3PVisry3PHLksBx6Mx1gnJ2YkOBxVa5Gx45oszK3mXpT
cExLb8DbttL+nR0xWDnugBbJeZ8APWBK7ywq7WHZzVqqfE73J7D+L0hTFfNBI/9E
miI9Z2szq6I+ngsuo4xoPcbPIS0MM8d6YtZespo7yfAJ9/FsBvpRctN9cuA/nrpM
KySS5jGFAgTuvjKIzDlk1Yxz+n8fSY8Ka+29ASIiaK2NgrsRyPDE8/SR8K4Hw6hy
kdmYPYgNZvCYoVJ3viZhWZduRhggQ3LoVh+YeEDoX2k8JNz2P4O6tpLIaScsAUXM
kBE85uvV2AsygzbDd1cEfnzAKAvknxLSJ7JoUreVJtWUm69+NLrbOdHE1xBV2Gvd
WdlSaS6yZRsgVM62kCMFg9VhUT4gLz0HSyfc31A016ebavC2xIvMRbrVqzKU4Oyr
zWgiRF+5hQCKfSZQ6MT8HdgJYrS0WDeGU6VZ8EKGqEaxojsShiiiTrWSgTxOcpa/
TB6WV1g+YFCKy7phCJX8bDZiDgQPpJvt/8SNqXxihNrbSpZd0FkNLs1Pm0lnyM8s
DuRxFVZRkNtyD5DlqY+ABMNwb2Lpf0OwzIcSB6ZHXOTyrDGecNPdGBl9uEs2gvxJ
YuZ9h+s0P43nNTMR6YKsbNbgD+2GkSsQDhL96+9KhpjtTN0DpdiLoKMLXao3w20F
mqE8juGYPl29209YUXa4hUUqibLVyFhELGItei4Q/IZqf87kyluUKoNAPRhlaIXh
t1yl+W8hpAwqTPYBAU7HPTfgkafllht5yGRBtJbTaG9LyYbJRVjYqI3vul2Z05Ok
ohaHgaoMDa4c/MWi1DkjAQx4/QgHvyuie7BV/xhZcncPEJyOZOTT5s5QTdzVywir
evX9y4ABHuiL1DGfMRjFCSYOOik9MBeu3S4z0puhSiJxv9ZLbSSE02EP3SUKL/zE
OiKaQQuBskLj4xPue0J5Gp/p+Tj7i1CB0ZamH5tIq2MclEKJaFN6wKHoFt8I4YqG
EG+dv7lWLivZyTEZAa4uxn3edj87f+kC3ZP2BE84hzdClYEvB0cFPKvc6rlMu6f0
EmYOeSoKcFe9RsphSmfOPQIK2QHNLfSaVmqeFUXYNFKjwfuGIcDxPlVoh64D10KF
yNF0alkAJo+bPxTqTa/5Kx/pXIOO62DTp55DmZMeLLAsb9EqKmn9/cFrVPAkCh1h
rrJe36Ucowtkoanbx1BN+Zfn6mPHCSsS25pujETLrD0Uo3m6wM2NCHXoguGJp+jp
2YUQn3fEiWY8/5p3slESffQnKt9P2CeEi+ACS7UxF20BAQrVOrdghcSxtWOPBLfu
Tl6dZZWdFW7xf6qc3jGUDCXBzqW2ufjwtd0XoFsCJrAr30WSLMBQKGCqkvJRiMsA
QvsNMk+UTuHf6qk3/Q2dGJRYVmYrinu2zZZqHP7dVKhECxnidLyllrAUx5avehd9
IS6303tdEdPLTyDwoZYLYSd4SqSX8OY9+UfWIuZ/TgMfXOzZt0yRMPdDvBbgQDY1
Nb8JBTCkBoAcWcgzuysE0MH7dm8d3cw3/Wk4xNclkcBfOholYuEYVbhl5SZfMeCD
YGkBoBx245KsN3uDI9giZMM5lqcDB2//8hQTcBHz4Gaxmt/L3GXnr8iQcF6QOstM
YvVV8SRg1NoP9gPmE0irxX8nUbnHeYCX196u1wXvkwtDqH7n/LlGJUwt3MDZ3n0v
LyWjgEJ/nBHcQQSDoyISbOqs1SwGrQ76VlBel8hPaDoS2XdW0tWPVvfrCKFXVvi6
Y9Uz5b5N/gBWzXUDaKPWMrLYrZiQVL9/2RUEGARs89KtpDlw/ewr5dqgzchasCY0
F+/bCE/mOpxtdUooVFyXT3/WMXzgzns0i4kCV4+D5w0KniUfiVbkBVtoFWDnld3f
fxQENUvhD7OEjaHGQ+b1NLbH0iPFEZJeQI+mtjlq8WGgbnYnI2cQJQjtCE8MQYiC
r3+KMKJ7dBcKOUauAxnL4E4+qr5W5oYeAbGEEvMdvesmat608HTdqCogp6zFFUmW
LpARG3FYhXQvSu8uCveobccTiYYRyb8yuX3hjA2iaPgyVQG07b9fWvqz4Ew90y5Y
MYIWNNwJ0dREDBqahvmAUPGOcdaqT10vEQtMjXFWe2CImRrOrLCNyhUTvGTC+EYH
h8zZMEbEZ9lK3bl6fFUZm2LJGD1368tpptLEv3z8vnuLMykA4DwwiC9vCDzB+25c
w/ZMTSdvVX32E4ErWGs05KBB17KTFdfCG7JdfSfw2pB+RwYZbExR9CCeNwcfGdD0
DRkmpnbQuxOBD2tfGqhfB1Vq4FY5sRA1NgxdhE4aquTJK8vqsP+gyk/q8eQqNGje
A4bs/kllprEs9hBO80cPiMMUCS3HOFc6NmAlF0JgpBP5G+IBh3ELsun4l+6BC/Ry
Q7Z0YnRNt0K3pk95gtaE9eHiv8DYiXp9P2o1UY20XkjF8NKevIUE+0KWsYDeO8bE
3gdlOFgIqDCwxJcDMytUjfC3MVbwr1Q4ZqyELaVi+0F5XSimlNMrX1zTCcb+IP/+
A0VEvpM2SoluuICYvKcA/t2nPXTFd2QnTui3pfMWDZwGge0nNCgtJY7QEJJLE0sj
w3Rgw6Pa5qhg1qTfwYXazD4Q8MzklanPBbqWWs7D3p5lz/6E02Ua88PfD7SnNFH5
ltaL/qmBpdwQj7YJmOnpas6blpfKVcjLJ3agPh5tXedrKVFBWIGb4klgDiZqnu8C
xrWMNW7vkNDDE04Ym2cFQiWjBY6kpJubaxdbNLzKHs2ux8eAcTLeDxM0LiH2sijA
b7k7BBaUGfLmVfe5bjCd1GfMkpg3Zwz+Ov7e9+DZPEutVpcic9daXOdAnJexIS11
RNGbWTRXGcsfxrOa+yyed7O99aw+Vy2qnT78zldLXNcMB8Zp2h5hFHdaChQkj6P6
PYUBipvF5+xojsnsaktOIos4BBJT0X5Jsey0UhrIN5ocIHp8ia0NHnCjUhAyjoP4
PPvag1NjHHbGXZxxS6Z9QcyBIiMDQeg6h+TBjS9aPORgxsQlSkKPFaEEZKcpHRs5
RZCKK4EgJLlh3K8Xl0x1/OVo4GewtEbmRAwUj1v4BZnHyfsxPieL5SqXJ0Kl9WTx
R7KYffYQy3Puw3jWFbugFFHMHBthvZg8YfilrusTJYHKdR6jRAyVPo7ThXeY29ur
HZLIkJ2OBE+87XzeCFMhoclpxOCOT37JLoLfeJ6AjgX4WwZs93LtOP/zbf3pz5Yg
zOyG8mw37+3DVfyO0wnvXj1Rt5x8NYjHXAGLJ+rsjWcz/QXgHiFuFFc2SEGD656E
smdPxH6CkAhl8eZ2m7WKLAYcDWibyVcgMgOBNM1ET+2t57WfwnD3qsKo1+Vtl+6f
AVZcFYwcBj2icMI48kSD6VPzWgcyMQHW4G6Vg1EwHEWWldEtxK//an0XuejoVSug
EaLEn4qkGBsFKTt1Hi4Sv5bXP0o1ZCvtMRPyPcXt5SWU60LZfIN5lyc8BJgB0WvP
Xl2bAgqhwH75lxhP63wOSTj1VY9B6GQmetMm6SuWddgXPOZ/pIhFYAgc6dkfQLGX
AAONfeN93X4k+Agef9zK6XGXZ7R5ex8ehpb2OFXtu0Ehq4afYph5LBDd1bJOznoV
Ivco9Um9KEHT3Uk6zu94uUGNdDqHIaw9vW/zw6FQ/c1jqCVCz7Io3/9fpaboZJqS
uZDQNtmwwKtJPizkXnsn/zi5KuzveVI+icRsXp96Bro2yZl87frffdPsWoIM6Mxb
SsjBMBIyXpRn/aJpdkFQH4XRJ0umSAUVzlDkyKgGv5nPIG/H32PwrzaE6y8dp5Sy
AoGUuHvglKp0EyUe16kmMuLgAQ/JYSOVBZJa+roOjn1Xmk2G6Ug405SG+LizkiNb
FmPZCVBWZEC0m4NHPSDIDVSI3C7/8vaSrOSYK+U+X9PcmdukUEamoaUi/2mOgZ4l
jRkcZE2KbwBOMdPOd23y1QwMPl2ViZ6B7cyRgYkOwFq2zBE6HoMOhLd5eGO0BaME
mLbstp56YzlfURshMEnWGoy2FgdO0s3NLuwm8IYBo3S/PBOfHxAtY2FvuI7apdsH
FQQQTBJnQ8+Wv+S0fiCkoVjqSJjofjE/u9ZXl3nAZkgbhDNri1G4fr46twCEBF/5
wPWqYj/ietuPv+Eqhh1R54IAojLoU/xYut1ISBr3ke6qlwIb4Ih3JBpOPHE0o7Da
5g/0517CqAhyvdqyQi5hsDSZUgThJ5J3iS8DPAD3MJxSwwPRzCiGM9vbz6WoQR9L
oaWm+u/2WbzN2ah0rJgfUD6Wzwn1WUb5pDe6VMaTeW5IvwadKaUxps9iKc38Wyib
H8ffa+bEwtpArrp56+V/T5rmfJNoFLRY4clXjalAqOW2Bi/qS0C6pMRzXEhBNNw5
boDTOC3pclF6e934IFZSHBClvMFPYK7ja0mO2xQlVgu67/UsS77AVZ/UCiV8raWK
qSHoL6i9Et8MPTUahYhWYvESFzPoZS80lQeX/uiiXqveyqnJ6mjD1tHWwpCDmJHl
5HceMTUOkPTPXD5JJNJslYsFzy+jxUPV1HCFGVIKbCSZjN/l6+UYZvWz9b5Lxx7U
b8RsOWyKei4oULBGjn5FYL6x6IyRtTJcpdvVpeUICafs9xouscZj1JpF/PMPr02p
yacT+b7tuW59EBbhxXtUN2+8YUg/GJcyIRLn7353R0da+enmRiSEL5gIND+va5Ec
Ffk5iKskO/ZU4tbObx5ByNi9Bi9vBVyUuuP37FRkPN3X+LNctNJzFI+a+Us6Yjfu
tQd2YmJLlAAKWMzgDlJabwaOZp7BBZ3+m9TochAZPKAICO7TVH5RoxYBMDB16Cwh
R+yrxJREQIM9EW776tE7dhuJW+Q9sUBBXfy4yHo4S2yBpcZZCBn0sKhCxrFXzbYA
91vftUChhc2fZ90vIF2CQXziqQFhfX6SLftQu/T+4TcWqtte2eU7p/SgbATTOab7
bJAAPB7NGgafU71enlpMwsVLbuhi/i7Zx7acf0xjAgA+zSprokAFXLEGUP6DXP72
yGFGbkZDd1Rob+CMud6Z9AxqPOnXjE/pN50vtcnFG2CAeD+z5MbzqaaBftECV+r9
K4qfvIIJZVP2jbDBa6tAty++BR9yk8QmsAMi96fHnJufMXW311GGqebv1Z3/mmuU
Mzl1ly0Bs9ZT1muIOO2LNygdT24nVq1a1ft64aBMerdHafUI3695C8eeJuzYC2bl
LQH0O4bu5lm36oltdAg9Aa7/NmDvyXCg5XpjeQHDo/te5O7cm0pmAQPae4my3BFV
g+sgvKFBJiSKI5KJKS0EhUtzUzHylNTs87iDKOlMbaE8I9u41HYLRV5obntnNWfM
xc1Bk3G3ysWy189LNSvZgsOYiDMGPZD7Y/rZ8Wyi1w0ZBFv1doksptjMigak/zbM
p0w27798PRI2IhVPKHXmbKSXVWHkM7GnfZdsGiCT17FB3EYhDJhbRAnfkmEuEoqc
g1qe8rxROIoxaboFp3ySRR6Nv6nuLAxw5qffjYurRYncCDoXKf3g/BpFEDY+Mv+x
wfmuE6VR4aQd+6j+mil+N/LNdz5Q7nVPVzxfXXJv3djd129E0UiTjkNhEDjyQoMk
gblkvF8Tg5uwk+lZf6i7SgIeFd6aK+VKyYc7niL1vey/s4PRvaqfyCRkC6OKj2RF
pHA+O25ubrcPiErQ01TsrfTCB/ZtQgR7rR3GdABJX7JW3sxkmjO5bD1Lz7RlUzd9
DLjSFAPQ4kkPJ1LlqgYhRIh5nJ0DWoMFY6hWqHNkRxdLrlzOt58m9xKT4hh7k17q
x2MuMN1JLbYmHLH509cE+O4sj0skC85aW64hAu+LMLpe9qmFncbUD6C+Gh2zfgMp
F5UFEYpr5HLa1NIrp9EOcEMl0Cc6zIXEIPKiiPWdFwnVmDkimTUp4dwZDIEaT94s
MUx4QMSXkguStJVYwhjud9AasHsrUvvdm5ZKyHyuwqa24cterng8vZyIdjwMqNtp
vqMxNYvDYn4/PmkeqFtAwHTHjHSZXGurN+c3BFbZxhvMci7sDCnaiWCcFWabBoaA
ybg25sA+V3CKjMPihccYUAG+qhpsH1rR8FghgGEWkXXQJAMFfYeKDVcpr5CxjsFZ
Y1dezg1iuqgPPGmrtTwxskA6Db3+97aIJ/TLDH+pb86gpvDsMbEV1ElrrcD3lVM5
2acWjgqYtIxk/E3G0rEmAa+JLFlHbaRKAodntDaC9fQR6dfWO99h2kHN22Tws1JY
FhcwlzBaN5L1Fus07cdLJmoHjmv+VFEb20cvkCVxhkf1TqAipDuzvz/kMWWSKP/R
hELokLs4yE9NMHpLXG4lrabbNJY7jfuc0nEkcgxFqfYBo48GAhiX1O8r+FAgA+JI
fQVXBi0nPpCrP7ZScnP0ZDdPZ5n8BREpPP6Nsbj6ZMHC4RSigW1E0awn/nv5viwa
GN4UdzIjTMjPCkES3mqpdIIrPag90OYb9fqfnlP90rMzuUQcuP4I6BlOwvIrMQSA
N3LgyYURLoPXrW9TaTjRvoPEibYjWVQ8d/d3O3kdxcS6DIwr717ckkTffxY2ilNc
k+mnAx0W5vpDpVHhbB9RLVU91wPbZt0h8AEFV8KcraBS8jU3RTuswBCITL9qKw97
9idhvPFl/7ujsr9Ljn2pZ+XLP5AatSwxdiuYMGZVeM+z7xvOkMJ+t6fzwdsWXcF3
EHiS41u1H2knAMLy8ske1EOlxJIDEH+darbZ3zoF6H09vSEmlPcCEFDdq6sbzElf
HZXzJULtK1nonpBayelxqbule7UpWiz+yU5yCmVaDpBQf0zpUvMR5R4ygj6P1M8Q
sN4PYgnE/cyGbVmaujw9OEm1kz7IMIxaVDBathf9OvcUhnbUUpgZVv1qDLqpBINN
pJfOJg6/FSq0hI2S4chn7A3Dsc6gn9f/fcnEOg08SMRcbP//SS/Rc/9jzC6A7gKE
xpWHl3AL0j64tpM7W5jt/qPWab/iFtE2k0IZEf+BKRuwMwYxQyVVfxKC/RVxuqTD
O1SDLhkggrG+iWf1T0wLLy9clZJJAtIngsUXIwfoNJTnMU5s6VQx3/8Euo9G4zUA
o6besypGBC56pwKcSS09C11kctfy3DL0LK43y+Zu5LAdPTdk9l+OlpcDAH0Z65DX
J9ADzPSH6c0OxUBjjSply6W98mjJISc8UGxTInxvO9Fq++DJ2CCZXK646cojiqvR
VeseFQbb01YA4c5PozDS29jD226svQ8evMqB5fYaFBztOlg9TAhP/trPizkSVl8K
2ihBd5WUOpqsiZwfXsbE92faOu28tXbkKrvF0Gaj1DrQb3BtKReujaELYIaBpI3a
5z0g9acOT6uwJYkX9REEehosYeLpEd4y5EzSBcmU/ohJKD6kn1M6JtyNdaD5/qnS
lREqZV0/8eWtLtqLVzR4jYnLpgjlHhyxeQAEt14FDM+COQ2zicIKgLqLGcN2HpJ2
sgcy08QLO7yEuyR3FaXv3aDSdnfgKvhCYMFbBe+bxGjH8YzumZOhEX8kHwV6voRG
MNfloPr2s1B4hkpdhU/joVOWcGGGfvET9B4rdTFfFHSwAxNL0is0+SS0cLWIzXC/
nAvV9Aw0UWdkM1sf3RbNWp1SjftlcY4CmucxhuaM8c/J2dWny6j3rKp81T62rFca
Kkg+Pj5IM3VY+yjRsF6WIMgG4bp6Xa45lchdd5gQoajIkObv/dDvLjuXXh29atgw
1JYsWiLKTPb7NUoAT9/WRsM6combHFVcov7U+8fT/o/up912bsQlzc8C0XvgIxPy
rr7gq1p86byh7HgKOgVb3qjBQRCi27dkDd6OKHNPLSCFYVDTYaTKuf+EeLyA8lEr
iZsHwbBvwBCFRopTd4NZie2DBMQNLmQdDLpP9dSC2e3hZFnefw2LvSynJMXLd2FR
sx8R+e1HjfxEJXNpGAfGpEWttgN9B8EAl8MqPg95VjiqznlyjnXkvzKCPLaflbZ9
j4+KrWWbKaD8Vjw7SZeh14Fhwx5rt3Pk6kqmEJMrE4qVPWovLIQ40IyDZ2r4KhJI
Ag2JnDho+y9pFMy6mCsQXxUz25N96x68cJAgmoFkUepR0xppZyo7JQWVIep1xbQ3
MGr78qQM5O2l3X+dGKIBoU2V/Q01dYUg0CLt1yagSjjuIlqsNgbS0V4pWdONT2hP
YIzC6juoXhzpMHQI8NRKZLJUuHiEHNBOo7YmmYoHrsZSss2whMinF7s36r5sbmCx
B1CM8nRgo00hJLJTV39PW1k6/JwEWpr+BNu7W33cz0wwkpZzSah6FBuAMQ/nC3P5
Pra4bEQWUnnSk2NQSxX9k2QQX+NbR6EueRZ9Mc6+1z5kctTG2j4HH0HUpEiQEwcX
f0a124RZ4b3/q1stP9m9BdWNIDk01z+rJLT8wgSN/Q3sdf1DRTJKPhlxQFZ52gcl
roBZoe7TfxPdujPVLP+P/ExCvIJ84OeF25lygF4ZnYUxI+E6zwgYnmt7y0+4vXUB
3Mc0rYuEGx6/9GAKXyEWPaeItq+gZMEjPhDN15KDglhvhh5cBkFBabrJ94vzJB1p
GC14xYafB6PRiEZLwSscnZQi39kBoML57f94VfigYly9+QxVlXEfTQE2GCennmcB
kIJAinOBp2gvt1ZjY8rXiBKZ+VH/zVy/2VVqc15P8Ud+pmaNHwq4DsEat5WuY10E
3FqWPlUpIaTdfbO8UAk4QQCXweoCUvBGd6ydAmEYVZNgtu1i8f598XD99EkgTz5V
/+Di4YVFGKqt6GorCBeCSU/WyGCHfX/dO9gcWCSYam2m2axKTwBETJ8hCqQjx76u
Vz4tlbxyRKj5Y1Fm7dmUkgX9W1GtL4dPIJnW3iOxYGERjG1avYDadgClhnTbSfS5
aqsdCAe9/Ly7jU7uvot+Ym+JWI493Ectl0wA5a7553sYWtjNtLlH7J4gH9Z+N7KM
IGRIL1lGmtaO8RUYlo3QJ1hruzIlimcdGrYQSwrInd6mxboLNKTr0z0iSNeTSdTu
rMz5htLxxUT/RCFSdXDB4vgl4yZd9sRxQijqWjecvZBIF4Ngzm/4obHlE+BrxfHm
uCJsQFW7D3fkTqVve9QM2GWBErr+zpWZH77XMUVOt4u2HySwZE9MFNDaDjiaYLCI
0ClOfKP5H5J224fzQmI1it33MuOt//6mr2ZAicNZjz4fLI8F80MR1Gnb+cEwDaYP
woLP1MIMv9QOED1KsuVb+3+mN+sB02xfUxUbyxZglsRWEHkGqvLTqTc90OCqtTbc
azoMwOFA9gDE5GmBHGBv0rx9vT70SPb+fBvpfaGlncMX6rR9LzkwdGBS5GemKxd3
bdDoIbVuQZMlSO9jl+m4sDviVwTj7bh0Gh745J3CcNNNlzu5q/MDA99xL8DQPFeC
sFrK7apNcd/JbKtQq7FPCpBcmsNFMtOwFEnUWFliLdbPTigOez811sNYHNEqP+YF
j9opCQwvtwEpAdxdKG13otEZ3OtHqjDUFnQZ09fRu7n26XYuohy0qgo+SiQBYbLK
yT/NtVkhnz0rmYbGlZEioSFYPA7gsSgjLBRVOTjk8V4I5SM/TDvL9TeTA1AUjzmn
xpCgVu2KZsgCsRsKqb49NiN8B+UUCsMSwPa5GHnAalXLdMJ12HrpqopDUeOjagFx
48AVwknvaaOdsyO78xJ8koJ945IiYfv3aL1PexDlRG6c3HH6pUSnoUfkgHa1WS4R
8p6HhGjmChSYMM4TJVni2yofnZw7Ysh+2RbYIgspVOU8LDmj8Mjs8y78tLY5tM+w
K5ynPVTPlEXvsQ0KujNyVfIQpGTKzb+LFRDmEzjsiyhJ1AlqDfUanAJS+kZ8dKX0
Nt+E6URu2iTRY/juJaMPbrv4Ldj3f5InyZlGoxdcmElXkpA2qpvY/Vnuucr3eAKn
fDhKIvoCEpGn5CYn6WR6JgK60ObCef1KPGjaSIf5I5rMdvRsAKGBmzeCNVi08T06
og4BKAdkw5JqHraXir54w4iY1OKVNfmJTIDRQSxITh0BZ6hjWbtiSHDdAdB3ajtu
Kb2j1msxL5GGOkHlSh5ujG3KP4n3kppymylEmbKbwqN7Qx/cvOlShgpDxAR2uhXt
sW9Zox24w7XHuhmD1YkYPQLXZbkYd7diHn73DJX4YfwCml8A/7yKFDn6owgLeD6E
DUYc8TPZ2Pf30lfAMUKVOdixFmI/8njDXztKx4jfFB4Eo0iQMkoifmFu9SavG/k+
eOJNBBBW3D9ZvJCo6XZoQuHVmFio9aKzHJRVFYbiPnCudFMeeRYeSaFPwCZgj59B
NX58Gqsu6LqAjkt6mBkXZSVxt2ZbSqkqIstGx2BqqTd/IzdNE0G7te6BkVyNiSrt
OlIyQOFvgwH0pw+3NHKpA5g6q8dIfge01jfRMt1mhWMSWUCCRgpHk0CUGg4eaFT4
BgTc7YNOQJEossFei2dRbgsPg8+bmJkp0EEu1esydb4X5wTXML4L5KTXyVym083L
6Sg+1dwHSEEvXVGBt7uAoe8eFqX293lFSirekRQrdY0fE0iADQXIUz2auQCdzrnE
6B7toFpwS5b/rYaEJDj4H0ZEP5Ed4oCFPOrOugytiSvIh4CZ6D1x8F+TNEN6Nbo+
6zrno51crOvL3BlDuu5fomdprr++YKGBIbdN6akz0KgzqXibSi0IldDJQQKlJ94C
knYiCSqe9M5sfvPC4MOwaVQvmI8gI6NG0SRFj4HA5ffy9JSRcgrmoL1aB6ZnwtpU
KFZY61K+VEsqMrDVTf6n8FOFVhaP9shaf1BEnpgC4e10FONmyBUQqKva9NdAZQXz
aC38Y6+Xy9mc6MsSO7M9WkWcF0W+lXzlBuhEtDI+2w5G2ad95WzWyYKmvsTQqcMG
Rk1Ba0iexlykZhfV5hOO0WOYSzBuJtgMLZ1giYSsutifre65RYxK3xdD+r3wg+c/
k591vBLoMHmkHP5YoeUasKVbezTMdthqatGrE8a63cpdSf6hyqSTztgdalBF+G+Y
s91GM1BYEa7XaFNIscducKR7378GcxXPRp5tKMNBhRn8itAmBWHjML2U+YkfKhz9
sfnzwU5OPjbBE6QQ+brkQpI3JI4hP5SJaGZ1eK9cB9saIpH1IGfIaiU6iW2W/gOy
QaIBvYHez0/GDTUi3RxFGfDYxQRVuLwhHVcDxkXuXhWRYS+b5vxspL+7a8a6ywbQ
egCUXGAoxpHTO8o/zdjXFnIi1gS/eSRPMe0qD3/xh443iz31jXr9ZlwYFIGPboPz
L6+dm5Hde+PhvkBxpd77SfmNUr1EiCM3FUjvqimObxL5IDO47X5gY2fm/CL1xTlH
2AOo8p9CoHdNBoJqCLZ+kovs0IrAhGlVPL71DIV4sv337Gi6DebYyydo0lJV+dmE
oGhh2z3IqI1vUpthuaI0IwFW6Le4X6U8v3vi5Ac2iy7wjfcc4okZ/gZ5QSIJZ+HA
OsyzrMYKSqY/fkDlUbXUI8Mqi3NS1k/8jo6V8FCjTnAsJ6ZcVIpqZDr8jJCzceKx
pEK1MHTk6JLVExekub9dJUgb4Cll0n1jGW9bEg/BZjrE9Z048Of2DRYIj42QoE+P
vo/mNyyBEM914oUe47A1Jm/gEQu5GX/4ZefBqBjkmXwVYrjjUUJDW9ZwNwK0jMA5
cf8OsfrekQeuHtfvd/RRFVEOqFUrxma0hxwK5u1DOnmfeZgjij68WYniSDFDt2Hi
ozvU+27jo2uCvE72y9m2KJPA6v3Z4GgleyWVy01U2jR4MFJL1wHNia7JOkeTcTc6
0rXicx1x1McZvsoPNZTzCgZLI0J73SCBPZHT80qdVb5cERBu0nlA/eSLYGDKXceA
Pk1Ek+DrEF2zzfKg7NwtIwlDme09Y9tGwIAvwPXjyAcIQL+0TCTTvCRLEccC7m6P
YLNvtHQX460ftz3akfgDCLZQBIXNcK2rx18DBNmQkGON9xu7ydbFl9Z6gqnTs2Bb
ySw3WRwvOZ3x/Qhr3N3MLOj4b0v8Z6VRhN2DDsHjxLoYU3/pnoZeBblUTKxJV6wL
PeXjqo4rUCOxdCdHYzosO6T1sG+TZPA+XtPw9vNoA7x4r40KC5Z/oPMAai8xS5oS
RAQV+BHDCsCNvSqIyXkJH/HpoYPNv1EA6ycH5bZ2LyWFaGwWm7whByK/9TG+mSl7
E3mPHIWijmTNgerYTcOZKFxgyCxMbtagUcSunnXy5wIFTI3uny4MkT23OXmjcp+j
2Rd9NjtYjqaiQ/wrKZtarjsx1Zi5WppFl3j4kNcaaM8m+7Y21d0TUZsEXvAhwCGE
i/7nG1L5Iz6CZH2SIW6p2F1jSlPCFh6TUVdMJVt89AH3NEo/Ev7crWXSC2YKoH97
YZ7LErLhYywRAU+cfx5eeWQYKL3xe+50FMM5nP451snBLRZstdCdf40L/gjCxg/4
T02pRTowgs47RA0p4upfa5oEh1zCqpI4VCVfp4jY6G8rgLx8KbvjIxcjvIMw6oai
SGrwlItzitv3n2TAUYw+Fpd5q+sX0LmIxv7XipMrGCoV/KdZ/DwyUKWsuPdoHPXz
B27nVIscg7xwKC1CVoM6nplI2p7IcUyGJEMNq1HPVV+ZYY9Rz6tLj45NV32/daT8
M5HSeiEqaOA1LX8nmxiWSoTuWJFQQ4mq/O1lQZb14BY9hdOgeRARhLu3xPhR92Ig
SHYcg9NsP0iOzmzrPf9BlNYyrGF9Nj/WcF9ul+2jrnAVtr2TZnuYzT/mQ8S04OYD
7SB+2rE+oeKqy//TZK3kDG/vuojhVsosTxDQpbWC0k0h44vsqt9tcZZIZLJcWiQf
i0XJbkTQuNyOrvoUd4z0XBulCXrkPei+WT9QdD4Hkryo7vivaAkYN53WzunKWafD
cL76IkRJdxg4PXMfhtLM8IxZ4T9C5nPyWJcineEu2+qROc69SvAYYmu34EQRBliA
M6SWEJfZGKeYPW2PGkw8PkAMF+B7f2Aiu1SESm7GSS0r+zpm1ssDhdUpvMv7RNAC
Eh4rU358rvcWC+D54NEp6jRXILmcaBs6hrwUvLnbKg9hxe7YaCpn29fXTpFBYZcH
olDGZ+2GvNsRMUlIc+NZX6xB3p2xA88grlTFRPB7s+cv2p+2KCZeDkjpDHTvInxq
rDorYMLDkMWbajMaKP2omkAgsGZ4rv10VJoqj/x7K16ph14hm55EEhGZkeAHCFOw
47q2lZDTaWSkkn5X5M9zwfVMs0SLnb/EF5bQGxptrRTQlkSuW523vc4GrCzRrOy2
B1Ym6H6jKr0ue1d8uiekU6bIJiUeWmt3RPuG9ea6JhcPD69eqHj4ou4yi8/uevQS
G4IeA73rlCKaEyYsROi4L/v+cL17nNpDZ2m6DGscUHBWzlFeYI81BbUwGMF14h1G
89FDwrWpRzXej7iOJBIUUerePtCdTa0182QR6A4GGW2e9AM+/TQBDsVmMnx3FJ2A
FCfE3/henISDWROjevVF8CPBBRzpbUK50s7ikGhSunkYn2MeQ1JfDPwBy65/Qdzq
jtvMfhVwCBkATufPwr53hKONswqL1XFvOMYKpw++MqZLMJ4yG7ByyswvPmKwoagC
+FJXhkiVCKFYywWU3XC1qUpT3Zj6m5HQ4lOgUepvBlARlv3DsfbmGm/78QyNYQ07
xH2JA1XoHHnOREevfXUkKYbesOXiK4VZnXBlL3b255sGMXKK3LC1Zfj6+yzLuUfs
H5kEYTau4DglJaOSGUFh+m3PNai4x6+2ZuO0HSnnJ9D2FXXCRHx7NcL0KkWEZzAb
DYdUjdPm8NUAUh2zvE+BQ4nEWrQBMbfcrB+ulL1JzFP9FeyBaa7SBNyPuid69ei2
orDnrCpxQm+JPNNDoF6nY2rr7DQbN3OE/L8UinezLx3YN9fjL4Mxk2T0t93aRWA0
H0sTxEvD7qCclxOKm8Hy9PSs8J+mTn/w/aPqaVTKbmx54b2SQoNpDYEcnrgZ/sg+
E5hYB4V6bDlgd3mQak0C8a9Uozs2oN0G+f1uRFDH7339IhRMaKvaHOaxta05EAKs
TjfBArT0N7HXoygIsgzZZhm8d82RKnaoQ+1MY0/JLMEmeUXWBlzlkXCpamqOHoYD
vT2snmsZgxMgE05WH9EWmJHc1trxiFO6sA3hChzyM1N5Vmfsr4eHGTQcw+6aB5Ju
KWxUc9wgliFMMovPI1C3nZRZ74nCrG4rbEnj7atYhY5ja8oZzvV+fQ9Z6kj9gNRv
IQ/wr7P5gMGmO2INXCcRX4gIgBhrxxAArC00r5Lgqv2SlOgcMvYz3GRLJqf9T92Z
lWRgIdbnr3fuXZY2UVpCE5TsHZH9++vuPOf5oYtnB+xH0BD4w4lHXAXNt+Uzn92k
8J//5IQGaSmQbRbEThdNryiy883AtG2JJY/Fqmy+Qt3Pt/fbsFxdvhg0P7tokZxh
UCx8y3s/9kGeyaKoB55r/iMdqNR5V0J09UwRNrkzmWaYJDzsrT1Rc7baXs8Tp/hk
y8a50J2eI6m/yaQrDzMcMTpDSQ+etY/NSlgIXFGe7mzcmflSNhqUmArgMDqyvMSx
5XOR4L5sM4ocqA4zR6KdnF95A5JXFSLm4a7sZiw15YUG04TVGrJzAPDzn3OVGlRG
HIJiETrvdlCUPK8I+XJ/tHSwU2157CQDyxdPSIBmwF/0uq6t0sSIDday9U14cSvH
U5D8sc6kY/3OZfGy8ftiKe6CAduTIMqRNb1kyeOVshIf6wu1YSN2SFMPJiAbnjKO
5NdoN9W6zGlUDGmsSIGdy9r8WdwcBJ4pmX55jCuTT6ryjeX6KzAtmvBLQBV3P2bK
Bj0WKDozoEFSSn12gf6B/9siUJhCvjbZqHcimD7J7K1h644n2Wuaez60oOg997TZ
RAmLaXxwsoOtFARwKJB5w8xK4/r2wk8mRJpbS6FIngLnXSJUO9QXeSOHsBr4+dOS
iIFpHEnVZQLo+M+dABxZxufVUc+0XGVczzOiIm+nnw6a89rkOo/n3klmSrhN3TMI
Cqt5+Kxhz+zHu1VtZ9LhUeumY5AiQKawHlKOW7mETcUgZgtUsre1dkNgzqcOAWqy
t6Kq+rzxscqqdIcpPW0KBLluDYGEnaOCHDmqxZ1KGKt9kzwuYDquNLO6D0UaWNWV
JYsEVLuixbpsUd6g6bYhnqU183U2cClWwjTfdMkHU4gKKm/ZWiG//4dhJ5DCKBub
lrxgcwj1zTdAUIRDjB47RkcKLscGz1ElJErAyuAZlL1HWLU25t2namH6bvvSGVqY
QonDZPalty68k4MV00McUO+5TNrOpvUNavEKiRWMRmJ5AT2c5NFJNR8jLhQ8osBZ
Icabnnv1CYHUwDsHgN7Y5BZ2xJVZpRbK2Zzl3MwCtzrSD1yY02vy0gFNiOHJDZ2o
b3D8JXlQMNVRX0Mx9WNFVOA67BImNX4IqYMXg+rot0IDmbLmBVecPxcEvuUYovxA
oNSc97I8tA0ehZq0IVD21JTene1vCM7WB35FkCHft62P7UlJsHF6eQRGgfu0W05a
QjQWfFwde9C7JfE0woZxMlUGYN3Zjh+GSxqYzmaBaa7M7t3t2HDxku/UIdoLI32l
ZIcPOuI0Z9nI5bDP0iFgTS/A1osQSchF21LbSenq+3L9I9wNWjgjZHTYBw9oEsk5
f/OIDUZfZwSdRAscQAds7vxugBj1gQJfYo0dXAHOXg2nu9h9i++nu8Io1I7/6KVj
ce69/0mD6+JgJvE17qAgA+Jxh5W8W+ejvo7oghwXEMFEGaom3xc28UpcjmUuzNqa
MnOq8OqjnfYAEIe6d4U/MdNcZcEE+XN0Onfx0Os4e6MydbOhSOgstvbwDh3cAEMh
b2j2hLWMXmW5svpdAP2YGwegn5qYpYx/q4ZD8emyh/33SoZraKL3cTF8zZqwheDW
VKafXGJDmTwFYMdjFj75yWikeBHooVHrrPwVDKdqRC8nTsE0CeOLYSFDDLACKwf3
Y7Y/tuCi/iSVVta/egswgQmNOWeYT0JNVQVQwEdcU24u+ixTOfq0EyR2+YsWx+Q3
Mphk3EehT9y/KvY1bIGdSC/mUXpg8esPTjNdnqtmW8fV3vohbTK1Rbf21eGvZEPx
kqToopF3cYy8BvX3de81SxsH8FpCDEHfl7IoQGPjyD90O0Lnnr/1TxD3SJlMSYw8
AD4HyarBt2ZDtAifxrCD9QOp2nVLAg0ExF71OWQjrNLIit6+ioKN3f7iN0cgRSkF
CJfFy9njWVJOmGpErPL9hMPp0CdNxQ+fH4upcEjLVER13NItbuufK/xvrhLarTHk
c70UpcZTwBt2GqA9OJR+6OsJKov8LmVEODzOeZ6rQV0fsnAgQnAPklVGFi+oMaZU
eckOv/629hFBUBhubwTPQTi25nqVqsFjZZe7SGzOcZqRFCyvbDu6Szn/ZGDZbNCl
K++maJX0SadsHDrX9BVsl4F4Jq4lJ7BagOknusVoP3Mlm12/oT50iPi9RRrvtmib
JCBkXA2yVhrUDwMpgOJODZi71JZZz1FM0QzleGrHkPHZVzrrIvW2hoxunez2xG5q
79PmrTqCyzOUO0ZGLPe4OfLQAVrgY5N6Ve+T7dhe6IAkkWvSR/lhUnz81y+f4g5e
WLhOR9Cr/MxZGWmyOY2MJFLkM7vPsXNhvBquvNKzHE3FsRVDktrX+2Bq7i01DBoi
Dci2ash4eoq00UnJ52ArDeUdYuzVSymODYDtyHg3Ao+xHmgDb8IVmJMJa6qcrgoq
dZGUOqDMKNiVVaaEnTUIBMB38T2+km8DZQEaPQBQ70taZW4Rr/N1+Zu/8vt38knI
M5HOq+AseNkOGjVZYFsB8NoaipzUc/d+rAE6P8j49ShFv67S6O6fR/cabrI9gPOb
e+DKFHVpPpUNzoyUyJCz7tSevwWT3zNTQZYQuqhjC0kU1H+37OrJ/K0RCJWMembi
UJ8x20G6ShFITwWfRrisI3Ww+hnmgtbY2RImylm3y3B3OB4yKThMHDKoKTnATmOV
5wh9HvOEvMEij1I+98K1Bw2A6/sDkHy2Q7fUJ6eYhTeNohNDWOsFU0h8h8D9Yeh/
uIns1ZTQjviPifv9e3IzUbyH2XCVzrPsV+J5Eg+UMYvLwGyIua4mTpsTRupeTHWp
/fTg3gCLI2ovAdfaINfPlH4UeiggpwxHsf08gQGzwfZ9SoJsyajsEMpooKVSL24K
79bw+h/poXQCs0+kcGBawjgPn8O5gTqJmOq3VNuqb9diofiU91YxRXIkLiOBnbud
cdYGmle56wgcPkUMhvaqWbDjeubKF8A1e3isj9NZmeGPpDx4aJiTmBloa5w0oESu
A47k7zrv6N0WuowJyEWSX/YVpCu4/Yg36lkFy/DMoxREQc+lLozL6+AXd2WrjoIT
G5OFYJQ8Kg7DZcGzRpIF51GttxGGtWAidBlbDJj6eRCd4lchxhBHiDPKR/zrF8LS
CJLWzYJgTPH7Y5WTXn4sEhTmICCPktJ8yna+p6IB/S1C32B/cjFml3XpWKNHMKuK
8o84cxlo3r9f4ofVEzjwqvYX4qMvDnOXt065OR2I7NRY10J4fVs+cnrshAcP2bst
eoPnFPNgXkc0yCaVyxMISE7w4u2A+59ZsOFO2yJlRMv6q0PJNJLFySMGmCxQ25O9
cr2KvFJrij8j7iUISuahJG5Y60fTECR42MJSEuwEJuXkMkIWXqRWYPuNAUoFerPN
foP2FLuv7eWy83JegLzdpW3LoDrX+yUQbq272XPNp5VIep0Qqf6LKMocO4B73uc/
NAsliTVKnuI1gZpMIaUT2xzOwajbobVCaCjW071SvWdXpi6llmW0cBcJ7EpFgdbL
pc4X4f729kpA4uouZbKhBNq31fMcnYkuf2uUHXU/VWFZBQVC/CgRQbZ5btkk6lf0
R/totGWsH+rMwvQbax0hPJ5GAB/S6fX0u76IMe4ZtnaHdhcBYu5WllNQNmQcJity
XfJTEiYOzFYLOftmwIPjjSBXURUt5b1UjxFiYBAn1Wt4eesGXsiVychYjQNZL6NM
UB9qx6SJP1r/fyXFsXzCFhpWuW27Ch+nE0+i9Yet631HH8DpnnqNMvjp0eEJKdys
zgL01Jc2wRCJFmRuCfRddEyVtQ3g5jZcgcAf+YLHWmRYVytwJHEYmSUL00pVh8Wf
8JxwuZNHur5/LGAnW+5ggJFq9THwpaSQM0rXlXPFee4osa1VzlXwe24cGKeNP9OD
ZLDoCRdv8lFV3Af8KVbtc79luLP8949vnJed5xPJH5haITnam2U7TlqnAq6rl0o6
1fTFMYS7aMjOAnaZ3lzu0WKKvtEtEu5O8R7KHRklgfmVlmbY0e5YCjKnarwvnnOR
XAsvhzc93Tx8m9rEmdwIei0gkqLP5jNHKBeP+5H+h3O3emurJocoYxuJQulbA21r
Ch13uGpI9tEDRH+HvzZgsR/tt128gNDKqobpv6o9FACPU9oU3jQbV/DNA621vmpj
Tmm2awaed2Egn04cwsU6pRnAvIfXNaOP9aIdQiUdCcYdQq5HcuUAEhfT3frJmW+l
G/TogiqPQMdQm6lhwUgJx2/Xc7kCtrBW6Twy3/jMvF5BJZzihXWUz2JyzQ1HPo+9
whj0wlqDJlsuB0y+4akifqdDjFz4IgPFavA0wIz0JWay3K66qVdmvBvQUE7gfzQ2
92ZyuWyZG0zll5VEkGlaU70KyKxZouATFzt5R2SkuaDPZrOVf94yKqu5h8NfHE0y
shnc7uIrJm9G8U1raUAXkeHypxH7/PG/SNY8yv7HkQlkl9bfSDiVDDKVETNQqx4j
Zu2nYg50ipwu4QChr2IqPgm1EdQ9PFV4X2yx1ATA/6bzw2OPRcYu6iWJJmZyD3lL
9ajSvasUwordSS2/kBVNxsAuBwnqZSpm0w+HE45UcSjxyck70xybnvLmpUewp656
1u5qI6y/Zo8KF38OGekd5KZ2Fh0PRIF6k8bmyfaj8awD9KQhkdQnDFnUHL6vKqLZ
Z+bzUYW76wDw2CsUUTB8n+EgpdaACJXB+vWh1S8QFySdrcEBIYK/8q1x4kXFFZAD
rl0IRMViL1874dmADK23qVALgI+dwtkbKFHGpU8JzwO3yW2YlUurZkExcztZIm6H
UlgZgOlX9JCTOehSpMzrATU37t0ybrbPxTQ5zYTMl5OlAdY7j9kA7Ow1FFUOdTp4
XkbYMCQaTwFK6xBe0pUKT7TKP+oA6AW+pzxFtc6XojuSNEnm1Z60m3+YyaX4c3kg
O68qiWxvIJDmBNiYMiUYQwYqn4iizm4bZjb5y5ilCpcWvfo3Ky1K0H7yd0Z5j4Xn
FMYZ9flpTRpg0vG5zAyG5PCY5xZxTXtye3l1IrYcy5hk9L4TNMwYFQJeaOtC5QIn
by6HXD8ZVROuEKXIRWHKyM07ikLjt9Koz+OFL11QRAxSEYsSFRrUEdfDeA6VisQp
O2wHeCwp9Pg8RqvU2Q494SQg3519tLJD3C44eum+VpImCiGpurSeQXGjBdOYRUrK
QLiM3T8CSDz0x1i36WjSBw4cTLNvkDsFh4hmarkXvzETKpaQkaXO6MFF65grLt2j
XnIJXJhgsf5OzSJITG+zcRdjwiot1/i7nIS/eKYbWWHHv7eRCWq9v8mX/bBmc7qh
tw0oOO8AyPJ3m8q5DEaUWMfJkOtViBvMo7uoYZ2ywKUo4yIFEyvbFMkRGrNwN2bT
s5S8iP44sQI9h0ebsZW33to0Dv0e1HYKEUbFO64HzKgZxTT1vfTTMCUaqnngyx/P
Wi2nvQviF1YjM2iLk9BVppLir7T+Ge0VCKNTmsHIK6rNrNIqUGAVhOFaq6IDI+9p
r+m2vagTY7AEGdOEPhCr83GJz/QS5SliezPB8fPIiDrY+zVSgPyCxShJFZ4Ga7IU
MjxbX20Wc+oxqyOMiYimNSvsoyQ9ZLIJtSHFGRtxEMeRQ+MOurhbZTHFIfjj/bkQ
OQqckyjbOFC2COZ5BDs8XRZzpImdGewgLkuCuBJkzuNEBJ42jyKGmvWs0A9+D2/4
a3uPsX9ta4Ekk7u9J9VyWGxU66PAmtJWMeaLziyygqL7226+sNJP7gTo+8s6wAOr
ZSRTkW/vhQX/B7LJe7FErEulpQquc5QRCI9O3IvDCxFAr+A8ED39gy2KvjzsQRs2
WXbDqUWay3VFFF8DXqs1Mu3TUnaKUszEVxWqKVi1Ib2q0JpC8BbQOyo4bcn9G+Ee
K4bcqjNqJV/DSQawD4V6V9q+1wZ9blbCNej0yycsN6TT7DXQKGEozlBpSIIu3qbP
DyrTlIn6c5DOXOUmLoDQlxAvPVDi5MnoNPvYe03B8ya3pPoAoftEBgbYSisT9+UL
H5z5FBIX1dN/tk0oClnpIVk1O3TDKenhf+TcnuI6EmR44JkNrraDzbgzEkSblzuQ
hTi1m4tQl8+WFtM33xOhU743QLQfgaCpKTtXat610VzgHT4h1VYMzSil7plNeSco
VjduPBwhvDT+cVmQ5ApjK/ROG2oIXgJVMORqp5S2MA2gi9YsMKrtrC+XevYbPZaV
e3yjNzFbBcA5cbry91japADGwjn37oJj2e53AMW5NrjXbc4mUO5PZO4DSX6YIZNZ
MXQ7miRiguhIT2/lTFb+aa+wr3MY4e6VGMoR/Kyx2Zp15WZAP1PiE9GqMgc8xZFW
oTEvB5jvU9tVhkIMw+SzjCLE+X4zfYHe3sV0XhGOYxOLvnYhhkQMiMdFGkTT+TiY
zEGev1w4rsioEQWHEOdzHjS595NJvLf52OKNnCgHVFK8alj/opsQ/pqLjKB3YQDi
3ahM9MhWNtI4SdFw+GHkQVHisNk60eqs74XBdKQ5d8+k2LIvSfsVzodDCevVxcKr
TPwEYc1cNfsMGgDWZctZNdkDo3e0Pdcd6jxIsoTvz5aALWLVrTstYDZAEzOKDHiX
39NfUlGRs/gADmd1DRholUD2SuwKI0iMJS45Up5ntvDUawJkWrG6vN2lnfcpbCpS
eufCI6RoRFAgz3gsZglSOUX5Ai6Yo9dfwnLUdSkBFtaPSd1pDus1+BTOJxAhQDhk
yOeFYNQEwSAhHmZEf57mb1n80tq+m9SDkoLIQPhXB0xS3OIFwDBe3vyPZZC8YK0G
0l/zTrJFxeR0QqkuKBUH+TijVye+5/lO28c4bruduXFVbIiaXk+WtyqtoCXWscdq
7MCfS1PuOLSWOhJGdedBoafa+Dy247baMzWZzuGYNffJVCFUwcoYLNwERf66aI3K
3VLLNLO23rzwii0wmCQpreio0YwKWJn2q7/Hv6LHsOr89GATAftKZ2526mBdHABJ
fEXoiCCcAfxpCixAFex1rumF9P3SS66baI7vNkEN85GqJU1J0vLRjMuw27GFEMae
ckwr8hPDjm/oC8/rHcal5RIQSrcww/BpxfPrW9RhoEN/2aATmeK2wvxmqk5KMKJ2
Eo6KPbcHNtHnomWLuXiu9LQ5EiIwCpNR0TGvklDE06pOAb84Ux2nsv1YvXTn3SsB
xd/+7uLpB14C7amkAHDL8g//Gm8DOq4zWB715knx578gNzyhQcRPmcT0wWLVx+GF
VlDWS1sPx3K5Ru1pXUBooDnXoi8LGfNN/YKgQ+QO33pwFJgnFhJbVmhfOnt8j1FZ
NuT69V32zjjpLnWARCEIoekZJUH/rCVF3jofhrZoV/dG5oY/s8KVTxGqbFveGnUK
QsHpYdGS2Ef7uuKYo0zFuVC7fWdLAuybMHR5bsaWNKQ+BXinvOFVuMeuTRUEiTHg
tqm4RJfEBN8YktUJQV3oj0JPcBKe4zyVN+DEkl0iev2vJpyOzT6vjMmpLgr3u01x
rgq0cPFApH8kFaief4NjsincxYVWvk6q3WxlGTJGZTKYiOjshs6e/wQnUtLiu2am
NfN7tGjRVPpqPV23UlrO7qjv3PEKMIRzTl3bc9wREixzalKIrGbT3IxwZ81q3jkS
kQIb3JIwXTJcobWT4szD5psAW1BVIs1q3IKwQpeT5KKxCHBkojDcWBmWOvTu+Jun
xHmMBRpQ/s+kSq841mhB5LfnI59qb6tgTnfAl30hoKO2Pq2fvuWO/OHbSO34rWts
X93mgIt8cLF02GBUArN2KgRtCCIAFki/tkFnC6iEjDM4aCqcv3FboAM/1cW4V604
9i6fDuG0S29SXl2C+qiIHPyn6+We08lZKJoXKLj+AAyZVR0fQ1ObvMsdPlztubCz
XRACW5t18R/uAxJK332Ui3x8TFCCQPwYB4FXjso0ByLEyHOE3efHw2CEcZABjhml
Fzp3C1KQbzKL6j7m13oduNAskk/zmT1H0zjCacVfFN1G30YUTZWhv/NM3rwi2WrW
3yaL1A2rqZvhGVAF9Esb8oEh6I8jBqJkkHLPP1pe2YfrApx0niOiDE6dqbfMAv/D
CkfkG5tFylYLuiPW0XzxBGrBa+Gs8yQiPfMwSQf+gPEfgpDpPSIxw2PO18B0BFrf
M4Ij8fqsSxdDRAgh+eFIkUVALNgkCt6nbAQTEYXFPAXyeGus5gs5JGa4Ky5YjMV9
Qep02TzRYdetnPB2TCNMbp9HuYOZdzqpcoOAr3GSjVVDWf+selP5xRtnnkJCqieL
poxtJ1A9Kt0qHb3wqoXOEmOY0f017pphCU5M9wZLF5Rw9UHiXBxbeSbHDKJrn3J5
h/28hyUD39ojKwJhPomdNJFsStCkM8L9KsBePBSBEeYWZ9M3b4sR9QiWW7JdQ9+Q
OKOIq0V+XmO0J2PvWRqF+S0UyO/0GheXFpJAf1+Vvooo4QjhH0XCEj35CXI4H0Tt
wmB4R8iAE2UiaqlWQ6v0MHGpqiKHLak9PpVa2/Y8F6cjXu22tBVTFsTQRKBp02X4
Np+Kx7LB4FtOhv6xGdMHDif8cmKLZSLdGLb5k4L+m5F8NQpCd3nThFKLVkCFxBgO
oJOLDxeg8ei8xKW+DM5wy7/w1NCkJ9RSq2D3+hierQ/S1Rf1HVUkIr6OTb7Jixkm
c+y/6bXlGrvywgup2oeBDEH1oolZElVyk+pLcVChDCYhNVJokFrE6VzWAOtv7TXB
qbF3mtdEJqPqSB4qOTthV8vI9DQjSH2sHSootb5rsFOAih1X/XL0+PX/CbvrYi4l
wQk5afOpPnvcRonM7SkmH5hPKxHQ61KEmIYU4l8sB6HJkfx7ofK8tSU1hCLliiwq
pxo1Qk6ZtpdZG+kNdNjfowvZePv+KaddGpai/H5RilluGWQ0jkK0tgoHYhv08Kgq
Z8tIzaZU9QRtBzePus92JMwVXmIBDI3kNCl6zHexxhM/879X9IhUSTzudjXH/nbO
LpD1JouZMVWw5YddMnxroCX2ksVjlz2d1fjvNlaBChL5/NYlBqISzXNx12m9H4P+
MWpCDEZLDZSirjJ7eYNOvh4c1RzmKHUlNoa8IBUBWw905fWrR6jMH+PpUwbqy39M
JL0yTDJHo3FdRP3tY9SDh/JZ2JPnlUCw6COmLoiGnE3Fuw9O5Ni91nI605/922HQ
vTbkMhDaIP/vWYXfD7wV/E9DFdCu7qZdY3bZTll60Btfnqj6tMv9agyAoMmVcNrZ
oQ+e7Eu6fgf/z/lwTIqV6aGIh9RNx6JTnzurtFdGlUVYfJ2aFJK7cQGKiKvM1ZoP
247OGkbAli9qfpbpi7+2nZjiMQFNI7a/2fG+UXI+e7uOhZg7dfU7DhGjQf7YMwZR
I0feOMJGLbvdpsrCmdTtjo1Z6Ujx4nae8s6N49QVj/ZiaUbShc5fKXyaiLZK6sm5
mBFRIFuYI+ilQ938Sq7KfjD7yWJxEpPHm2LTIA3jXiTmgeUP6Ioyv059rYXHzf6P
SJTSbVyCM+3dDHxFZKOOx0ZWQCc44/r1RHzJ0IiRurUXjXwwqrTcHF2eUN5rrH3U
orK+w/NfcBuOyvvMk/+WxhjMwPDK3HQ/WCJ7GSJ6sUvZ6Q3wS7nmwrwIIer3b58L
SnBvcHKlVFWSQUjjgkGEC+1+tVEHQYC2QD89Z71MGi/ebJfqW0EZKFh/BjOCEObL
xNv+P/6tCNzs/8jQZWJhXqNKf9T7i8PPFqbGB26WO58ZakFSWSeAGxSS1zhAImQw
`pragma protect end_protected
