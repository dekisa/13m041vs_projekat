// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tKIutyDGnY7g20kdS4tMiE3QtlGQre7u4SxpBJpBHuTRARhnzyP2+Cck1iSVlrbD4N85cleC0SgQ
KT6zWo278cbLVDaeFWfYeOnsUGkdWK+toXQfqiGfR/bqIWuXS1S7r/t5GzaZxDF8QyGw+i9BdOfJ
n3m3Q+orR8vW0URJBDQ/5Cs5l9b9KG1vnYfIAqICtLx4qSY3HTgiZrcB3sMqbd/A9scsezeEFuIE
HoCSWPgqDZul9CQQJ853UHRsUKwPSevGsccq3SrfJqkAtNt/khdPKHSdTsYvuL/FFRv4ucahUQ6A
ASEnuvIqSe9Kt2cKTV3Aq62YYU4GBIgbnluP/w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 39472)
qGIb7by7j9PqKvfkXdwVyCvmgB1H8mLPAcsOF3WGf+H0KR+mQpRCSf1V+jFNEOdiWY4XD6cv7X1N
KcPJn31XdC5UAmBuJxbMhu4WMsNsxyjwmxQdhSd9Liu+JpgoTngZRX10H8FdqS9dboiWjxUug2EF
hLKSVFmqoBJ+Xs4TdBrc0PHZmgMjGzuSBg1HQ/PHtsKJ/tWIEt9MVlfu2tpoFP19UKaktMbmklwu
qbDiSHXapLw8OT79d8Nx+hMC9D3k0W2HKmLs927sbTTY13BDN3lLZDbCaKi4tSho8IFQoK/8IEEO
3Uc/BotSAsBMaKtw6khB7aOEbw/UgVAQ1nyoUdOwtkDMh7/frzdadFtPIk1fXJ/MYDDZR14EOC2X
M6ZTTvMGHgRFHLl1yWL85ui5d4fZ+eWHlUPgafr1UlRNiUu/uZZf0pCA8IzQieexA0+nEJ2t0E6z
jy+Q5vgkFcDHLS8w2rdz4dggmsbQwKnpsbhg+4bF1yJAzjIADDi4E7BV8xHLUqCW6I120VwMi9a+
Zt4LzdIAHHuQM/HUrRFuruCApijrKAy89tcJa3d5SjH822zJQHNWgs9OGE7+v+UpUdr4K318z5oq
9czR8cyV7LSOYEwVsx2XOE6il6oIrQJgcL7DbbjsOtX1aXnRZ3OGMYVHx9fkt1nODHzALtc07Hsc
yj5E8eWv5qdbAuxrfwkG4s+Y5xHFvReftA/uWwzC7IR8dmCH+IP2BmtLlUNTk79L3RqRmPwZYiBf
esTprRd9QUQ5M/yNlVrqEX1XdQHU46nXeAfh/UIBpIFxnrh3dyrNIF7l+1vdcObKDRBb3oPIbJUu
FcIcGI1FUNd2AuC7nzD6JVHFG5BijKsdlufdB5g3St1Oyk1qSb1bjCUbGDGjdv4ow9iWCRgZ8fLw
ouZMIxgV1QYu0OBsaEX+8UQJ10migLyYCm54qpYDfFokG+c71naSHDbFK9dKlV67iN7jNfql3T4d
Edl4E37KTO8hMkzDm9nk89opTRYlPs/mMTa06IiDjpHfCluhlBqb5dL4KbETvqcHpOlGzTf5ZuqL
uIyEhJ7JSqUatFrKKg+Bu2okONC/uuiMP/OyhwYk6le7mhYRe0xbjzB2g8Uc5ST0+UCa5Imr+7xi
ijgqxYjWZdZqT3Nr6HLPvjWjWYyaxvFZmm14HxwhnUvXQ1cm8ofEj/IBethUsQuCRb2G7C64ZDMW
5HGT7DEM5Q2xP3D85IE3E+55k1OXeRCsfXH+0AqfzHj5SAklC0Hk++aez6kgsh/yBe7Wv5WyyWIa
6jcfkFea4RopFvZaswipQnGSNcESmGhwKeJ3Qk9pO7Ipq/7c8RroDQfdeSwO1OgPuFSuRm69RXdc
tzsCfOpdgGf5iotpGIrBgTpwNsea2LoANME+raD5evlRs3Sq76tpt+5E5kLEf8qif05xpC1vAkNB
SbyvB3qH7drWb3YhPJS+pK1KpMma+vZ+Ar8nTTzsk+H/FdKMgrDiuhduE1JiCybZNBpNUMfl/oLT
/DrFFViwoXLmNMp0YKoHt5yMEqSuNh+dW50E6occ7Tez3ycwc7LJoZJy2kADnkz3z+ZBEyxvqnHQ
gECa+6eQy/XyPkIqIYCqnFhSS1UOpS+MvsA69bph6C9JkyALX5O+qxwnR2/TGJeQEVRGysivKmrs
7Q+YZR2q+pbsVL0043+NHUf2LaAyskui1R79G1HKlpxOjhhcfBUabYzYc/vJ0ZR2nZJA7YeYX9CG
Hb7bZL2l04V0x/tx6o49eCGZ5JxlzMocyonJun/kNPyvUh411mHcv/crqhk7e07G1XrDqOYh3Vj0
Ko3Opwi42qcrFDPp1L95f+80+m6oqNTCtvW472c+PRkvocALDS5a90v2tpkbvDQhLv/Qaik945BG
EiELY9k5817u0RI32+JjS6ZXNeKJxGCWYIC6JowNNlb2HA4zo2z4E3zdfxOYYZAYbIL7IbvKnHI1
VbiTObNZ3M9vtDuaxutmBoii8WqUcmIU1JUxTIGELWgR3uVY+6FKgh2gTIvKBvk+hbKg1znmAd6k
dAgtbvAIfZ2qUR1AyQbyIFZi+0CnGqJBVbn8UBWIiWMi4YGn/F9uUM7sM/RwHnyVyIX1XEuJTsrE
eBoMeV+wsaTShkJQImOGfxEmuEnV4oOprh3WQKzgSw7gpjilB0Q95eh7hylLZYTXofigTDLcAT1c
NakK6kMECKHyZ8Ee/jUAJoEInfmNa/bMfQBWL68O/prh5h5GjB4shmpqgKSE7v2atNRdPyQ5i6uT
Q+eODNCBf6pAz6c401lmkJIehEPUn88fuZZAoqXEjiYDqdXZU/EhC5pNdgVMK94gliLLO/vW80rL
q7PWfxbZDjvCOVn00tYQ3zHY4GDRoZD9B1RdEHHznFaVZpg+xVY3gnZH8/rBVRZZYhJIjzTJKtww
43yYwtD/UXY1AKSjM92zqbmC8HPUsM6MEFqkgsD7jJHKjF1oo7g1Z13uL19SqgDIYWGutqahgUv7
b+kbofkcGdVprHMuA9z+DbMKmkAPalC6Tw9V47W63kiOr/In4Cook+0azSyZopA9nCLpBFg4SYa7
x4LYAA/ybCUMkfUlu7F7/F3xIaR+kpWWbmt7tsg9uNHohxWQFbnSFveLos9RyPYAyvoPq7S6Sikl
mMi/elfwsCsyxypKHXlqgMJ8A8ryGQPMCNd/X8vzApthdRzHPtvlfF3qliCdN4wuFm2jJ+lbvZuu
bTAwwOtYrzdyJb0YhDZzl80Jz0idYKDeNs7EDHpK9JEDih+6SQqt6iZt/qMTxDeQpAO9bQljHwpu
nDr/CrA5E7JzeCFQOY8Lnj+kbfLmhOjN/aaPz6GPIUWM3dzgYuCjl6kTJSVyLhYNGTExTL4A4N6T
yWtoNMqfADIzqGrNHnR7gaF8omntJJQHDQhrGNkSrXY+RlTr9j9gRz/YyQqqCt9g4sU5AVYVaseQ
6VfND++RZaAWSiQnL5oW0Rr9pbdR5qFwfq4XO4BzOxBPYYHMuyTyV5Fq11XzOyD6a3d6Hdm91YYW
UTuB08hva4ckk4x1xc9EI/ieYasE05VhBWlRhbeiGG1XBQzuAQ7zpLZNcBeHnLIzq6ciMk9DH22m
4ErSLvE+hE+0VBAkh5EMVGy3oCSfPInzTWK53Y7FrIDIwLlvAaw4csIMsZmQyu+P3+4zDrPiZ/8E
jnVgGuv17uq60al6yxiQfvQgwOS6PXos+sbOhqS1z6wRCKqIeZ/syp7sa3czcVn5XWCYnm4C/Uyb
GPb5AimMcyx/NLDeKi2+PidpQh6/10AmCdM9/DRFx+ZATSNlvE/Bz5l0ooTC29l2ynudLT8bpup7
zxG6W9Skq3jMXGk9VPP1ACL6flxqQxNanhY912yaBk+hPzq/xnEzqQrM5eq7+3SMBZfgVG1SgeS5
o6rEkJc7lWsVRU0dXrVyDwsn0Opagb6xVq904d7Nfh/uiqKIDZ7bHA0WlTcL2LP3hBWTCl5GmIAn
xGTCCwt+G3xoeCYRtVgDv6hjhDy1KXAt6MgwZCe6F3ee/TbEoME4Zyft1LZVyq1pY1UOIyWEUhrA
JE2nvClep/AQTPrvj9cIH7aOgcDBn+6vICzi7eB8+Tp/GIo/vzh0kzOCt13byefX0uYd1zLY4lxS
cbHgvbDVig3jwhbj8kfo819VQkLNCHSZFkswRpanmBwe6KZ01mllqx6ypMjRcF0YgaUSnODRsXLW
mTFhajEuUr0L0PbwptYzNSNWCCtiT40cLgZRcUe4ieyZCIcAOlM5dzDimAATUpvDPjBOsdKqsfdv
ZX4vRKXDYFB2CCBSVgj7RlQgoLGw8s/NO36xFEaN1wO+GsRC75AJvBsTWkwNuJJ2sE44ERZ0TWUr
ylYW3zZXFd/VCcHaai0dFKRG3v4khA3bQq7E+F64pSGwawWui8SXfResQxLwzfzImXxcmkPCudlf
cjX3tYZ1o+G0J23ADs+k0tuBJ3nALwVv7d4hfoLNj9UXwT3A8Uuvr0zaBFSxCA2jvrxLf0tUND3Z
F+Hl7MaAYXppqorKil6o5BtrQS80S7+dhBD4oSt18fsBw96WSjGssePKdgKO/iZS25nhAFcKF2Kv
iLWuQwUdtXe+zat4KsD241Bz5gRfQi+pJe8O11w0M4G48f0ZiBcfXO01Ly3JtalvnGd5RP+psouf
pJ951vjHhIrtXV+kXn8PpljZkVIPB+Xp5ybcSOwglMdzeUod3foWovhjG6MFdpAxv5aqKB7FgOXs
iIv2mwYBaHWcw4w8LH/QRoPOkrjRpNqNoW/IVI7WsJFU/GxO+m3lCz69Wan84VEc+W+PcEvln1wv
loO372LK4ES0oCgoM+r2mG6bDzz7H40kvi5uAUvJ1n+neTWTNMUH+BhcyLvE17TA/BFco8uDwt5K
KWZUeinAEGUuy/I0mLWs1nDAQywvXsoia3tporKqsSsZ8HBAb7XVlFUoYo9PRsPhCSxpaT53jK6H
+H/hDU7IYEZCRUJo6NoiUmcYDR0sop1hLBs8NbK+2RFLFtc3oXoQetBT0Tu1VaE7OFwlMZjT4FQX
gju5YfxQYLiQ0FaFTLXjtXV/Dw705PovFl/GCvwqJX/dIT+OEKaE7LAhrS7KY/RV6o6DoUIPy8F1
rjU7VFLasaBZZMexZgwBAzR41sdN+F94OUr16DgiTWpQqUu8tgeaY8BXSUZx7Iaxz2UHH4sYNJNC
+6wGNyXY8F7AiXgSufEfx3shin064dDhUrbDmSFtQaQWeRHZet096EPlZLUttgZNhiGQ33tUISM5
ljnXnVFAHgwen/DVBTj5vWRsKmnEjH3eLMgx9CBsLkse8lxZldrXf35f9uLx2+6pVHLuqhDvybO0
BQfpr03RdRE/K/nKmeoFxSbwE6WfjfFR1LujY3nykPlqd4wof6aSDeYSyz0oyrF7DZy0Yn0IEiUn
DL5Sizt0c2optkkQftMBa3V3R2nhOmjuzmZUILhT+hRvg1+2b/KdsgHmPLGw7DWF9AFRVxNMgrsz
W3tyqMj5NowFZzdfFRzJNIF6Ea14vZgAFca1sY9ff0kyWbNcB97fryGBFgRsnDOb1m103mYxImZH
tBH1UxxMhUmHCvaDuk5Wz4HXVzrqdKIbQTxvfI/9IJUuoLFDYHG+HOkJn/9iECakLK3IkhzuDyZA
oaxwns43svapHeHOsKsOKZ80NVf9p+85EhtnaUQITESbLptzKzHOQ2RfjGIO052NDqz5osrssmSt
QJMDrel7/4I3Hn1sp8FY7WEJZdyxxOEQNzAFWwTxMj9h+tvyllXuyOFF6TM0PBJ+H5GYxVev9Xc/
mQCWC31nug9WR4KzeW9beOLsyxeveD8TbyDgdyzid6gofCqlRyCkIvi//MwdIfX3j9S3lTbFfB7a
2d3XYIM61efOCuf2kufk5hrEjbwzM25jQZ2NYD4/Nu9DAKblJ+889AgoD+kS/kz+Zpx9/gYqp3sh
3xMi7sSec4dlmIgmKh9kejoovWiD6Ar2+hF4Xx++2D7R+l8bSqJnekQctZBVZWOvCEDVzK1kUpD3
UULFMLndXvRXcoW0NiQVjwXgmrDtADEYVfkvK7E69TfGwbcDj+zHPmqqSKjHXgOo878iD92ljkoV
PvfpjjmjbC/pI8QcrJnJUhJ1HhvBe7cQJzesOvd8QjQ6S+NSJYq5N/43ZMahwDfnqh0yJFZAX9dl
p9c/jfrRO0IfG/qoUS0OchKZv0qWqpmVu3ALjKgY1l/PKXyQOaQL0w6ZLP6eofYKvKaDJRn0dVkh
cJE6xvLTPHQ+IER8UP4Fb+oD3fVJRf4Nqn/LMpgXJrFA9oFGhranBChoEqpUWXJvf2l3MgFArEtV
aG3myJcjTBCj5wQXOeG5fFTWEdUOclL5+B5apUDSbJHv9wItCLi0eUdIx582o60ATomi0efYe50w
dis5MUwQ04VUNypDdmTLJeIMb6E5Kj/RE7b83wm75DcElC/pHXeVbYaIQMzROtjDC9q9Y3aD2bnC
1SkodB4Wua8XgD/nBrLiXO0gOVRWWS03IgICCJJlkGW7WRnbPGEcKr0qNjkWHIsuRFow+UmfUCVy
y4lUuoVGHpnT3bXTMEXZbzPqOarSzrmLMYo7FDFECfqvnErP9l0YsMjU+GRx6qUK+oMwq6Rh8ulM
Hb+vh5RcksBw7qJ1E/ZDcNrO5ulIXbHRnFohKrz95lWfO70VC4EdyN+zp6UuU9PG8DTV0RJhQ8SL
xHr+OEYrMBZFWRCKIQ4p/gXgtaqAB4Inme/10/fgEo3TdhFXb1GJGYF/is9REJ/2omDwThbXG8fm
IEK44cnf07Hc2qsIQ5CNX3k/Y2nWo0hCDjiktPm2RsDbmM4VEgB0OANib1xo4xJvxyLvsyXtYnR3
G1bJ36rM3YL9Ubz8reevwJyxEPw4fQhcLJDY4AIYMeBg08t92fgohbGvngqsQpk5FfawFpTJcsgi
XtJuilDT031O7IBAztHcZ56+I7KNvmuiPypdDCtICnXNkYVzV8bqQESH4/tn0cGUvRvOdQJZtfii
ZBxrbY0qoyLaKOsxOqERUuD0qHu5aGgOb5BS/+bKEj/bJGS4HiZjDRhp1PthFwFFQ45EpCiS9tMY
fcoRkRcaEE/TbdkwEHNNISQDU6oTEn+cwjg7zyHDtUM1N9Y0sNHaareXP4ZP0+HSQJRxJ7FymdDk
/y1y51g62AS9YqKFCX9eJSE70SobgMhGkmRTWvHiiwVGjF9Ik+bENuYOnFvEd5Wbm1BaG5HPgXMp
pdWUGT0TNrhHJxboaWYQeJekt/cSikTatRdn4SzLLipl2VZb24Lvb/7Ax6FjQdeQPFyzAe6AVjqL
UbAoXUnRHgvobMAyNkM2+eO32DG8+NCjfaUBsZzgs9/qJ84Wa1Pw/BiytZJNSPIZ1cDsIzOua91K
eMytTrkqcaPFsFaZ8EahBZTIm58LJqlRejwnYSSNQT3Yoc7L0RGTvG6XAe2OH1tPn4viP9K/YUXk
xCMqbJ5vSF7a3e9gJFlecFoZVBz3sNEXn40zr3D0YpSY14BHnisnb5zjWvGT3Dd7e9+7WlBiGEkj
L+zs2FaREk8HccWcagOXMX/Hkmg+rCAN0GZn8yetOZm7BEY2gyNqi53DSbVVPjEtxU28Rf0nrLyM
vuYJbCIXmrI5Bpmkhn5UcamcSBWkaW9TTD/Mwy+v0PeX+R5LV3gllfU/ZllEhfR8QYxwr+SbQSGj
BwaK8fzyv8VVA8xCmWE9Cch8G7AD706DOo/i+MrK6dDrTt0T+yQ6TIK/1FwUWD6xPq9ZesdYyopD
Pia8mZtH18zOyfHZ5b5IaTechGLbkaY3SMtPbgDIijDg1i+gAq08O0+Gue2pGHyPnCqHeVAQnTwd
HFwDWzMVEqfX756QZrWzw1oCADrA2TzSGe9C4G/QVyWe84JFeXBgg5f1PtrOvDPOBXArmmlN69Nq
plV7z6TxtyHYjM47TyNVTB1lOhQ5bSQyYQzQHQVUBGEbsyp8Or0lIX8KheGtsudmsRcJjjWBB6JT
p6gNXqGw8prQRbn8mMGqeKZ8BaCwNvLAqTDxil5MNIAGHuCCYrtDEAKVnGg7+cPCb2pQ0ymoo2kN
LJdH8zoPdYdOdo9/wcVnqy6c0UHHPHNv8gS0+tWQv7aAEfuCAOzZMK8NjieQ9jkxJsQ9WazY1xak
FGjk5/1XVOuJTYLTkQt/EZKKg0gtmh1dS5JhnOIoMy1wzZcsY8vE3fcPiFkBcS7a9LqJwFWnNRkr
+AaLsIC9VYbFkwyHUciN61OeC33aDqxdOvKU3p/dmwzdKxr6O3xv7Ix2k/ophkPVEPllu7hRpdWb
or0K36vbPmuk9KoX+fAr2ZmJHLJc92zhdphXW/rf5TKJTaOQgQ/ppGzDiKOOrkMF0UQCH5TxqDJF
FbS5Rqdz+VeXuktJNocALywEJDAleJbKwtClbVKVjgaEY0ZuXw6YFAFxCbPf7Xsb4/WK88JJocrF
Hpinrvu1bGMKVC+2aCq/Y387fV+luRU+8hNqfJmk1ohUljbAsxfIMzgDDyTBNUkqP2lIWwuQwVqr
1sMCiFCTcU7pnanTemLoPc3i6m/Bc1PbPw7IFXzMv/M1g2kW24yHRPAMP2FfumWWirBPG3sFlzKq
4yYcxScxmPnochL9SPjY4aBq3cMOa4qNNWYAmBgc4XINmOIrowRd7KYcJbiLXcjlz+YfDhixe1Yt
o5RTE1cfhM1+sVoz+dzvra5ss8X4YmWz/04ro+G86o1kXnm+mvKsKJTcjfW/REQlvDC1tWoa5QP5
PSy9kiJ4LJAEwUG3nTxpgWKFJBVUVL0lZQL70ip1nvFtkAW6N6eU1ZYhsuhznZhWcBk6CY/nFdSP
rLeS8znREk5M7ZoqdcMQIlvq4g3pBvxNuTRsGY7L1PrcQQe/iExkLi4IxqWa85k31by66r2AWQgb
eD6smR86q5QGF9/C5e9W80C4D5tbNFnSR2P7l/TnKSsi6V867OOVdIcBZMAuMjN3aPmg6u9DXabt
yYqDFLDnd8At1COHCCyTfzIlFDuKqatuprQrsidg1LUcH5OpIB7Jz+nknrLfod/uTJ02uF0ChZrF
50GPWYkxycgEHW7JTHI4Fx0rKWGThH2HYXd4N9hh1v43PYvsRZntsWrMxJUdEX+Advxm/e/bC7y7
YZQpNPRcY09MSLuIXRYPKAze9q5IcfDUnZyc/kGGfBrgyP5A2xNaAyEZ2yHKS5hfbsnB8Kd96MPF
q1LhWURb17bcC5Tne1saARt7BMgY3AD1cpi7sDkt6E17mmKeO+JfT7vGttMZCJrmK3PQU8juDHiA
gwNqsbUv99l5tNvwm8I/sMBqG302Nqy2DPL43F7HDlgCF6HxOf6jWF3BEH9CDY02VDP+G4/vQc8a
miil7lKRreCgrutoQ9xkYeapOj70ch9VzO2Sq7ogPTZEblxYpbEZ5XZCMAAlXqh1vlMqOUUowjDv
ZwPVjq1TataWCwoN2zVT1WfjGnZYcJK7tb+ai7nu+X0f/gcrCs1uHigZHrK6j7WWF8fYo7qhmsgC
79DMUWmBj3RmVbJpZL7O812bBvrBlhCBsaaCJbjZvXqZ9URQEUdxb24VwTmKIt6Le4M1GGgyRkIj
7yVom07Em/g6+m54wfWyK2iyF6ohU8bgyFotw04J+XrYa9xeEWyXufY6gj+LYZZ31SkyvK8MOz01
MrPtZi/OtrM42lGV/cDxIvoPkMIZPTKep2YRRHtP/6WF5vdpnLva8RlEpglLe/hd/IGgM5CepiHR
Xp+u94Xb2fkATvXcBTyeZJg4m1e2WUsYpDAIvnDGbgkZ2o8kXmIddyzsuWnM3UGBZinKq0pH0zmk
8TUNuMsEKzKmRKSgbbZBC+BJLYXazSdgDX1gvlp8Hdiha2V0wcC+FT6sQ2a6la8emWuvH6QL42p0
bBMXsFt+rtnKku6gS29R5ukL1tMAvFkRsvmDrBlo318I+f7G8kPPLyKxo6XMiZM4bqMI5qnlh2C1
R56TKeBJvqcS3UQM0sshv1R+pGr6R9D/aNy/k8Ho9dxp5l1hdoKxWEuBMH9FIJVeUEJg9YQnCRoY
Q3/9B6MWQXy/s1jz2r5vxaNDYrrE2pPbETRm2OnWEj7pnDBLsch5w/GEfjV9NR0F3IQ7AZvNaaU5
J5JzdZBJPmFUFAEFXGhmz/PLjGMbmJvYZXW+lXbgSKyoeoE6NK2/+yk41TN/qkM83jrUSsG6Es1L
MhuFtdncDCwXOEW9yxxeV+u5UMOuh2B47fdAaOkOnCNVJzX2QchP3/wqONYRGWdeZ8UbX7CGOczf
EbcYJQmEQVU/kjGNHNbDSYGNJeKcLV5yWvKEBjFMpZ47zPOrZiOWgCHNO75mekeOu75DzIkH3znp
gZbCL0bOZSxaxu3wewQ0M8w0UnldXSn3yEfJwx6hBYIx6pHsdsAmpM+4HqV0LSHRVqta7CfdbM3l
gJBm5Kur5mk3VkfYiqWpjiifiwmuz0G0VMbjY6cM7fDkBuU6A8+Pp8zaLZ45gIPbiFHpyVGhg3U+
1PNF9T+75Fw2wbpCLt1qog4FW4xHaOKqW26yeO1L+GkWEzg36UiidvzVkQIIY/bTr4xWaMXYmmFx
jTztQrDQ/pNGPZn1z+8Ay5wEV89Px0HtnTIllJUz/sy9CKf/v0VYdgi0JKU8RCGr8jOLDq0+dK/2
Rg/09Gk37NslRKcGu6zKjmYbfZQRocmtlrYn6Xfq5pnN87rx72pZ6XcgS7/yeyH/1ZlrfDVOdPbG
drI78dfwxgWw9Zf8gaKTHqBBYguZ3fgTeS75Z4XPNFosK12iA93ZF+mtq4SJ/R7U9mOCB39p8hYc
eRDSW+bP/1at1mARlA78yp7S/j4nbEXsUEoYLYkowX9wxM2N523uK+doXPho3yrUdCchuSNvkhhq
YN8UpMXzZrcYHrt4E47wN2PbzmiVD6ZOIKfujp1n+zUcqRvXeE24BuVZ+rCjOPFy5MQ1MHSyt2XY
OTjJUSekwyqtJKL1Bwmt/c65fU75LD8+hdThw8HZ2X1ifMA+SNCTvPc2VZODJH6RSWpuGT/zt56I
RqD/kgGYifRROcP7D2fVdfdWIsaqjhpArVT8lhX2dpkl9xomVpqL2ae9+64VvVCw/aQ4prr08xdc
tegAXDKXW8X1jKBW/3BliAvSeW/uOq4b6lRW8aPzil6ZXJVh1Jm9lKeQUpjOqQ35cvsiPkRnFzQo
6+/W/MNFTZzsm0p/SA2YfRI2oDrqXktQOBH+wqlWSgRnPkrq05M3fmd9F6F4ZBq8TanQZUvQLXoF
KocoUgJJrjj3SMX6sjsfMlN1aAp4vR8HaFAFgDnRjVlRQ01SU4TKTv87pXbGnPFJ6ZPrqi3BT10l
88RZLUqtYoC2reWxS5K0WuB7Xa7v0gvS9Q9ups4HllACJf2YD+koNgvqFPvw5khDKox8pSNjB9WW
2v9ZjA9xNiEhSHevsD5fd527stobDmAecjwV7YcBRHLTOcDAqg+4d8EWW7yJxMzTQRRtGDL9Zy0y
D5dYW8UTVuPXtjXq28Ha5UT1o0RA4ZW6wtvsxqhR86tNSCEWZZjItbPU6+qtEoCi+5oIGXeK+n+S
2bltV0hD24CMHIIJHjMaEWFecMTRn3zNDVUVbIdLe//VRXMAaad6DRNadjz1h5P1wdixG7M9Kn0D
DJpD2CZCNO9Z0B2wrwlnDXkEpzA6Zl/6SkqJAL9MjB4hAKudBFkDInPVv3wIV0qEDZceXDw9EYhZ
xskNs9Mxg0Xv/ayhQ0Bz4XhpxhAKZhAQl1ls6NSphs3rN4T6gGtcYYfsOwpDjohRCeECpWiHyycM
ED5CdihVdU8rO8s4m2+xU45+7bSiCTfa8R5KEEfMdWN/FIjsSothJY2r9Q2L0kC9QKrfTCRr6oQu
RFhpMncFPNqZwz5LSJe613LGw3Fgdk6RFMmDMqitiUJcshTgNELf9mk5GAryATz2JU9Ubq3TK4YH
+FQQCYDX7ucKVZJDzJbfiHPAZr7t6/bv6Hd0Z2r+RHwTXqymUYmRUuOGvJbHusJxr9jTkVUSKr91
2IxyR3iiLlnO3lrdje2MBvTySXzkpdecMRPYOCLehLw5PYZ4q1e2cYwrm3vaTQ29OLit8lIC6RKF
7bO4im9vV3W+vHfuJ3eTlM82U4WV0MI5WBU5vL7//eB64s8BjTkof5+Zzuwt/jev77KNayDNFBX/
Nu62RZzwnJk1ZrwMox/rZN3q7lTYkJjgDLRihau2wPUUescWzZgcFhZ2MUVIJ3S4QYdMOX4Jy35G
kRinUtSkkl6u0aCZPJPachmzeB9D8wsmt8bMT+A+t+1nDYNwLL8m5s0lm91/uh7eELefW0VSue0/
5IoB3gYMswyelH7S44DXJBeZVqbCPAxWvJdJMhlL/q9WWvCB6RKR+9kiPO90i/yUvwzN4DNtLWKH
u368iMNhPFvQMnkzjRGZpHDbdNfzyzVlqjOIGq7ixpwluQ5YA6JiM00o4QyaI5OxFS59lJsOCrLr
9WW6eFfv6rfjHSYDg/gt+H2NhYSqLQfbLNxmAzA0cDAgLMh5LA4mhR4A0NPuxxQywUoFhXcIIB8j
L01Lb05GtbLSfEcUNworJgT6TOZAc1CaT7GyzxTR0q5KZrqrXqWKBap9HACZ7YNEEEgu4PqBPEp8
IEuXDqscUIW7kJZhqkWcNpxi/xf/iIel64Ik8hv2CxmHMDDNm5LNF41+POR8PJ1Uh7uKyOm1RQ6O
mwDF1nOXCzzcMi7/0QPOAOmKCKKyYpqd5AmY4AIHDXA56v2eAekMuceCZIyesC3TobbkzX9nqGln
r+y61WXRhPGL8wCzPPdxT8JxVjG6vmZ2Bd+kKc1CSh6U0OFz+8w/YsPd4izQwbeSXbFmqEaRBoia
i7XhsAuRDtJNVC5rwCJEsAZR7D8OmsXLs2AEC8FipeH9gXZx/R5Y0PA/FESj6i6nkZQ4dHDAX524
4i2d+x6EYMPId9DF1jpDQNJUN6HcSV2L8HCjq3KmiNqRx7gN924k0pr0EejjVnQZZGCQbDhVe5dm
cR4izwU0cjQ92Z9IvRHYl+BXn9rtCYSMF43QRxSLFUBhNG4lX/V9LWLUGUdVDbKe+x5sUp6cUN+I
d19dgqjcNoyKdVMAPAxoAq3uzNEwigvBjXX1/NiFYJnodjZp7ann57U+MDZleA3YchmcChIqZJDP
daUeRpj2cDYzJF/QVhW+UpVQFUFGPuibQ/zEAITlEZnWQ9CO2rb8A4Gt8FoBakj5gLqrwTsaaj1x
4Nz8Hf4phzBpUJE16VNGAquiwFRGYzp72xaPOYrghATG/6ieV3oKwwG/6cERXnNQo5xD0NnQFaNa
fMY1F6EF6IBaLqueWg2rehSziFJNEqZ3mfkh/Tb9k/y5CKO+xfwt0IfvFymzS8fzBeM6WcDoUHuk
OvbcNsCIK2NaeHTaVqRNCVC8oSTENr4r/NJKoaItmxvCkNojPKfBaGGNqx//xhaCqLtag2vwxYbJ
4FwnKvE+kit9fEQEWxn8ANsFq2ui7MutwEBF6YYVQJf6xLJzHdlc/aTkRLNB2edtGoArMGyocQqv
rzjEgAZpiyH46VHAlsbqpiP4Y23tPQNyRpsxHQuQizk1vRpbLF7lmSeRAJt7vCgqA0dM2V3yZAKG
PmzVk6ljCFFCRDq3e69GovX6zEtVp/dgnwc6B9J50t2SRdu69NDkuloKDtjNU0dgJdzrLDxpAsKO
Mq5jdPTllmX8vV+L98RO8b26L9JgTiqOC6dGe7gNSs/cNtoRPSZ06e0wibWe0ClRTdBplaR1x3xR
h5oS0FSRKkvlsuTB61qQz1p8CsCpY/73Y5kAfQjAlNlQtPL31dpVtWcE2TZ8cQY6imR1SS9VI2Q4
lFrYm8tInFUTdgGjiwjgNwS7gncROWNH/l4+VloQAwolkCe/8iWBFM5UTIoaEKfTsSsYCuY1LZoT
WkImO31ki9QO900rgkC+GRFBNjFXRgQ0ZDuVpYRdokqXpPeMYB+OloM5s5rOq76RkPnMEzSdeLpW
zZCTNXjMGHDDhvUYLkv9GMHfuLPdIb8pEkIxCsvR0Kz49/KwvylY92fV1ec9+9wi36XBe58lx/BI
x1s2gCBORB9qT8EYYPUIeKjD3w64l4d4vP9InQs3uH3ZhRId5O9VvM43TW+mroFOCETcqqmsR9i4
Nsm2azj1ozMYPuKpmONr5v/BfM5N7jBuGMRKm8+h7tbNUF/xhwhADh7BiDOzDp4emLZhoHNFGt3t
s+EFdhYejGpxTC5/OZ9O0xMmZFYGG6HjbRGqYtNoq5pE9B7ETT8Sfpgsy+Ww7lTvmUbpbRdG3VIB
/0/dDid+KnCSLFRKT3EHJPqb8wt2RKamuLNoFTacsUG4Tdc/L/g6AVfu8TGFMyRPsueSgeX/q8I0
yTYEdIukEcwDNyK9skH4J1+kF31p8WBvxAktTGiPsgz59ZCJJnYZs2PwyuYn108Tp0wyhgMVFdo/
eXhJidu5sxNfCP5BjV0ubVe/JkmMTPjtDe3TUlxfzmMvs/p413oOQa8wuIjhlLp0xNWdn9j3/kwj
y/g6vC7Mvg1cFBFUDAHb/HxE/ybBuNZgxrl6uGnM3vmcFV6xVNHr2faibCewLO+NAMJdVXMmQ0e4
IJ+L8oXMsAxIzLh8HkRtF6xefy5whvUHSMVmirrt73YY9ougrTPq7MuWphJSPdxfmm6VWSkb5dBI
KxJ6WmMYc0E7eiDxiQpMtcS0+BKWyV+d8nYw4pmpAAIMMH0ljmdnWXXTy7ty06yD8uiSvVPviezi
1hTuDJiRe0FBrAKVqnOogA3d1UJuDmiup4mm5Po8g5wOXXOHMb/QC0/isDuaZLmXevGoviHh5gKX
iSw3lAfUzVtRtEL4r/h4z1zc7fiZdawY+O5us6wfUxJDCJC+xY4Oxd9L4YhN7K9T3Q1rXwRjAwQq
7vZcSa2fiRSRzUadFHl8OSo4SJWjlaQtvFzjARiO/sIRnrHB31FIxWYuUfSHvV/PIZhDPQ1aHQ+N
uQ+zkCg2Lk6ncaIuezJ9KW4OmuYTCK36DANu6rWNfd77yDrotFlKuoPBJH1CaafEJ0F34A74R9qG
uCLDjhNQ1jJhlJanRxPJYG66zS4WP87vECJAl/DliVpkx4UBURXlieXV3OBX+W0Ciu044gq3Nawg
RhW83emduKlgDjFczODayE6W6aUwBXd3TWDJsLZeYKQxEdvGROD/CM44QCq2r7ZpMDon9ojAVzP7
w9Hv3bbpP3YmLWMaJFZg2ShDJiH1PI9NHEqNGCCuT5WFwVcBDf1eJzmtnvQRcbul1L1DZSHrxC8Z
ryhJvY5TKzDkHMAU9qqrtDS/wiz1XfeKpG36h0mbi3ERHUhLqw50TLotRRQVPX5HeD3FDdsx6aNo
whylPrkp3+U2VGnpXgW2af8F5gpjyeYN/DLHKJXfzUCAGlTzq/ncWVQ+wBZtoPbceFtRY9M/WobG
cUNMvKoOYor0t7rLdMzDpF/KqPMkwgHWRmmfILt0LtFbYjkTRjTU5FgPyztqNMQNfpwmiG1GixIR
rBMOBnPv2ptJcxdvL9T3oD3n45Mm341HpaFeAcisN6iMmzs9iDy6vrrLAFQc+fSvbFKf+1XDGIS6
7dkU3rNEXdmuUcYkaF9ygI9WSdqtj01/+FtodjDr6OOP04PaejURzABmIc92gCr1GOgwZlA4J8wh
bCo65tPX4qkTdvfIQ+nGz5cg1YoJVESxbfyIBqhKlp+J7l9Vul8C2aHXMtT54igx/lmutOOc/zbg
r0E/ImmztHnAotNv6KYQUl3KVJClvTjqBvK4pAyEGMAkgdM+o7w7wcvy5uyBvc6lJqSjQ06+hqGD
YK6oNr+AnPUWGC4qkBin14WpwhAZU6GsF3OKGFzpNkQVlYlh7kvBWAtHzlwlnjXL/aN+XPl2XZye
/4T19ZuFeoDznrbtdUIybwxao8fZONxurw1XD9t4I3LBUNwW17cuJWIBrVMnjBMmk/HSxxu44dQN
IKg2NmT25zObFT8iryxV1cr11u/LfgqwjryWCsU3K2jhp/zdQ4k/0SoEkF3k9i/ANBSKsw04GF0Z
zXpThlXYKP5eOAtaFyGCLMBIEFPkZinGrmDFadY6pAGHHJzI/JNg1botZOYflIGst8ziCMbxhXqG
YUQ/b8SedxRXED+G76jnaOL9SoL3NJc0I92KB8JZ3VuGUGG7Nd1sO4Uty7cYxxsmbI0rtDb50EBO
vGCj5ZWFbeBOHm7WUMjgqPqN7OibJlHqQuv8Ta5Q0mI7Qji9lfuTcfjm2ik3eE3p3SixrvbNhDon
9xEOMlsHVpSvkJeCemjMEsYMsuBBZAk/GU7myLyWKN9T8rAxiE7RJCyHOVPZ43iDStadsciwc57X
LDbc4wZqRgdnaCC1zf1W5w9n7pFaRUMKyOw5sLOddrnRUr/B+163poYLzVGshE1XbVwf1R+d1U4B
k+tP1LGWFdPVEWUEI+J7I/rjbZTZDavUOBtr029zgJ7xeQqVRSGJlCPNz5x7djytQFeK59tt5RZy
mqTkHnds/f8MSoEAWM7KYpqzaG43eLz8u8MRQXMhIgRZEMmUBbI0u0Q3GLnQh2ZO7u6Q3pqryufF
DQCRSgD9YP759+v7gK6zgdl+BgCrjUTvYWwacB+ayULrZ04LbBOCxOz1HcPcJhO/DdoAj93DgLAP
h8YMRJrFIeIp1qxnXcFswzzAqKp0YOGK9/oRhN4+TeyEjcqRG3ZZyzQVUWqSz1LLPMsaqv9dI+Z3
3FFzINAWehLQyLgcRmtVntTrPip9qQZpiFRBxr+rP8c69wzWMVvDFkadWQ/PvdblqFjL/JN9wTy1
+54VUERYhKcYImJkBBXCaxTwj/SE95ZDrEdgb5A1VynU2rEvVK5OG475ragsqKRN4g5ead4tUDy2
W9/Zsd/jQYPRQ323uGa9rXIokfGB3MbgM3NQHPPJ8cit4hgG6wxzMmNj0fRal25U+Y8RXZ+zzMK8
LHsZ0gHhFX457EbEsA1xzQVDZUUCz5X+U7YbVsXqqDYpRX5Hy0jWoScjiKhL8VKMeWV9vbIrw0ZE
8z38diqWGv/aHsfCA7L4k4+ClMuJ42s0LB6WR89hI6jsw13l3fyru7/r+uPucq2oTC229q0B6HB2
1qQkIDYp+Nz0VHxmZScbMtWQlC5tGNrfCuLj246JtJq63hJeAw2ysONYXQhjaD/Uj0991UVPXYnM
EplLlxCOBEqOZy9NoLj/mQSBTLUr/CdZ+p+vKhYj6TkOWdADx+UEsm0kqXYzN5j4j0Ez4JA1Ueyk
h/qu3Tdm1SkJoJLynz1pdtYQuU3KGGGg5TCb7910hy3KvxILrynRdQUcck6otZGCTgwUr/n2HHWY
NlACEoFgNIplbJ5w9xHzGvmEpGCPX05p3v8kBFgFqYyoQ0BTSeIkU1aZj15hAamMVQZSOZFe+ba7
Srd1mlS+IHrbJhWXORiEvmMAXt8hjUrgXi4V2S3EMPut5dne6yQwMZwAq4vQFZz/TSS9CRootWiL
SpkirARcBNBbKYB64hdfwYHCrDoLbcJMxEIKUAS+AS3hTcHWhdh/2ATnT5onKsyZVqq8IEs409Qe
77zXNNECBm6SvzhzMMr4UzPpkB/q9XMBJhrA7BiUFxCASiIz1+/a7ykSdz2LxZ0nMLiVlH6fDWJE
5HvWdLZR6tjvPoC4FIOQ7xwu09Pzo0i4vvYp49k768/YtvI1VPZVtgb7Rdpzcc+FZsr0LE59JNZd
tTuk2GCZ8EWEE8Dm15TXlqYeMrFp0uj1djZ+2jdOkt3ABYDvzMYYdc/LHI+E6DHe6n4fvAfi+Gcv
Ousg2JDcc24EYdU/qjrRQOFZNHpT3RPa6UVXz6P6KY75wyGo0KwB6QWTeZ8GPC51V0wNik6C70ut
Ki06yMR47Sm/rnPRQ7wv47jOHjeTP82luDPrYR4JcdUgLVx2dZjuctmR3uRjGXow5zA9E4LEw9nE
WHPZIzJeAP4XnjO0SZ5vgs9u0B2Ws0fwQ6GBw/yqjIDFST6Npj/eazAYvyfjTzQf9Zej8oeuPaOa
O4gxdTDxiGaqxfvRriHW88qsaEeEe1qtzElJ1aQEbQH+L/bJxecl1kQc60eRbmoP88rKCaJb5TZr
1cFa2weCyL1UupoCvXQ6BWfYVonQYmqjVOjIpE125iw67iMuGWNA/E+ZAeMyu7OaqGfnAxQOq0ZM
TOzs9+CBDey2vA54MRG4AHih2oDYhp7KD3mSFRCSstgooeO2bjxrnD9IhgLBji1xY1Af5PE/dV0a
FXnfNLms2lIHEfTATKdt+VeOJjWZsV5wss2YTMJOtYRPPjOx6v4hysjAW5gu5VeLKX8X5FSciyjr
JmrDpdYnGGQwGPyhU91DBblTldiZ8AeWBLPXZT693gLyvvB4q2u6QB1YNffJGxDdsaCGLGIv4ZUA
4N+bvKl6xtfA5H8IPoOhKs9x7DVuqznZpUsb6+rC0uFf+lf4KL1zDkUNR6eHKdaI5KdMW/hU4MxG
G/BqwlP783rK/VII7vdCiVj3ni/U2T/Aa4f5D6zx7g2zcOqlKRb3so69IXG3HZWQ/Zr4SlD64O3c
E/VbiKr2Eo3hkeAouIAG6dGOm8LJRCwkn21N/tP58XIvQKsa6+f7yCLRKX+UK1zTBe/GEiJFL/e5
aw7mKd0bo4A4a9eJq6xHjGS4whNRBpu/ZzuDRcSo+bmglFe2xYCcL5iwD1u1Bcll9yaWlkJWGjs+
yuj4v2lDTDWhQLMWMAperjDFGvUyQOcuQ2HXZ4QRoIoyXrNN2pwZAvyAh/UHPCEXy35Oojk65gVC
wd6Tay/kb1Uu6bOKhlTJxKngVaLHm84xcXuY6iWFbIbA9H67CcKaqZRxKuG33LOl9Gh6sLQNYn8/
I1AGNTJgcXN1xNiXI0A74mfbZfQ9V2TBYwTrh+lgyOT1r91xKtykmLgiaI4qHve4Ui9ozjGyZWkW
QPZuJGS0nA+bSwEAI2KMZb6IDDOSc0CHlZ65p19hzWa6hcSgbFqcBVD2Rq26pfQtBaSo0tId983Y
iXCrfA+FgS7BOCO9mAA/pxsbAAPHjWjwu+O42crD3rSLkC/syC4fZoEQcJFwMZY00KSle3xu/IEF
qB4Uz9DGOsaIxi4/KzQXw9hnDHjI6t3qhjs2vXTHwOphDiq4rsvVz6B+jvER7C67KcSRWQeG91MG
/haHvzFd2RSLAgh+DQKZxtsO+Tlqhyj79rg44SlErl6yq2Ijjsa6u8xsbSEmmvJsfqKafWg0DmJz
yJO9kCdZ/ryItEWpxZQUTejl7+i6pXp+qb+TOAU+0G4vaqvsTKuETEPj/UXhmZREk7+R0iP/zEiW
+ApzlHOYAXdEIFrErrGofQLJ3BZ5Tlh/Z7hS4HQGPTVFtIeBxuh4spNQj/BG+vX93W6VDg1xpzHJ
SAGkoYvYLOmx3ZhxbVyJZ5sMO2mpT4bx6LhLhIOiIddH8SQwcZOmL1O8MYaBQPd2nS7pzNYqBh1e
7JPfvFXWY25IZWVrHxiSWLr2cgDzxEcyZiIRnuqUDDyEiG+LTHmYKKqh9HiJlAOSAXTPosEMz9j7
aDxPgOXmMrArHgjB4bZPEvjd9iO71ujqTq/9uQ7kF8RCd/N4MER7WfkSOA5Q9eMJlDpUtkJ7GSeb
Pc23Wg4V4jnAPLBq3WNUvQgaW7mIyF1Af+HuYywWHMV9AvQgYPrtPLkmKTEJKvLdMuFZVvKLQekk
q+e9HGvq69KaEkCgYjGx8lRgD3oNJttDCyEpxlMhmZ1WP5DVvBIdYFcqaHGDyjVXP5IENaVYhAQZ
fFQk1fN+IZpGFi1raqdYyhLVtm7ilAMLMLof+HNJYYpz8Ay2EkZcAej5359zOqacFLXZvIzS2GOR
i29dKoW0D2I6oTJYVcjQbMDrCNH5ZPtXOMlAtyB/h+vqf8T0xN+gA1hFXifOQJ1UWhIhg04k8vD+
bSDphcpKn6zcn6SjzEVWfYroQ16hI6e64PLutZH7ptssLSEHThMglXNVNpP+rGrizov5B/jwiJLW
3Ks53BcWkYfOADVs40366D0QArOLi5+AAJXq2i7qlPybAFJnMugSeb0x7E2PJ9Hhxw74K2iDuCWW
fo4VWGx/2TucxLkDus15YKI7HpUvrnjeuoJDlynV/JlGtQxSBgSgUSWkgn1m5D5/Zixpg8TRP0Zs
Sa9AOAzqJCZFCPU7/cxQT2zq4nEEqAQK2zDN/gUFGwT1GnU39j+Ifn4lAFriMA2TYHNlvSBoefdF
usAfhEalo9GPc6FU98fyQK1ZtN9WxNgNbW5kOh4pM/rQ0kw+43lz8cWvGsyUDiEJc787I9TdbWQ2
QXEmE3bIbbp4BHXrvZI9kaAmUE4QBSxj6ZgeR6jgKxfIg0d0szdY0v8MWcdLJbBOKO531mck1ajM
t9jHE9L24X4mGOi/x5MeuV8G9+rTG3/KYjnei+T1YWig+f88iVzOsn9lVlrzkHbK6Uibmseq6h+b
wre/QCX7DYQVjXdUUFlSSmfyRIVScmhn5OvLY6LVzMRrqgzEOny/XLR51vLJfCvW1PJiP8Vex17x
vZmBHjdjON7L4OmDKAXj9GpTnfx4F0F/cjuOybzfTJqLy/0WdfFMpOiJUBq6TsVqU/EmJyphw9LJ
95vv6XtTNVMC13x8ImZMaV7rY1i/mKXMSHrI1F1MzxmBVKKQiOpA1ztJJ5lF8t6+wD1NPqbsmqbB
k9Jy2aCpk3Kqx3rOTcgYUu58Z2Lil8wghaifFtwLTEPxWrVH5rTtJQPYqikKKeAF3rzJradkecxh
VJr7e2A0OHvfCQNnanNlZYcTZOPsRGxmeHB0L59d9EY3DojNJcYAsnkMVm4UUisGR38wEdoZv4Yw
Ri/enCurotVJ71YLMFoQQ5mxfMBzjgVgi/RX/3VTEmJostWiY8+PMPtLdl3rO6BtdRi0C0b/3b+Q
y+5yqIQvpnEatSB0GP1MkVJZLNbWML1jLFePbj8Nc5ukxPqZDe8YJ3qq329ePgBQpGKmlvQWnIby
InZYJv9Uyvj8L6zbiHcmalpSeu4EIySEZY2n4BF8+dbbp4g3esm5mQJzjESBf6idtrOU5+7kgJzF
yppwuaXzuHVJnQpQR7To6pvVu9bJJixnZlVEQ8H37a/AWxtnY+mYfOe8T8mRVqiN4Z0T3enfnrtM
/yYF4zGX0446j6CGCvv/ejfdyky3Jue2cWO5IxUDoDTEP2wXV1AHhXfitBynhyCEHgQRk8XUienA
9/AniTQB+H9AI76DByN4wytDFMS3iy5BcBjjl2yVnlrWxBdmB8agBxbCDkU1Bxl27QWQ4WWCWk+6
bnAT/yut84ExULXbhn5Zg438gDsXxg3WiNKx9sDljjZOt8EGBSlBh6YuVtMWaTZnzQzYabs1Hr2b
il2YdxQj2Nzl1GRtGWPfUeThJT5vCnYuvDtq91GXRVtoh8bOLYxuFYdmkJYnLggNvw6lI5SnDcm3
Bfb60T5Y/DTEtjTFtl+2+lgAAaqENuje+QMb2Nxx0pxm8w3ojYcyCm5GwJPte9ia9RnCXtl43HvK
vO01zWZSsm9ATInkT9B2LTRk3NsYQ9invQ+9PEObVppMb6pqATYW/Dj3U0T3yg6Ry6tjkVsiYPEY
79Rse0IdR1bmDSUKhA53eXNOhjrqDEFbVZcq24t/wYvWugVli+IOaOTtwQBGWlNhr1kxlFU9Ow6i
5KXw3W9K8AbaDbz/CTh0E2it2GRz5iok9U99D5e0Dc3mLlsDtQfUwGDjjAaVA0nIJviW15HYzbGI
fDrD5dUeQJOe0V0BhLFQKt1yqjz5jsj1Tvqshmffxhvu+oyBSEnzev2o3/HW7hO5nY/QIpdBG4pt
pBktmexDYwuLtBso9Etx6oo5YPl3E8+SuXuJncyk3THn60sUe+p6dpjUhvok2ZB2eSayU5PZ9Gms
KKHOP0w7xaA2sO9B7fMieHQeeJAad/TYJG7pEOZT7J0e5tAdjkkJtXWffFTnZaAFPLDVGFVnAezC
XMXCWi3FWUOMmfk3ehTxZZf9XNd9qoCZd/4Qld7U7uhKM110f2JC3qT85dzOUBaD4JJvi3iSC4Bz
kVWULeHLJ3iJRmsL3wzneH6kGF0Y5hmlxnJ/aObl6GNyyuBiya4aKOMfp92iwqu3LwjiAm1ghZie
x7jwFjyqC6u+VSJYCf2r5w16EUgfLGrV5B5LrQ8TfgfjKb1yH2sdcW88vdhvUWIA/Str4RLN6Rof
KIZlCLSGhYX9ZTO1r9uh+qwQM+3uxwzCEyhUDld7WlPPyUWj+mWNAFX1au03+f07tJ5IJHfpblDY
x9dO6SIQl8v+tebZctjivjDcdg8Ip5DBU/JxiUgZKnguuu00faK5XVDBx5nbhUKAnHlYMHx3euJR
P1ajJ71vqTCTWgVJ6D+dMN7BcscjfUI5gQX9kmQ6PkZ9fZoUpM7uGxLsN29WwjinhpyWQyBaIAOE
jZJNL0WZHhEkQuGA/8lO+6R+zm9Y65z52L5P12/yYobl3RjN5UoSRSM9VYhLWSFaBtsFWXutSqOW
Dd49DiNT3jrUnnusJa4E5rxFUgZrjnZAZrW8NgQUNEnRIYP3VjybpfmkR1DOxEz4IzGE4Pjtp7wo
mJhwVLnM3dzisFLRIpqg+WRlAb5joRLhjmjglKDOT79K3uh1VI1Ybz30HqCkVGfGLvvBrP5SgFBK
h5aANILbp7XgHSwz1xCL5+NsgbqAQUCViQ1ujW2FSLg8JGf2RypBIH3vPjdL7UGWbykpZBgeAWY0
6BetfAGfCvHRFQOpcI5RZjORK2lEVZV6cqDnJea2vuOL1igP73FSoIy6hU45DsbQQqKEphwENNT7
RouyXtKHXb3CZm7PK/F3oJrlpiypR9YgbYQFu2tKw+a4IKYRg+QbOVMHeqR86aRQIGTRfxAHyiO/
LTW4UtVNF46kI6KsS8zqWqUIgXczQyXCtx6ihnqmiEnrRRWhRiKWU8K4+fPMoatXcARAXno5eKuZ
XS6Lb1YW5jl8SCJ2o17/dpFDoDYRwARtf7PbDocG28zw0JCoXC7W1sGh5VUAahycL8qy8veDalWq
Z9PAsyJCI2lNo4qAiP/o8g9SX/DlqRe6XYvBYJG8M1QSIW/Pd7F7+GxFzjND/+92+ZE2Nd2xNRfB
TZ2BAHkXkchI7em2V18dS3TL0STtXwSHVsAU6SdojktL0MvwgvfeJVytzk0AZSkaY1gbA/5KyVzx
S8f5M6WFE0DmE1OG8p+1HM/4sKWSzweLEzYuCX4FP6Kioi685ZCQT36GkfH+6RqV0A1jhqZZPHth
FQAmP588u9cNwfPaZyreWoSvcPL38jwrbCKgICLeALAHrR2oFECz6FVWFh5pi6r5GwettspJtad/
ZZNEQ5vhlGzhxz9B4MX0bP7I4SDUmQNoHbV9GEjEMgeausSGJ1tjzOHlVbi1JY2PjbZ7cgk5D9F3
utM54z92NrpCHaiSYcXo1w+3MPEHldMgMp28IBGMpnayed7pIwQ01oPEAz5T9AqxN9/QaM1PbScb
xMy1V0THsNfok/J2pUI0cWL5e40CxF8eTUGwODBJROecGpCxb3Lz5RiDmaIyO4FQ/6mfUFK3ndgH
nUzrrY3VWGpNrBpZy8KQNLI9S5LrK91aCAvRKOybvhKqEocPUKIUhM65GPNQjk5yixJa2r2lyLL2
bUyhRWfuuqU3XxP+nR5nGLE/8OYFGVysZ0wCdbnVmqXBedHn1TungGRbkZq5VMw9vyksk3tcC+N0
n91dZP00ej3f/fo4Q2HJYSQIRk9aLGcZ7w3dLlzZ4EdI7MHlRk/8Tjcgh/lncAD7tfb+xU4z1uSm
kWT+XO/rNx02lrMAjM52JLlc597LpbUO5Ig0VHyCkjTFv1/xuwchM9dXGrm/BkV2WHOKlaKDPnji
EXtfECquz1wd7f7GkfRlVvBsBU2v+83bf7ggMahhXCBNoDHUt4zJIDuoPcBEKNGqqbeEP/tYeGQh
Nt4MiRKwcXLix05CyTr8QamMuCSUPwZgxovUlY4gPEVv/ZVP7y7WhG0U6rNsIeN1+zaPRsnwLYga
o2yH3ufw60aKQbSQmh8uLN180Ctf5nmiPUo9QsQYWDcAYPzd44YlKl8d5VaqfFwdOftHEKEoiQRR
6rcyU1UMlkSn58q4DCdxbsnx609N92X0RDMRP+1vEl/NtKJttmJl7peycsIvGF3eHOLt6nZjCewO
d3MyBi3vNwdnGyMVGta/vXrPvySojPFw+Jm+Be7Y8K+tmlEUu7TNh3rqskRjltEfxULIR3hE3l3k
EOLcSYYu1ot3VE6Go9OZ/Qq8ZYfikYHR7JCo3vsPBtgotXh7JbqumrQNuj8Psrnm6MwAgkRa/B9R
s7Dn9rmFSBCwRYQ0v3BTdSJoiRBPYZvj332ZM9GzvNJsFyaKAVd+0TYlzsCHMX3+nhfoX5Owygy4
oXe4kC5p3DD+OW7j4fYZ5Ei8VlYyLhxa5MYeMgV/MOyKU5tdOXlEk2Mi9aV63u79kAF4hmr+ummT
FEHhUkPBh0nKUUktRd7n2kM5PI9YmzFLV1XtTgVGOLZPE3xPPBNL4cJ0jexxMA78a52qKeGVSJou
zIxzYpzRFER7L7G38cu9tLXh3agDdM2wp3lfBCs+V8eLGICoEcd1dMH/5uNA54xe3m533FIu/ob3
ptVbkzC9T1jQt3V5Z8Dm1SEUU++QnwFlJyU57gNWIkFCZdgMbQ3ZlFL2ZdigMbYwRbii6AEl3E55
sDQjR3KdPCa/unViJ9eXg4wazmTaq2EcObg4gzi2JFb+YH6z8f3rYPnt9Fs4QXDfR2M15nsM8Au/
9W3QteeRcYEdwbOdAOHqj3NVdinCtpQ756UyuPnvDJKM16KQ75nI/fXhMYJm93bX6RafwxpIvRpf
WacR6yWa7YyEWDxyecFN3sYh8oXbh2ZV0/DQPOovw2ONrxvhw/QGoKagejgXk6oKQbL+ODXm9zuR
3+fhG3tu7T3fgV7UefA587binCfGOCKjcxPZnCMMSpv3hP4KEmDd2tmWt9af2w9GKLldUyalYvb0
YrIKKkV9LJBkiFlaScfcIUhwINM66WCLei7UvrbLWq5ljeNnRYPDfC2J3vSikmgBEf1qx6fBCGbh
V5wcVghdgwPuvYkSmohASUO+06ICo9u69gmVNs8xl1K0X1k+l8/8cb6xMgS3iIxzrCK+Fufg3yz3
SzBq9tEGvuvmBLTIFO8QoqYmJQFxjbdvStjKfUhA04mDeCQT80ecOPTe7AGCYvIkY7G67uDGAHY7
HSKh6LFy1sygwV0bjbsIO5tDghVnHg1QGhbeTQbnw0Mrvl2brwlRNARKQ2b0ZSk+D51WlBlza4F0
rgv+GI9e9ZfmlvtCbnlvpfTzeFLmolApQocwFpuOcnCTogKJdKarfnXyXOv+6KIBqS4NkJ8E4bv3
lfNKqz2Yya3E57hM6E8L9hVIolavXkKbNc7RhERZWgsa1YHKfH/GNKLe9Bs9t6EFdHcda0Hh9z9P
wzMyQpP10r44CEixKVKqWvpjMuiVe6c2lOD3+7JMmDmCL0dx7hgeit+CSnCvl6w+8J86Xqwz4kb+
KHd/uwZRbUrQolieI15FgWW1n5ZcXiNj1Vk0TjMW2aHB9/ky/1mLoG3YOUcxCZMjJY0n4fiMAJrl
SXzTh53f6Wfl8KQ8lppO4l2nHKLy1jR1gv+RZoFTdkFtHhBrwyPG2Q1MVpcuHkQo3Z7/z1UTfQtf
MgLLxsW97Wcqrez7BprplPrcNi327R5chKD0JSo/JxRjPzhwmNoBoVChrvy0G67A+r0JhkukNcEa
gslTXWwp228xGL9s4QxgnxBXSHrBybRnWrl1tDoCFtxKND5L4hKTQ5K43TesQkHrqyPFvAvEoB69
rOFqUi0kawQijiq5gV15mODzGrej3WRayiiOcGGXpNrS4vaWEss3QpnMpzwjMOCFVvMvGJnrKFBM
mVHbJkmBKSKqyPSs+3L9kAZo4u0h9hfAg30cFF3vNwo8boebB9KsSne3loVqrAKw/EcrC88IwQJp
0uvEPkUNnjFjqizl24KKoN6ggfY6pIp0ZrRTQW5/HNE+wZtWJcQ+2aOq7/8GZV4WKgNrqJ/J2kkM
ft2hsKsHlzyhnX7WluDuFSvn3ACR013l12+5yn3OsatH1WN/dcO3c7kMKTLJCXgRk3cfQExY6FDg
9SbEXKmjDE7Hk8YLb02ss3HJhk+UiP8ic21YRYus60MnBJEKIKn8iX+qlINjr4doGxICEDRBhHcQ
iiemsg0qV5YfnQmsTbQ+b8DH2Bw+JT6QsvcEr/tQosHo2MEpm7dmu99MBbu+NuBRL+Uqb6SLou/S
/fJ9a5o40XxXdPcaHs3OC1CdfghzuxQLyb6oYgIOMs81/Aho+vYHTrKa6rpJmjbLggFMp8FE425A
TCyS4Jh2N9YMpIOH/Kw4WcED9HG5ZHKqV+AQJd+33Nw45lGEqNYQoYlInoyFFJLSVSqD2Uc+GTl+
99ODov2TSTnA43WMOm9hiRq6W/8rgzV+J2w10HbQjgGw156QnPE4H27fXR9GaMi4xORgJMMAEidb
JYOU+r64K+8kJO4zx0jqory+YvRgAGjnbaGVbS0MhX6inxFJwUt6/h6yPF3ZjMgJbdsDS2oDGTfL
2uBYyaJe1nGFj+B7nYCIVQehDGzZGrIR7WCcypyypdPOEfGAEKeMgu7NnogOu5MScS+ELFGTwlVX
IbgeUlC9hwqu95AxifGTJbK1whFyVYNmZc0yarHl/+d5HQKFL5RmhyVOhiSZaBkZFKcWsDuJ5IbB
gnuIMzwMD51+JadUPTQDUVwX4kMMMio47vTfxEWaLpAM8KJNOVRNT8mNVeJ55wVo3JatD/ngYwhN
lEJTaB42mDU01OXB1VvkBcp4LNtNFN1CiL0RXnT9K10YRLPo9x35K3EDFXxSvYkvE6/es1Uo3AXp
Q8dy00o2RcAVuyPpvdHPEun1N6Kut108Gsn1Z6EeW/AuZAYT4AOnVgMaL8J/sZEDPcQWJO8EcMwf
W80/FySMH7jr7ZWiE5STQVmWQ/FrBPE3e1ju7Dps1MfYDT+zXgVNWSyaO1UEsW7rwXby8Sj/sPNN
40vont/f0y6kCpH9Cei/8r+LeKbPT3BKBb/JXjiZtNZtQ54nOpt6lhsj7bhtoqip0xEg/Pu/MKNi
Ns2N2aZvN8/BjeiM6aFpJPrb8ofEDWT2sPeDdO5v8/ExqgHVPvqiBQqThOW+Or7RkVLZOSJDq3oB
YfbbR7AouJUAuQGXOfaMcuDbADs7LunXnkbW8/Sa8t+e8RgGFbQp3/s2bqeUg6bwYnzuxQDa0iCH
rj1KzDfm5WXczpqZWui7GnPTvSwZ8R8Q8QbGxB8xm8tSQuD73WWF+NuhDGWWFbgAGd2iBHZDKcq7
6LPnlhORg0X7JAJWWbbWlF2Jv0oqXZBh+8aL/0ptNEyhzZdRkZP1cKCcxOEtTovgpkMCyG4Qo/58
y456E3edBT4854sVwuOGMa5q4IcptMGkEVe70Qj0HfxvROaNedlYcZRmAPPwNf1+a0tWgJnkKnE8
RS8EckdWnuz26RMsr1eaTopjrMPRohOfxHrT3Xwe1TLrSDNTEMXhpzz9U2s9owfFH8+iv6Ncc/ZD
itcaL6Msl5tGhr/djfvw5ZNwoRxj2bbzSIRHNA606An5TIZ6lJfX33cKPFEJV2LwyhA7/3iHusTY
ACmDbzWqbZi0s0Hf+9iYfDx7ErvU5XhZjaiFE8m8EVGMPGu+kbtOy8jE4qDCab2TsdepjceqfMOK
pTzfOLKHStZifdUrcGryybAXNeDPPIfiR/tKc13bBMX2b73lbuQBQL4tRnqRt8CMm9iVGloSeOpz
c+0dRO73pDJMGw5uvzCGHPAAT+Q2zO3EtAqwt7gwJNz/Jtl2WbUe5mEKmrcNgM0NwURUZBE0BO8W
x14jG4i7FwcXxVR4vqgg42pxze+HIiOTAE/nxx5+HBsk5DesK1EcAQTbWLwkayPn4igU13jFHBzx
aQE6D/1m3MmueK0BSALGUTzyMBfjrw6VxwU0q2bWEQRm14yLoYZerecyx1LfszoCzutgHhgX81MO
mOGL7yT7prkVHspms4peGLg5jBA+uL17FVkqVdlgF78Phj8LaUiAcLLoznY0b/yg7eoBkfCMi1h8
Bwtu2XoaS7OrG4KwIqbc957Yg1gkY6tn9X1RTQnj0G+jqOWIkHrS8ugZY9qKir9/d2MxXdnS4+yX
JmiTSP3ScNKhMnCQNT5PfzdFYtx28HeOnmAqJmrWcCVZ29u6V2LK0qryYoMgOR8T9KhOFYgkPLFk
XQQlBysrT54KUIsbHwTm+B/ZPr4/LQPHGi5BFSZXAhFJoLl0XyIRAhv/G81SBejIvcE/90leuUnB
tA7FZBdPB3ZYtentcsDq8RKmeoUcoBDkYXuO1ScbNLztef5Ren16kbcJ460Y4qodWFk3ZmXK6Mcl
7iBG8zLsTnefgp9/ykJt2RjAbgXyMwqcbwK7DvJUeI1l+84VbYZKrvMvGfJgshSHT6OMoH/QwBFT
txf7OKdd/78G9bWJn2MswszGDtyq0CBEjuTnLgryejs9bCFR8V4EScdVW4TcqLeVla8vAMaOdW6J
q2eBJBXvCeyRUbvfLkOh5jallyNHOjmKi+1SyiUg61hSkr1IA+CPL5wfePVcZbaZFGJ85VdDlZ4D
VncavHjDGIqTvoWle51c2cPfz8zrIn7WssMUIL/EAqsUOzJ9qtAvu0dgFKj9yJsYDVDCL1FJ0K+j
sENnZgrvv8Hmiw4UHDdWwd0XNn1WLI2+cLuzVhgEKIe7uzV2Hyme2ztIxb0+mG6+xv1Yz9SVj/pO
wLwPWPfcMwxjbyJXywokdCkEdsGMNtn+soC6EEGqUKa+idH8aksETUKYOSlr7+1itC5QYOQhskK7
DoaUbjAZ/IC1ZwlOYE15Vh3uJXfCwuF3cg1Sb5Wczv3Irm4UpXW0dYJtRR0DBFnju8UhFKFKvVSd
l5clYHTJdus/kzQAvNJiltXqh2jCrsqLUmBSeeAJPErzIouSweRxjcpD1NzPygL6oLYzFjdHcTQj
e/Cz3Fw1VDgkPRaOTBlVXk62dwBC27VlNPUbeO6KFRRh4ULFWpcHNwUDOaoVtcbz5Zb49iqLOtEx
2HkWn8Q3Xrc6h37rD03icV2HfAK5F1pfRgcbtnxBQrJOmutP1TQgaHjigllpR8/mu3P6FvTiSad2
Wu0aAL3SnkFuC/9Yj/vGdFSLwYd7yCDVDfJJUsFKSedBypfFdpfAaOiyaYn+zlT5lD8NOmkUdF+h
g80eOcRytsWdzFLC0xmsWx3WwpoNVIgAwCthFZTktRggnlTy1qT1zYfaw7OeLqLHwfYWnxUNw2p/
tiGA1+PHcH8vmTMlrr/R4HWuqCaHFi35gmJi2tt+GbFtytgQNsM/WWQCcCMaSBggNtFlCSmX9JzR
X3HoZPX92om04cGelTtSCL7GAa3QF2UfUbgHaHfyALQnwPrbz/OBiqe3ItddD9ihHIjDpl5dGJI8
imj2IC/HXW4NwZXTZWfmkIJkP5J4YXm4F8NeSVS6lh0lTb4TMSz1ApYxVudF3ZSgqmOAQgpoIDCp
FfXBIcxLXM9Ec8XSk9ykanwxJH9D7d/jLErP5FsdL4/32Bo72gDwu7tYnvSOLY81COPzUZE6WBcD
XyvTEFC1fMvGkxZN4HlJvKssz+MZ1WjVxuMpGMxqMZucu6d8IDWj94v5o6GFRyOAahyddZUmQuYH
o5M3Y56TvEyEYE7fNrWj2FFYaEukaq9JLJAmfDQ20mk8bkpvv4Nnr6hqnXqqshPq2SMIAo/Tu4Be
ruauJktKOuLLagS6Gxno/7O8qLA5Tp4KweWYDKFJe20rnzPuZO0cT7PdPBHt2oW5H41w3idd53wz
ozVXfEAMUjfcpMif3zscaPudrhkw3Zm8z4plf1L+Da8qKjROhcLoJXuZ7U7CBWP/XzIrbBe3zMiJ
1w+eDqIx/hVWwsHeNIEdazSCHrgBjK0rHImkvJeSIdrP+RfNCSU86ceD7YvSvofguc0HUHC4Zisa
ygXNJimufh3H4MopIwec16ddDB5Jn+QryQr7t3OXvsWXGROkSQnavf9PUfAkRC66wS8KNWjQ01dz
e1aQNeCHUJ6wJ7tCnk8B7walcVq/xXgM7Uazbrd6ZUmPBO+NfUKdxUE6mlMiEb3OEFm4hzOjVCeG
sce7OB+9oEchcCnZc/AInApDJ0zbt6nMUUa1TpAbsAFdkUydBkJI4vG/c2m/x6BHxeTPhgeS00Hb
fAZ0WKJmlznkmVKT9BN/DCLky6TkgqK6407Ixdc36jwCX4JiBf0BCyZjP5jxTAFlb2o9gEOSrc8B
R3iPkwWyfR6Cre1qVcEDSaMgLc4P8m6Ptty/lY5jpo54mBN6V73WZ5ymSJvqD/xd0+IC+6CskIQR
z7UKrfdJdFd7VAKd+D7AP7Z5v3l2qYbeX8qTVQXxJdd76QOXHaBJTbbhrWJ/5s5a5kRBIdJuR8an
DbzR1xgTXwHJDez4sr7RRZWcz1Xvrhl8zgNxAfFSxfQLjOiGdlmyCXlfg5f9tsyzAXCv2gAq7oe4
Kq/S606wmaW4l1RTbU1da2n03ijxkHqYUn4UWdNFru7SloaCW+bHua6CBT7azTphs6rMdSjC/5Ux
O/9u0tck9DL2csH1YMEkbQzqJUUGaHnvAecfNkVzxn+jmaMtZ0fF/eIJR3h2xcdDX6gb6T1veK42
qOggH3dfxr6l7CUwKLO8eYXGCLJkTJpQrzAt6AGas68sDahOn/vR9kPgnXuaKxFJrzGyOMc54nF5
xwrjzioJiqzMredndbwnCxABpswE97RydRgU4ubSzukbuy3224UhabrtL64yYoIvyRD25Zx+v2A2
sFnpi+XW7nwM5YhMdexDNHB9EBfjjdo2fv4jK5STlc/d7c5IsX/fem1OOAaE3hPHOnVG33MHAzRO
+nIwDg2VKGCfrUpNRPRS7wGxhseqL2JtKbvHuuVfXi+p2hL144Aq/BqK95MSvi9Lnu4UPt9Q4LKT
5MqKzKO2FYIWkAJfRtkqidzoQXdQp75j6FCZunnT/4D11S584cL0bUvEt/aY9cdpiN4wC8hdVM/p
jTAHqn7o1XAk9Ssfz/ub6ggOshyTeeciwc4kaE3BHy353vNPSpK3nWEUvMAv6pcUhfmzSOVryaUv
q9p13X4ugnUxVDgRDKb8w1LIdxGpWyTXVpxUKrozRXmr80W3H/Gk0Wj6OU1y2CFNFACavP6QwqTl
UaAqkpnPCjx6ik24v6ZXdhRUUUUDGmNu6emwrR7gjdFY+mnoHEEE8m1pTyZzSHtz3dt1ugN53laF
94PHylgFWPlNw8lsOKSS9kdzEd1Vkz5f5nl+JUb1bINA0veGdx8F1lhZaTBLU+T9Ppb3Me6gFJiu
uYPy6aP1iCkhC1hK/NribJXsIbVVpT9PX1ezb3affZ4D7iXU6XNhueRr/jS0QWGWSUfquN9+eSvX
XK+hftS85oRPhtEWRlADQxY3z0HNG5ccObM9+K0oOW6YParYl24rXko98n2oMlhNNVFmNwaPubKZ
ZenQthyBJysB6L1+pIrW68wzWCwLXtPhzWQgHQkF8N3imVVG6jqrGEMx+sgaxemCw/7H8hUcUCFC
w5X86nvVR1kznZBa3+b2GjCvy7FbJA5MiqgQlzb+kacLnbKuWiQ173YZCCJrSpT8+Bwwk3r93JKF
DJpEVsd8AXeTtc7sMevWHIbaa2MBaAHFH3kY/nmPC4MhSaNr9CYVOi1DiFt/ZI0B3RmE0FZ5hRHE
bINZMkK3UFvs2qLnaA8wIplnijmz++L5kIkHBmQ19MGGzU4GkAAUM5AmDYiJmJpJelHEoTG3j1/M
BP9b2v4xmPeEbCgPUxSJoQursMjoW7fjV8oq3kr3iCGokUojgX0B8mnuHvUZ5FmKX0r2a5K1giKP
IHyvAulsL/6UK5XKzV3QI/TljHovOOoSM/cr+CWkmcqFC/FBF9xyh9vlXBH81+3gzT+4zjQf5hUi
yaBhBK/fCqOX/PTx985lGeiqklz/XmuRn++b1vMor6n0DFs49dO2/UXol8Qf2kfExx1s61+2wfud
HFeyucakU3r6hSjWS4V6mkN6jANywdubcTAbuAFIB31VdNFRaOQVEyDoOOKIAeRdhAHEPG3aSM1r
0Zg0VVMMDWrUU5Ol6K+D4lBf4z1/vedoddvyut9+UxJthEhAkhTCMiI/++v60PsHENtj/rSNzaDu
mw0ZftnCFGlENJnrC2QOv07cXLCHvi5mmEBqe1dnfschnZGcQ5o5LYxDWJvsHRIrPe4HdFTZ52H8
QNAofo833eRB072oiNZszsci6grCTi1tmaAB1297Y9XlkmQW7xyIAeNf9ALoiugRoWqBOcXA0sG8
bOM8FreCpIm/CxtovTLius33zuowc7NIj6XY62XdZE6R+cCUYMjGbbqumNnNUoL5IYyutCWMIqj3
Rx/eir2p41mOsQmhvy46hpsB7Enw4yCAA5XtBuV/0r0EJQjw84s+7Et87KcFP7Ad07O/kMG3M7VE
SKCgmHCwozkY1OebPUaWylPwww/ykcRTBS8pAigwP9LV0OAh8CVlOkMUl5TkoScdFONBfwYqtFcF
x2rJlQ+7kVqfgo8hHNymc6Ikoj0XO5EfECI6PyrQPdvC7VBZ5ii98gARG2jdihNjK8/H8Lqq1D70
WxgkPlz+z3CFAUSLHsL3bi/KRHOenwVTVJd+9bliGYbjFuMiYZmPvsrl7zbHQis+UVrcqd7qClr6
G7EkSaLkhlQ34OgiC9WovhtCmpm0JhMvuC5geSWKMTly+6rNr/Bo5eQ/BT84dmpjD5Ieutsd7JPv
rXRGgW7kIhTcCniO5Wsej3gyVygEvroWT2wJuEXjykFxrZCD8yTvzZMXl9f+Ch3tWT58hPQ2G8zn
HwmG6TFr0yWkS48anF6t/kr7RcOXHXlJpAwEro4rod8OGIJJ+b48hydlpOdPK/rVu4T/u+aopOhJ
h4mrnW/nPQnxorVeNSNi5cjyjt7CYQ2XpYL/2lHYBV9mvX/qPErO1c0H5kkvwA4IImCsM2IASgHh
2XWKYLf7casYt0sd6tUELGSQ9K5AzjLtJwCTKcAmZkIAXSzF7UeZPyh9t1nTil2wA0GyCSR+LYjl
5AZG8t1UIfT2m66hkQJlqy03e88Ocus7+Tj6yU3MCU/a00QVW6rOE48S2zc3apkARlimigcK/rGi
Gi8Hc8anzUOQRr9EPEZLALOi6n6JrMlPFn97YIN3e7VvyzzqON920HDJteeopqRwgQITSzzanrjQ
R6Mq98/4xzxxzy+SPABXxL0REBS/IRamPdoR8T4sIPsZL5xcKHIY5GtdOzo0hKb7FmuMN2a9nGwq
9MVQtfcx2CflY4BpX5tQ0Dk6LzV7vB1CFzGoTbRbXXzhXsf1qpztskfIZv8HS8OgqUrH84Sh+PDu
uDkdNc5h1TCBBDkumF/ebRJtR5tY/JUNAuFVC/MIdIPn8tpXiGVH+0f/p1i92/Om7snwWiIGQvxa
5Cv1aFaQukSGuAc18NBRUhGYeTZOSt6mblB2f3ZdXtxzSARirpx/ViDi9Rbb62ZCblXvIODvVwv6
O4JZwYhX8uiVD6vRNpdiIcBgN7lyBUaLwLVrENvNZy1aRMQsythe8q98J6Ht+SlOrhRN8r8/kKvL
Z9dH4tV4oV8VbQ0/6LoZWxUUv+6qDbLHsimxT9mOoWPmeFxGTnvfLpNq0E+cbYEUwWgCV5krlbV7
+8EIPDsNfIurVYWi3FB4fmuBOVVhAFtLIOXaV+sqKJo98QA8crnAkRaByV/kMnYrz4CKfCMqMNtO
MLX21qgSGGFfRdiZ2CuU90EnwcUom1vLxcQtax45foD08DGXFlo2/NE1mttfq8IrXpldY72jNHb5
ZfrukovC5grEpp03Qu31WlxhuZV8tUc0pGINZ9GyKLSSwA8Sdb32ghsDS2UjDrx1ABMlOhXFyAxX
etbpvqr87IatViZYIbmEYH4iG9RNJOUMqUCzrsOyRrcKpC3p4UEEX1H43ddiIh7sSGEYkWi68RHb
Ra7UrOQPSgTagFxD0q4wHogilDpG0S/MHsLgUPfMc8Mb5jsdIfdWuv4w7ZbOMXhjYqFBZZSvxrHz
+rNcfY20RFON9yNZACDH7aOqjPu1kRuGJWDS8verTAHjQ4K2PCCQl90mOoK1nlUcLEU7BGuzoxCe
o/wPd3+aDMx/IbDUBS9nyhRxNvHJ955LJ45D0MIS/9f0zawcEwHOWtwZuTPExgTDKhNccYj++os/
KKc8+k6mxSp0z8/mntYj+q4xjAj6MFA1Egf3cfMFRZ4MOoZjm8Kib9StlMIH7zw9/tK1ib/KoTJD
hLUp4jQR3jesDvQSAnxxnu6EI47CNMSTlqfYh3+xdiGA4TzraUCLsn4nHd1K40UNSQ26I32gNtJl
ln0cDbn1ySKOEcpR+pFKjIwQw4Z8537bT48BF8WsH+OoTWj1NXvTEsB4+PrPVcP6oaXzT2EfaVqc
RLZW25eDG7ZDnYYOYyd+SV1k8tx3Xr4IXrdTS63jAuLNKdXY73hcail7l/bI4dGlp+agVZ+njUaM
+DWuCJsH7pYu4Mnm90c2tVX2Tuhhv3RaaOw26vSFVQWTpGBR57oochknn+JX8mQj/szhyCYfpmFt
8K0vCj3DR95mAXKYV7CyEuv/4/c3jL9HxmQGVVY1ejnjjGZb2+oZnA99O1aw3KFTQat9iN95F3rW
Ksd6BqVX5u/Ecsotklplnln7rORyYHDIFjJw/2Y2zB27uFZ3KR7zFJA1dxbuyJuYl26ERRnRMZrc
bUG3ySebAfY3rg86/rNpvfRutwD107hVi1UuOIuIuIWzSUi03K5N/kQ/Ofga+pA0uiYwMVjnM9hN
h2Qqu+p1AgWorV+7WFrViY1pkTKtfaDExxFC3IDbXEvnEYcQg1nVafyuOb65nMXRd1oD8JdTvEK8
Z/g5BgIeGXeWcAKSz88iSRzGJoghwtgmwHA3uP8Pyxw0u6SacdnNm6JaaBno+EFG1lzOKTB7aqlI
MyH4hQMkWjtrFNs/DmeQQk0yIpmCRPtpt+mJ2Ay/TWbfme3q2nKpo40yetK/SaXy/XhsdN8oy6nB
iapcwuCFA5AmcsKGefyzlngRXqTQYVJHqQY6J5zEv+2i1kPAIdl8DKdoX5rEJsBLWcxaA6or3Ydv
Z49qxkZwMRPPphv01psV8QI5y0UwkuhMTP7DlEzejcNidrWNxj0+lpeKqU8Ox+nSGpY9i4gknDN7
fnrswx8uYofbOpADby5mJhlghuO2CV3NEKIW2upt4+U2v7+JOaKh+A++RhfChWh580YMZM2swPfY
ML9Z+fRqMI/YM2QWydO90tYiKJ/rEZMvf0Qzx5WO9JU7WPfg09qzDzGmFFlbJiOPukeRMJrDBgow
N6Ng+4iw0drg/8Tx174rgH3j/YLDtP4QuFUxLX0JsguE909zZGFYETp/d9tIykyw8OV+H86eLv6c
WnmjnAK9ODjhPf52hrDXWOvDpJrF7OcTq/YMQqVWAr+XF69qxvToQvsL19gSTvcSK2qiwIntvqy+
GiPk7LfnUzBZ0YXSkdJGjwfmAFZGRDZQrSBdn/2jQkvtDpnqR0iHU5mhMnLnTZe4OELt1KiYTnL+
dned9fgabSc8/gxDyWeugH5cmtPz3SKtpBoCJaGU3IgU9GMjZLsBiC0DDIRNDT7Ra7E0El7P/JgJ
cON5hSu2A2n/HR6sF6KFisILAlEPSyDZ4fV7GEvwyUpL8yIde/VLM1TJjjlxUN+ubtB3PtwZRTRb
WRA4DlulAEkbzks/fMEAGtZx+c1bEdSeaaGHBPQtO1JO8Mt38Kx3En9Zsm1HiJv44IvnK7wvDFkX
K/n8YK2JCk59qu8+9kA25z9d0EcqC5/FQsqJEGDtmEch6mfGsIQBRfl8alLyzRX3JF3aWiM1hU34
TzEcyaBC/CHTqpZxLq5G+WNH7MuyaxvW8X6XI0dsq9w41vUa98oQFHF6PTDOuFmqTGoDeZvsIXDy
LtnQkM3n4RytMze2OsqPqZLVyWjJMVs4UQX27T0iOmR9JUq7+R6Z4nyBtB73vc+uuZTF4Jx48Aq4
qlm/wGYRR9yNagzF0LKymYuEhAuqIig4bgK9C7czpahdDYL0xvJfikXnihzT8Nm3yK2tiZK0Wxw2
Y1wSvO7J6gEMTtm97fPg6NGRglFrXrZuC9ClkbkHJTi9qx9VWLUNoNfiUEEmV3XSP5SZSHWIg90N
KRGoN/EgGvRFN33oamq25+evh25Q7pW2fRSlok7OYQkxIL4AMlhMme42RJb1gf4BG2QtZUTxjrxn
px0G4V/qE2rkXJlSLkqhZ9CLnG6pkky2eGrAst7Ee9EZ4yg+WbwWUsuAKjY+QnG4slODaja+BMf9
fNimi3+cRyyx6NrUAYFjtmkYnv2WEEEcu2J5g/v3VpNe3c7GuKuJRMUE/0Gn3yTtkuIPASWZ917y
5mgLrHoLe7khhkrph6f8zo9zjSpCmPwwpwP2H4SAJXoj+ne1C6dWFFMc+Z4YYWUly2E6z1iCJXhv
srH1gGCjy6ZtqA8IyBcARFzHKtvNq95Ygze60s+pZaF/+rqiG5pWw1k7bBvLMpEJfuzCib7p20x6
/oBGzBQj7kCvWha8b+W3dWkJ9JTVzYOd+xPYN6cgPd8jIglqLZv1JizlwAkGwygPV5qbSWZUIQjR
CPFlI/YzaiiGWT1x5NJq+KJf8Dv9a4YdEA/mn5kFVNP70k2FnT5ye2aMy83KEQ5uJxDXkX3w1tsx
D70r7mXlFYfzILbO1Q+05ZK/miV6+m7qrqz/2/PS71af9XNOCzJ5yQ6ATp5brqBYhQ1kx8Du2YKU
Nyp8aoMsLlSzbgVK6jtIbAotvH4IGKI6+O1lcK256ey+ioEuwcPHVaL4JxQs9aYXOaeMckEdYaHW
hRqy/HRjmLO3zxxxGDAWbAKSh5XowALea607BGt2SrdfXbEBoisx5qxYO40F5g/GpYxL6kJpizja
reQgkjdA6DtBuX+CUlEANhrzNWu9dtds6AsB8IPYkiZHS2zY90H/r5IWS+nrP5+kmQM36MRpCW+6
a1jjPDOMBFsFjj9NVxY1UdfaW5e1JT5Oeln3w3T4JKoo5Ck+IRqE99rerviHHDHzoP1bdEWximkX
R/Px9rnoE5ESryvBfwlxAqLMuYgFW9dVmiR4sAcRhIjuJaZp0QnLLfa30vFlHg0NPedirAa5/1dK
9jt1+zMMMV6vUnBws1QJkIKmn0kushA0pCu8VS9icR9/BYc9FmN5qHQ64g3xG4VK+C+emOFxmiuf
8pin/40k7ilpWQsHSOqPWFQzK7xZA51sOljpm7AZt5yjNDk25ovdLSstI3GZ1UCI6vsZpjLIbxKH
M81DLjH3MZLP5nLm6gC8WmC8ZfxleMO8kw0RdfIpbiYgfjQNnrq8pPh7L5enjGrrk7ND5B+FzhLq
OvUWsdYc/ZUGWV0yCEjX1wscrV7cl5cE+33SPOG3FRA8sRK2oTIPt/2+pr3V7ui6QaJfVMhSzdeP
//SzPj1xbqL4P363A8LKmVtwl5iA1U4YTJUPkcfWUtH1PBYPRbe8IZyhWKdc+E4+K3zAsI2bWsLF
qN8MYVYrHT2tXnBf1ARdN1hMXVU3+gzAcAiDp8XA0H1QmP7mPHRakC1Vmss6pMpFJ2oYo5JUhkUR
iZynNj5b58fKoIEQNf+q7zf3QmPpd8xa5Xa7idGhnY9eL1nYIPDDTm8k7mzJa0Wob4CjLgxKbIRV
EQsq6b5eDxGf0xaX0al3DU7IYwSo7KUH4DbmS757GoDc046duek1OId7GZ3yHOBMhVHSDQrhrJKt
8WfXJRLML8B0Tth7tamnD1v14tTFqYbkG+W5/wYWCmAPxgpXZlt6FSyqVg5lsoibElacq8uM/CzA
e0XDMM8eovGXF/zDe6LgbAUNuBJu3MrVxJnL7HxC0iD2jdxt1RBNDWRhkYO4Q+RZ/BE7UDWrGBEg
/05ImpVrxdBFb5zA9O39G3lZRxi06BrYO2Njtgxd+uiLhIuoQ9/WArY0UCckeYqyfoq8d5dhKj5G
mJqruDgKiIuFdYOvRk0gJPfSsV972mnI9RP6blLe1ijvKHtm3ftSUwvnAz0f1i3sxAnsgq3MZh1h
uxzSpgDgFBgFmf5ixzoispbB2ZH2FQvp3YxikDoBYZGioyOJmDQGSVhoJSqcmbU31GBsfVOmH7vp
ZtcyzVejSRNr7f84+1xBwMxkypay+Bfqg9gEo/BvBhx2MK45MOn9iNHE8awok4sHvopprFhlCDfN
UHVFlWk6x6jl+zcB2gR13AjdpwP24aRI2GSl6gJl9jiimxIpzH1zOVgLrLWbe0A3T1FlE7QFSrS/
bxJcccWOZxM8y3A40mI9rP1TsbdHeONTsHe6tK3agFWZRGblxzzrG/EBlam5mPV0OHcm5Q6x1hZh
eR66RzyO28IIXGsieFTgbjHBs/N4M+8nz+FchSYTxkblqAj225A6y9y+GK4bdh2U8l9mp4TjRUMq
DBcYF0X6ytezZxBnRlCiIkBsYnvpmSlK6TzDDZSnlnHEdJxj7D+zaCozW+XYO4dgIQoDJ06KMbeB
6Xzmm9KOKD5iw7LZYhi8B8FA3BTlRmWjbYeNsuFi38OINyNUw1AameqmAtFDmqRU0ixKU90Js/IU
paeLxDI6sWZi2ji7WCFgZnFJUJLeyF5/qMmCoAKYlpbvSkSpKOtutDEtPgnVfUdyIZ0g6rmDhpad
xmZLvEkkvCZJOiGSVnUc/gUB9CsaM8YcuKf7qoigZZR6YNs+15avAq8QN0P+iwYl53fzOYxuySwx
23Rr+C9YSBMwxSsvmiAzcG3f45/L81GSo6j8FnsDR3l6d0jqJ3Bb3EFOqH9qMStmkatjskZmTcpI
APK8pWxu3GQ9kKg0anxuTVBD8HC0ZKBMeBR5r+r2u0gzuRtP4OxDv2G405Ms2uG8WncNpBYAJdfr
lDAQB6lfYwHuw/HKm9j971vHquUaj4KoyicYgDdxhd2wMwiVDWkLjmgo5WV8Rb8ozHLYLfXJPtu1
oDpGekyMoeZlDu09SX4eKx/VMVCZ78gBJ+Ji2c3qaKu97BaWdENrxwu2sOSVLa9er1+MM4zI2TdF
lCtuVCiuKkLcZ2lhMS/dSxr8AVFT/oUdek4p37idnwWX3BNJ3HSXjxvo3wlDXX6Fu77/lmsvEnzG
yafQ1kghLlipWnFbPEKVheTVYr/QMCeHn9DiHEa/41/aQ1HNbii7OPwCyAyZGo2yCHEM/3lViVsQ
NjpXoD20SnDmnDHD+0hQ5hRUwBASTN3aLOFTPTcTPDcNfoAjDquNhpRXwXCQyBxtoDoXPrQ58zBX
YG2K3RZpywPJm4Y65UayPSzNf9IOTqMDAGprmP0wVT6lvO7PreE7R768pQBOhoH5dzbjlRvZs/3J
Bn3M1CWgL43kooPg7UCHQm9asFDFsyqHeWmTxpQ7ZYz2QZFessu5+Iqqsi0ZmJG2ZBjDqbl7vULz
JwB7fkvj2z5XW7hG91wznZtMGJmjFJR2xWUZzQoa3qCUHMle5ZzySvPOu6rUAdlJr9LombUkvL7K
T/1SzhqAPffJus3tQMpJOpODv3x1mnXNnw0qz+yrNM60l0MlySKHbPknLvhzKC55E9Ck1rkilWjD
DzULgDqcoLGqDsopoY15STmTs/gbdzoxN+xpbR5+XJIaCW29kgKXXv6pNaVl+FIbO8fF2fN1xjCk
udOvPZKTaGO7MIzoIbyyXXJPOWmVzH2Cbief7sZC7YERiS87UhsvaEGkN//ZKzt3bnvXooK/h7HI
p9/Do0RRp1G2VNKP9WOwQDGpDYxDYT/XyWBD6kpUob8iCKqiKSj+ww+MiUhk3OpewCiOjq4fqyjq
5So8BhH1Hl8ZUVX7imwyVfn3pP2mg+cSZnEqTAVYanb/eQqjrWC/qG+9U+YmRfGSedBn2BO37twN
veyOhn8bWhb5HgN4j1hgllFLzrz81YsvADAqK5NQmhRbjd86dPIG4BeJBu49hoCRu12TVbrVMFvp
EhoaSJYXMNDwxjWaiRtrghRq+uhEb/8QjbkoJhAixRxOyECA0NF6gsuDMPh16CtY4xBIJnUKpLhD
ej5JxOwlL2bTjkKHKcYUQ5FTfpxblP9zrYhoBvQud/sWloBlXgyIonoxpjVemNINu7Q/ujBEiNXy
Z6yEz3gWHZAS3oH8Eo8tBcADJrHCeZfCN753z8wLaWRmoBDv1pwIdJc443ci+40+qyXw9lWgb04c
GuAx9yNg5fJ8LGPYjZmH067T5cQneApgCpqYz5911+VVI0HkLZUAAugb10ML9MPSUKtDsyIKcW+k
ZT+TRXWVcLnzhgehp2zaQGRiakFjIW8utjXYZb3idnUFI3MpUiEV7+TwXEICHzeZeHWmNj6pTxDm
8dhdf1+LmZXxKj0B9X3lc88kUSlhCWFfcOvfgFs6/OrcCOvtquyRiz71ma3kdp0gjdyKla6RmZ6O
AAH+T7db7pptU+ynhELpVXo2UBHdeOYiSnNt6S4MOMO6TKfm8ekB6lCrxi9sFmR+4k6unfJCE0k8
oh6UiquiI3drdSi3KbPx1fO/H6JRRtIsYOV9FFp7fYm5/VijBswrkadD9N/vme/VUSXqcHScoCcH
9yyDAPnxZ2G8n0XvgbnqjnQ/qUZNTa53Z/6S+qO2kbM7mD3PNec8uAP+RWnBUSkp9wV3uMkQrmMC
8RitmDLB5Oy8jqUVSbs2d8muAtNb85vTKA7pE/E8le1tId8Gzfi5M6s9DR1QP1BkAc9JEd1EKazT
efecGIXFBKUHDa81drgsAb1c+OZsnPxMK14q/3v74RIh3P3IaMq4PG99xHcwURLwEWu4Vm3//r5B
0edcsMLNL5zbzCcW7nPlbTAUwzkVpJCdPnRRxKW8ztruwnS8Gb+1R3WFowsjLbpbVeQ1cZ8uO0ft
G+NNgEqxg/LS9XK7e8pfc1ezVIS/ihRiPvvQnHmML+uY7NUljOE6P8y3ljxsXqxDauCom7nDDi8G
EVfSwL08L7RipF41+RfNgFbyZOr4T7iSbq89Cm9CGwLjytrNXAAErdnsRKVL0nrd6o9OLFKzp3ly
jM20QvuIINbO/P/+p/Nh3JPHYrk4dyi+VkX78INQsXiEiNBnvQF7i2KJHCcrSK8j89U+bIRwD14x
C7pEqZjRohTUsJyMf5H9tM+espH+OyYmCvZN01+NJ4S1KOidynjz2+QPfODXxZPthHe3cd65XCyB
bVaZyOlp3rxlalrX8p2HJjhYjEQQW51kve03X0a3oQn3ux/xjcyGOnCDo9aPhVx/vNxi71w5N62l
KM1Nv/tfvVZujkRVLAxTqSfl3XITH2PQy6l2YA8hWSNmKKtPcdy2nGE5iy/bzqKvZKHGL8Bz1SGs
zoir94gisOEWAVVgp2e9gAnBKPGOQaId6+SSNlvSWAWkvHMiZeHbq1Wt7slHyW6cUZGuogZyi3Fv
+dZ4SArg3HhPiv4ZZ68U0++gya6bThinEml8Gys2r/J9qyBbYHz7XcicOT2Ic7j2vcFcNQ2yPqL6
S2wjuryiDiDiCxQeDIEuK30wk3rJGJp6+Ig7PWO8ZTrPLkhTKHIqUKr/i7zdogW5DRjGAoy9MaDC
Q42vYLuocWbGEqQW3pwNk0mnravt1KOLSgAHXDzYoL3RR5BkoMcmJ3GzLgWdaDqxE4h8tuemrnjL
SDxecmJTFQpNZ/zX7UxHR48jN8aq/+l+5QOKNr/UgeG9bNvDsMdWyF17WddkVC8hii35xUiJ1ZW3
kUjj7zGqgAGxQMEjNy/PBhCZSIU0lI7BXfDpFKCOqsU3ZStpD2nGqOOeFJsuJT/1m/pFzJs5ljfE
T/tcdtTqVptNPqVPEA9x3/CzaFKKa33RC+QKib2uJvXfZt/gp27ESKwneWH1Q2HBGOmnYyKAyzk+
CYUMCnrW52Gu2upmg1yy0Fqkw0nZMr77fZfP06xl093WU+u8yCwjlFhXqZpUSm5v9i+QPZSrL0HK
SJIwItk852F4VUwsmjfWdA7809qsNcZJmEZn8lqoouCQlpNQ+DU2+OxxflMBdmIRETpFeyh+2H0o
+AzvgjKzfPtgoLIdvkq3/RAhJycS4YZxl2sfL4np3RRvngN1ajQDVo3hQuQ7oYrE0rCoEvcgw0wQ
bl1KCu7CqNDP42BwkQ5uAmZCh/QDN0ZzIhvVyTrPxEFTGs4Bhx/3gvfJgRP5+wt6f2ZWP+4tYh0e
pn0Xg53oO8pnXo2EtKoV21RdjSFqM8yN9RUqvmk/WJyU0fI0ycL6E+95gZZgvjVHTdXcAbxSaej4
a6SFja28VCeTnmivpG8b5VTvtN7zbk3fJcSWhcViJAdRa0MzjjrLYk5UhqFtrjDeLEXtQZEKuTkY
NsvgB5HTDLGNKtOid7fKVupgyvA47VqFt3LiG/9LyU2A6xXG3oKjSRSbYLgZiHOW1vTPCAtOqCyd
Vm+JCCcucmxKWSr4kh26YnZmVVHdMz8nOXmYvMi1m76Ra2FXnZkJM9yH8RDkF0fPAilRLAGr/SVO
t4tAnmwsskm7B5cCDv/XhmcRS9oq87m/eiT1ADGdLfjf6XzE9oEJ73JDEDOCbVtNIT+SixySvoRS
4HjtRAEM3W1y6jBu0sEQnM4yBXnP2GqzRG0nbxo0DbywGgzsfBi9MyPedNRImNdRxQJcJRqpUdJu
+1VyUotmZX69Rv4/FvW26liK0LhOe6Wa32IBI6UrPvYda8pao55ps1ypTrwDhRazeIsxRYXRqNwX
Z8iQ/KP/ljIZEIr0Oj74A6Zk9o7vX1XTLSLtlOjGoLER+R5zkln9j5lclAHmVatbbIF+KhB9aHNd
ndblQXHsnkdf6qsGmx41RQ3K9w8KPwxcemkegC5raPvYRsgJp6/+2cAyYoB0O447BmF6JVMw8GuI
L609ylDTcGmPZRob4QZX7MDOc+ATtT+LTnSNWhyAhpz7+xj7e4dXyd9KeWQl5uhG66z+1DxPCslw
COJvc/vN/b+lsXM/AqbyoQDN0LeuBAd8m/VhK5dMs4mrHtG80Yd+R/zpvCZmAAfdc8xUvN3xGO58
BtLCDr/60i8qkCxUEHryN5GPfF+y0R0tGWSKjBxm36eq/r23wviGIc1uYGoXyC6VJS5jixva99Gz
PG4+322yCfjXv1GRjrqZuViapXVZpu4McNj1DmO4N6VJyYqnK7eZRWw3a/i4ZAB27O1F9gKzASkL
FMq/yhqMtJNz4ADSVcdrH/ulAieH7MwVKt+tHiDATM1h5sBsBIDgV9ySC9bKhjS4/HJPYzKKgdE1
GNI3rfBkc3dN8lXJfVuvkN6bLzY+Zkn1AY0wnY7ohv91KIDeZ/0xSzKfaP9pwbjACkgyeE6fpb2e
iUzYNB+E6aeazF+jbkCbnphZdNV4e9891kOY3GoBDOl+qYV8CBn6reZrDEG8dM8HIj2ElsFm+jwL
gambshABJ1MJsBTrLPHlym0IGAHXOt48Mgjaywebvk6FM07SRVKsBuZ7r/9xG5Wey0qSvm7Ff7Eb
EGoU7TSyaMX6y8YGSSH5Arq9w3Cw+rfYxGKRTVpMyB3EAx2sXWGJ1RJEZt8GteOTmKTo/QlGnCys
s/tpdaolx9E7801FcjBi5NVF8Q68kXmx3hBo3YYJXeOqNexDCPC6+jy2ZqexrlKjVd8Muu/m1rLE
prYzQyOC+VLTP/17198X9dwDHY9PTzZiZSsCwiMoTXRegZ54eK1QP8kuRMuuFndfHTVqRAZN/PF0
XEJ9FovqbOV7OCffVhTdzNpp+R+DTpjO8GlQ+2PtbZQhAdpGEo0HNLUi4e2kOizo1EAreUNcR5Oo
ZY/nxDmDA/W2FkVQnfaOPeWNeTITswF1wq2GebbfKi7/cc542/RJu+vpOF0qd4EYcLOYMJrWX720
G5QpHMY5umdmk25TLJIQdcJX/FYznnm6X2d+KewuZCRucIlQkNg7IrtqQvVitT62ixnRE/eIf6yI
9rjvKM3WvKhvovIWcVZYesDMe/GbpAh2RPpSpXBmwjSzGa3VuunqyXpnDeoK9g5y2qmtYZyK00VU
3CW2Y0sOWbQayOVdDa9kdzYOQKCGKtejXLn2OOHNBNfpgqnfGgnONV91dwlUlI1OdfyqD3popaJU
TI5Qa3KMGMl8NlCnmbG/9TIS0vrP6F403BpLv9tJ5N8VtxatCfOsa4RFcQYst4jcustvw+t9/ude
afo4+D2J8yOxfJiF5nHZE9wtoQFGD0hir8h0vVlAlRpq++cd/3D5/a2xRaPEElrdTkbJlXNAd5Cr
n3oFqyhd2QxntpZ5wd+9ajyZiZ5/nFKDb7gmiWQACbZVatH0C2OROj+QR6+U874lZf/xy3mRhMTW
aRJjGeXyf1JvtDT6ELiXcF/ZBfyvpssX1Yb3bg0vV5cZNnZhwjweLWRZenyR3V7HvnNTE+RFC/pD
pElIHxD+V2sV7mzdgy8OJ9dkQXUhb8sk8ajvPICBhLigVAP3aGb4etrr4BM0oElvnr5g9dCw/OSK
ts1OK4yI9HVjFqydTVyRcpgamukaYPjEATIGjCwHdnOusI4JpwvRvsZaC7HgQiZn8fs5tK6o8Qu9
i/x9BaVPL7L9xsl6o3iWwsAGoHCpcHb9a/jv10qIl0ZNzUYQ2PXzYnzTp0M0yonM1MCHoTjQ3rM0
OlQLVCgZM2QYBIztJvTWwUsfazc/gDZ53nUehWdWxuDYtG4DJJ9r+rNNgnp5AgrqJYd6kO2L2Yx+
4f3NQY3pWt+pFPZsc0EREv2NcWyv6O4UO85jfFRs/l4xZGXyBrOJBXvnAegux9DVxsgRJj7L+A9d
zGza+U96vRSR4WygcXlQr0iozR2FxfAGx5Jua27pfyEyqHpz+0oDns9D/RguhgGMV7e1yONqkBHB
dV1d3XAGSYvYyLUUsqeAcST+ni9eWwGcM/eBVBdkLMiIBggOhJNR368NDmbZV5LuPJLiPZwXPlzO
dyW1dixd9dD7U79RrbONJozEEZWHcHMqy2wyup+oGnxAW+Pc1bW2AEiRcjDRbrHzPcVMatbjtjtq
ojzEfeaR3C3myMBAQjb26TkV2zDjxOr7TBIGKRtCB866/pGf9MNdpfoUU8YWy65QEROdH+1J2rq/
XevQ06AW6suAuzoRJJM8NYXqzbYvv4BaPM6hnnw8RJLuIEUgKRCtrTZYr21c8FEnKVxsMmLp09BX
2NaiEoAm/PhevEBb09xjl9/X/k8yBcNgPEOtTtOYtux0/qSiHpAOfuQJAiDObIazs7wNAjhWs9O2
RZFW2FjAtxr8P4LJ/o+aI+R0gaTSLWDjz/DawW1VsGvIshEnYftFonvsuVUXRmcONVtHD13AqvIS
BpcKQAJy+xGP31lb9hInYIHcWKBqNBbPWh0Wam3o/h3Qfl//c7aXPASojQsGMEiuxtmxeogNO96m
n42NgRYUWLTMfme1ln8XMs/zV5tQNoE2yE0yaeMEZdE8Z+8omozpJ8OCh24CS50W6vT6dgoDtsA9
cK1zWtyFgikxo6yxhCYlAO4+TA2l59pAjvySS6693bCnqySqH4SCXvq0DxzWKYOoO3LkHLC+qEis
tCdS5YSZ8OFQEQK3gFxckjxDtgHr2aa7mO/3lJSe3XBno9gIk6nR1f9yuV9EYPHZjYJkLryTWHo7
Atc6oEQdpuCMCU8JQjxOqCaNA8Ls5d7+JW8sAVyaCUPu3MHfjSULkhzx4i3N5MesaIcK9dK7opUM
nUD1hH+4OnWhvb9hsO9/Yi7sufPPpTiOxhcN8E/IXUpGwlEKpqsSAlEqxbgERg3LrFZht+JVm2XU
ueX/BERe6pTT7x7tKXIlhEKxrFgdlrROfoD0lMXpJC63Wg4hjLpIweJEIveeViJBbf+qMI7FEQaz
xja/OLCghec54sadAxQ0Q336zhPagOshSs07N52JPn63Uneu2vwxkUzUjX9XkYSw0ODtCAPZ7pjo
CTsyg59Of2niSxNX5bJqRJcAxfJdthBPIQIqg9qQXvJxf8ZDl49zg5aMzTtQWnKNdSIHy8rfZDbV
yvypR4vkfMh1wREJps+Kd4dYdlq8upF077voS/NKjkjKo20T2V9T+qsZsqFJ6zGy2o43j3Aizx6W
qb78j3r1Gkols8rCOeMaNSerXVZBg4cdWS1M4rIxif+hG9qIIaD9G+yaDXDeMB67a6EFgVAQszv2
9nvXw3e/mq0w5WRvkExtySllIN9MwMXH8wRzQeovZPH6v2+GiZSEe8lo7DduYJE3I6NKjxVoQ125
qEdSoTWlBH4hqZNnckI4N1szhX5Mf8DnbjnqQpG7+bz0UeIKXXQYYy9JQ5b+8dAPkuIXrJHNTHBV
v+wQ++qvS/VasXNeGoHCAA7+Mqa16jR/3d5dw2kUzt+kOhFMXWngjhNZ8YbZITPlpzA3od6I+2rY
fJVivwDLHPi2YaLdRB1xY6egLx3HTapUhUJLb2VshlmlUs2Q54ID8d3pF33dD0kdd/EVaxn13dxq
jAlinwOfOEQShUyMmcx82uzYZUulSIwoJKW8VpzEcb/qd/U7HCEfQMcjZkzu5KV1ATRg2fckaLS7
lW8AkFHvPaQUbVd0LvU4X60piipW7Az3DlISMEy6PLgBvwoZ2yKZndS/bHxUaFRH9YQVPpw82vr3
PO6ZlBxSxRKoktPTcqNBg1mpAITpQo2YObHwue52Ats9yLyUmWt27Nf/rF54Ul/E0ESGr3Zkyb/i
WxpIOxegMntiv7STFWBNNAWN7vPZFTvkVQGwx4nljpqOmvbQjImKRjMZjDatuElOWRVpeUMNEam6
ub8F5MFSbJVSsPQZ8/ejNfEBtkYlLC6THW+6Xd+dytahCL8Fcg+L/f/E6rZ7oNFr0abd+/Y3rPb+
NlDq17GskH84/IbMziLsotbNf/BkToEq9Dav7DBd11LzSmfQW2yL7iggiJ9OENVeRy1v0Nq+6nq2
FsmmRT4fFwQG/yHPV3Oj858UVmqpeeeQobE3lYhLJJOD5CHll7de3nTc1pR1C9nRhoCEunTIddlL
TQ63107O/FgqTHwIljNCp3BJVGs1HGCeM6e0q0g5xKlp/he3mXWWvkjoEcSue054ciN7nSLCAGai
/5zHAdIpEVENc9FgrHqCGDJ9i4g3PNkgZ+h7OAsz9VlhPqImk7kgjLY+ucuaqCBkMFf11Uyuj4vA
AiQu4gomE/TjTfQ0pb6S3OPyfAt1mB2+w8bGovfLL6d2PlrTos6P3czGktVdcBuFA4/jNo0jr/0a
ik4Et1bVY6Mrs/oeUCN6p1DWI59De/tneHON4ICHJtthhElp9+IQqspXZ5CP+Mt7b4aQsL+hBVnh
xYjMTQqarmIVyYXGpU3CM4w342aRdWUvBVEKIUFrHE6FHukB2ocibjjDMgylJuD+ndke85krdxFw
lvjqXjfHDzBVstYCVtqMdPxhMZB+rZM7FkZiAkfkxIYx88wcFGFq8vuqZu3M5MQ+JaBMyyP8tO+p
x7lQWYn0FdMBY9BKg38D54781t5h8X+V15SL2ZXd+98VvtWWf5PSc0bdkxzR/WcaPl2ptQkcDxtb
NNIvqzRY8vAh4JAb124sD0lKC/PLzmdb2QR7jx/BkW4cnwfphGW2neFLA9K4mTPOXUHx+ZNh6OAw
K3nIZ/o9dhKnVSO+sgCxD/qXq2bWRn7kBRwjoIN8VNpVex/NbPR/YRRbZavW847owJf0uFhdhBl/
agzGM5AyDRxkEhi9EKcaef/4Sv2fKkvE+WjufN90huLvyhmk8t+AV7a5KBiPyZjJK2ieb5mT4ZAL
qmLMuZsRnEMgkCLp13nCoAKjkVQ4iIv4PBJUSr5HbmP60/95fxjynWEB0K/zLnaF+SzJDWY0zKn0
qrbFZMK1CxY2YVN6wKyM5kkmpLdEotqjKkAvnYP71qJCERVAfuhIDPDvfrphdDj+t7ydDZU7se9L
znBVSnsIXOrNQUxU+lRlcdCTHDAwiiBbQnLZ9HbJg+IQ3nu2TBkR62JUFhIkY1jxFinIECQnVcl1
m7ThYxWwLKflxG56YMScf9FAvMyoeVPy2D/orBbyD9pPErGjc1vfFFLXXUC+3BwNH0X/UE7HZ/7E
8H1qVUwlrUVrwb45EGD9a1V+VA4sWR2RXlSwePLVQnoq3U2/0bc0+zk+qFGznfwELGXdHTExTDsp
FLnjYLZ8KkEIx29Bm+FhULJU1sWoeI3a91vhPVIPcKpfz4nTmf3BNXV582e/yICHbiH8JhnaMxry
nvNVmk1ZddVb+6hpECO6Z/I5O7ByLNjV7N2a4Znqny7k2+RnmMR2CRpDuA9IrnlotbKYoxxJPdMo
ZnhuPw+c8mgn9LzXQqmj4055EzGAwIKjkw0mKGBsCQ5AMnK2j8QivxslUYa/oV75Qma5Ksk4jbfL
n3tVTyEGiJImflVaQskRR5wOdj4/7KU0z9O6PHT4ei7KUx0jm5vRtqjMIx1JKWHKhWDt4Pv+8iJM
R8PvxtMkfHnoqOap6LajOD7opZffnS8vcYAZ5wCDoI7YsDCTVqhUtl04MGgzZEdUaK3tSjtY3VxI
XTFtjhKFCwYv4g8fxMcCly8blCcb76k3qRzZX7LqLUuXzjb2lfuHmYrR2g7FFVkfqAjNg/eef3sX
Z4McmDbNi+YyLq1LYc0laVY1oR8Dfx3GuETlFM8PRi+pw8K48YRXoMu6hX72Bqoo01+9IvHZwu48
2Y9BymTrRt7mktheCqycPMqKy1kY7undPm7DspHfDOXzc1VJ7enmucSrkEb2sJdvF/4qjw/d6C8q
Y+YG1ZcAN6Lo8JlnFT91JPK59app5g89D33RImZ3c/maDw0UK4vkeHengTBfYFJDIRzilKqkgzDQ
zgrS86OWLx5UG1msDUp+cvcTWnugpAxvijaidw7+DW4AvRvya0MWv9hdHUxhvFiJpxRtIfkm22Qs
kfn8HNDycrPJNtDf7hzVaeFDfWzwM/x8PyJiwi3gM0y0DvRn33V060ejJ+bUdqAxCfHre2UkUGIV
wCLUvn8fUqBEdbckFwEd9a8+66t66gDyZpY8EQKwiYa0yC64K05XuzGEsjqENOm0hDuJGeKpRZDp
ExUVKKOYuLCYCt/h4j/yEeNL41OXdOUSQ+iSzkTBqUyJmSgTA/zeo1xW852W2Mjx4GxAM7oPVJvp
UjoHAMYzrLg1DdHXoygx/KIc5jeidU+hoeYszW2NOp2vChfNZDwfRA87VKfU4FG/W4oecs++z++R
eUFmqw4/Th91WNNBHsXdizj61kCj4HoJASiEIjr0FIfTNFYdyPjD3yLibePfL9z6tqd13Vm94kYJ
e1kmXzLmrI71JQ+LONnkIDOGXF6siBrMMeGxcil1Q3AKO1+yKyNzcQ9whsBjOnkVvc1ow+I08Sro
+2aQUIzf2eXcZ7jWuQZT21u6fO+UB4ZsDHbA+qrKoi3lC+GzSZanX3OiZ2f13zMV7NIBpy4SoJPf
4UPT8tGTcsxoStNFv033sLp1HNfx+oh58x+j6LeK0X69nfewzjutfsHlz8DoIgpnntVbX7rLdBp9
dvRJaYFoehtv+iCwUPH7ZbKbbUT5vtQMtfw535bzS93tuQXEOBfDsbTYj1lZwShxZvMzP373BQsy
+PD0mddkrLSmzZ2ZJ2zXIMXtlWUjc+Zxdo181c8RzlGyH06YKlRgk3hTvbVwNGUNEoxJKtR3bdro
QA3c/PlqYh1WGe9dKlN7raFkB9p5pfE7qN5NIkof+RtNq4n/Libk7JFp2KlmkUPRnSD+6Ak0nK+Y
zijqLsEoWNmjT+xY5Mp3xFaS0DtNn//u6/03u5ZBmxzrMDUgGmbSYFWnPWH/hKUSBZJ8EIvv5kLs
xHK4hOpXqP7zk9C0stjFZjWEbkoz/RKgaY4zBeeQOJVBpuxOaSo3qbawvHp3MOZgXh8uKbw/wPdn
lGl5M6gV3AOA7qelPNDNoVMFuYlUTye6efzGOk/M9dQYkHDZcwHA4jjgQ7bqbLGGmXsG3bDexDPO
G8+YIqkFaPRhg8wb4ylf6npeIYCfQpyiaQkJRsFfa8RsvFM9tWrT2I6vkYAelW2j8VGUzAKVUYfv
goeWJ8FzIcgDDOlxI7cdiFHsvccr7lF211jkISr/qEx1UvmNCLltnuCTls+k1bqSJSTZj2DK+unh
WW1vvL0GKjpwHXOp4W/KuTcOPWYeNUEgUD4PpYwDU5X9zt3HfkcCRAoxs7K4sb+cZfiGpTNbbOlN
PFF2VEDqJs4Gnx3qznvYql6JXWctzNvFxlvQEw5tWuefBEtLllzCsRlUcLiRLmio9r+9eJmUOpG3
G3aA5fGN5T0KNoqzgmsKuuLhGhZXiX195t0TG6/ov0MS+9JwiAld8WziqizPoPvQsLps2SdyJDFz
+Srm5xxpj/Nb5yixy5U9vvYb2HCZ3DySQC3x0JhfHgevhL3/a+yJR9ExC/P4nAEhESdxzL+kV1cr
C6wu/1zjvyFIp+Ua1HLSB3KnsS74edARHi8YcP6ZvS6qGmCZCO1ma8wlyGwpS+tlWSfaQfJ8OCZY
A7gruzYJezldZh9Zwcl9WUmI8GzBl+E0Ta1zvKKDTxJwb+3PRmIzdJNXG7lJjWuDlBMiz73Tn5uD
06vA96rksw3nXtceiaZEOFuIY9285G4Nn4xOxTreksR4ZJ8Iv/ETyxsNzxW60Mg8eOX/yj6aMvwn
DbPV3h2xALVSAulVvqE4/P38yrM150T38Kw/6M8X54V1dAbj0+gVUTWcUpA7kxV+rM/JAVAEKBSU
qJsGKTtrXmF4YZWZI8VSbXR9U1EdjifWXxxeFlSBy+w6AemjHfZm2riJM+sxF0Qu89zjSgAJYe8C
fy/E2PL84Yfbe0NSBEY6XmsMLZJZi/+JTb9aFAM8NL60GoAighIl48nM1NxJu4f8S08DG2oWC9au
yOVmUrVO4PL2sSreY+VNgpfJdskjWOZO9+22YSPkeloBBgCSF4XAs5/hu+EMwxPngi/WYJqqrq9d
OPdonqavTnICHKXF4LhffADoQHU0Vyk/Mhf/htMVwZgfEwU0pEql1G4W1kXqgga4OIgbKhj8wEjH
UudEseIvV4sEN9LTVhMENViMs1e3z/6kB6JV7MBv9i7r/rYta9SVtQoYOyHj8lBW8YzA5HXHs211
Vb3PqwrN/xiV+aDDPbSj1ysZOUnMFnYfk5E+DVU6JUKkGttt5uaXd01X0sCGywZjQstm9CQiYxOy
tAyckXpIlz6z3S+nj1T+QZclg0Utviexz7JzOY3W2Ch0S2iaGjD+o2Ll8Lpm2j0o+P/1Omh61hd+
P20zfucd0jnBUqPaF1WiPIMBIp5NeSYxZ5J0IPyxL11U4Jxaapt1aYXkYjJ+j6q0mopo1q21wX0K
rSDu+ZdmrL1IafYfPEaNeFpwi4p3caMEpbDINvo5Y3JYKQH3FyavAqIf6YXj95Q7MmhnUO5wkU+g
d7MDErlxvFqwoWJtdi+YmLmi4rSwP5B/pRTZ9BBpbJjcwcsoE1Y1i4Li+DoX6PHNUt4VJQuiDMi7
nlPVsbR5fw21+HHO/Jo0aMvnzSs+TXsbAEdb5UiX6yPFz7jb5aUSKnTGBgdRztgeSheKSHPnFAFF
ZQ9OT42WI88jn9HS7r0Zq8oZ3f9STtCAi3tJfJWxwgFPKl5QoGuwmJ8nqeeIryfXxwaA9YzH66YX
ayOpYAotPgrhYQW2ld4iandwerq6PNI6kgzLRV6cNtbi5deV5FFAmDqGTCQNnepk2DfiLooiyPNA
gWM6kbjj8aqobNxEfzpp77odDwCpRE+518Kodpc7kya8Om1iQDWejzu3emA2qK38w/By0YqGJZNV
gqurWCv3WAQ2GZe01qGnoRgSbnRkKxl2z6rwEdoOjWdxhyvqEeqhoIEMwqLVjmYxkJLpd/KqYJRO
sB/hjTikme10JTSAXEyHyXjzZCFi29Ww0qYOOGVeJ3lM17wHkN/nSUZh3gXPGFZd/i2OJj4PJThZ
TkpJZCxrTJkUHELEhplMz2KWb3QkJhAW7owkwQwp5HCoXUOyIMHHzL77dP+qv7cAmk8ak6O+iQrz
c5CPPGcQOOqWNjtBIvoBtOgOYonwavjDk5sf2F7G/soIGIt+QLmoCFLrpjT+ariH0j0IELRLP4JM
aD7xQiOD0jLOxBL8q/FYy+3MpbRc56eekGRGAmpSE86PV5z2suKKt9CPA97H2bRp9KnwKuvRLlKI
q37bWPfgCJnDDUTetKuLRSOyvj2hZYZgLAaNnldIgJUKRcUeyvBJ2E4HA0KXpxVXm6tRH6mMKNPI
LJU9lFch4qtn6CumCpUzMfMTIV4CEh+KIQjwknb1/AYvrL6YdsEpG/RoTSTgq51bEccPWoghRu6c
3rb1f+n4OitxDNkAoyZTOrk3L/L03FPaJMhrpqsh3S5x9frjZHCglcDH6CAAClLSeC+JYzUSD1kK
k4hPdQ+5WvXvhxgSiq2gDJ7wNMuW4XWPkmrXbgnPObRfcM5Hzvwctoqvs5gwOls8WhLMzUBq3zyb
JnQ6SGqsvXCZssQaNxf7DAW8w8QZeQ29ctabT4ZbvgvO2MFvHIWzMZSqrehZP9D70DUedlwdM9kH
m2g8VOHTG66ujm5TIvtxGRpdWDGaAKc6u+Zrvdhnew3agDa1/FndCuI3TMAdRadplPKV47DYUco2
81neTtqI9wrS5Ojv8+6GyshaqvDXqEozVxnv5AYjTsM9tFqlCgIYpDu8GQ7nOsSEBb5Lp3MzyS99
S1vMHdWnJJz+mzzJR76rlLNdN97wxi4rqn9UqHAA8jvBZhoPnpViPfd8dRxW/prNamu/OnB8hDKE
n0lLYLbUQrhZPSrp8wapCa/R0ccvvSeGqCPrTDEaxRwrdUZ2ApqQXhvRkz30CLPc+jPjLRVvbc31
27jk2ywthSGGJ2Ae8iBtuyPN8uAXomA1qJE5yeYV2KXXI/bm6jDlqBLITXtfFMz/e6mo3vjF4L0F
P1XE0rICFpyI8pM4nt8OMIpwBNaSO9rPqf6V74ug01gvLo6yXd8a9hJN+3ICK7ejn6csY8La0k5m
zezsUTzcF+i4J4QVm2Y4b6LyDGn/Mg2Fhak52A==
`pragma protect end_protected
