// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
EwGa3uOGpOm/xvDZuq7gEHhc8+2cR+7eMuSjGgv7i/orGGrX7gMj/qJXFktK2pf6/1lbm81f3dlN
h4wYPaM2uj5JtigCWb9/kyFxf2ExwGpmYQYQlnD7QfIrPUsqX/22HEpQw6DWpF5ug8628MjdUzF3
5Se+s89yyYTWYg2mE8KjFaEoLG/a4xkh2iEIhqbuCTpakMgDYv/7rozJC56IXGjb0gc670OFw+R7
MQz27rbSfVeriVtSai3T6vxMZSiE9V/SgLysYenuY90O8EX4joPc1feziCSiHvl309bQ3AhuZOcy
CLsws275WJ5CbO3uxGXoHEKF2pA89GuWEVBmag==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8512)
rtCg1yGdZgYT78OsIv9pG6znP7Q+LqVSXtt9LA1uBgselScmaQ3ohUWflyAo8NL/X5wyVu4Kj7II
2qbYmcvYjzsDFhje1/24h3EK63lToiTyI2+ijrptqqyLuznecMMS6XLBGiZKeNMet8SK3DFOiwap
/MyLebMa0xTOEAlFKdec99QrzSDjiPBTZgY0c3+VidDv9JPfCXhoKoByOq8IPTnoh+DUymSLBqE5
BFpEtgfEAkP635iF5Pq0dPvOm9kern5EWAxxgoBTkWuOEBZY+QXbab7lBsNBFZkxhMr1R8f1Cr9H
jqL3MAXGRNgqfs4iZoedE+ZOJIunR3aI5vFWLSD+Jd9AeuGvxKLzweacOM9D/OruubbifcyXFJ9E
BGYY6FqT0IAXd2rDHysFa2lVr/0a7tWDbtGrTsZcknGJaLHFcsJrJQEme0UV/X1CfJgEH5FhwQRe
W+II5FycdOeY/FL8Ufn6+e5FVdDSNjf59231mkFIl2465S9juTweDd/1f/7i0eZsCSp9UNsn7zJo
eEOxYijtUKtts6oMCXWdSVD6tNolbTeDmpQ/tCbEkdDGOreoN34xQd1ppW9vaIpph9giZw+dxVYs
1NXX8KT7zUjuDIphTqn3wFOCUd1z182E2plfdBVkvLKHxgpy7sCBfn62mtCY7qlzZTWDEcEjmR99
Lw0Dy3e2gMGt4JoXLjLDWi8p0eS5f7Lt8nlafXKN+Nt6KcNHbaHTXQ/0nCigzcavtdAT49qg/s/4
p8ddMsO0o5vIUt9JripHwQZfctxYJEG/mZvSColB7CwoDIU4zIMUpQUbudQ7bUwZoMLyjqZooWWC
72F2Ddq0XuXnZbIoUVUh/FRRCy5aiezrRHEssOhKNTWcGc2vI49NJKpIifSkXM7FGwDVXUDiRS+K
HiX+FG0tjyP15ZR/UCTToCAxyd41PELzptyK6AFzlRdi0CVZVWaV0nzljGzcB+RemTHAKSIEmHok
v3OV57LRrk802mUrxm0BaWHX8sMx6PMUIDquoMkb0vgIPyn8lyoSIIy+Lzrtrdp+U6VZb0mSYhXC
+2nTgjkCLGNqGSPq4GZnG4JVOCrCGXTFqWaKAQwstVtMNLdgpSeXo9tDI/HvDDWck434CVzokwuM
oAgDYLJ1C1uhV5iA/Wu4NcW9Y4o3w65AR2dy2BJsdWl6DzfzHg3FCbrMCR42ksoRS6BdpvH1vfht
0f7wS8FpLtRMjgV03d8B3jaVfBymjGHSs/ZPJW8/iyRBHmS0LXi+fO+UZo9G6xnhf9S3lWxKFPcZ
c13WY0wV13vwkVmde7014CFfRVo2pcfBrGrPqJhW+pj65JrbkEuMrNJMzYQl+M7z+wrsxYqUONgl
lzXAj/gVrrVKVlnuCRUJMjBncpC3sdOUwt08p3qDjSyPclldJRrUvRjs1xHiFRKYecIXXg02wvwt
OniMVg2ZvlnPabxV8zPEWikC/eQ9h57wq6zcOixTUaSzLSOI2KP83WsoM4JpjQw8RuLQxRdtd9In
ftF8BYNIK/VzdK9Wdu7HF06E4+T2KS+NAbKCiIk7KTqaqhUa/nWkRTZj3zcmdiiwn4XsTrL8juRr
gxtyHSZ9zAUYC1KCmyob03g0KhqPlHAdbJxuSPXi+ugp91WkwEfzxwbacGdPZE0AbXoJ7R2La93L
4D0GkHHgl+UytVajDLdMT1fkvnoONJfEjJwK+qNTDUaqx15g89gBGLq/2Jt9thzfDagGr8FyJjq5
ZWm+9VpPV1fXLZMvrPSEZTyDQak80hxp9D4zzMw1Q/5oUiisp2Dm5JhVAJJSmG7iHGAozWplCKBv
Y7GHr3s3+tJ+ysJsCSUcHn/VFatzxqTorX8ltH1f260UyQHoe8ZmZ7NgG/tvXLDBJ+ThCisywKo3
zAbmAERPBBULMq1uwS5Lrq1b4zVtzECuHzL9NOL7P0aR8JWDw0jleJm0wHvb2ejuvStvjR+CEWMl
OON28hXmLyBLnDj4HthXGpoNpbK8qN6ypjCVncvAYQIdPrKlVK/vqsP1MduwGdAKf0Rnn1xZSOZg
1meSqufSaQ38WnMh6kt6G60Slwzbz55KsGvHJVYMPMOoDlbBkXPyKqr77U/htWPl1psoliU9PfJe
2hj1/bhHvqS2gonXn1cRviLKqL1B11JEBmiPnPk4vCdMM3dfLuCwI+jweiZfg8qxnCnRJbJ/5FfB
tvraImj+ocsIwI3SfAfp9kgZ1LPFBP1rM2HnsnqkHN8aGoU3old+ZxKvIiz+si5US3zImlB1rN5h
ihkQP5sb5WePv09hli0vBq2Pxd5r68iXbl4Rhwzpwl/wFalr/gabDN/fOV5h+WsKfWGoB1SlzFqW
7U9RZbpIY8PiY7Fs27ZAUrZlJQ+xd/iEJYghUCsdDrYhiJzlXj9MQ1Tz20KYa5R+rh/3C+3WV95h
DGT5AFPpai1qjnqmjtdFqpexbIqUA9ngkQMw/W08+C4sVksuWY6l8bfOheBHm/CbHHOo+gvjseWC
TsFSmIk2H/FkCReXXs+dnz77owKpvH1/NKYcrIwuiVfTh0+11/+YGQwoFemnHHM+tNJH8WxfZsz1
IKpDxMNgmxMfz0YFxKN87BCuhqo7qLa0A8dOWB7u0cvJfg/nRlyreO2xrfhbKdjIG1qCTrN9BNNb
8FSTNuY81VrqfJByQyRVYhMGOaFN532+ReICM0n3gk2LpPmYbspf/eX7zQf4KgX5SfKlteG9PzFH
EJuADh3NUVloTgieeOeIbcvL4WkcaLZK9/oP4FbB9lOXiDK/C0klr3yWmNpV47TkXk4M+v5Yck1s
Nku3Exwjx7ZvnFbF7pSNDdXNHbtp5Nz7WIJ2IlvtQE0XlGSJPnJovH/S/8oNH0RnPhdqx/o5O/Nc
/CcAqEmhHU8WfGMO7CN2iU7FkT/RkOEXMWsLGQ1LbEG/HOI9hhrjFBirAleoeJBVY2KJSEeMa/qm
LhN0Ioy6a691OIrf7ZfaadnCHVKhLElB+SfuYVXtFISVzQctuZ/Ag3FWSHkkaYstoJQwIR6kCgb8
94QJbscUi+JF0fb0JO02lCmz9+x9/fB/x4YEx6gS50v40QkdP9ldCIsgOhf4q9d/7D2T1l97ztBu
knXnc6PeWGS0hR875gwmvVg3Cyc1FCwSWQyZfWGcRiBgecGU4JkNyw4GbU6uaEAVneeDucxYeXV9
ZiBuX+ugX9NA5Enkb4hfI/+7noZtCXYeAoVVgRUSJJRTOARE/HZbatQidsZVakTmBjgAmwiHl1BS
r2eqlqB1GMF84GzSfzMQNkhsGdkgCsfgbE7VxalEjH8E6GlB5bdyJWjgrRxOlbiHuvsX/jrIGiMo
8MAvmsrJ7PSNrJ/u1CNt7S3Ze0um1AzBEPuLqgjXrNxR0dxNltja6NaujTuoASaEqn5bB5rhYduJ
F4tRZijfZ9+bG1sfzcvuwXBz1GuoiFb/JB2v9bkY6sdW8JnE268hSfrEPGBNHYDyaEXzDSW7yKVV
lkElAns+KnLc15kHc3mhe4IlGJF1cw3Tjhi6g/1MKOzmBF9FyGM56+ca+/q3PO8yi6FkTChm9aG6
xzARLdZ/Ak42HK2c5Jb/e/RpGvChE+bIt9m6LH62uo1vsDGNTwXTMW4WxXxlRH8/lafUz1aCLoaW
7wzHOkW+52NmGC0I0mgo7sMq6lsYqQacFkMbP8dAj8QI+6LxarmaYo2vhNY0kof10VA/vHNF5IJb
Fox1CjYvRxJth9YCqSsiM9q1pRkYXw8EvPCAFOFXdzk1WF/RoD3WAkI2BLZD8ej7k7J84K5PppJo
GLnv3b+OqYa/54JyQ+DQIbNl7Gf03sERrkabCTYywAQyz2jQen9g+sHcGhKzAZlja67a6SzwztUF
qZjW64E8Umc3Z/tzo6Iqv//+LQgnMN981EWFtmDyEs/xujrSPGlwHJbuJ3uz9xRdpTE9xXu/g2lB
1WIPLEEVAGVLIw7KdOkifjFxhqtz8rAy/fczTJlFiVaf/G7So/TrLEedmnMGqvtw0FdoLzoyLLRm
Epsk7fNDfl4y7+jcZx6NK8AiiU2OmJNYVwuOkQCe29oG1smmiz7Wag1DnGKFLVDcg7PF+7OUW6qJ
kSbNZ26D7b5W32j/zAE2OjocGfYAtZTxd3IFK9Gcw9LtSyKjEyCA2NjYpXUKS1CJBBAw18G22mx1
dOE40bEddxbWwVV4jfzbCRbrWrfvcAAp6TDluLFtWKqKo9PQvMT2eOdRBRGXPOlGxrTAEHE04n6e
ucqDJflUdlD60L4+SOY+Cm/Y9xgUHNFgq7oQQwA9m7NGXIwlneJe6QSO0ZlE0A/8QtaLAa5DDIt/
g5p1qNlYzt6LxbTIsLmQEreVno39avj/ob5rPfMK7qDNbBQvbn7ke1kPQHEwhkFUX5Z4gzPh9gRw
KXA8PxqeHbxf/Cmqox7Wyn6j0cW7wjlt2pQ1fNF3Q1vpQMjcukAjYkQEqjTczyVOeIkalY1Dp6hq
wx0rN/k9MNuRTrcTNz1anUPUxbcV+zudjRRKzPlfhCxLg2ITlUFo22qWIRFGJ1eb399K0JsmYp1r
rzEAc/NSxgLwnQ7kN8OHotkJ6bUjqgcF0Ry21jTVK4JiU1DO91JQzPgCIh0IUXq2pkGKLLB3m4ZV
EZkWxIWBVoeI6UpflZV+Fun8bgOINIknTt1yBb0wI98clph6zNvb2LsZwgIvhuIMTDEZW8Y3jFIf
lHvhHphvw+oTllhv9H0L+Raxvg59I7z7lB4yCVJb1aYjupWemUwB7e7dz3fXwJ3l1j/6gu2sptFj
BPJRqiqum3r5X5380BdlSISTbvLnkx9Lki1PfaRaQ20KrpfxZGoJ2W2mEXjFftjWSfj4NzVf7Lmd
AXl/liLdJ8kFeWKU54JRdSVFxJaijFaHvfqXy4ZtlC0JaBi1qWolJ7WqYs6qgT6cjleyFsMU/Qlb
Yq4eFVgCGJWfjvr98sPXx8qsLzMJXnLioj37QObds/Yr9oGkIT//zMupFNpO4tNRP1dnXdiVHmwQ
3grmJuS9Rj7jHC6Qk5UbKk4C0dtKF1xwlZJLnu8M15zYXOtVMcGCpxMftpszR3j9FTR7kLVsyZe+
/mSb9uvDqEOjNN+th7EB6k0l2qCy05DYK/9/tlABoOH3Dff91PgKNjMDOft2r7IvjGgCITwfxX88
B7CAFCQu6wqBcCTISRyXomLOSMg9fF87Pe+kigYQnT1yj11t8aYVTRVo8ZBLdyGkaKObWJKvqFIW
MUKxqJBbOuXd4jRNPBhMhwZVCEWW0o1bo7fk82erAzcjTgI05483OkoCjFfgnHeiWkMZZc7QlW2k
kd0hkw5eZHclJVUpXlxZasz5IMAoYJepJ/3m+QZ9bn7G+yQH5RjG2q/IkibVgHKdwuCAVW3qNXiF
yxRRiJsvbWzPph7YGOZtP3h72QIO/rsI4AuTRDNjMX7rMbfIOYP3UikGxOGl8mHKpBhEznlsu9t/
Km94xNA/IUsYQt3rstJA0JA9eWwwh4cd93IDlOeo6GLcEcCEzK6Zsj3hoc+ZwSurWT2Q2lnLveIA
uD1Q1vT5Zq5fpDtSFER0JvJLL4MVIgXaFiPy9cgR+cb6wyqdedtOXxOof7L1jVrskQHtfFBdiHQF
7LAt/Xsjj6HzJxFrVaLyF72kMoCqXbF+y7Jvu7vm62cIm7EHUWkNo1VTVtRyQH5uHCU2UJ89a137
6ZxILUlVBSlXQIenRUcsgnLkYmuB5mvsM1FL9DzlWzd3pkBv6+wlzwhrisqlcLGdbeKq1sY5bAO3
y9xGq7HF7DSzhSI/JtRdeBct6Lsz1/BwhK4mHuVbkTQPnN6c05v6lpsotQctAe/zzmiuBIWcbwxI
2vaTD4d7Oac/ALgFgXKG2d8eXH6cuEP2tggYkFdsmW3t3yxNW2mPZL3mD17WzNvbEo/uglq1NiQA
E1PqwHCpKMlYhksxeVrAo0vnKqeLxqyZmMEy/gNkJzWvBiXjo3RC17RONYw3lV4L+0eQ9elSX7Hq
jy7ZPXH7/oU1F+qo/DFl5+iHuN4isHWryoSj11+IYcYcOCXxJw6HdR/cMTtF4iJf0evOti9ShcOK
EpiVPBqPnGm79LvpmLgPAlWGCw+y7M1EXUxuEnSP54Tfp/CyyJ7WfTeggFZKw9t6XlDk6Ox1MhzZ
mqsIjZ8RqaDgImVzDVVLoAbOGntjgfrEnTEjmCOjf/rr60UKvuj7m3ckeSOjZx38PJb72ufkI0kq
S/Ovu7P75Q8OPLdC+sQYnC+Y40Lg3NfUR+ogHWQVCruTLHh5AQl/2oFrOfobFvpoA3v0yFbJ9jrR
18wbt665D+WoXQta8+YSBSJXLGQyQqVfdDCYoq2JW7uAlb3Ytg8KiX83ZIsH7/eDhkRAmw4hgn5w
zzGSte0fcrRBvrJ9JxVOX5mXzSRg7lX9NpwAvCDHv/xUtpDWKuYTwJc23pSAIVIGzNhCTtJPkIIq
xzRUvc2ahMf4pBcYZixCLgtj5xOQw08tGtsyawfV+FPvF/sHpkMZCvqG1uhWJl3f4HYxgkYOGt0E
k2MbjerJi9OukwwooJp5sLg3qRPZMP5m11pyeeGjVh17v/V3Il5Ak1UjrRAOaMy1ihSY+/pN+/he
VWCWBSNQAU5Zj1U+6sAfO61D5XhVwN6a9RDtvuRN2bHYwLfT16wJGZMTmEj8zfrmwNHMXs21FGoR
LZSVT9STDp1IsYLBNWsHJUHDqxnRT1NfBYtGlnqW+nXfdV6+J8HLxlG8aIltRRI+z/1j0Jl2IXK/
wuu97PmOQHxVTZioSFJzEA9xfNN9uc7kKQQ/9V/+K4xp6cYRUZDM3vimAgAC5sMKLE7wRTLk+7Xt
KXng/L+ox5A2JFtvAxURiKOnQw6fCoMnbo//4CE7t2W8eY2gFt3knPh5SYqIZS9V+zdjJZIMU7N5
H4Va7vCimAMXLEblej/tdfVBpXFQRxHOmTHAiSXHtf7J4Oll2ujiun/AE4yuOnnDHpvfs6IhyhhT
hQtsTbwwjshKq1qEe45FvRRAjkbzqZS85Aj7Y5DEPkTD3sA5zfa7kiHO9VgVc2EHSi+uOygKvQey
dvzNVmBUyRC2JHemgXaoFDf1MdJhLtxMSfNEtt8WciJ8JYXxILySVu8WyNtM6jUs6y2XxxGpqbkS
KqVNJJTI97cUSS2r1sXM6D3PV8zjsUdikeFuMRnKg4uoCJ3VzS7Vc+alDZIPijRzf8Urre3Cqjza
IBUb8M+Bqb3rlmmHBg4A2g4f8VW5hlpQqxggxSExn16xjtWrq+knC56xesVQVvMODK4oygOviJcM
CygxS3oFMHMY/gurfHxRFUoD7n55G7dmhWiztasQWWqqCf4ANQcX8zRmEpAsYi6FKASFlnShj7Fu
2xTknm2WITnWwWXobqIyhy/G4Vi5UXxU4I/6R+lDzFDxMqqaIvKjzv5S0MfqdZjx23T1DBOeRiV9
10mP4WfBqUurXc88gN90YE12DdR3sjelRmJtx5pxZ2lFnA/nYVidW9F+anTXtQ7qZaCuq4IyJefL
NZ06rXO9VaTI8ZEu1drLGfWFSmZ6opcO8WmFfUw+zQfa0GmqVMaInuS+AfubpZIPNWufeZetJNRT
miorAT0pC0tocQe2RKRkAwCcTDSUGJ21rbS/tNXaZWCcfc4EFG0tzZQC8E3yUdCgaBzbI7Ncxyf0
IB0/iaZilts3wDtP7PcyLB2KtRJZzlxPM3JYvpIKlXEbjZhnT6RFYdScmIuizU7BsQ85FwCgJtNg
eoF/Hnhh8dGM9OzGwrZC1Iaff7hfAnHsaRlUmSp36QgQPr63asTuL5/16oVXtbtMHS5bes3ZuI1n
xBINjIZuGK6s6B/+9q2ynYkT1+XQKP0CxD9OFamb7GJq6uBGY7TiXjChTqLGGdHf6Yn3h2BnwOiT
hkzzaRO3LU+oxDl+MO5b43gaPLTZMdtbJ/PDdlC4n4nH/h61hDldHH5Cow6VCHlaiJVHDdiyqUcs
Zv0wg2e5ttt2sWqw3uJuuPBE+0uhtpJmoUdWKmNZvMU3hHCFoziN1WhJTtE58w+roa305QpVGeSw
8OBexiMn1U6wZ8YWnNLk1M4jDS5HD1JiYApPlZ+xvyGQ01uX+/NwL0clL8BFTdAtR2mK2pA7xfQD
55Q2O2BOdb22riok4H7z/AfvyowHU8UdlsSp0sMLilx/7JnKfZn2GLuzm7uhhOV9Q436OmpFk82c
82BjhKs9vjOtQKOw2vrQkIJY3u/07doG5CyZiE2wRz2wdbpeeyd4nwlglRBKy3DE9IHl8RxLUCuT
Zwn5Bfu6mHZbNb9yvuNaDYM1LvJKWwzYhNPjnt/IE4J23oh7VgYEm8F5C8jDJq9JrgoeCdyTvdw8
EhbE0dnLYbFctz699/LYghfbGgxFpnsUIn5in/7nlkNlQv6upG2VZN9rUApYXHJiwkZNxm3Fe/G2
vl0tmcFN8VSlb9PY3ogisBKvMHnaNPcWNQn+OHN+rBDvSuG9+HKeCzYhN+ltyC4J2LrFApTPk7Yx
qdkVGMFy/51Kbdb18S7YA5oATpZemmH1YGCg22J0s2Z8ejRFmCOm8wb7BHmuA1XSpXL2ETPlxmKV
U6ucfBMxWyHq8N3ONT7+VJGgO8+lRVJei1KkCyzsh+xAA3S2P5yd0EUCBf6qqR+bX1mPhsp4PBpe
CcvTxEnL2XeDL5JBvcIVJ1HT5YsqYLhs/RTWjN18kaIoEpKfYyUqNoqZ3nNgn1YxHAQ1L5V3JBg+
yUmtZjqpUMXA79AGGPnmq3qMl/CyXWCuZ3QzlodwS0JhmCbCXSUTzFhH0lmbdyQvUCcYJBxrFYKH
Hz3vpJLEyy05Piy+eVdkg4lEXnzgrqhHdfvCN2snHEvXZOvRUzUN1OBSa27noAq2hqfmNsqFWTp1
3n1FEWw7YwvoZtzN6ywlLhu8i13gGnqDWLe/Q3jP7V4i5/LTSr6HM180FD4uAv4gVVoMkGbK5wiM
/2xET97kk6Ro8Efp1gb1BPFLyYP1oXQ6ctd5NJS4JP42SYmpcQiXEmFd4XNyv4i/exG3gc56iGfA
NknNSCygGoX+1HKhOEZOK9GDXfrg2hvtZt6QrYoQLS659Q9Mc445SrnuisIIBzakGjqhRnoC61lZ
i/NfX479VjLOnvuuHTPrPJYQg9LQczt1TnAQ3Gi3xAWUWfyo5RjkaL0JhXdcv6EYay35/svg8en2
DahgZlXte6tmLwZ7+TOnlUld8KIh/t1W+NLksGG3ZJ+SsS2dh9kRoSYi6tK9Ar2j5BM9SesCn6H9
hFRfVvbSHJtFnB/y5z+Gu+4Y2Z8X3eTSc7WdaEdCxhgOYRo4n+7gOE/fr+gQhc/ftz9Z3Wfim+F6
jdSi7j8iZpUHr36/uEhYFUpPgIobM3sm6nHrsNIlgoceiDfOhYiJ5iC/mn8+Cq3EJidEkw3sKEKu
6ZlUrjlmDkwsY/noOlBYLwDm9Kcmq4yMapIRa1hu3QSegZwhr3pHzRual7u5eE9SV2OwrwNlK5Nm
haW+bftdE2Z1XfQHqJBwaKJg/zpDFOQmNCHuURJ4gthtmcA/chvT0nouuDzKc6MGcC6H9RbktPts
usJMkKuNYLNpWeO3i+2waR2pfTvtZYj91uK0M55tnKQoFLyJiR7g6sFrsGJLsLRfOBEK0ZYXiYfL
P7bB+aSm7H+mhBayN9fmXJDTXAyclxR50hSkWYSMuTonuNIYd9UqPDnanVWbjTFMG7DptQ5+ISS/
SMkMGxbEaPiOCkWq5jNY4BPU2tAxrE6EVqF1sfto5UU8UoJPmsRuM1cDxoa2QA9NvO6a2T2wh3hL
VEZjC+MtiU5uqH1mokG3r2rXvyWwjo+0DCIDXrMnAWD2aBQ0h9Spr0GiiWr8rDtZyaJghv+QUM30
uDQjWbEMX06Est6wv4hS8S1otPFKVM+5ptcJsljFYEPGVxARfz7Nmv+3MsqGc/rEYZ0+veQxqHQi
Myi6dhSyeltDb8xNCIyoH/Jxhp9ULAVhG5DMyHqIK3JlOCfiG6B+p3cR+MIfjC28EpuAZMh/hRnw
97i+7pDfPGn63WmvVb6Vb8kqb4M3Xb0sYZUINdA1e0XFawZpKvCxYHy+ckBliCz6h3GRBsBRIMyM
52aUxzAYuYSLA2YvwRV10d4bUnAWE/wyl1cofuJzrsp6DGAhmNM2bQDu6roGRdx6N99h99ZONXru
Oh3J7yaHVPj2XNh6vGu5VQqTtkM7aJUThMcBhGdDfb7qhMvRtmOrBIgDVZcIah9CGnBtwi7t5Txo
ITkvnwCW+NviQeUvx+nPCE1zU1geJ9A7RWKmboUniTGQ9Ulvo6edwcnTZmzHOvj+n3Q7Nb3C3Z6b
X1oZ/AE7HwsTer9R+tTOYeE3iAIb1/iCfIpJt1By7IuTAXLwXtkuI753lS9VJpGaDNDpPun+3PgI
YTIY6WttcB7PmYHYp7WmXQujTfJ2a+WcVUtM1M5ML6dK9NBI0j49YwXWALKlJFqxBqGGV65pIV8Y
Nrti/L9mYl1faB2UtUa9kLK7aQ+BzGxyCwWpHBDGaq1oXdl18f4UTnmVuCuTHG6BpvtwVwhnmuM+
HJv7gU8GBzN8oAUHbcFDeG4Y6VxZkg8keU5Pyu8KuDTZQ1a8UWH+J1Lai09QZ5Ba6KKhHDlJX/+E
LTMoV3XI6Hxc8uvmXUlIMwCgOJvMkPTb92tXXpJ7RJg16fQN7UYcIPmZwBjvLf+TX0T1DHrDSA5O
bswfxZiNxw3YRxJ9Xnc3QGpAzbbSWqleWzY9dkZgiH0MAnJCnFMkgCDNB93vYUDIaepTIwGnfw01
rrlW3dJolWivz0T9eFtxJTj+x4gllXFJBEkq3LL7Wx5FMerH6uj5VsNorDYlVB8m5aOC3UwDnjHq
JItS6EbLNalNQUkyyT7jlwvYPDhK9Bq2g0kbkf14+PjNw7XMsVHvHPjtUXwjsxD75+tlfVz8k60M
a22HFtus2rxarJ4uMLwPVH3pxRh7Vmyd+lEaxaGL/q73jDeuM2GyNRMQmoRWhbDKSfqz1TsuZcT6
8Vnsvg5Rm0WUJTPVLUPjhuN+wpjOg5TAYaaiYcGj0hqmTx2iXEyVoc4Q+g6dfhi1waBK4zrwXo0A
FkUEahZn2VAdPci/gGhYaBe64TAjGBR0jFvyj8DSVPpaKTpjHfUh30udvImKs0jiTQewSXSMFIdI
KW8RDHA0YuGZYFAju56Fg1xTr6FbFo48lGz4xE07trhTyxvNXSLe2z3XsWo9CN5gL1PMrzjvXQ7U
EnjaSKvcA+mLWIoa8RU3FEhtXV58VXenSAhZ9R4+AF4ZgC3Gw0JQMtLKy6CpYqmueDH3fNHg8vSL
sd39c33XJjdN7AaJwZlyc8lNAg==
`pragma protect end_protected
