// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
PWyBJKAd4MsgKEdPbVGHViYyylR5lMipQTemWa9NcBRXTOaUjl3GS01Vs7Fp36uYdBfsA1vfrEET
KH8/QwGo3uKIP4C7mwx8CR7S55AJ0epH5P6kFEjXp2bdZt1ChQkvHEmios93uXjgBCYqGPfziDXP
kafQoix/yMPjXFFbo5DCj8pBWtRMPwde3EZ9PjNsN9qYKysXJRhSE+Zc75USzsnY8vzZ1KcEi/g+
u1p61BTkEZrVyhVzLajvZWlOMP6wP9lotniUKNId6aeH7TGmx+RwKejnoafuOF9upCAewgbvr281
yOlg7d4E2HVZqpJWTSJIKpSsKqSx4gOs8B47KQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10640)
88vag8Uq65mLPheil6gKKzIbhdBK4lSw9mZTh/tp2WFLJWAW7EPUtRHP1ACPBR+qTA7zPWVD10ox
06DmgwA2L8MFYcYZPik+E4ROCbDZE666r64AsH8q28Lq0vfAar6vnkI9KVT5f5g0LdV6d9ncukNR
TNDjdRXu29jMF2MpmPwbVU9zRjWA7QVn+E+xQi3fVRSSVPI5R/ajL7rzD7ji4yaBe+3ceF72YXaR
1bY9uSuDCLbySusdyf1gFYUWnNGm8U0+QPSCTool43+BCw897uoLjPk85jMfayPJgvnUT86mj0uB
UAOwEViSNDzlbRnQgrO58Ncbj/zDZt3Gv6i0d4UO4O/kIzXJ5FMq1ZPaOK6fu/QhRIbjPElKJX8/
SDMqkERO7PdmKlYUpBTr+NesQYnk3Op/Lvf/AQ8l15JELjj/AJhqVLiP1sUCsmvYEGcWM5TeM2Lh
lkAL64LCH5ifvBN4w5og8olR6yt0uwVN4+sEiw2Y0dMj7/t1aDNqwFFtzsnuulzODF3TVFiCiWsL
px6S2ww/eOeOC9m6vcpA2S6elFPL3AzuZJ4qIhVjuDVvhzYEIJzGVMZQ+tYMjZEdWL++NO60fu94
lv0uXft8RzE7/nRPsDpmw/+idEje5vAp31JFTD+F4c5w01lOg2PpgDouOuHfSfIAwaaZo/i47YVO
VBBCQLPNmV95LtHifPZxCtnDWIoiAc9v9ZWsI8Zb+QgwTHEPg06qwgZeI1NTL14mjGetVIDqJ6re
CUvtrPAv9Z7lHgxaw88e1qz3anHMhnJn6Nu8+mdyS6s5AK/nMbz34wHTT683CQDqjleCA1BEj43+
X5iBRcoSAn9dmg9Ts/sLV40d7xUQbWYBdqVJA9xJV3Wn5H+6fg5sykqKmsmLIz7Q/MjbYBRrLptL
0IY7soFU9aGW42oOa20BpqAN+5JNHMMn8EwvsvszbejMAKzXqsuaUsMzUP3tZiPAttOUYdl3UnUw
ruBqBZaoT/aoU3G3rLcFgytSOgowXl5cPpO5lTRWuj//tl7GgdqDUc/tME7RM46IiZnunb/PzvXx
lbnfElVLEfQPqRuG8ruh0WfjSWwmBo1Fj+v9RB7GNUTnqBctZeMitAaHsIjg8GubrqSY5SitPwi6
Oa3+/K8qQEinZccncXkB/Skk0/O2xgSVm3LOfmRJ+5uBj/u/eYGuzehmo0X7YSR8SkZXabGOhtzP
+Qlzn/urxGmg5/FVA3PT7wnXsmhWCKSBSWnxJUCVcNdiNX95JmqXBuGC6BP++j1kcm6vLG4E59y6
jBuIX23UXHzJfBVlKIpms+VdY4ncnZzQ6IS1yFEgC5Ma/f3/BG3Be6XXvFF+N7fz5nPIjKjJZnkF
tKC+KFnutAGKKWD52GptUc9PBYXtJv9opnaEVlIO5jPsRhgEm9iKsXXel9TUXGJYn9bqucKMS5Ow
5an1UtPd/iKUKGlVWuv4xfc0iznUQq7eFHic4dpM133ju9aDgCatVxk4hGk7HlXNd//24vhncMSP
veyYuL1BwZkhkxHS9zZGMq+02lNyC0elmbK0Xk+3UXJeXInLAduWwYljO9B25eoMpyWWyz2fFXiL
8blkZtIExe3udLKFSONFfI50HcONZ8mT2BCFx6TSDl4uJ98Dmjmd8AZqgjz40DjWrlgYgLfuXlpx
X9mKNFTuIspeV/YcXdZkjy0FjDdGoqStxgwhGNZUUlsUtOclBa8BYbSaGU/R7XSAqvSFQU5E7syv
3X9XA7a4LQU6gKFtxS3oIJ02YBApvHXSjmJoffa6OpWBN5Jsq37BFiN4JmOfrK3hidbY2j7YLCsi
k+i11oih6kXQeIdUPk6/gjjNUEoPcgVSEATO/CGNDgSNe4rDTGL1CvxQeQ7FtPEjzg3UHJA/G9wX
hLVvnrX/sLKSKZ6Z4IYkap4HKzrWt5k43waCbf9OMCHMhgkMfGN/GEn4a29USyCkKQ1uN6SkBPWx
M/0mvRWlx6G69O56GanLqWibQEfa0nZVbBooNDtVPl24bCBNuZlm/96DLvsL1gaCxnzbFSoEDdXy
LHVsuDBAjKdHygbQMgaVr6A5PG9ua+GFJGUlfkKyDyvPr56z8N6rcAh3SnPhdwgMAzmMwRGl1k3n
8g74DBDbgE6J6kl97Wpf4mNekyOhbgpR4w+O1z6uRouNtRRsmW6yYtM0m2m7tl4mLdpNfFb43KU/
KBA3bn//pCzCYVqX9upiddlVBcrEFRL+YcoGa7LxjPrNvdbdqKV02XCQecB29q8m6Gn9Bu1IkfKY
gzbTvomq8BElCZI0yZgnFT1arWRCDZoTOJIC/0qqibWPUfHF/c81smWZ+kL2BiixyY5UsGT6Dwe9
U2+orzr3QEV0wQOuz09d5D8bfxiQtup4RObcr3Q4wnK3ZNdybx0DU813Wkyt/UBAvAAWusvdby85
qk5xve+dhyAB7Q5uPa45Qn6sKUKDj6ZwN96Sj9XMtm3ckZDzwerZacR459AsdK+72YLfSgyBirNK
4WKqFgrFs96VmXNNdqwQ4YoB9w/65v5ixhM5F5bt1PCgAwfEbQS8K+30b05Tr1OMt7gsG3mAFoqj
tRrGcvQAg6EkUuiigK1ArRcJDbGS2iwIlagfYuw3jRyV9jyWCnlQg9G8EJ/SePwN+dQtKWeApAc4
OAFivXtt8IP4pmWPMzaKGIIIrB8tiYVvfncCEyHje9LVcu4jaQNM8+2Y8/5NOUiufnfQ41XKzsHH
2XuDoQNGdJBgkPEAvC0+ixPc1zRYnUZ7oUcR4qIVkWziUUDf5Dn3PAlRIy4Em0lEiMOL1J83dwzi
9qBDzNSJLMmc0eCDTcVeiYHnob7Xj7fThT3abp8pED8WcFmWwrBl54ihMJgyrd9TjCFYGWll0NI6
GMsPii+xt9c9VaefAgyUWyta5cGS3HitZzcweapzUU5vm/wUdI6v6Tw/nMuKfpDb/fOdBRo0JTcJ
KYOIU1xnUrpPiP1Ua+XtV0MZ5UaKqkVHE5JVels9TVkcmW7UgfbCJ0xrdxfZb+uRTdaFV1dZffAm
iELCr14wR4GESyWwnMhrMPjDsEYtYc+XrdavgwnjYfHuFzi8/Aqcv9V9eN4I3d8LaBBmJGlpf64T
YQ83L+DbU2OZt/CzS3LlbPbeX6LGj7rDP9UMf+XZqTYtuChVKO34xAneGb8VquX+Z14cTyTpzCOn
wVgSBNIUxCn5WvCOYDdM9OXX0qscb/bE9G0aDIafj16UxZhEPpW2CWwh9P/IfxqvIue04M2E3KJP
1o5IqzgoWyr8Y1wVenjJdlshhY748fYpaB9rDWOnzDGPvA9+Ppkb5Mwsj9KiAKJhznubS4+zlOBW
EKxLNPCP+fsJetFdQusF1o0SgOSEhk3Q/y1oDEUx/VWtmt0HFRKf/Vl83nHveOuZcq+6/Lph5dm+
DkUTeqVYh1zRUkJHsP79pvpm+xvZ+pP0k69vmDmQGM3+Bjv/giHSPM1srj+2XBUDiZyWbBbKQYY4
slaqp8pzW6ZpDg6TbfYgnaMDlU/HozRQRYdURWaItoLY/OJva8ltyP+vKEwcaTsIn04bx2d6fXJg
xhxYsFF6v0ceFrJ9havyMxwfs8NegYSNydxhZWnIXzky/xu7mz2pqERdw9kn3XfxKcPajiVjx750
aoVcfML9yD/cJpwqs5dLpYMoPtgIXNqgZd9l1YAhqzGlwRY147398N42hQh3lAO5duL+6LDhq2Km
+8U3+YBkc9gXor0RAWDDflA2TVQLwTMffvzu6YiobOFJYIk1btZwSLOX566c+KsxiGc0BQqMWNJG
d7nJR825wSOGLMoQTmC2K4ehSKcOYyESGNkVow/HFlpK4PAm22A6gHMZIC3nqHv93Wp23M7S5J3o
j/ghxG8F+iKKZ5mIyMeYl/NtlHrC+u9+Xp3oghJVHWNhTH7c5dyikDk8MTV07yJmo5of4oMw5quc
f2dwBYzHOFseAsoW03q0QXncV/K5uRSGzt2S0nnKiGi+Q13sDrLHRHzEvq4nRJU0qD0R9A8tIn9v
yBXi6L9lzLPSfdSGEQXdIAAmkpglRPNAKtqDGsk3O4Gw3phGn3Q5JUdTK5PT1fzPiLTXZOlAK0BF
7VDiwzra/oxkJQmeXxLgOMscNmxjFnjruqUWkwdWYPD4+r9+tPSgBjSOoUu8rTqwx9sgOIQVq/Do
jRD3MGwuf5yQo5fGjKWu8jBrlH1vwutaNI+NkwtycPJFMf2dA021L7n+g9W5xfWLpjws2AF7Qf40
EcsVCH/eccdcfCpGRhHsqlQLTrwONju2Eo5tmSpWyucTl4MTvT/Dx6BkKyoRGsMu4DWn4XOalKlK
EF4Y3aOk54qrSOSyB1QTWrHBS7YMvuVDyibNapxd6b3WchBYb59QY3Kk9QZFUhKQ90zTMh4jwFvD
/qRcUwgjc6EfHpzfkKKEoPk6uxdxwvxH/LTRHk05t2mAseXQfxhRJJ25UZkVb8IXV7yplBN8SDiZ
1iuG4YVpQQj4Nqms5RmQMWw03/0DU0+QJFP4YfeHcBygNLB5Ujpcn6tkaJOhfoXgWg9LyzYvtPcI
EyQPP5Pjy8bKpIjaTTRyMenBfWLukMQDbCzJdvMsmpnf74HOsx7TPZy5xBazQ3WlkEE22ZlTzlFt
lzs+1A6s6T9MQfCmk9xHhHlHA+sPGrroTQEXRKO0S4RSqvqsjvSPCETH/s+lYl29uljnSB2iq2Bh
K1UatZW51DTkuFUV4WtMQbHHAiMlkWn7QaqGhDC7rh3vu3R6AUocASlZH51I5D2DGnWTKQc9d4jN
CzaTbi+ipnKgdQkn0TrXcPnVeR7sO0RSmWeldfi0EPaNVq/UVkoDNTRpqgvmnfc91Ou1SgFe0ccx
YVYwS0ktOPBL4ZkbAPHKvHPdIKQ8hsI3733T9A5Jq52iLP9WdsI0rINVnom+dMq+y5HUNDbaYzJz
UVIVUeJoBbN0h7xj/jQ7IEQoWhJNAahI8VXTR0O6+1n+R+AUO1GZ9wcgAK+Kf+nJtWLreCbNZhMl
gwJb95DnCyQMLuZpXC3e3jkq/kGfRX/agVzq4NpEQCfjsoz7aekIVJrf+trC7g+tV2YV40TNaUx8
pupBNvrdecXS343UzLFKqz7TpKrvW0uPyhvwqjwehsM8ImJs6w5oErqqw9Qc3Zd16HAPmR89ps2H
Hjmwiv4Huqht0eGoKwIgEaqNQrY2Jn7BOWFvWLc+A/jAWKTfkY/QFGq76HjmBoNZGVn3xf6OBOKo
g5pGdikCxRraVh3gwLb25uKy8Y7GtPh6BVpnGC8Sv+TEN9roldkpMfXBz2qojwYjAq808LPLdTUk
Kglh0eQT9iVVXDqcPOk5aEaes5VvWpFEwRmtcu1Y+mZ2UUF2UhMIjndvBu+bfEHJ/y/TetDzU1fG
bvYy/UYKxMGMSM+DaXTebnbsnHucKcSv77bQFd7aZW1Q8Z4vMACGboFbRoPZkJIBivJGs+DNG+25
/9PjyA1cKo+IDQL+KSLo+ql0NR5Or5AmBRC1A9NE+M72TGvdSxZPQz+hH00HyXVSQ2gkHpVaC6OD
UJTvUx/UzugDVkwUZUoKI8qGof9srqXTS2UvmdWPScR3TUa1kiZp8GzDdFHbLyLOwSDu+7Kcv0q0
SP3T6e3Zk505vwJcRQfFHHxbnoBYOvwPNDCb2LA0EhBdTNpp6qe5Fy/djwiWbO5gIvBp8K/8BlOD
7uUS6//D6CkVkn/VD6bEDdEkJb5Hkr0FKUUVMg24YIAPSMR8SyOXAfzMTw4nk8J2ZAG+c7g3TZzh
GnZAbEyBwgup6k3uZKRNPXJagFUlClKh4vqx27vkW6btSwFmul7vEXj5shWofkpp8rcLCMgMMx6C
V9mzWHqP62foFHHLEemKMifHH/a3kRBZ5cJSg3ZiRbMNpTnuZc8VF85LTJex3+QjM2zMAHojOck+
zQ0CNTiP3QnkZ0jspLqwHRSvuYGoO3fyleo4x0o15u2Eo3N+qhxQZpaPhvQKzr9403DUFc3kps1O
pUuMzHiNieVP4n7ITuydGWz35z2IuYhvQ22zGFH40Dlzty5LmYk0Qs+fmUOzm4T/LHJj+3gc+HiM
rQoJshOVnG1DZ+z2x/dAS8tpcf89MY4iOL3IjGhTRVp5jZE6AstemSMukKtvIAcaT6eSisIwDEOy
DAg4U/45rg2b8KCqHImNrCo62Y6hcZc8vQa/6BRB/iCKqdIMdjdVkRTFtATWEFFFu2e45chYNz9f
fT3ndjHQIXHoc6gXmcYawihw5H7bSwpXFg9AlMS/vh/p1evCy+s/rrJYLNbuqUmyZ/N5It9MHqpV
oN5h8paJAv/qhLvqnJCaaKNGNTJa1juIi0OJlpOAdH/PwJ04x38Vkf/3Q9Glft4P7DvB0YqgiP7k
sJhCz/vZfUggQhsO7sarpwRR8FXCqDfLheuV29XExZGGX+gG2DLmXr4Pbz9C+Gh5YCjUiKkApq/j
hg2n0fNvhN/l+L0DQK83dFVUYRZpJyrV+d32yaubIA8fppxXJps+/bzI0L4WTZ33L1nuLB0p75au
bFN8yJ+YEMVlX6ymRlZAQaWpJekHo9DL+2gEvGpzEWPlaAIZdODrl8JGfg7ak17wLzbaIXnvi2hx
2r/a7teSOsQwxRZyYn2RZRvSpgvZ3lkaQOcVmvYLhPLQ4iTuom0GvYCIL9hos49TprE3VCwgG2ky
NWNivdp5QoVJPRtUQm2jR9BCllMMF6cCMK2HU5aE4vJWWHW5nLgBMCf6WDKevFpxFuvFuTiHVK4E
ZBMmVIr1r67nCNepe4yp+EFKAUQbMMoDqk0xc+nYiyPxRGzMRimAdBognzyrtVfCcRv5CXkDMsFm
QcFcpxp/bAfFh8PmZKbMn2Hnc1zAK95aMb3gE1Af8B11og1zevjBY4r1qkstw8DWtldUq8MIZgck
O7fHJG81I0WYjCT620bC2UTsVfH7/isbRTV1fKLgiYt3p6o+54+D+7nJnnVkXdfZbE0YXvCKk4k+
AghbEE6sXGySa9Otj0V44efROicmPxwTPU97q1T/nNgvZjuxO6KuSkA5iebx1S4Mwp4WkzZwWErO
v9m6XaSjNiU9WrTOrlDUNDMub2JVP941dDPeYWEJhV/8j5i3MeKHjb26plzvWqXFtZxDFxg/Nd8W
t9YNwkabHCJhRcqYqEbtX+GYcMc8oqVxgZaFSAvcl/c3EtYB7katV4Osrbx1vXlY/PiMo9tzfhde
jV++Gezs44wdr2TQBOzCHPUc2joFP6pQwvW8MxwkB/8xpE8B/+ZulDLh7aXxXv3kgTlfgIkz9pI9
IBSKTQ+WiIHHjeY1a17PaekGQaQLGwsFXp2quaECiTykkzum6ZMpVTAuz5rgxHKoN4Kx2Bk+0i63
+jSAr8MrmLjORaLQqGTKlh4+9jDPH/0BtOAXuXvVUxpuKSq3tfjWnR/ELcr/AjweGYLdbNTd94aX
aDgndTI+lASFDGkU5nrRmsbuxTyU+r2ebji1n0BCiP9ai9DMDOvLpg1d4LGVBxlC3h8XoYmSPztB
1Hh/ziuQ+epo53hD9XcBKXdPq/xMQLJi2J6clQquJnMiCJ2RqSqp/gd6QCSXCMbOCbvLXMxsYGEe
rLKe7m6cYRSl85SLDIp6ZehZ09Ken7RtEl0sDX3SK64QyYXdil4c8uKlZKhL9bs1QusktU5Uwku+
77TsaSH9dW9D2Qmzu5XTYXL3QBGsjjFHC+h30GGaRUAln/hmJRhWSlT+0BFX2KB8rhW+hNOiDxjH
WjXYUKyUg8oEkDDQkznzeSOgp9ofXIxP3U0HRySe9lm42v43SoZw4UcLxlLwb7m0Y/ggX1CwSkiQ
XvLfbIyGjkclWe8f6KDtVMENJXz5kGqGTQAIxArMKJ/LpOoG9zGitF5c6UCLM6ipLLuDmyGqgu3l
zFe8EHnqcUhrcXwWlpHWxUk5sFs9s1gyAnAGUuCP3MYB5BPLntdM/mhJMl3AOGR0oPGQzcjzq4wr
cFeU67e9IMTzQO0rehah/oq2QNgiVZOmD6z5cYmo0rejB2xkCEwhuegKybapA6zTyfn1TyLjQAnw
wd38uZ9SssKRi77CaQ6/xd1LuI/yX09b2KIpZwKxe6R8eisAchxUw687tgWZIMvycAWg46puH+bo
cVD1j38YyHaL3cRuCZymt0iDlNQ2XcMkxuft+lavMSRTtBottXSBl1cNxAu5BFN63HnAmyCmIhDH
scB19dWCxkatjmPe+rPcPNkJY3FocU+9hyJIVyFQP55YctfM2WjIsWAOcskuo5Uu1O982g1rTCIS
g8g+cbZPny+CwIDLlMRCMjqKo4n3FSoIW9mIdiUcmKZSx+1CzZlPucOIJgMQbMOceFVDrPYOQbO4
tsab3r9xC8aVzWCPr72o7HyysK26ekTcp+jU5dDXXTqj5qMqF9g7DULPYO1XH+jQKzmd4oDw+7vV
UZ58r49CVsQ1AlPTD3P1w3O5idCUf5ajdXDr8/qk2OVo24NIeqOTY7o59k3ORIZ3uIvmHYHpUxMK
tASlVz0XnIHW4wzSRpIbh/6QncpOkCzpZSdNBudNH/Uc529EZ7a8+4ZmtQqx+S4CfzXHxoMqe+z/
krdGiVwx/wcls73D+HEDXUMf3heGMA0uNWOUHk9KHLDQRg4dPTzzpRLetoT3m1swzJa4/TirK6Sa
Ca21eWzjyWm6ESntFveSZJqSXDeWFds0n54zceqF+sHpUiXZPd79I6wHcZjYROXvEP3gFT/Trcsi
0ey0Y/MM4aQH0Zml9j32So0tD4IzUQc1sycb3eN8tjHHaO7dG1De3X/ugR6WqYvtQ6obuNh+TMrn
r/USqKxS78KF/ef6dtqbgU4QDfBHQJ04VtgMKQH7nSy8iI01K5lpn6YcjPs6heZFrsNLFvP/x2ze
0DZzoWiBN/bG1spNbiDH7XWtL4qbOtSdvnVgeZ+9Jz2bz1/f3c07E/diOyGykpNBGywTfJjbSZTA
o9ssqLfWz1WqCyt8POY6vSkbtdviLTHYj+9qiBg6QgthZz38MKwnMgjlxxZGfMyyR7Bdq/MYGuYt
8IdYSJPJIYxqKVF9KB+11qeeZmAXWJ4rnKZRGqffNf//FKVtv1KYV50vvs/HI4TxPrIOKLGu/443
aCuOh7x31239NjQVCKMUiNWwlYsYUH7l4rg+HD8kDmqJ936ZoyV0WJ8W/ev7izJavg8sR6JdR/Ry
pDOAWlLWJWY3bNUP3tQaqC+M89FWssUTafkCe76me3bXemwaZK5jrMySncGkkR2UxX56NKz22kCx
tYMPkSYHAQlJXfF3OXm8yG2S7Zifz5INJiTuFQPSFseNDJCNWnRq5+0cewo5e4EZ1bmOjuu0M21p
t3ii5KYpmVR4+Fma2I2wf8Z2zN08eiJc2AaV/oAb5huMQbq4S54dKRtTs+L4gm9hPudoxGHz+4YC
pcNoYx7XLxkMWY/fN6pWxllzRVkmpafqiDdxJPFItS7CP38qlpjiHHKjecBgGMtP5sUxwjrXinUO
1hVVZJGd+OmwUH7jOjsUninh01PMf8k4bR8DR1KYXrWbUmNyZz0r2nmlQjnPGORKRqsPCffDZ16P
xM5+atQnxMCJ5s5f76hparB7VHllkqiIkqpteOWbsSIV/M0V2VvoA8H0+SdqFah7IReBDBHCPTlb
JYkTJJzvTxnpH2F8exj1D/6Y1O9BHY//dOGQ2NWvrhIcKvvXRqt+wek30RJAkMgXE/CewpVbF3rH
xGl3lXhuJ7z0L5wUNKNs3lFk/+vo59HK+fgPzrZsAQMdFMr9KUze1SBJtWzmFYwdB65CeNE3YNFb
4AUuNtOTua96CPtfWjDQiHwx4iDjFBy+3VCDCRPDWQKKfqCzmKl39TDkUpw4dDxRtKBDQ/M+gM/6
M7rUKYDiOvf082uik7MYICA+3JSy5/NZ00f9HMDmfarDtDffSse0etCDE3HF/hmiBDDH9E3z6hsO
PC7mx0LzT1+NMkhkqf0bUU1VqBDLPTN6NOj4tcDI80LsSGE175xNG73PydL0HXcxj6/OI8a1tLzr
2pMWn8/IuJMBXFZa0hEICnNhlSgvHdk5zGStRTO7g/waottw+rbIA26OPFOtWh8PVUeULWYnPyPN
78OXNZ+ybmxNyHTQAhPSzF5Z8lLhv/36+7YYVSiDls2gFTwmWj2bvlJJV8lNEoReNK1Fr4hXfOIV
p3seUtb7+LiUYvP6dhq3tOk1wRsSDJW/A6yMRzwXR4s57Ld5ScKc8wP1o1tGLeVOf/C872O3N5PO
7HT9YWKdNUX8TRYjTz2wUQtIz4Is8tMLpIxC+eFnttDhErniiGk7jOnHzUt9sg2D6lD4JbtCXh5d
jn8pf3aYBtOqDwkT+tIMsL9ODD8/6fAjcComB54o0DCmtdoELoByY23cwQ3gjJCYF9l3tBGl2RZd
JcPVF9U7dONVvxtqOyT2fdBGQwte1UYrXpxuM3zF4W0yYra4cJZGIQtXkUS903QkGfGQWanVHuQb
jqE5ecMVxJtWsM8cydTEVCuYf7ESKa2/doO+QCGwQrKHUolEQrxg4cAOz1cX3tbn+6OmC985vQIY
UUtqRJuDNp6InuguaubjmMCqo0qstQ0gen9aZ9X2YFZnKXOs8fLFLxfa8EepRLSwugZOZ9DDZ0fi
aGqs431SJID2C8umCM8Bt2gMdWEOjkgn0AeiyYyEIzXiylRLML16un2bLcKJlR9PccfzSijYaCKB
NbmhVbL9ds2IPE7VtK7K+7NrqUc2z4KzhY/iipXgOZ566C/MEdNUWcEt7/FHxK0v/Xuh96r5E1T3
VbynefzRqBvrPAz7QXYBTRZThGo9yzhu6dz4ykMMCQQmgvzy8VpscuiBp8/uPOxJu2LI9m9qC+KW
RqF2Zjk/vXD8USycxOjbVxndwX9g23Pq8kxOQC0YkWZabBqhL/5eKT+hSIY30KMb5J/Jnb0aarOk
dCsS9EJjZnsodNtSvn+wgWGgQdb/NnjxBAtm9KB1TEflF+DX/Z+N8ANW96pZP/O2sn6M+PveHYRN
LJnycrKGMd9N41juyne6w5sz97RGjskg4UdqGGKba4Slz5F26DragJOUOZKCpiCLr1d38Cv9ZQyY
5P49Q5BcJbogLaUDyp03gBN7s2DXmmAE/gV6wcrU0Ux9jAYNLJX/MNClu2G7eg/lNtyWEjRDvwep
xUIV4pIDH/JDi2u5m4ljbqE+x6PyZJOyz158DEEIjZvy5SZUH5tqFGgHUAoRuwSbXptRwXfCXVUC
H/9x42HR4DQJaOtKhPKLUaJ9MnZA5Yb/7OQRU49k7EiYokclihWEnlZS6xX0va+9D272ZnVkTdBY
tB4QqyH3+Zry5IzGl3n5fnuINOHobQdltW8Qu2onfRCI9KlGn2yY+ewwDpSvzodCruGAfLczug4/
0yLAvitssRiJ/ZgfyBOgj64qmxBboYRaI3Bu5agD5B4MDfD+Di8Ern+inZR664KD/OsbVX84l6c1
DE+h7meZpCTzE8OWfgRqt1rKFGcgEMpBuZpNzG6MQA5k60P0yd5zs0FNCUCpREMhGJntlGKnogqs
3D6cKXol7YSQWnBw7zJi7zF514wLeTxOUJwALRfX9nulP5FwsQZPJkS8pMMGzgefopqWRWq9I7eW
BYDiW/Z635BUUHRz3TaQDqbCqCvqWk1jHG3z53UfBOw2miepag2A2GZL81gehHwYxXN6v5Su16TJ
3QLCLjObWaSzbzLFrsd8XS0RWoBJmtNDQgJsyeRzFeH+ybxNePgLJt3ZFCBZFWTCEwwMFNJaTAbp
36w774EPYac5Q1G7aTSUNNGO7TxpKmp4tTq11+aiZZBSgBq/6zo1OhyKyFM5Wt/0+NyTXfL5OHnv
xm/AvG5BoExNd2gvCcQTArDCX6ZNaod0jtQMtfvqwfXDCFNsR3sNIyNVOTirk+qWn7+O236pBMlR
5igdRj2bSFDmD5UY4u/BJjc0sV/HzNorwewbd/zSUyUFWBI1quDDLPKq5IqKxDZuBQomwoKqmzDe
z0oM+yVpMKt1gK/tJi60MESeuPCDwHPpaMNO0bVkpRr6p3j8PmKsBSc/LUP2K2xO4lrNztJiU/pz
gN52PVKxxN5VDq8jo9W4Akjmj7DfoWDSekk9LBx2JvJK5COxpmQhUipqvOGIJu9gf2gMpxnepCex
4wIXxcAdTiBHqHyemDqPfuHyZYbVTEz3CgyCp78l1DBB4iroIc9ANPrkCRkAiCENHtxr/4GmYk7v
+1O0evR9W4Jwdi6FT9QQDzQ0evnPX6+5Z3RPrwU+/OBY0o9+AABS/90WXllxPkgTWFdjnBphrpK1
bJk0h5OoX5MaxkDSP35NZoRDDchH+6kI34HGly+U7flXXrr536JcdFnmvUNwdMIk3sZQu1izQdbp
4xRdx6W6mF82YROFZfjDi6gVem8pDC+EepN7mIN/dHgF5IFVQdbaGjLJVSpBHzYUUwUXP51FBusT
5tjwUK+t97Pb7TUkUehPTD2Simy9I1+M7hy1fkcQLsQXVzUajhGJXHanpBKy/Arq64ZjzWp6ytfr
+KljeMjwQOlruOIpb4LYeMI0KYUU3Kt0AXgyfqiuT3VS0otTXLdcLZyvfV+tj2pnwtL9iv3ZbLkY
PBvPwXhGcG1QoNpZf0tV77of9LA2H6Fi3/ar51KTJZjXiKEp6r4nAER0Bqtginu3axW501RlGEAh
GsYP/e6GdstsyftHm9wQHAMhlecaXzkmYoyGg5McSIQQ6CrdqkCZwRQQLWo/wEZMy8DudeLoGDvO
HSByK+KzAAZMJk8i2y4h1TO87LguscJ38QLa0A7JH6dFUhaCb7m4+q6R9fBpqyWttAyp6+ci+Thn
Dz7+91oLhUyYGsYp+272ry16VWKRd06CSLRrSz8PqpQ4grYuLyiVrFWZY4dwvsFtfDCya821fAaO
WPmmuAn5Btv5cq+MmZC5ui1VwvzVlgc8+vRv2u9c819ycyuTc+dON8cVRiXFoLrWKxEi28u0WDQI
oKiktBIVPa2OReTKMwE4ZMgJmhNSZfwgC2Xi2wzWlsmPoX15uHIFmDOAU7qQ3JeQjg0jVJbtYpWF
K0yth0xX9pPwbhHu0zctmYzRVfQSLbPnPeypBdqRR7j+YzparGLJoLhru/2GVzrsxjatENonFhbO
lG0jKoHlpOJGdHJzVRNue3XmhlsiwChOLbEcSZOYbn2R8kV8yWox9N/1l1/qu5/tdaDdz/+vkuzV
0fIGjbthBAQHpszEaRXGREk2Mfo//MuBAT9UQU1IeCK1JwMM/hsjY359gtDbXvAmMhPvzRTC5CUC
re13Rz3PWG+syzBKWq/boNJd4Rrm7YpRxoHHH+TcaxyBNCB3bPdieo3ykHu8T4+277MlKhjRYp1D
Le3bhAMcLXLh3akgKX/xk3QQJsFTr/bwSGP+iYzoOJzcrz1kHBvQKVxKSNYhUeMg/30Lgr0q9eRy
RmWXIf69eI73+FPicDVyRxDeit5gX8e41VRep85I6wA9RToD/wTFxVyClUC9LzPIdpClIw6ttCLR
UNu5XmoSMkIwwKQSAHZeFGKzF9iww5NbOJ8g6iH+N4IoXcABNYsr0wVA4eMb3vilbuipndDswylK
TLR5SDfHxCqjxIQMi/09M7KAGqNp6OFuEdEv+Q4Sn3hXTVEzdJ34mroCCRsUgzpOqoB/qxv5zx1B
XdoRDU7Dn5+ZGZHbvNh8sfTGhnAZACeayrVVLu9yV+V/lbGgHN+MGNf1VdpgyPWTQQ/KmDSJqSmi
lw8VSp+jlowLPHpGQxIcci9gA7MM4YSihcPuJrRhDnQc69ETHO7GklAMS0veH8d04BOjrMCEpifG
BQggsuJQCFoef1EbUr0g2ZGydRbv1vb0wPOawIg0RdpXTjuR9P09fB6NRtMNMu9mAjhI+bvkMqXo
JZPGlrL9oYY1cG3A5hyXRC7EpZvJ7IYmVnbKIyweg5jduRzvfldB39ySLObwFiHxoEFXZRBOFAi3
KyMLhpFM8elUPp5pKMq8B72Y0MjtVVvC7SHHW9DiV5VTrJUceXYwvHfvECanmbDInWxKE4F0BhRA
pOf4tE4/WD5VkTOCrSXM3C3EuZvyzYK3xxfyUQq/PGL50005+Di35CFb0p1093VO7yaFzPLmGITA
hG7nlGqMEgK0V+KC3DupVNBCCmqrAipw0B2/ah2FxZh/+aFdjTM=
`pragma protect end_protected
