// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
RS5MMNCi9BZiVeTBH2AL3cGY9sLCFbGxL3lt3LRLNUr6KioFD9m2Ok/J7WMKI775lTrLGtyFCDSm
XqdFvdQN0Y4AOUjRjc99QOFT3p5+2LiI+3go4m3awQR7eIv+jZEI1BOkfOtcBowfLkfwLDCchash
ZH8CVPZBOmQuwaw/NaCaeqXS64lghRciaqJWbNo7DPznMl7/gE1VImDrD5UmrI+eJ1AzoilYrtmR
a4RizK+Gh+Z1y2cp2TvepWJ128KvMj2s77loto0IUNENBWNfZ84UNqogHBXiBhZovEg1jkgfWS2V
U/BLGAeSVaN7sweESPNxM7QqxoLmlIY2JOAHPw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 31536)
93v8Gdfa4Q9m7WdQoPmeW7kWt0SdjfaVldW72Qdyhi0x0W8thcjrrCQIVCxLgLeO9uTjTmwUELme
e6kfSxmuNDCSpv7Xzib42iy0ieBhGNkwGChxJfXF+5He+0fh+0SXSXY0/yvfJya8gwaqV5Sp9Rk8
kr5Ee9/P9SzsZUzt+gJqn4K809B37+JMQDxiXLyxw6Dj1OQAF1dgkF717vovOATpIAg5lnsMsKbw
Ce+MaaG7HzDmo0nQ+KmzBOGHRLXBT3b4GAkI4Gf+S2Okw9oiBwMqhgLeLabnQ5zH/DpTdTiY2QTH
Dq149fgea+KqyBLRVsOQ/c1amjg5DCP+I2cm/L2aqHff4WHS9GZw3c4EYOODzSyyJVjxHpjnmmL9
CusDSQlXGtwvniQBB634XpB/Nd0sKbSEW5KiktET8YdM4wh4lwTijCHWtWc5jSsEg/2tKdTqgLp6
kRaC5LFkNKpeysFie/yi8uzvP8Udat5ByvqkVISQU+0Ck+EdxnJecihd3ZLLrFRmYzx6rTa3MSiK
MMlBK1qpzoU/0l+MVC21nQgBDlI1V63PkTLoSWQ8kFtyeoSPHo9n0N3VaUrtDxGt45yHnms06cJu
wOoTqiqYMWzvlUsqfqgjMcC55W1lwAyXBL8v7g3LFWF50OAOFBRWcvGXcbv0NwTa84IebXuzof4v
gEFtsg2gEF72IAdcG/CCNLY1Bz7C0xYfgDS7AAWGFq479rMUYwPgBKKm2hnv5/YNGX9ivkTieU7a
kxIbUtRm4vTWh+A+/q+z+e0yR5TVKJWZUogzBwzPklWI6/I6tARaPYh+PeTuCyfZaI1aFtmmgmXG
3T/IBKwHKLs0S61ukipHmoFSWiOGppivNz5SnfKvqi40f54+2bV5hMRHAB2/D5CJHu0tbMK6TjyC
epvD60hXnIcCVDwBrDV0bqjbYgWYj3DdfBNdL5VKnmMVoR5Vd2mOD+XtolClBb0g2aLfQc+bKjiL
229avzKy0XGXgay6C61PiZntjqSl7IjwZ8HnkcE9/9K6FbQBcf4GKX+rJ/MenyrkXNK66KnEqDrV
AU9qlP3caR5lJSIHDDb9/fXk0VqUkKkBf8EfbAcs1PWMLQPUtWChrOJCUfv1lE3EOByajTOOTOSU
7Z7bWPd+cyqHXHrOQ7sgEgFF0DNACrDdOyzLGPWkRh/vQuR9yLJLIzTf+LK0fJcu1N+xYZSaao/d
l7ewHmRbnn0jOSqR6qBifLMBLXk91gBPwcf3i1l01CQt9rhV8L+MasctWM4b4EvKVbnSVRUB2QzF
p+ko/Sa04Xk0u5UQuyZKrIpo/iR31jJU6LVe7w1HOj2gUzcA27wb0CaHYX75Wf4dcD3PArX/ehsq
cEWCMeUTgF0QdDsI1XpE6tmQd291090Rd1Uym26W3L/tQ8KbGTGPsb77VerCFZhzmDr1wGQpk8QB
omNIGlI52alL81BanjROe4WDNLOZ2ja+Utid4//Bx4s2LjGn3cYcZNevnLPpjHqLpZr0jfBsyGIW
ZG1Rv6caaAqY/5ewMOrvL7oUMRBffpLNBl86UurKQkavCN74SrNzPSuQcxK9XnCHPEbqGdkbyppv
Lwxedy2+MXFYEyF/RaYw/RuxW5gM7MFg+NlZ+K8tkps16pY/ziAp9rGST8/1LVEG3fvI7P9MbTGg
ZN23O4IK9nacDByK8qcQnsjs7BOLWrYhqyKAp2K6o4mVVY5t3X4NC2G18Ss6eKA+XjsNW42FNfsz
MtfBD0tbLowx00zAsMiV7WNjTpZnCLfkgKgXoZPyuzhrGWIklZrrmtsN7tCh6632eC9HOLa/ilpR
v8k50ye4ekYhLUm6AaCJxgO3WypLiNwRVUup8FOaAzQQQaFllPaZP6KH85nXfqnxzgxzAvPY0vO0
iHaTUhXAktDDYvFy8xlrLf2Fwy3+fr9AVjxzvvDG2Z0exXFRHhVvxoIFCU1ezElLCDCjy1tK2I3O
ct45arCc7SfDXFAdNOeq2ne0Pc7ibZgChgdY3b9lc52zbJ4+9XzYwQKSGmsKB68o+1A0WuFXTH4b
CnVKVX7VhMTALLMuzlliVFs0Ol+XbMo2u2qxLI7KR/zcZKO4tpAG4tK4547y5XDrk7v0AKTnPsk8
V7DxQpXNWCS5tgc1/tEiqg//x/Rk253PlSw9f9CuJZdz/CynoOXcQjsdVFBBkS+Q/I0Kq7IDz4hh
OVHEd6fHB8kSN3FH5Twgr+Ho4nZTWIeQEOW21r6UWbZkS/8cqKtytAscD2uwwIBfvfPgA/RoCKOx
K7YndheV9ox5SKEgZ2Ht7qh7675L1gTeSe8YkyMR0nRNfzNqJOkbb9yaa4BhblGI6kNctYuXEgEG
TBVEXqKs7Y9WTqjaSsIWuc3gBMm8PYvRLpRWXcz5AKG8CtUlgesT7X94hGbZsSOLLmO3CnbU36z0
XRpjJ0PuN6o1W0DX+1BeSDTCByw5+a8DuTWNpWo08nmY+L6YPJshDa7A7I6JzLg0TMa+hinLLKvZ
rcUjWVaB8S2p9Q7G6/Udkrdcr9DS/S1V943MDK8P9H9aXmo8vokno5gpVU6NAzeoHAXnmIA9awpU
VKa12p4sinrhSzwJSZg+Vk7MBETvqQDWgI79BUfNfbtU8c4f/QWYVp+R8ljzg+8HFEY3cfKYU2uD
5Wol+51OtdYbZQuPRVLvKLL1xX9bUwTeLuH2Glrloa3x1kj+VO8X/BGdDMqS2mRSu9nU5aUoyZCw
x5PEaZZuaIVEyWQw5Tkn9qPYPtT+LW9/R1YoJVoZ3VqLMaml1OFfYQ01NoZP8C7mpYwnwomc8ftz
DbkEvReJtQ8Ck1kh4MOl3sYn4q2XzkrReAE/i85CzeDtYz8jkZEgMX9K63p1ZXjAWOewCfUGbZIP
QSH2qOBTOQxxB29dSbcN3yqjpW87Bqtvk2WpyuVmxnD2LLVb8kOxoOXK6L6l+Kv7cpbiBtmjUkFZ
/SRaMA4AZoT3Tn1F10WicY6+Luq/kWjsxOSTdBC9lF3z5/pxYrHXOlFLta7dQkQ1ZD3tvSkahqOJ
IWl2TyRatOzexoVnnC0IbUp/AkI9AiwZ0/IyIN0zhPjSHbIhNpUKKkiyZ0yjxRdqYMX8f1gMEhMC
6leAhA6PID6nF1g+DQ+f5Gmm78TmlI5FfLmS7Nfw1ruaZ/NntWg+BVTQe9/pkUR/55m3wCoaVj4j
d8QL+3A6N98Z6hG4MWs6Ovcx3DEGYj2negbZyDzZl2eNpiYKRBJqCvm5KgAoG2O35BE29jbkWICz
xToRv+nwPCFQrwoNbsumzKFV7V9x/RlgDRRJ1Ccua0/lALul4TJ/CIZ+dqE+0tTBUxj9SafeP+OO
OLqrKY3VsOGHbH+xf5gHxjfOZ0vTt1gSZjtIkFeZnAlL5Gg5zuB3VaTMUcZOTYyqdg4A0f+VqgwD
m/MoFD7YkJIQ1l2+aQI9ZQnJL8HD5A4Q+VeHIRb6Gh4/XDL2fO+YGPBdUUMuNU/1Ty35As5AC60m
OuGCF+xnfSnwetNwMlpiptAqypHpvI4N7XG3cdDLo//9we7WjJFczlgPtuR+F/WJhOJ7IPStrJnS
ywQ2HGqr43nO0sJzZ6gNT1lpCz8k87O2ueQ9VM+prOouDfkUgDrHErfs9ewYL7EyGzOUzx2zo9L+
VaI+SNf1yRaW/+laJMfzMRak74y07Q1NJkygHmMuybLqtpzWCs14e2xjUWrVWbMuyusM84R1xVMc
H0gLhvSCzILZ+tfWmi7jFPOlTkQU4h9DgsMqrUIBQKPdsif+DvHG4/faCFAYIiOtjYxFUaN4U68l
2J9eQjUY6FnvQebdX46qh5NaN64V6wnPsd6X3j9rmVaciWYlnl+EwCbwbW7y0upI0D/uaDgnxgvJ
NfTsZZ1b2TTN+iskDUwjwc+hgp/SBT4NhRDyvibJY8FgAFg1GajHVr4hRCNA/qLugzqfWoNbWCVS
uN4juJRt46L4Tmbhdw5H8K7V54VX8AT3MmI8B8PXGNS0g3NCepZd0gLmgbH7lzz28izoZQ2v1X5Y
0p9uGEG8PnlKslVD6pF3ys4QJNVEi8jb0J3CfngDgQUhXSlG2WFWql3FsQ4VOpb1rAbvb/E5bZyW
DjUPag9ioLTwsbYjDL/iFLnHSVH4qZ3TqO/RX4lCYpN/Jw1qGxIQGMsRI3Bm7gDL3xvu8RLpmX3V
+8MpTJVKNMV7prmhshIkFMDYUutpdPFuA1mQTAEgNWFyrbzHeiQlCFCJwEvTv0WfuSbHyOAF90Kq
P6UiwxAS562X1tJL0EAEmBiHVISDKJDpPMDVGEMCmQAI6tvIe033uEuXzM6MaVHYPgmJ6PKhATll
BWooT9FKjrMkJU4BDXzv5auxAQY4JmZ//GWhFfyIzbmEOvbmGZ/5X6ccexbYRHvYELoGqFmW7c+e
HULpCdeeNtTrN4AKj9NXubv6QsuifX8NN0lM08QcTu35Y5ep1VKEjkhOgbpbfYhKtLb+28G6B8fR
tzuHvfWjN5IXnUwj1/7LOq4zYmxsYUshyvkVOEfE/fvOpmldugVWKpDwlZoF7VGd4HAUU+ujci7R
cpVXHisWkd26PFri89EqcqhX6mGA3ttxbuHSH272xWK9OatKOKA+96911wEQXhNyDKVVzDRpxBAP
4V+AnhHwhN+CJwAquQTmtz1qz7/P0F4kv/QithkqqHZG42K7Z7fNqE2D9vkbkapwiICTmVMWQ+IW
0vggcaKJfst5FgdhKqQpDSNHjWCUWS4AvFV46UHUZCYYfbC5epvJvg9B0C11NMctBrQd+A1TzQ2l
28dm2cdQRPcmQLIkOceUU15zXdwn3jwKauFmkf9oK2aLtXhp+0X1BQAYsGNB60kSijVdWUKcWImK
NpD8U8fe9W/LmkIie8Qva2LsydZJ0YJ7IU+v4uL3Z085sRoniunTsuRMi//fdMdQun8WdlaN6G3z
kxZSeb/x8F0yUsQIb2dFF4WLDPBRwyyqyeyBe/Q0eLyIhQhGLE0nP+9dlp/pbBHMVLFq/5EP/cpb
fwYEctjJO5XCeQj18sqlWWJzoMnRtANdh8oQymTISe0Tui0GXMX69d3RHX8wxD9+chGkooXZmnG7
h36W/5aq2v17N2rXqHn4WdejTX8Ra92+1M4IcOhzjTgRlgQeuljys4gSSHeQ8JH8Ufg2ZejODenf
9P5EY0MtOuBi164ns9ummBVIY9RflCN/FP8HXVnSWPgHiVdoCxRN/lTsOlznR4cUsQr3ko+yrumK
K/Z0S9aCYMn4WCsTutcghJYQIF97UERewQRQOrt8oLumAkvgFTdOrFSv7XOx6X4QqzRm5n3TSaYP
rFIUKEsXaMCzqtP3pi0DTOTwf9bvBPLPwT9TnVmM2mo3jFbJ5zzZOH4Omh33SuQIBObiO6o++TpZ
t4FX7v+Jr4xYfGHGP5jkdaK5gtsaY8eh5sRoXI/zM4UJ4nl8XN4Xm7SNt/uIRw5lGPLTHH+OysS3
2jjq3Znvg8oUCUzVx9N5MCq49iA1jyF6sn8iaVK9N8WdzsH5YbIA338WB5rjl5M3i5TX51nYUuHi
SPTRSsysKwgUaWBRqchUUIkVn9UGLzi/RN5zEbMg2HQpOdkypidJWrT6YMlpp3zWgrLwlEWz/4Xn
2RGiAOxLagpW2j0YwCtSpDyAcAlsJQBYCTkPsiBihMi1FzZEKq31cilplbvdhesbyZzOxxXfQTUT
HR4FVbprh2u/lop6RcGQBTXn83Mz+8nPEkllcIJ1P7YFW6mJdQIqbIi6AG3TSoOhHpO18iY39TwG
eFV300fmfDezhYQ5CN8fLwOj7hSKe5GrHchmyToUOps7AEpT8xb9RY4+st52FL+SMFiRLt6eqav1
kYUZf/S9orhCdqu97KJDDN5r9+SOnX5A68ZL2APqF6C2vg0T+AbNEJDIUffcAn7tDWwzxcEzG5f8
4h0lEOk62I65fVIz0v5gI/X4EMHGa1eLGkM332ypJGB0qlruJq9ckZppB4Ol4DK1OfJN2xeICK9m
nnbG+KnSWDGnHt00VwaTeHHHEo9hcyQ/BYL8hov4GhR+IJ8z/d6+U+quLFmojNH6VcV1zwq6R/u1
xOPmDVRPgLLZPvPtl+yDClCuXWuyZuqSMqXOuLPOcV8D2FChg9MnulLZkaz/lkw57vCHn5p9BsgH
yu0NVDBzLKJdw9NSY6h4d5R2YjhWspUcZXj/hXaxR7s0OLNPudI1Txf+7Rhb3hgaEebGk1BdJziw
XecJFYWLadH6BLCjKtUo5HsoNpfQv2vckmgO9aotHfNsA7Gc15LKrc0JVJxI6epCBSAK1UyB2U2l
M1KhJW9a2ZmOzwID5gJmjR1uW2LFqe+vNRpHc+964WmarEQqpx+wWW8nxzFNl+nWKbFdc6PJvIv8
8Z55N9sAOSoP97L4DKsD16Eb98MsUXnG0SS3UEs9X+7aVeYQN2J3/HnOO22FvvABndMogr6gSdMD
pyx951wTGP/1fUlQycBM7BU2aNS+DHle/YFvDchRxwhjYEwcuUhGfMyapZGFG5V+WFfiZXtO3wNV
tsWRuLSAEg4WJehf2BHUj1svKBZETZfQ1J2Z3l2oBsnDz3Jp9BCDqRbUcTON6gKGdgp2SqDQMM0V
5ZJLxWYhwqNNYtMG5TcSLvAe5LccswjiDwixyDE3PJKjSNu7/hWDtbYDiVuQBHalUoPTJ2khGWVU
TzCRmMe97hJv8pLhXztWh2HybSeTyn+JEdZWMYhruU/ylBs8okCEEmJjdm3Oj8fF5miAdxGOdtia
b10M2OhbEcJPJ3YPwzRB+sONdvvBdTbVtSHieYYz990X10EsFlvvEvDTS/bnMUDKB0m2lV2rCgFq
XLnSNqUZixQNKbDeyRj925DS+tCVPbkCzb8VAFhCUKWMsN/wbm2ACW7aFV+59bwl5Fwemts5lvij
E9+Dx1Ybv9GMvlKIuW/4+/6UIUHS6gidbknUhe+cYBjr9spkqoB36GeSHSW0SsSzwYVmjEwcQpOA
NHHS5eeFlabSzZAAwAhSsl+WtXQ8D6/9JsdsPZRSvDL5LBRpsXqceomdnQ6KzHnA7/QdJCpfCkeK
GbkDRsm/ZJluebeQxDyJ4Fh03EJ1k1QxJinKy5EN6V3bKhyuj2Ze+2Oyh2zNTLUAOh13jOa25Xme
2Ia/9XzIIIQ5U5PoVcAYR4y/etxZzXqd9Qu5XyroU3Ux4cnkUu6qoYEV7gOWFKuNongcmnJfKFuZ
xoallkyBlHo0LkqiioJFReER0k+dzDtD37zAwQ3yB41SUoKLBdB0ubmIYCKJ50OFHOgpAwaJbil6
pQIUrLSlvoG3J0tLfyxief8SV83OOjxg9jc7jyUU54saKI8gK8bf0iW6/R5O2Qz7h7xSJbljv2MX
bOcQGWK9q5uCIpsPcJ6pCvjaWYx8eP8lF/zLOD7isqzxA24s3Jp6IocsyNkXCqFA3ueGDR/9Cgm5
abYAWWF7RzTQQ7WeF0WiSssLeOXBeQbJYWtot/zXror6lVuVX/om7n9zdG6Yfbt6keucza/XpozO
aoC0yZlXvq6o1mGCo9I3scuThtKJqc9286k1ud/C3xutyek65upMhw8VEQKPfBS0RZ1Rd2wDM8ho
aheqvePAucd63YgNxIrB1IvIXpo83FEnoUgOuOFyL7BHmvtKMPW5ImWkaWf5MxC8mah4EmUKMqAC
0naWODrMT0xKhF+kRB+v8lOoEch+PIyOY8XavTCaoBLQySSzQbgeA6hHH4Ci9kJen48tteLrD3HR
NzqDXN8x13Ii2KPNy52qEIavTOYJSGbR4bgdnbkYHbXuwNVncyqnQwR+79UMVdPTHSRHNavcTiu+
wdvraPbdLrb4fGIifwKSN6fXm0xMBTWLJgFzOPZy1xuWNpcrGbO7wfmxHVoBU+JsHLZPcWakyCmc
DimJ1sScWORlbtooQ9rAvIzUuvlL4TXQ3XTeM5z85svhPWRD40Xa0gUKIIJPIuV9sS0LgVvSP/kV
za17sEM5MjPKvd/t5+6um5xIhOAQvOmYAmlZvUcQ1BWQ7/uhihESjP3TbfhyyM7E1kr5lUBz4eNN
UOmWQ7Z9DsAFRrG92+lhR5HD0fqiifywqDMVQ++/+5GMYis0uQ+qyHobzjzXFMECGNb9CoKJyYoT
8EI97fNs7xUmugttVD4cOk49GwDPYvZnP2oGrsG4BgZ1bGGpfwRBHAQxD5K/emH6/YrgEMg/gg3c
aKQGXao8njSSz1gWef3qFcFeZAnJqUdpiSNwqFGubvc479AgS6VksgCYjYN/3Foa6JQIugRq+ihV
PXD3yohDm+434rkYrfEE7iX/r2zzKERkWGbqEZnRwpMGHMVIV/1tIH2K+GSCakPa5C/snZJ8A376
l5KEedFSUbsd0uyNgNjFOa1wvZswT31PnGSRLj3BNjT9mJZsLPFyBK2d+uDWl7j9ms3+7F0mj48q
/b18VzvKovlK/8EGHew1tgpJKmfXA9wuJxk7PipzqGSYAcwpED4033Df13pK++RzbFJ/6YjsiTUo
nKaZYWrZU5tU315u/3WWsjF1t0G0nzeuYru9SQBPn2V7FwSkp0P597D0DlW++G12km9hryf8VhLW
OoLqUzuySF/KHr7bhwKYcpcHQdwryit6KT6XjlembwI4A9UuV9lE/Ptlwm2kIRArZaN//ExKBDcu
ZXGFYWIlkTE072FrT9ZE3d6WWg9xqlzKtGtOUAW1QmTtrEoaAmIa3pxgeEo1sFFadNp/4HIexbu8
y/tIgXQbEIxFFEUAmAHbq1Kh2K52AVMCqzX9d3hBJMW9q2gX3iEk31E4sEQ9NEOSEw8PrzTBs5cL
/R6vgRyvPPZ8dgsLlH11LKOgJ2+FizKewMdZOVAmzzBNi7r3LakxPtjBKZc/01cG3poT3kGtSegf
cT+90cJwdBduS1PTSSDMMddje3GmJRQihyZIBOE+/qhlLIhTf0x8+wJdqrC7H5E8n4wyY/FMzPXi
QTbxAcYFXamE0Jf96OB+tz81l9FCJsNqlsgVdIzp47VYZjqiiDAPfNJktAhcPl5eOf/NlwwizjSA
QvWg4Xx0aYGAHdhjq6DQXLd8j1JbXHSII8CVPTozcRUCJn6xnX1u8hfD/QCWIrVtL+PglwdWe6Q+
Ho5oi5fNzKmoNPJjuJbaUql9OstHhdDDLPAKJEnRrL9Es6Gu43jrqcpVS0rvWYcmBPsvjAr3mQ1x
VMS2e1sFIDM2uQ+FhUz1CVUCxCtSNpdmBaCuCY7xLVtu1Y4EQKF/xtgfBvg773ImVSZPqdvRDHrn
RO7KH2M3qmqe5MQ1Jafh/dse3fQS5gGJoEP7p2lsF9mWfLXPnwYgXZWlfttS7Uy1l2aS7cbTCgBX
1U+NNCAW4HF/pBrKhOyrhl30UCCN8ND/Qf6cepG+/DtlOYTJsE4NS4scFwLB9e22PPB0VmHpPvgR
Zr2+YWWZ2OhF7PSoDf8tneQkEjeRgQwJTuZpvbW7ti3toTeRzfu4EtCy1z8nqNfo1KSPna148XtK
ULIorK0ACrJWC/KpfVlxw871lkCfSjyou20T51x9zpC5qYpFK03nnWQZjXEpTEUS/0zuJnI5qsT2
64Ww8NSmU/tqn2gbM94VeiLOyJWW9kft11T00hpTgQHwTe5Ii+G6tlHcsj5UttW+gRco+ZpCUaFB
g+y8S/2rDIvHqW11a8GmhnsITzAOtCdX461rk5F5f/42yWD4dc1/kFw6A/LOqAeYKjKazWkxjr3w
1UBLB32zE8h5pVjH6zulqTYP/T+B9hI0muZ8d6BdywhQjipz2C5m5g8RNiTiosUrZNL1t/5MVIO3
asIBK7EE+4LW//NUbE9PLJnyhIdeqACzyaOqj6/J7xi52dWnI9DDsBB4v21fzlyhlYr1EdZYnbe5
czPZANZPas46RiUcQYxJSTto9+50XJUKwhpm7VJhILW2t0215nCVEWyfb5arYvbXICl71nX5JQ79
b8Dl5cWIA8lUqDi9kSgPFuGgIHcfdNwRqTTtCHWk+YpMB+gp1H5GJhDAsWeyWeaFwan4BtFLylnP
ulFGMTGixOHCS8UJz4bGwyaXtxCNm7OluGWDe2ZyTrQTXloLkPumMRByoMNF1X1HHQGzKkFjgO6h
wmejLGTsAFEgCdMmxzGG3hsL12ftGHJYd5x2pCkYj+BaoYb4V4ZdoTZOikoJ+eTCrX46eO/qKM31
01EVhJ8TowxPjK+OSxQnOQkzPtLbeYB1hXc22HPOk3CVX5GRTiAEUv9QZIjndc7uyaBtvYvqQWU7
v2MevVXgj7pHj7QtKbk/I1NesEY6mHkVqF2rIeqoX//kFoGS7Y2OB4E//nFv9IYgR1zIbzUTukyq
SSSearzUzPMc8E1gDd6/+78lBlgoHNkHLamKXD5JlFQV1VLIReWfdQTCKoesVV5U2m5oPS9lHKum
KHgQM4YZ3+7eIn8ZlMBnObFi3Sb633RcuKWDqm6W1ksfk3uFpXPoXsmVMq+QNHqivsVDvWAlkGVA
P7VsCJghX8rexy30KIPM8Crcjl/exayGJf9MdbpuI5EQngT2tEXuvLu+2Ru6A3eMC4O1cZxe1sax
Jnp2OkrAFNMNsYrritSwTXdGO66jnIhIePorDdHrqrICciiCuoN+3AMPR5LeMZhGH3O2gTxDHMhC
1f7/ULX7jSdgKV90QK7voUzkDOr7/7BcvmMoZL4bJRjNQHmfZc/Rv29nf9rmJ7J/1V2b/DkVDvAw
YcUhjp8mfGCUwJZ47TZaTEYtAhVL0mfiFNVf1fEuf77VB56qxciKK1ETwgksf5a8dR68akE/sP/x
/zOlMGTGAo0mClU3EGwSIXU66RaJYmdkuMFQ8LYg7uFiRlml15QZA6nHqhBKk7OX/CVM0QEF6HgA
HRm8P9JaxLxPtlxr9TasuJ3UVJA36zllGK/K8vrgmTAYu0MZbpRf5yiYwNPEjHhYVWk8SilNr/+F
I1+4cki84UasRjhKqVbbECiGrEUlENTXCqChJzldhLwra6jKoRjjauEKL+6Y/y6vj9E5/I/tPCN2
6pJWL5JqIWt2I12uBlGaBsAOg4hbdbdpjLB7M2TVbPUmdLqev3aQkIgOqfgIypg8PTlRWTTF8GN2
e/9C+rtulQYfMYB2MKstv4NxCIdj27YX94iQ5La+ZtZXtwWu3wiyz3mYrzb1QFMpZ7Pi3OjsKrBS
WIIFM6I3npzpdi2ntwQn71lvb1WZOUMKhif9DxopQtzuzUiJes8FbZj4tqV0dRzLUKWMqvvQkgmt
kJFB7sp8jFH5AHRUD1PyF3H45UP3jDAALrMHzXHQ0x/qRxhuT0jUvaKHXS9qMwda2zDxc9pip5gM
tmZYcmvCCLuOgVFmgwXMxDTTWu9379ySz6cQWy56mg9Q5RPWglqGNqTKYr/1CNtzPeWpb6BwHYpf
S8mERUC+HCCV/TODb+zi2tKSGJcdKboTz5V28XXga4x4gALYW/3IK/oMkm946XGon9RLaZyrK1lt
8eXadKiWE4lHjAk4fLxcQ/7Y4GcEfgB7STnTK5Ly+pbYbstx07wqCOsuR7fUxWd704OtN9meWwa7
dn3+QTRjI7amRJ+a9/Y/c+7O0M/+7AgoLAoCTB8fZtKU3+QFA96aF5sAWd9UlaJGUZ+T+JFcjYtK
bm2SfSaqM3sC0fNK4x/1/duKu2DKezhQS9zd8A54PUbA83JCkgYhG6offbZbuO79gy8JM58o+rCo
Ukc+8OSQo6vTcA8jmQgq+XHwIaOh8xHc1vhwah2PeqJg63PB0lAaQHcAPzoGDTEaFq/zG7g00ZUs
9QEw69Mpqp6l/uz5J/iYrmS5EnTRM7I+0jqFItj05up8kbpbg/0y73JhVa7Cz8bextSk0aRmEzku
Z9Hud077/HpM4GXF5bWczYEy//zkM6c9b9AwEt44uhf1up4VmLSEZkCq2l1Zo/yqzv7H4/57lR6C
Ku1hL5CNXqYdGoZ+yzYmwsu+UpBWxPE8rPh0z0+3XVnR6OZ1wHtv6Xkkqdkytkg6NawZF75sXQxb
njibpk7blGEW9I4gKb833pMAuMhGURtZNsMqg9u5KJZ7P51JWLLPu/m85jIkruxRZXcUA7L3NI6m
8u4KFjqDEKXgTBlmMHiWjAlprgWxVFr49mKc4/VVsZzPYSPRl5rtARklnPxW6sFvwdVpqnP3lRYF
v9eqmKGsAmyy7MbdR1elOQcRv+0Nf5WvE0cj49RKWKQIbBYjr3Hv6uZnDvkuY38PwGyRd4QvYXww
/q2cazFcIRvH0yejaTszmetvNKGsF9Pp7aUNqKVjYHAwS/CTdm1UgsFwoTO4S/4ejDhTxWR1phen
IBwwKUWz4vdzDZBuwz6mPvZFhto7Z7EL4h5qyWQ4326zGAwKYZKAUAw430CWDcxrgdnlkXMRdDuX
qaQV8IsJXaYIc8p0fyrQNzqyt23BRKBmUULUg8kxVv+rkrSAxiuxmNbTBO0zwuwBnsuIJd5qxpKW
WdKGS8peDruLRsei8UQNT/CuZECenQTxS7V6YNMIwYtrSDvxim6+ou5cz2G8iVLuKII/h4M4F9p2
Lc3XUxpcZ1AD5RBaKRkYQesoF7lC1SXstV2vrpLGUX64pUCSjEodQvgwDB1cn+s9+tSIB7pMxFTm
dx3YMS2N7eWhSQ5YcciuDyOwELmFLMEbMzJ/Zi6y3jiokcMJMLL2qcnb8yPDmjfahhluHctXm0bU
BdvexXxAL8IXWf2hAUhxDGYNraatGAzsPt0VfAqfavgroKrOWD0JfYztPV0jvJpLuT4Drq+iv/7g
z7C+4CYGj1OCM3/rW7n9z5G2ixh1s4F7ryldo7agrWAwxfnAHXtnmPcs6Lo+KfgksEi22QOZydE6
jFxXktiFnnDEaLVxEmPYx57xDJOXE6wNuphYlz+6OpxVDDhvwJpp2chxHMuMI+F8O6jB8EAZzE9d
ewSjUSY9kxabhRJv2xfVAfiEE6KquHyX5Pl1GRpeuEtZOmT/HoO4CNjAg3WBMLEerb1H5+7ceLZY
xGGq8tK3TdTdJd0mFhPI7lGFMoRMg0mp4iXYeTPKQRGH7R1l/tuBCV7ZvfRWmGPoAKPb3WIFufeV
jG/Xk3vjzm2W7L9hPBzKrfzABjCCeSPUJoDhRDOtg7SPMfFOJW9WTH1j5eqW0dMhidONbxAX0ZfT
VB7GQFwKqQQDiffm5U2J+vGyS1Vn8R/W6xDdiGeFoefSBQCsIy4aNd26WVkpHvPwtVf16pMXEiv/
AbJQ2+cMHu+DfbJirMPL6zn0iC5Xb2upr3ZNLAgzTmbNu+DeE/xBbYXxoLX+6xD5fmb+5AKXtW/N
IN1zGtD24jrr+6V5gG6Bttqo8e3k/1WtZ1uZX/pjqYeggCKzRDZlHHWmANIe4vOj06y+gLbjWC6z
ZhIx/YdIURLXJ5ymT55UH9Tg0wZqFC1modifw2OqKk20Ezpk3Vq2tUjAtTh8NVNW71uArwaBNuDK
02jfnlzwRQkbyUSplxcgN+vuM3frwUX1EJRg+n8V997h8Q8jWaS5Erj7Jq/rpxkXlkPBkPgmbwFG
P5t7YbnCCLOmH7QmVN0K5RIfIkzPEhMpjawgTDqf5CoKylmfeZAczeoKWM0BR8bcIby2f9vrD13/
K/ix2FjEKIsNOdQlDe+7uZ1MPeREU4a+Ch7BN6nzjz44Y0QHfTc1HE5wRffonH3mnwVvJQiaviLm
DD2lAJ+75sxEZ7OWz+CZl8+Xw/Cwt+Jeaiy8hyu5JjLOmIlhUjIQq8+mIGE8MC4MQ1bQ0abhGQ66
jUHgZVNqGaIHJNmUlQJ1AS5twtcdRuo6PxKaEFiGVFu6ihPHk0YVMNSrDTV4rpj607WCAg/ZGpQk
N/mCEWfu3xJ09hGDYSBBMFjgF1fQl8IboUQnaSugBpQVIFmqD/5M9TO21YNwUyHvTDA+p5YXZjGR
wgyeaDyvqkB6YJe5ravg27kiK/d5oJXQ3NARY7yXUYXKClZfGdOIQKpixg7GNVv+/B3H/hXKFa3w
Eog/MLs+L4SRCkzp5G/2PJ1e//20quFpK8cGGm+4LIP7BcFyjBYDAYZ9dg1ILPfRO0uIlL+b5z3m
kJEOH62indWu1lyUnVkl9Hm9S5sU3QGo/FUMP6JiY6VW8zDj7kN+OzHQwF/WLt1gFGiXmNWWZdUr
z5qUvs6lhpCOsTd1DI7/UY/dQunBYxfEhWhLzftOVXjJfYvj7r4QY93bZTj+edbdlXcBqsN8VlEu
IPBz+Iwj1AANJLaJ5ZCKPiS2dPq6THIxl6e07+P7JR2P9YN5cBPPpbb0SYk0QAfSmITxefbMVuWa
mmTVFrTEc2CBt5jt5q6T8RMdzDSXmhwh4I8e5ehcJpv3xvCTC7ChZTsfngOQ7ri7sDjMy4B2wtD6
pIUWfDTNZVlXeLb0uW86pqoShAfNh3sM9Ob/KPYNRD1Oewe0GOQTc2eRLronx67re+MgsEsUvwHh
LarH32pVyWZpDUGZ0u6bxC+h00Pho/+LrdF32mz9ofgxcd1vaUzCaZPvB5COCaDR61dDKb6cfCno
6hNPgSiPZk8audhJ940aithdXpwVDjJLjFsrtR9PndA65AkoVub9xZjEkQliIPMPlVSKNKYelJN8
dIkVJOxvr1smAwctVArmUcdWkIl75YLl53KmahCE+6m2Y41UYxqmsHNlPmDtn8aDgk+WZsMeCzKw
h6oDHsGsPM0gT0fCG+Nd7A8rfRCXacGJtRLY95B75MXlDc+cE7ekPRwPe1mZcO60pz92t4MzJh5E
CGe2bgcjBg0dbvvqk9sbdbZALq4MQycSGFesCYrhyeoudUG7GcFmEdaRqKl/9+RQYtYd50Uju8Rj
690VnZ6CKZtTH1oaH/bHSaKIZ6lyelfRTj8BJp4jyRWlJ5EO3Zj+cYSL2qjuOcIkww0vW67RPtSA
7BC9eiuP00Wh6ozYPYdX/zErAhSKJFW+txnwzGGHYkjkOEZ4ydT08poV2OKOC9FghadSQKOzZsVp
1ttGkeHI04iB7LW5IMrF2gE/tET7/+haFSFZqbOkQOUQGl9QLZfDvh28f6AidJrDYlzxms9toE7d
B0GRLMQa1pxhHmal8AMY0gpwXoldk31t4at/m2uE7ioZ2R+/FbJXkiR4WUsYq46UV0k7Mjc3PIPB
yDKTDKXMZRrkkDLFV/IvABRhrtrPYCTh/7DggsFGl+ctKajFQTD01yCZKl3VBmBwTQ+nRPt4qR7y
SlDFtRIqCEmPI9bhEsAzlUqhU6pLqjthQ1KcXcflA2FeMw0zl8d8rFt8s/shQwoMiR1oaluwEuqj
DFak2QEfJXpdnZpEP+davs5MC7vph2LTOHiUCC/mgsJGxU8Rzg7FNO0CLf8mS1AIpzG5/lDdOf3V
xlw93lVG4IAR/lqrPlBotA5KZP7oNoklNLhBGWd/Q+tNMd/qSacZqO6DpnezJl/7brFQSFf/rVMk
s6pls28s6AJfo/yZmwiNqnMmr/acQqh8g3RKGAkdVn4Hn7xtWRO21PY8TTYC+5GuhBTqxbwkX++y
wQOsyJhNaTdfqQX3iGIwg7P580zUA3xeMONu7Q/z+5CMnFQnPuSOeLZpqGkDfGcwUUUYsPrrSPlX
zY2W0H1aO06IpuqNDq+Fn3jiJsZNudFD75FKAYPkbpi6IfHnkD0Ujsk9Pe1LtdIRl9AqHztp11p9
FXCSsN7PlRwl3Td5FXVHUTzZgN+Hj/NmMRCVUJaG9x6n1mK9YvJEtp9C1nGwHqIYriM1F8moB1kE
9gqDj135eCa+lijxg1jJWTQQGCYMJb4eWQuEXBdm7EIqUCmObiiEp6Z3gXhbmIonVWl+e1L4Bm42
pWGzKnmByX1EMYstPXaHhyhlT+Ad5FZfg49kK15xtTAORJblX8YNqkv6/HeaWUNhy+1nAMnJVbuz
lpCEzGxHpF1yIcBYZVIprrPuzEiGNieZaGJxPzeVRDE3TSNM0JAe2BuFJsbB8dy2gFU/Teylao7U
w5LVneFvCtpreH570pq6SO/UYnFPc5ueSairy/s7zwHrtveYPKsOcJL4GHqRHc47JXi34e3hTH+m
G0oUjhN1yO+4W5cdTzJGHjSPKWRNJf/FJ15A0KTSaWgT3pB4dDC5wAzQ58yqwl1EbL3x1NOy95Hm
j89PsTRZXQi+etMN4LrKB1Tp9kMRgAqg603EIhn4F9bJAw9SNJEa5yCjwdfmoMtR/NF6NGlhUuC0
tgjcmW7PfRK+3vqYnSLzgJlftvu4SWuOe12qppjJXp+DdURpVWv6rJov+JVwpW2yHDS05lxUC8un
iddifRHuLsmvmHAO1arkaJOa6Scdzbwcle96LlxS8Gs8pxa2gt2D11eRaoqv8rh+8q7M1RuePrnG
0Gz00Lv+IGwyZ5ljqffxdVne31lcUWwWElnnX//v+FblotrlQOAH6wwHosyCcr/bsROvfO4fO1NF
jhxXE62fNgCbyn6EpcBQ/INJoIrCOb7sMWG3wQwMSFFy92l2Y5P/4khKAxjAjIoANaztFu1JB0UD
sC4Dpo/rtCEiQ8p6eTj9/8nVXmJw7Kts4FH8Gd7V2oOJllDIl1TXfSpopAbQiYuBQ74nj7UV0LPa
9L6v+fHdLRCbdMV4nU6hic4gHBBClzjsr/fgTWot1afv1zOCWBW2ggnMSzpQrjp+LMrS8+N12aO6
BO++hOV3bG3RTcj1xCkd5jHm5Be8NwLS0n6jteyiiIjIO5sFUn4AIZs4K6o5tdxpum1RPN5S3w1W
+on7RgcLrUXeIqLUXwlLL+MsE9Qo51yJtRScdBt+4r4y7AqC5MFtITUJXHDcL8Ks74pGUgzV0FhW
lXKQID3rRhELF5JIVHAIllFqkrCe6NOWniwmvOcMinaBX6+aXlk1ZmU2pXBqU4wCDpV3l0slF30h
n74k2+HHmf/marhiv8XyTCUyGIxYEEG2yjYrFdyzJYw0kYu1k2uaavIkbCDhWA0IdSQBJPFMD5NV
GP43ZIEyU9x8Kwq4/Mx4Bj28thYISl3ZxhUBgX1v23UDhzff1epvFauTnULVOHYgy/TIbgImSMoQ
Gcij6FL7Ligpbchoag5AfkEW7bKoRujNupYoiqgTEATDt7N1f/LLr64J6dpR104/n3jj9wBOqZhK
4aUtfmUuu/pbXKCw8HXlE8zaz3D4GZ/U0O3XY1McMxOI8fX1SbciaCif9Xg9127xDxF0cknFpNZZ
aNyrQtKRzSzNvc4EKZbyJneN5FNafmOMS6Lkm+ADZkngd51gZclefm+BMKqV5p6haCTpzfloi5WA
7mrvvdZjai8bOmSE28cHjlD8i/V/QClOGxosqiVamiYuGN6SDNsD/AUi4qUEEtFNafZZvBGFcxCK
DvMf70S1ytxnxogVkhd/SyD+KYYHfNhkKpYQuhwyQjZ17ZeuPshdP4fXFVpDvtrC81bfR7+FrvVj
YTOQZ77a4lUUMj1DN/IozCaSBErJXrgbBOBd8lNf4nVeVL2Hu1hWc/Bblnw1+rhv+WVkJUrRvVf1
mdU7fer8WCiunASH5FWb96d6qqScrf6f46fJXPLsBEhMhVQEiD3hReBAVtQhOQrnCBhXpuSCjtxF
lpE2FAPiivJvvvqtRhd2+lDxQOvvS93xe6c1+nAHgNzw+IVRQKADI5siOheUizxHF4IptEdbGJUs
oRqoqQA2QqBcgV/wuiSx0EIUIhv88HWy8dRXkiPRIeJkCX66w2ga8lRMg1WAuYN+hI5+tAwFUpE+
xA5MGPpP1DsAlPyKnzQ0rAEHx9LfwE0EDG2Udpcuu+smxsJh1uZrOUjM6tKz/7BZb2WHGRBCb2bc
l9b8cINQjrQMm0d8rac8Zz++d8A2eBVDwY9jWoUBYCz64qS6Sh3TrHwzJnW7gzHD55UiUKjp3sbI
QytaF34mtiN8qzA7poo9s1o0OAabpMcA0r+2XJo5UE5ah0Ii3DgdfkRvElwJB+cPCO5H04sK1HPJ
O6VcoedkPKplFqoWXRjLMFTuAmKQg9rk/+tgqmks7F72RVcCexsaigV/RUpxL03P3FYrXVLeMcfq
NIIVgWddvvwLL/DPEpxOkCeUyRTr5iUF1qrUJQjDMHaMKX+EmJ4rjuaKEeHQcq5KndJB4LshL1p9
Wl+LrnftatQAcATlQybm8yoJ+U3RFaOvhtjr+slhmosx8NRW8ylMUH/IY8lm8iAmpplL322/UvMH
7sDIlDPM03XOl6P1uqpB1tndkDH6widb+ezLb3s4qqmKfd5kb4ttDmYdhnshfh/UhGRptH3P7kNS
jGhv1zsIc4pl8Wj2QQWEz78Q0oV5gaQFsqNqjKVFfCGRaQBsGYplW2TI5UIhwYijVE5IvomtLhp2
CCZgCzVdRvtnaBXOkgTkDSIZleBfbPSExDjODqDf4abkVX1+5z1mwit/uluK0sYQcH9+MmYsBolf
ieEpa6hY05rXYt4Up3lsmxxgfm5Mh6X6V5p9wBEKuc2dTLMYJxCExUrxC2AZXwrDOpLh6hHjaeRs
EbqJXVCbmZz4nJFLpa0A+A8UpKdM4TyXZCKETQOR0hnMXbPRLbc4u65Arw0zULtvW/U+B3ZFy8bw
OlciSk3ZAsyYl9/TWONNRkVk8twcRe2woI8E8/qShX2rT42U489dyaEaUpuyu7CZ+QxhdN+lEGqs
hUO687tRuoffN696dP6s4H2BVU4ZihKGn7JP2jARjJYYolXDCZB+MEishL3ZTAG3et8WgCxMESS1
fsZxkkxSUzMLs1hmEQx4NPbr1WEZL8J/63IMtpYcTokAmtId1/Sg1cpfh4dZMP43DThYgcglm3Yy
PQQXUS4p5YUdEEWHrF0RszRHl2xiKBWdMJ3Wh6e9clckPt3a5X8qn5lFzniq0Lvigidi/6xjJtvX
QrOA4s35xjhAwuEOCdlbP/lINXUaIil15hJVgFz8ciJu22UUVzl3LAGZbi3RRVUoXWHQkL4S9NTI
1I52ibOaQZnYx6unziHd4jIaAANCG4FZVAc7GzSOeM5OL8KCQxtdaT8oaFrmeapxqKqT2wFyxAJq
0xBI+J6wd2KYc/mUwaCnmvTStWATeWFTb+YknLjoD2uWxCWxkNHhbfXOcv7efB4g5SWfJewGEVC0
u+riBuywBrdZbnPW+2+FrOwcc4GN0C/RQRTJprXQ05FfWnaIjXr4CwdxWt0jiT1DJodYIVCL6edU
tp/MMfoOhJMFkVzPNvIO3i9iYCGxOf4sVHvIZwiGv9XqRz8LxIoo+zepN/Y3UYxWZxLWT5iFskg4
gPdYrUCkVYdR/HZDECqHTvidCscE1qI59yeOoqKwG3yrFalv/H9hK/JPhj9QwI9zex5IgFVe2rbm
zh+eolIgH8hJysmmGF50eAU45QMJkLIseSUiH/HGLSUUpQQE75EkwFIhh1sTaYZAZ6PnUCo9F5we
Z5rEHQiCUv6XAPDczNGrw93GnOxlS9sId0SoJYDwdgNehgDnAAlfWEEDFBw1fZcQUi0PKaRR7RaK
l4dHYIyCO32jiAUuVPzFqnxKAOJbEgGCzekCXqukhWZqjFXPaJbTFh4KALzr8nYPx2PgiAOlMZqm
0DX//pV2IYURQEz0zSY7HfDNMf0jWDB3n5A1TnYn/PgbWb77LU4ULFbxeZVpevx/yh9VaNhPdHMe
BFPMQ1FQCYhxbNPOZ+stCO+0abhsKvWFwblczFuWOv87aRdk7vso78ol2bZazi0yMRk+2XUh0+MU
hAH5Fa+l55J/2NHnsGYZswa2jE9d4HEb8MBOYd0Lu9s1OQnfVjOKRUzbYEhiQdlp2W4NrsdRgLyf
q8vP4odTrFIPM2dJNQcfLdIZk1fs07R2PfNwDrqG42Tdne6XC6ZwaBXXepeEUX5KWqqPYC8Is8IF
p9qtXCwdxJ1GG/Y3ULk61kfbisGwUMbfC4svACthO9ZyYxp1PntgYf6IBbSGWiTkq4HzgtZg9TiV
UdS2gNIpyBOwd09PY/OXvKjjjKPbC4VS2lhzsTe05Mc3Wy6gB1EmM7ScugLdOGKIxeWpv4ZPRN/+
2HXnSuI1R9oBJ3tJhXACUVHngeQxBHGVeagv72Zq8n3+J7VlzNYBQVUm2/SUSv9SuBdVfAIms9sC
50V6EIrQ/plEtkk7JNRoHfnKm13ZwLfyVbaKah1PXy64APeVA2jSl8NRZm7AeYt+k3NGDDX3qYXv
G1xDF/NZAb/74DZwnLj801GpUwEnLayIvfIoZgyDXQ4dizueJLOh5bw9I2lRcR9+kOfsJrQzaUTJ
ssvfW1fr0g6fMK7ooYAgbfycK44bbpz1YS9CaqQiTh//SX9bQg8rm1TYhq72aUwFIWbHuDJkXHle
y21m6HLZGTQTbfs/An8flw6d/t5ZIl/4I3dLoctkQ85jJQpkj12shi3gVZa4XRd9Vo+0gd9K/Q4J
c/btelp4RwdqUvm3Ky47a9LtnHh7oswXtX7kNMfKlcfGHvIMWIlKClhf7upu9NKWB+P/2RNB/CvH
2vsb4Ozgfr5MjA0sKASgqdaKiNUYjjnaYyF5MNxZSGHiaJCwymHSzuTkboduM7QgDZl6RkU/1ggK
ZLtPToxMuYbMWZ3wYSUKFCr30AqYTrn2uT961PpP8WvVvj033qscubf0f3oNZbJTd+ddLsWiDOWF
UaJl6O/yV5+ax5NmEH5Z1i+zCCKQ7f8u0Z05DOFxW8mY0OJF2vnreMGOxa0JusyT5VUd9rqzKV0V
Bl5CPqw/1NHf1ir3V9yOG8oEGB9ChGmlj3fIEK32CU8WtAePqa7M6g5KbsLaCMatHRrDfRfMH8aC
547sAe3b8linIyn1QKQtt9PmFRrB/ujCkXP/vTARszng/088b5HpXuWPTnHy49HmmvAzgpO7UqhJ
sOLeaefHe9ew+4VhMlaJKrjh8k+rY5vagPosHYkbdUGjrkR88plPvQdGI44VqVuQ594i15NSqSMW
7RMk9zGQiy5HXQHtgCN05n0v1CVjGBvSYxB77lJKFkovmLQis4bENwZh93Olg1y0ET0LKwnxM/b1
VmRAo2oKkhdp10qdkVSaWWM9avUtkguegTDK0npI7mkF/ev/lBaPGIOGefY7UE47730Sed4K4mLg
dxOW2dGERZ9tRWE/BR/QSGa3flDKd/UjIz2jonWsBkXH/6lSgpYdsaFdeixxYMYlMNffu1YlDRkx
dPBPM1oJOtByJwRvyN2cYsrrmGspOhrwFQztt6rciGbGh7nl/0vOS0gvIjT4p7Ek7Jc6oa19rcW9
Vx6Nc+J7T1G+0fMmM6emZja4AiNxgzDlVKLq+4xQP6jjuL1jfAcH7+TrsABAV/v5OV+mL3WfQd1X
EOUo0Iz6U349v07eIXGNdgpOdDEm8NmDVxi0+LjWSN7bS7K4TQORR/872D9JdNfI5LyDtjt/gbBO
d8Geqe6VG0gAS/AcFicILaGc2ktU7mubNDEtyWIHZrHVGdYA7NeKxiy9gDOY03yzGS5TA7nOC1gd
7IzqaeX4RYrVS+FC9jYshgPZeOdVC4xM2YQm8/wffBGbT4pMlcTDZixCR0DmeUyWoHESQUkqdja6
RjHqC2NRSVQa4djVV6GDr9LOSydZQMzt0xOTR4SDSPOGVGdUtyIO8E5yQOoSD2zrmTWpwewNGi+Y
eyhgCm4oKV/2laQ2UUYkY17AFO0lVVgGW0MkYJClSN+sfC4K7ojxZUU/NfMYcfjZ2VnXrkHyaKLS
ASbFO1Y2yj45R4X0jUH87sYlO6OhL5EEAYo53WIw1JRUPzEz4zIxL15b96fxMn7dCKGlqxvqRN+n
EI57eTfb/5Hlt9r3BiS2/+h0lH/FoT/BOpRa3fl9hjN7f5QHhpeO6qpAw1ms2MYDgEXXmAgB08WC
yEoPnNvTi8d/1vZtW6GYPChFIJ8DpXaqjcquhW2NUZQkAFVRWMq1O1Z4R50fppccauBv74yrELlf
DpSfP2JyVI9qXXJ0zWRPLFWSMgiS3HYb0vM4c3FeTCodpofzeQrD1ipXEycPYY74tX0TCcPRZCA8
f1+oIEZMFbg/wvRWjaxZeEgkSuhPQblb4JFe1if+uMvsrWAywbkYFf7yqBKwMxJha3TiZ9wbyIWX
nfCSSWZ3DgBZYE0eME4C8s4dbu1e99PXugWyjdA+k3hZkDTyZxVQ5ssAWelu0eJWTKKAAagMgAvb
lBXH1iSPgn5v5tzgKvgzdvvobgj4Bs2bPW8IKkROta3Fi9dJzi7UYjwZHaStlC/BTFwmUGAhoh/g
JfOt99ppYLsQwe8dlpRXw0hcW9nDPyh1mvKM3q0j+TdT3poQe91dqFnJ78zi5oJcSnGotsuTjLP9
2Vq9YIdbgsVWXUIqIfv5SG1cR7GiOccpxf2RaNC/6EHw6jm9oO4le9oCiDmrj29xDIA+/6Jaoa3S
F1MokKDSo7gYBlTwHVSa2X/DSQSNW+2o7SJgncDrBfM1uYkKzzf7IG6jbWxBfqDCaAdpX4KBtnxg
oShjGvkF/dt/pHBpNfn4USIOvDFRJ1IJZSvAW7JfEgh28IcITXHhq5hht6U1u7pLg6P7M9mmjZBl
BKSHUbGSULXVVeghalp40onuZAq6i22jxb0tKTxNXGIutle75Vqj6ngf8e+zR6H6vDq/iNHTUj8q
+IKx0+w6vV3k2wHBaRodjQINz0nIzlM9+5d/lha7iwdcwr5NQEWCRRkDSc2pdMaC18KBnSSg2Njn
dNd5vbW4hyiqSWiID1wOMoXq8UkvEdtTwkWQTJHtBq626lwDhicQoO8TGzsRIgQ86W7WfAg7GUay
GfcjAfqxvWG1HzouOnvpKTt18i/1g/LRqUsdh2d4RgOp9fG/24I5xPhIfQ9y+jAVIT+lCLtmBB94
tJUwVO4FlqM0HFMt3/6uClvZTFsgwvGLhJnRgE6y9JAi24oEUAwHDHPRAvL78rHBusdJc3pKZspK
tVJdCamfDbxkFfw8LjJe246k5Y2s9V78jcqNubRD65S94gehl37S96zx5aFHZjpuAqqpwcAcLGpw
72YLUSU2quUinIJ5w7x0Zxa0i8Mw5jyijdzPgW+YNLMpfrAiFNbWHdV3jzol/W1vsIeS4ioLcXfs
PXVFdtJNPyiS4CvjdQY/bUr62equDj6z/Qlrh79eHMYI3879FTA679tXqTiQuAe4jrdujyus9SNk
gdqrbN3Gq+t1BctZdfIbm14YCxEIkOFIlb+4Rz2BcvzP63w2OA/nwLaWy23E0RYr8xNfJMXbo1ud
12e3hvzH5wlgTFGHkH18sGZ3RYcLF7+Q+Vy6igQUa8qPZIz7IEDJpnnVUEJGyFNdtj6l/wYqWUmK
yKX4w4A8EgW6sXw05LoN9Un2zgqUpO9/0tbvN6A67mVA+OL0p2Ao4aySv4laK7Tr700S7EM/yue2
W9X5PNvyj1oXcPegSHcmSGvFDxv3IAffhj3PzkzPzoOKyDaMA5/2z3fL/7wyznAGwiCq1pH+k7vX
+X93ZGWfQx8ZrioM+iYtJLQilnibDM0gpzHk7k+oWZpNnKjmWiaax3H0enZHwUulxJG2jpy4X8l/
cM1UW961xM+YjjgqC6tW7+28AdOtN4MkSvch5QkBYkFPrLZokb7YXM9v7Qz9wmlK1xE0MDks7Vc1
349i7TqIM7UhEy/3UjfgpNnycdeT6ZO+6AXe7c0ViDHOmHhlAogixozZvBHebiT3l0CeabEPANS1
gsyuf0IK8s/W6/YokswU9BG2zj7l2G5o9EL06P17gK+FlJuiKG0hHLzRZSkQMsHZWPF46DrQ40Hw
G8QgfBpL5cIr7dp6jqkwg7CWy8oB0uMPoKI11Srq6HCuISNn45+PoWvvSXox1MzB2eMKGEjQ2hyo
Pg9aMHb13hPI7AU9spSaXzypim4BxuXS2KFnFmwDIDjn3nJWjhKCls98alSUzp5DotJ06Teyn5k8
eSYiBcnpj9tssfKrevK/l1eLkJimUkRjnoBoPig4PLrbt5tWsqWt05usklU2ItJ0FLsE2BN1zqVE
/kjWLFE2yfE1zZBHxy72g22Lx+cn1/GerwtJ73J1AyT5Z8K8K1g8baI3eNA1BSW5VzvC4+ctyvSc
vMWGDc8o6oF2PTw53q3/dJWkzjV1NqYLA0CvjacCQE61v9Pf6z6pvjq9bGGVsaH4VGGceYXwYFLR
QStDSO0QhCYdY8wZYas8P1SmyBzIESyXOBqSmy21o9PG1yPheRRX6YR3BFYSrz5BCgWJWe2vtm+F
ebb+J7+omIHpP23lIs3oDpdwQko3qFykP/8tw9Dwpa7ByUMeAXZ7HusEBSfSz8DwKD1mICyGfXf9
BJIaIBAZ+ewuEbPAhC372DRnUKYM8WJYdIPBdyyVWNMoyd602j0jIb6NCeSh/Jp6Qw9eHIWnPjg/
uIadFpKQETTKLGx3Ma0uJgIeS3kHNVu9cC7JBMk5ScpHvJBUF5sA/Po4TP/1jBH4gXzgHlSj9hMn
qf2h39UOd9lFDqFjDBBQ2oMmoEJ7YC1P8RHkY+NwwhaEjsaNaWpj04hj/vLKfoj63mDVFshsXjqf
DMTssl8xDClPYLgWhpSYO+69awTgaDrpPDHoKGkpDIErVwkLxxam1XMKcfzhirnCC08KRYEWAUmt
C3tSekn/SGE1qQHzUd0b+sWMq/rqG7EwCqYliQm9oWMPW9qetp9jvw+OO2DvHrcHZLi3tf71Ua/4
yP1LTa4mzZq3CQ2RDVrQk7eSSelUd0pY6xYVnUE3/56l6HEMdHwgF6rFE5jjvP8oWOS6oSGuhYK0
YbaA7hSNMQCGHRVZ91JDpW7RK4x13kd7/m2Yx7s/qP6mKtp9HRTuBV3sFAF3aXCAAKwSqVOc/ii9
jbXG8HlQcOj4yMxz87LnRwxhTb5J6QQxYnzriri/IITnNtL1tBIbXWaO+FX0ZhVtJ5qaTe/L2QdB
csALIgpwcGPfTAdKdTJsyaHRzNfxnj/JUAcM6zlmQKaFp/uS1QZl2yhHKcqHA3Bd2yaqKtGzyKtn
WZpKnwqJUwBgMsX0nLUgF5h8QJwW/ctzrd3dLv6gAKBc+jz0x47WqeiyL8unomb6A0AydUgGrg1G
6RVHsAtZdTlkbk1ZVsx4GKcqZYKGgqvurYM0Rb7dvuiekb6vJG88CrTsKICldTDN2+UGtegRxHRY
OK141S9L2o9igc7ASxEfRCNG9htFlCRo/B3QSkh8v4CUE65SOT4ibXGGhqqQX7U4C4VjqNRF9tJX
Lezt6kxJ8XUgYsY5hf24dID0BkF2OjIgri7B2Djwe7DbygqxL+Pf0gEyDMwjin8DchMsq/zAdx2B
L0RdSlg9ARr7GVQrPa9+4yyIPM1cmlxXg08tkkbfDQmkyvsGgn/ru43Qe3OnMrKkUfsFlwHXxPoP
AXjRYwH6A6xVRgY7ViefLglnwMdUTSdHM+WZlugYSPAZ10rllI9OQTuImVE2CGfiEHxa5GElkWtP
7Ejy4xdJEW+7nScua5Y4/7zTOfjjmPcQQuqlHrHYDXfSEeFMpzYM6OXPRqwZnnAWGwDReibOX0ir
niHx2C96eY2YOz9fnmLIBkAQKCFreos1xE7k95+U5ufQMTTqK7yUvn7xzaN6QqH3ryuXVOBvwswe
vVAuygBANgQGxqgD1bj0AX9kfXTFlPNnGaxLsvVWQVbMMjbB84tx2470XgQq2ZszLjtdOXhNN+cZ
kMH96hQiptp/XcUeBIZe7El3emjKW51Vcn2oLILHsPzgrX4myAnBteGjkmO1hVTRNqP2nAP5uCIt
2OScD5XUBX+w6xqdKLxbLyQ8g/pPf0xojpWSLShxqVubeKbRMyMNUlWv0QDSwdI+0x4BWQN+eMjc
a8gukuMoqCp4qoXZ976FGP7zUTo018BLXn/RseXtfW8TlJ2cYi5PZfP/xNqOdt0dw3B0J9e8ICPC
2MQUg07DX0dmDKUFZ7msWEUyWQLzqosS8cVGvSfqKEe8V8Q8k/6GmlH23QZnkHuqXMWzAt4RY3j0
fQCVFJqfbg2wYzH+8ZZN9U87AD1iJzOvmvae8nHh1pdP4mzqP4Iu0C5FKbsmbn4IVACd2gkT0uYA
EqnMQcyJp/5Df7nYBAF4aYaQ+usMzCalTLdy/csqYs9aZfq8B9Vc+D4B73KArjDo25cSTQUh1Xvg
4DPuyTiDE/+v6iuX2ZFk+xoMCNejqqPT0cBRnhHEkcu+AKfkVolAwhc0SnWOC+WnUH2PyLzTPG5w
jzp1Jz+nMAqJreOlFQRCqktAn5DW2mA/DDwS+HBwMjpjTaN5SJ3bRZOeoPLJnarcgNOvHg62H78j
Q7n0kNTOOe+thQyGV40XisTCcl23RSTVzWtYdt24TRMyJPgY8In5sXmBCEuylGtOQ2OgeG2fuDa1
WuoDNJjruvDBfXrHazkviSw68nSIqz8QvlAJc0OlwWn2Z1gVNpoI/7d/36dG4kuIW2EAhA61TjH9
bhQVvdfbZasJS3jMZQAsZF5gMkWG3X7w/ScmDfig6ziNSxriMeDwpB8bcHpQ+PvO/C67pGCTT/od
340Z7L7eAlQaaR2YW2aGoylM3Sg5jOrbqNaMtCFvop2VyWEg5fNHQvBH1Nsj4t2CUuoAZxDp/mbq
26P5vJ+bLOet1mLbrB1asg7n1OE+92Jf9mg0+uq8ko3oUMD5MCcXyNYdsVnzXklq5XrsPhc0o+uf
986/pS/no498v/xxV9Csvx4vOoI3CdiwnRkrtHDMJGGrIfrD+Wud4ropRNj4XVnfxCJtYKLptCYg
jEQmFyQJcHjjNPlTC4O5Faj+JWHVUNfMRYfnmpVxCZ2dktoj/BRNj8ZNNmMswAXLnXYuj4Ru8HKg
43YKJ6rXtcYzFkaV5heaUxLeJqwhzVWm15RciK39dN3rEsIt6hGC5EnUftmsjTOCU9g8pCECCvaV
2ojMBQ9NBtF7FlAXqgGRbC59Gdo5PqpQ/B+1F2s+sxYjthwSN/iMEf3QGZFqmKLaoWI+9UVUfsnZ
yhVhBjzovsRNSI3d55TaeN5se8pZfvg+rRLf7MwMFHtzYDfYVSF7DzuqfnSW88CKqmbEFqpnNHau
MCpxogEXPUlFWLrz6aDJ3KLfZ8jD+zcysGz80/wp4ej0ooZxuKLrF1iqszYsNlxC99DxWU0vYmuN
leGnsPOS5Wdoe/TsQDVXgrUnvEzZC8LgT7fNXdJ5ZK1okA+v7pknCTLepRkRNqFSpthDIO51QxrJ
gucQ/nhnljvexZr8NH4j3scVtb6upFjqrjHV4JM9jvn4wnEUVOSzboRUDEmXZmtc+CYLcQsnBA/m
Y+4lPFUUP7w2vGjVqIegx5TsCkABFeTVRQ2wWMRTdeHSlfeD1BzseBijzNzVmqeQqvGMXfCT7oB7
toklUkk+oxfo7ILqW3YhkyUk4Hcn4jnZ62Xzk45M1ODv2OXf7dgbeHjj7IPy/TRLeicz4CShcizM
94hT2Bx7by2ch8SXLGWpew0rO6drl/SJVuLLT/x/PASIMmiRiipe79PAneXoMUNXzUkBpRDS8MCt
pVjfn+0/OJ4qyZ2HGcaepfBpMBAc1rswX0HUwBDYW4tvyBGH3vGiCxlQp6CL5UnQRWeJLmHPhnjE
TPbl8ZleKaNzljuClW5nVsxB+GV97PjaWuyOdKGdstS0db3AEeUMDMCLmLnLaFc+qeuWfrP5UjRC
zkaOslWZ+oI0fMGiqvg38En1OEi+6yhLmOSPoEZhiP7eppfG0DZERcJ8kbnM86ok5n7emZz4gFiz
BaRDBnuYy2aDsgSuydgymJu3dz1UV3lLRJweSjV4EKLiQpb+nIK69cIe4tWKWmDs7rEoFYrQrnvj
27WKftfBIKQSURVUqMbjCzOTW9Ymgbfwg2iHmV4MiVIWBBhnT5nrudlnUm1YOM27l1BOoyciZ2TD
a9YZUbsyTvnozuvKVbcaIIo3vJFtvMq6hWLWKZiJ7BuE3PuIDfMhLQjMpo2NmI35sqP3A9nj00Yu
X8y7wG1fZ5ZI8RBJo6vmoIGYYpHbK5ZBV2qlXgtfL4SQaNw4lHX4wp0XaOHpbLvExPn9r0gVC18a
Jajs8zI2qFRPLqwxCVEob4acWFWbgKag4U/IJQvlp9NkY1vD3DUKIG1Kb31F0Z1ERiJ2YRmOOiOh
L2k8NqwDknjR3Oqn6VArmneiQff/mZwbPNgPqD4GNzZKp/aaib5NAS5dmnx+aDxi1xOQ95QZVBFf
nNlSgE8jRj4sUGP2sW9welmMl1MmhY77+GYtOHuZLCVS2i23dZW7qXFb704aQ5N02rZtkKhdzlzO
PmmCLODX7qUXjH+20exiscK3cxcSuz1bOl/TlRylbWs9zDgGOEnBjmQIWZdkE7fJZfL977GBFBY1
ba0hCKUgfz6EKi0v7PgLiv06RrH8IY6QSQGXsuONvslqbh6+FJQ0Y0A9MyDKB9pX2YSYRHexakNp
2PI6B/F4/iZv6B+eQ585HsMAw7CEfjMH4AOjanlMjAzdnKk+Gsox4jyBXJuKzvO5KMu+OQN0VIL6
EZwJdVjGJKSaMVmvP9BM1SGWkTxqLmng00jvr77OuIPheewITmPZ0gzY1fXZ0RcDzr55uVp0y7vX
8qIHPhJcQ00CnMeFieJ4QZ1vBKfJr9U3w48qEUR+xVnIHgIxg3SbrSQuknWi6KE4YmfaEnT8/ZNj
BAEd2UlvCspn4hhhSJGukiBn+MAKlorrdxg+3eF3XkVinE4Yodu7f3afkJu/YC4+hLF+E80pEMTD
Fd4Y7ITufDg0gE+/n7DS00MWnB6LDYffrEA3ycLdWfTEecHsw/mqwh5wiOODAXOtQkXEwpM3x7wu
OOjFeOnCqZPMoQYNGwz9YzCwe+XdORy27C/LJzb1Ba6eI+QFPqDzz3Ia1zMRoWJstoXLmc/OXcao
GSHqCmSivfBS1Bx+w6Hu7fr5eRU+8RLKiwtjKVj3VunkkSS/NtIgjPZEEWgrEXO3LqfECGopG6k7
OdT3veiGLr9b1M/CMaUosX1cdm1NtUcrIv+oGXRDBPPiP7Qepjgf2a8jWpOi6GMpPPFweqFZIdG/
xLDj+5Ch5sN5/35rpzD4BkiM7+15shyk62tyBw+/AcoAp3Ho8WD+3L6RikXkyUFXjF8Ubs0/r+G1
c4ud5jIRhascdCvk2fyzQNsr0n+7gfP/00bEf+BHHjaXjd2LFL52bN893wCmQepoN2soU8eBmF1w
zYtImXvoCSj0sbA+zZpYffLpilOxwUdnmzIpslHNKYFrksBjETPvz04OqSXnzST0sBEiKIKw+AT2
WTElhpHHauV1vjKxIV93KxPvO5usCbt03jF1kN9u3h8RQufJBfWth7evY1a+pgYlcmeUKwSBMTll
C361q21kXWYiN2RP1Xmq9aOJS6pUwKV5hXW12Lst8GvUnxiEl9uNm/P7H84dfKqYDdr/O+0EVoaA
R1DewCa9GczHegNLTAmlsR4t/im7Q0sZvfOf6+/HdEMB+80dfvsohgjMB4UEd3wKYOGZSGWBrQiK
stMgdZStOdvZrSwvyDiEhbRYx0kzsreMPrcudZYUoF7FYOGhkkVP52kaeVcduANJ9k3COVnL6DDW
6w6LvUJ58vUrvTVaI1gUAsQ7baTuYImLtgIglFsWfL2QIaUsXYvvycn6UqwE39UgtLM3vN7o4GW7
n00U1/CWLtX5HYxEB5wDpY+qH2ukUq1PgT70QbMomvDYlhvBMaOiPobBNqhPdm+WzRfSxMDGGo1n
K21rlh/GAysmFlEJ8C091Y3CueMQjulm6FSJ7BA7e5hSO1bcFgMvytHNSYq9RERaxCet6TtvGwG1
PbRVQPpVZnAcIVcNrwD6qKX66dZIeiCT//9i0f8VTdv5x3jHvJk0sCBbdPR9btDFDJPQQeb0469Q
cRZXLilhqWTar+mSB3IDgKcNMtEM+N5RoCGSTScgqHIm5LaM7EFwiIL9NG47wZVa8obctDQP3n2R
PnuBpCo3lcvLjIU6eyL0rwAlcePXIGazWdZDAJm0u6v/iAqaCqFhcYP2wxI1rrHG7xgx4J5KNVEk
LhxVgkSsbUU/6xsY4/D97DoZEjdIKrz1ca9602AxnoW9uNC+L1vbH1yR8Gzsx/MkGm4//Lht6pZ4
UjVgCkwd/xnIQFYNZ6b3q184qKLURgZHugPjAf2NesWbvngbQ+hTA50k6ZgjbTxiy47GDhzWt8ro
cFKwsUPAL3lNKJFWUs6z5SrQDlKltg9G6l5KgddxWm5xUkFbHeHeaYECPAcEHiX3faHNH3+rCAd/
rG2zV0xZiOKEQfY1POIBs5SO6A4zgt85iXo9ojOczQsTNK9fToBP5yjPdw94X4GD1anVEHHBL3tf
BvR4Q1qQ/0r5a/67+4OuTqJ7b/96yzR3RcSS2bRzS4Y2GvOrLcXsNsX9dTQVGKXhzW9RcZCZJly2
ug7ck9gcWB1s0FnnzRQfCd9GvartM7xrGL71coNBfuuqgUIyRqscDekFk7hnf1UuMr9l1hFXfjed
2fVgmit2gB0kh+YE3giDnMSRU8Bbxzbr+DDdqDTeUD3TmP24JASJw9/ahcPsIkYdBA+GQnzz1lBC
8r/P6eOELVpaEpcbVbnjMqbO3sHjBI5OnaadCttCpJgZCqY8eFOMmIwfkRPe42NUEtDkLjKX10ZV
miBpdxCNru84fh6fFvP5EvgttaC3ZzC4+BFRmttflyxhi+ktIdHdKTK9vv+0nONuXCG+r34l/Xfc
wcdXivynl53yhYNy+EPRDPXr7pgBCUPrORUvEVu8NhYREgXmB82tjYdVpioRttai71washpvCz+3
mBlm4S6pbGgAO8Stb4bGvs1ukonRvnWX+vDRQvbotTRV+YeRhUvn8zo5pKtG5FDHdrDY2HPYI3W2
3OwySepwy/sGrfSPQk75Kx9TX+zz+csIZm8GTBGGbTNAd3XG9VmJMsenwm2KEeiHgvXL0XohbUQN
ufzYOZqmU3NoO5QstLyFF5jmYfRcWWLdgQVFbGFXWK9LcKTsPCLBSYr89Sk7iaYfR5Vjy1QGsf+y
fe2Fhz4HB0rNapS4E6hVebeTcQbJBQmn32UtHMb8sG3dFJrtXdqnPtiqQtmxNTSlr2CLCpbFn2u4
JAerz5hX1qJX88+9BYNBsOTHs17qKGGgJJkmvJXYQXKHhqvmFBAO8beEFGKbprURmXilePRbcl8A
TwGfoVclM5ZqjO7G+2HdXAWh4bLHa+VinXbHaKG8gpiP3BVxyqrEAcyfs0L4ewSbqLQ+wZeA4kyM
7tGRG8jxTYXHpJkv9Y2s4yVuvF+uV6xUgABtiuSi/aIK9DBhAusPpinkI8H94/B+T6vwgcv7V8RZ
3whNbr/SgjynYSJecD8OQQUtyBKtl2qeEAZgsSNq80IoWQz5fuee/hLyZYhDiCoapGIcsFdQJqTr
O3onMohAap1pzmZqZfiI8r7r5Kx3b9sUARnMTH+ia4onKzivcHu+3kf166yZhC77K4dXmL5Ev9iz
IeYKX9HE7TwAZtzsswhgrvUUWUJ8+NjyMSEIEmmJL5fVo1hm5NLzSXdpvMu+3mqNsoHrucyvii8B
N2TCB2F+udH5gATbfEFZnfvQS4XDDURQQwsoFyaKmdzRnQskW8qcftRdXLngAGaiJrNdMB2ZPN3R
ofPgDIVcx5hfnYhhYeBChAvvqP/aZwZjgvZ8NrMjJ3pykNDG+szYDW5DtkeU/QFESafdq1CBNy9f
3cCLwgpSnz2xliEsaZEdok5MifXQfySh2A62PbXyoMSzQkKYjbJ5vuuxvd/lyL4EzHQCSHVrxaiZ
bmGNATBHoyhavtXw6li73SmZPL1DcfNeEoCzasoCbeHKjC/gD5pLqsVGC0ScGGLwBA+YU60flP2S
O//j7ievswG+MK92k81fKsXPTm6T2H7YeFAGU59Fag6s53XJx8ucg484pJXwN7BaJht4mh6RqoSj
oBBCJnQLBdZOdVbcAsaRUsaIbNGsTBY+yNe57uYOXaUomGoD2Fhn8koxOBo+TA0N+rvzRbf9sQSj
GVgd5xD/AtNSsEWptgzp8CeROX73FXxRpQ51S3KAaVNgMSyqaF21Sb4vbBiFmkqQ8BhYHFwdaZns
Bs6yclh8FcX/cgiVcZfUkNCBxjsmeMyO7HVj5EpoeHd/ITUmJgHeYa1NYeCya20PtybfQPX+HfPz
SLCaMUNMcsYt/x7jJPJA9R2dy5Z08gRkaNu9M7+GnQZZidrVuHDr8jrLJg0Q9V3gOm7KrS+jrEVY
VTyDyulox73x1wJNpELeBvSIhUCIFTL4vA0ThL/o8koLyLHQYjl5BA5zErM0f40bG0AHGkdRZO6N
ogg6qgDGQNElffEuHC+dVWxaCHZPo9LJGTicBnpEBVKRDi6r9ZlUS6HoNrTXIhjubLplk2u9Gbx9
8eSDLYyY8KziUhq5hNhwQVPEAo/BAlzWJIbnfI4W3sTzcte5GLBcGj9INqHlbgOk4aVxNv6Xo48a
HekNA7xxlk0vn0abb20tIIkKbvzDJIyoa9G78odwooxxdTkJ8Jm9RNVklFuMw6RyXEk6461fdxWh
f3EI20cNEc5IsHSxcDTpDVVH/9qeqQ03PE7LcxExt2mn2oBEosH9fgxWqaLyexHzcHVeWVuGR+DK
Klh7GxalwrdbXIpP+RfapI9hOdEu2+b85nHru2HoC1Z6pGAYfgVZZIZyT9nDYs3DyJehTRUB93e5
enX/UI+rP1meG6NXlchfZvdHsiyzgwKPM35wB0HI21mxzZzTLIB/YTeJKQNTBwc5OXcmDYSv40Bg
lOPfq8OwKlJR0gSkWl/IQ5KsVkz3EMPREXrzko8smSNOd4gbzpKbgP0tptI0q8XJOngRbSxYDLDe
xk4v4vZN+vZlE3JRdDO0mHZLxGoqMzDwWOmeUc/cX9zJ4zI/qVbVopJSaxlfcTj/8qHhYmMaLusq
yDu+mo2OLJGsdhBi6eTR/OsIQDqOyUCiQy0VUZMqTX58+hpqBKYw/wR899TFdhoshypvVF8tWmUV
G7WvQmfkORLI2Bcwf/5FG39edhLgc4qdli2y7tOndjK7SKEor0aQn/GK3j6ZyCaKNzADguVAcasH
V8tgz0rhd4IcfR799kGjd3PhlmA8bopNjNBciVCmJEOXX4/WzS6MTlxJzWgaVD5Snl1YoQwXEzyR
5sm8eubzLEjQiwPDU5yQWETS8MRsBev7xgD7UC6Hp9nLyz0osAv2i0JH84AsexvSDblBlCSTpS/C
fYNwveAa1Fw7sSWIkDLQ/h7+hcp9rihGTznXUjt31YSTTM0KBdXXgZ45gHJg/Rd8UEXZ+GmRq6Gx
GF6FB5K5gOGXBwWmFLWn/LpjHGcqiK3Tfr1u/Y0gXnNn/eYrM69+4GZk4GdUVO7FjfOBMMO4HO6s
5yUNq/jcfYBapS8JNieRyZoML9vwKcxA5niYgmJQHokuNXHs1BStbThn75yK5Svl/o/zngqUwAxl
y0p0saHEgyA7gxhEXm26ohUBD4TJNigJij4NUF2Z5f3aNWJSOYRvmGi5OObJaYv9/uc/WG0hSVAS
DwIkt4fCucnGSYxdJu3rXQhdTuJFjjEKhYNGMK5CHl168SrdgWm5Z9JUHLjNbBI9AFWqAl9mE2zt
FU2GECNpf3hbfEOCwhZT9MwyWEhsccQ7NUw642P6mkHVGZbbG2ZQbvIntZImQsAEBN5lGQrnL6M3
ayP40rX0FY1UjwPMX/7j9vnfQqCd3/cwOJUnn6u9GaNZivb1PEjyD2rY5pLjDoj8Nr1mJLKpS/68
nddGOdmK5OMvy/NJcshon3tZ6KWYu+Nk2cHLzXBqT9xgl9Wm+GkR1u92bVvsdLSffycns2aLqa6p
twY6M8KbdrX79FG3bXFuNpF7rwJh5uDZOFYj579WS+fL9bpkJPv2wA3RTbZrbGNXZKnaOuCkVf/Y
OuV8q6HOOlGmdJVBMQPapW1HK4br5JBOZ3BMcIMoeSPlCPpNzaOLHCEtiSCriDn13qvay+Wq8Z5M
QlpTk5QZAQXEjM4uRENqW7VUmsY9qowL2bynoOv2A9n0ccA0VuVSkRbsqP35aOdJirkjJdOg0No2
wj/UE30aTJv/ysWH8PlwAg0a5EJcY9o+EkC0yRzOsT4vmhJhCXYGYyUckDTlW9M4cZOkAp3HOe5W
YhD1mDGvbfJ2AIEZ1SrqEdPKklfNzsRL7jPfrGvuUmDzqdNoc0ugpZeWYxVuUuI6LhUX5l8V0h52
f2OAnOIo09y/cDHroVASd7R3tokY3vhBfyrduoOCigY73MLnvVZGQDYu8ePdP3B9zAXole0wsvqA
RCGgNR9PsRiX7Xx63xdf0b7FIi6GumSJ85mhoOtX6kPRuQ69jFgL/IVMZMdNoyXaujm9VMgXB+XB
lpeHoxrnUt2/89FBpumtldD3ey/hXNPwdgEwuLgwUh/u9myf8V/NfjOuO9UKpnqC6g6voJLNgMvl
cETo+0JkLmee2a8IRhnKkgvyhuEq7zinv9jbmQP7eeZyPgQYnPMx5+4mJKP2dB/Bz371Fb0eFj63
7UKMbA5Sw9P3T4VY77g0odJsgwzGYRPVbCEnxFtk6nHiMyy/bB+O1mlVw2doW7R1ub9CzXi4Ye1s
o3+gb2hbahH2YjHclvs9IHZvlwD4YhhYuGuhqvRsfZVHq+tgnnOlMZPQmDMitXuREzZJxsd5CIVc
4HT/Y+VhuC4sZYDjXD1st/4kXDbd8KP0HucW8+2MPsVu43u5qJL4A9OOOMr8vf2/GiOKs3dJdMMQ
reOzRiDu7Xn5x8QRisjPEpXhjAKgoB71rpa6yjf6jyqm0HHc2g//Yo37XlBlx/kszFMCPSlJfQEF
coFI8yEJf6bGUkqKbezw+uvJ7rGLq4G84ZQvqokUq0TfICHN3wgoA3vM3bLAZbqOOc0lVQxMRxQL
viYmo/hhPf4jsagP+mty2VKs7djFqxGb0GuknEY+I3UhgsZ6v2xCMTsi/Ql5ySHywqtXy7aoy/ok
zAA5tNQZIg6mDkGRpfg2YHl1Dufv+7LUKlb0loNjIACckpBr1zMJv7IjNla9TTPJlT7F66d0Zuxu
xpYg09SuyOJXvs/UHUNBqL58Zj4o0TI2SlsWlfD8DwuIkBGqtk+HqGoTUJXQqi/PSzCxmr7z1i10
L4AFUNalehO1c9APnn5HDTDgcaqKfT/QIh4IRDC8twS9u4fWOm261ytW8j14ffo3bXf2/uNL5Tnc
gQwAVexsxZs9hz+A4e8Se9GscvTHRDUxyptlPOdK7BsCVqRBq0lFDCUaj9QpNpPj+Is/uCITJa7d
3OV7gjCuBUB4yLvCemLxGidnyB5W9j4i/xwdp58zoqhXVGHsThRs00icvlxfe6lg+A/ki5C6oRbu
hUl9rtkqfiYKga6V6VGFG8HgsBtnjK93Gq0aqlEhoFQxtNmxRGntknV4kpF9Ybn7VlZkpThFvz6d
lJq7ve3AXh585J9Qv1ThbhcUgh0L3eYyZTlppGkf/R6ercEmlnR1y0byf1eCiv75R3GkcfOsRONj
hlfJWXlBI5h3xBvcP6zfolm0Q8vPRDGE3swUCQVLYP4wrrNNUoo7tINzYdFYN932LnDLi6a5IyO7
0XdXqZbI11f8PBDHbJSyQ/yuO/jjg9EBoRoDhE2HunuzOHurDjiWiaJKhhPQG/a+JqBfLpZGsYYO
M1BXrcgvMPnaS1JMefXFFOro1iQBigIzoycn66tyLKEP4ZhJ4czSLRcKAyenS1OaMLYB9Cr5I0YW
vTJIIKh3kE7xf3occuMHDzeVRRAhnkBdDsYGXiEC/5LZE02bdtWQVSNEpdRhRYiB9TsOkOMRblLq
ycSN7BC8FJYwgaOxKjxfTn+2wNWSqVkvbd4DxXYnvR6S2rYbrqEd+EkK2IRK5Eh0dH9GXkjoB8Dx
CVUnBWzUQawbLMMgVSaDf+cxm/iJT+TRHrDLUkuu/OKCHu6xEcXDK3Lu6Le1cVPN4hfcsTQ+EZa1
m7Xd9t7zGeso1kXjxOvPB3ql5jPfEIRqW/Cdjdoa006EqHcHfzNCWG12XKe1r5/0WSmsT4AqTwvV
zmrNnVgvlF1xwHk9FCig4ithfMTTb8Y/BXa7G32XDUFRta3yhssD4ULx/eCDnKJKkH/xkmUK954y
YmCLKamb9+CisA3yx/G41O7EKt+Dzy7fEUgaw2OPtqmW9fZzbI1CcGExRyGn8SkaKK4J6VyfzpmJ
vJroo0Iky/a3EVcz18lk8eNqgmOOhH37CLdrv1Bt3v4WZvc6JKfqYrs8JckyQkb6a+2X57NR0Aka
qAdtxNfA61oljwUpDd3YrB3uV2A2Id8lmoZaWX2pPB/C+u7HjDzR8i8fXnNyt7deJZtv8VAtjISm
z7dJk9PTg+DFzPKC3j5UkFcKupNWCk8rlGEA/Q0xK4ClteQ8pQSvEpONYLnQBlGROQBld1g7H6uT
lPAAI+BHTnPVvsJ4o4CI/TTrBm58HcqqapTDs/EQjmOpw0NKaLzY4+6CT8Vfwsohdq+/orjjxJnr
QvrWYRk6nvVI86+NfdUyqqafGaofpNHi8hkxqV+MA92nbtvXiG4vCyEMg4YkIfxPV0IAXiNpHtUC
+XGBCAOM5Ab0RGuYnpYVgZszttWv5coiApxOHKO7oIBoQfrGLJn/zWDlVHSvdaRyz1XLH1Vk6ToU
z9l28UY515S0NxktCQ6bHRHyIS4Y4PhPvJPB6Uj1e9MRdJe5IOfz2N9YOoQvsUxVFVCRrZuAQ92z
bicdnUFu2muGKozDrhqY0/kwn4aZuuBd8TNq0dtsJTIKrc5lTQ4uQ7q5/KVZFDmaq1fURE9L9pg0
0tSJTqkO8UBtcNF6WpJKBxQOgOxOYs5w1ovE7Qslf0fIhM15LsNnoIgE7+Ptpts+ZXyQzblkD9gf
oOnlKUOJWtoN61ykF77IL00t70W7DnOw2g15uZxC6ss0wDRYjATyIO4rFkpKyYEvDO+FC9rDiFvF
FW98O0TerLiFGBIKOrgtDelKT7KF7kx1ndRP1hyLl+BBGzFziqw6rt21KnmoD384FFzNoM8D81eB
PtACBta2gUr5qR5ko4ANcaiacmC1bMy/isGx49bV+Ki77NIbhfOoXR/sNg4QAlKmJ7LnE5tzzk9b
fiMXsnHzBlKP2QgOmoTxEmN0eF9PM+Owjt6R48lTsh6gEnQ84eHIhrTf9aO5xsBxlbwTJ155i9hK
zqcBzVAWyZwEHPb2A+SxaZ1YOcgOV1xQFmkGrkMqVCM19Vuww44Bg3mT1KS24OApoZcwReLyORsn
Q1vMEeNdsHhn512ibLGDsFUDTno4e0FDchwh/8PovexO2JQFSSGfIWaKGnH7rNikQycROn3JzAlB
W08KryjPUoUjJGFdtXi13w8lO6YSzY11ItAANqNzmItv++RygNrtv35gu63K77h69zyKDBI2SDOq
+0EQVDWVnzKJ6a4qmxG742YEt4hRSw4eUVY8UBKKIxRM95q7lVh7qUxYooDeSC6Too4p1anzB1QV
cMewyoZ6B0+4qsVBA/1abNaph3LRiR/T3vh/wRRSWmZIfvJWm4Q/kYyVynqfmI3MEcxJoVO94Pft
m25L3rWnZ0zoxcDab1JMf8mElqpKMVTE5a+/IusLMU63j/XzNu5hW61HD2guq5r8nJPZ4B5FyPJA
96TwyLiwhUilBO6UrbkGfWAUl39jLfhtw+yuAZ4xLaII/KY57IuaB4Q1qW23KDiYYjadb6f3P7tL
kdZO2yGsw107xqPSbu25dyYqVhzpNFN1M3Fz0m1xLF+DAKTr2rSYopiB32zR6DghzYxn7jnzHnXq
SYZDemdwewBVUR4nh9h3hqntzgboie5l0qqcu9ncx8baxXCZsuzw57u+3m/M7e8zXAEtGKZj6taV
mVh+F/h1aqnThfs2v8YVkT5ct0Z0yZxhd/f6aBza86j7xpemjPt6YPiVVvhlpjaEdCDoe806TaRy
QTimGSbNVyRzP+jcCl1avL00P0MsB9RhfiE1RDSH6hdvN8p+ouZJLZNAl+jLUgZwP8YD0WeMWTuK
4FAan15FRNuGgvDaGX1ywwlSRSAbE15mI2lyMy/qrn7cfdymYE3DgcvrIfA+rVoeE+YRoWfEHsn8
GzjPmxYjbuXcSPCMO7tbYwPGyBwGt7ZKxzL1jikwIlRfRGkcyLxD6Zos5ps1MJk+lscQDSoxgSkh
qjyF4oXmimy/iFrdoqJP3ydWldYbRErwCAtRJAIbwJmkVU7hwuO179a0zHX/Vj6pItSoqKR/sP63
/6nnbAyu+Ii7zahObVhDasVmbLqe8iD60oxibLv44SNJ0gI/IsNL4vnHLlJnaHa2VhayxRxzUw6Y
bdY8GDJi+CSRZlphqV2dh9JDIcldWett8s849tBlms9/RnPaTd9kxWirr2LbTwaTBbb3lr0rrtxo
gihDdI30WsIkj/8uVY0KDhm3opn/qiDOPHSTIOqRrvyeVlX7tkNcnSdvRcBEFttWSw7ob5CWgPxl
fJqkolNBlADVrEz4tUXhFNrB+bhpp+4Bm8PyGe0WqrJpitSWByqnPMPPJ8WUeHGJIZ0RPqd2ENFG
lCTuGXUsFvvtol6oKTc+YFAr5I2TMd1WfUwY/picPPkoLAssJGa72HdlZ1J7YiNDXao2AYgX7KD4
UkGmASmffT2KBp1Vg2yFnQuM3ZYAlpjaBWSXaadUbu26ioeUueKewmA//Z1h/CyDxpuyMfTsisa/
pblCWVblvngiVr97aQL79Nxkhs08ffiTjmVNUgzO7XLNPSZWm0N3P1s6i7bhz0wabTuUMucbmAOv
mjj8P9VqC4ltE2FlbYlSL0kEpAUf8rRyoqY/JJv8GnA0NzT8D18Yvvvu+8SovCuoE5urprjiq7FL
nf4BxAUWYLyL1Vrc7RjJjhn0Lp+7kCLqeL5omDZWl0iznjqwaGe9UdbePdyVIWHDm4cFz1Uc3nob
YWaP0WkOzxmzkx43hOu+6PZ8ZlvP+Sxx/g3UEfsNv9dtbqJSOOnhamnQAzqsneYJ2bcPdgcqAm2U
bBhLRVR1oVrde0i+T38/jI+pLY44O1GP+8tv3SHmBcRnVKZo2C44ETE5O2yKPyqSUlUd6iSaZ13A
0VL7uTkEAlErFEDY/Zacv+j/XH7O7Q1COBbzYkabQUs2Jmnl+yLCcch+YMWJDpOOfyUFskI966gn
Zdk++WRM3KVnvOyb05nCJSlbijyanqYgUTJ3Hi9r4zZHXXz/bg8O8MfZ+yYdZkiGmdXtWQOrHXmf
nuVbC3+XeWa2NNz6QQ7IH+bxL75sLLnoa+Iyh5XtadM+fK/6upvm9n7J1EQaeBYV9DrtFbTHoqQQ
/Yfrz+hS7mwmk+DIH62fsHvIChS5YPs9B8Chij/5eHQA3M1D2f+ck+RoBYOnx5QmeZ89iyrDFBe1
q/eJwlcFW+PJbhru+Chw9EGrCc+OqRZTAvUwyYZVBF/7TGcZwZxjfFIQ/b4XKlOFlwv6elrrTEqb
5j8IWctu2W2nx4e+yepItW23yJEAF9LaKEmKN2oxPAUx9W6hzXp1A9vNhBpZ/bf4UkSCg3cv3lQl
YJGqBTspUAd6qSbheO7wYGIPeAlc+8y8vXPxAIZxSabhNkjLbhOda3lrYT9pFR3m5F6DQVH0zj2V
KmlFGsivfw9+0iiQb6pxcb1aVwQNi+27Zu+y3YHXQOABVjK2kmmLFSWSyZSpjeih6nvOGlpgPNKW
EngvOcuOTFkqfUfNS4VfK+8IgWn671dH1xRRXC6E4xSOKvqzWQnXwK51Yf9xO1Ok5yWzW6vJ+MYk
TFpz81fDHruJb0L5d1EKpj+9hpYC/XehJLZuet+sqz8Xjm+IKY7bsQUqqZ7XfPRbNCFBaI4kokiF
aw6QES4X5AQuT3ecVV+EG5Gc8+22u1CqoIsbxp71gcIrr6MYoK5uIXFpgviURr0OYKZYl2vkWr2t
6+iAS0uGj3ZsbaLc3F8IHp1KcBj+q3wcK9S9170jD9NFkgfgXFZG1a9Tr/KJDpuV+JaoItHeFSpb
OgoYUH4rPEWChg58B8piKZUIRafcVz3SffwuWeqYXMcUs1v2cGTsLhqRIQPMgihRIsts6cAQqwjN
+k5Zk3rfmfN1sJozvifMxsQXE8EoI/GLMBjIzfup2RGDum4adkvxz2QAuSJSbPf2tU+2toqSPDgS
YN0g/75Y3tRm0R9BbdYTxwrBjpn0BUHMK2eJIO65pRApTSmCbR77n3Jw6tzVWANM1hNx1hggbX17
dAgLcbRzcpKWP0U4YufTVZfp/XOfNEcpcTJtjEgJTcK5Amsr70LXlzVkqYqcEMZfWxrucVf/kEVE
29OXzyPDFEiwfT0KWd2qFsUq8JWQ5n+frcDajWRA7sM9dEj/SFeVCZlaqI0sG3uoxZ2PTTqBaTD4
J5Mmg1oIAjmsYZ83Lm9hUf6TYJuzYBQYgnJ0gHYWIhvdYMSyfogNCwrDbkuEvoHN4uvt5jPkteeS
79f5UuIcOl/Tyw+ZixOVZMm+NMytiCkQmjoz55NTzm1uIiEvh9sqvMBV/ixDqH9o//ZAev+ZgZw2
i4vSSsNDf9qoC3zl7enCVL/6qoEiUQ744FMfNdA3NBAEQk6LpnR4PETFpDu4Y8O0p7SciyhHQaMK
DQgk1oHE8id+ECDiwYcyqPFocasaxjG6dM9JlBKrDuHoiO6tNEul72TYeYlGn7CiKuTa1LM6vxBT
ZNnK735s8XS1p9vEliLMKXwzHOb7NEk1XjnwUnYa3y8XKXlZ39PfRvZkqRyCToUt/s5i0jUDMTCo
kxOwUpWbn0f/kRvq4mS5SBcO16IU7+poJo5jU76kw7AfAJu45I//QEb6YQTgBu7/lf9o7P4c9ERr
VyJASnd184SqcoewCR3nyh3VCxdpq532Ho1WzAzw0KIW/kH20NIlWNb3gaNfri4lO4j2JwdMgsuN
geHsTp9M61oKJGfZdQqzaTj4Rhi5byTPWSO5zAVodJZOONZEHzYAFuZqL76HP9XjDGskvXZgqUXD
DXJkVHNwf6lzUpChW3KT2Y6UMFG5IbIoZOeG68o1VPWdz5VTT0CEXjWlfgTcmehls7z4unmswGDF
5zFr3Pp2fKf3bfYWuV6w32Bc+d6vq3baDyGx0xHQAEbh5GmyNzkOfpq36BZZZCMoHB2njCoegjLO
s6/XrZh3s5xU3bZ4XS+MoIrqCTbPA08wnBxWAPaLpObWGKoiG1g4jZiZgZPc84KbLy2b7caOhJmv
4KVBha0llGQIbUmswze1wJDkr9fffwVzqfeRx4UOVaTQjjX+56xkvqTQFJplHSRGDuzP9plLFHdS
OnsKANEOo5MHBftCZMXrKO6wYLIdw+aHqOBqGd2/AY7DfVm6yRadUAJCxEW0CWjjqbuCy/NU+7Vf
AwN6z+l8QW1qE+DLV1AQkYgFvpk37Bf6vqRhbYS7Ljp9HvSjSpSVdQszB22V6VAZGUt6zop8nuKy
mmdOvKHVzp0M4CzJ0QSYJ3hJddLhCRKzs9KCF48iLjFmVp6A8bC8Y0uxuuPeYPK/FYu4Qnomn8i1
ZAvQKeAkETX4M1f6twl+2nhsDaO2jmaslJ96ZWkjD917x5EdvCIVCpXfxo/omx1BaxGM7Z4ViRxv
Tlg3gzCqSb1T1CiuL2V1iZfTprVpDH7SzuuHpHz9VsLF5r+sKke93FoYxCfIVyQRYsq3FeXWCv4y
X24XRhesEr7nvLxujdeY1/j8SVAFeAJ+qJVEGqRPmIZE2AKwUDkqGzBgJOD6mLtuEFq+DO+H5nIT
rsRdDAtiiflqnI3KfByNoEqJtr3DqM5zhgyD9iZvxQO8yz32AI4zT8TaEp9mWM4CtGSlUbpFTZjO
VQh2c/ri8rfbCI2Bek/BZa3BCD3ck81TWpW2sQcCnGzNonUZ8LJuO3OnOGC91hGm4ZGipiBpKye2
fH78ELjqHhvoR/UL5/2wYR2nJEjcdzOpPD56VrAd6/LoRhcBufCxcroaDNTk8rxPuzwMV73NLyTO
HLplpIDhNBcFDQFLwIhk2nF3YuP5Oz1V14qKqoTxRrscYcc45DMP0HWDb7aU+NDqGNgaBxn6mtld
2xaeNdYJElFfMZti9CFaZGR+EcWdIGPFWDFDx6dpqsCQ9ahp0nbN1xm289OzSNr47AZu+Za1PtzJ
sKVBUxyE+NvMDbMF2xhS
`pragma protect end_protected
