// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:56 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PTeeh9+F/QkSitxSp+ajeRBDnTBNH+ikKsSjnO5X3+wU/iiz9qMNX5jf7jlc15bW
j0XncS37jvf/oZIyx85dPoY/Kt+bqVgVhCd1NByVUS2HmmqXjnZxzGK+Lnx7w/YL
nWg5rDuR8jaZz7hQkZc+c+0q0ls60CyUQtjH5onvFzk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 124784)
T3n0mKgGyxGEpObhz1JeAFNUnvn0xSBH6tJ796jIWRppx4URXU5DQhqHudP8qoaM
wTM+DURe/j6nEF+QfmdmWO/UJnWwPl/RnMY57MZ1xTL/trrvKnnDMSUiVNDNg2SU
8rhfFHaCjkmF8qhZLe/0Tbr/tEE/RDxZQJvhqOVhsiEGzevE1ginBFE/4i/bKyyz
yEuSlIOdg8p4435eS/rQ+EfdQ2VWIu0UJLgn/uP/iuf0xFe3Vv8Co7mApfu9KWyJ
aicQRASc774TmEEOkjD6Xfya3jnPPWq9SO3GSp8fXMnB6RsI82GWJi5P7eEkkBzY
kXrNyQIxqQlegGY0WXFd1LgUzbaqR760N/ATkillowGZ0NSmgDCMq3j8zV1LT/Ix
/I0nSwXi+XZeT5PVPGbA7OxXZ8j3Iky6/V0AK4RkGVaSaTX8T+N8UzcDze+/MIT5
NaO3bERyJad1nHPWRGE0smieZiz5BzyHF89D7l008wEU77ONOyhWWYJqzI+LkX4J
+OUWKYkSwYYnCXnGSFN6zmNai1P4p75ot/jz9DF/FidW8i1NkOn3S4Joadf2U/eM
KKVvhhIUF5PnS2J5FFARRroX8VaRUPerpEUt/GHxtR7xGrdKjmkotjPygJsMvgF4
zWDNHfZVNddL3jlOrd/94PXTZokKnxYpcevUl1lhKmgkOmFFYgqxzBr5bv6eQz8G
bPmQkYmrkTsKMiYN2gZX5AptF9DBRfCLD0nrk4pbZQKRqcaS8k442DSJp4g/2Bxq
1H5LodbLf0Vngieowp9L9ZMICAnZ1SnuMQYnLXfqBdaDKPKUDwyhCpFO8VbGQHl4
An9QFnreuwB0VjV3rXxIjHiJHvh9a7z5p3x+BHVB58hPhFNieoky0WZMC7BGqi1u
OvoWOMV9oXwvv8M20oe5kyUa9VLKWYPntG1vdp3oPOiZG+pHFDahh0uQd+vPj50t
O7LS0knHjHv6oFMLYQ3H5QX8MNeR9szDokKHYAq/lInohsPPRreY9QqijBOszukc
dk8YLLKCou62NcbkZzLU6eu1HtfeZBwk53sOoxeBccUhNu/+O0TOKoWQVQn/nrpi
UjrSFuRTRLjP2yJ5G0jV7d41Rt656yDRQs8iVlSxpu1AAgUPZ7V/7qhC4iex6Fa2
fO+W+3klxYVGVtbg4/H+le8KYQNgJw3LSUdekhduh4mpsh5er2K+sd4QVHyIW86j
Czz1O+bLTh2ZUdCjzZ97JLPTJ4kznyFE8ypUfgFE7+kbgjyg92J3XUTq2CuwPN+X
HZ8WTSyVGai7K+miwPqwuTBMT2kdOw6TySF919QAj0PN5TxGpcio/AP8xEtAWQaw
5fTLa2cXbO8vOQJ0TapmI9r0cesvC+KWZBeDyUEIA3WDshoSQzNvDDG2JieSuHv1
bbxl/ZfkfH6XK6KZLNOhjCvDH2CQanLVp4ydKrBtrcyHwohqtb/GDyG7isp5lE9v
F6v+tjzpnZxJpEA/zWdELV/e59KLpYzld0D8I/u+rKxBLDViS+78LD+4dTO8/HqP
/sgYQPC1Bs7pQUhVy6s9GZ6wNeK3+O+DH+u12GUN1LPNtFizZCNnP3i7k6gFpPEX
xMfQvgWjXpUXYLPMYmJk/EfQZt0IX4rs+gpwNE2KqU3GU+P/V7rc8iUAR94Kbjxp
IVhluw9jmyYEg/fwsKzwp66h/4vVwwV71eFDlHFlm7oPjR0yu1+oVfiSxk7FQJPu
9aJN1Mp//IoRNtBCeSGsflLDEBc2NJGXsT0AB8DX8EmMeamcAIvskbv6dHRMQ+68
OKLuoPqmGNF66RHHxJJ12+N0j+ro8WDb6/mrYVNhdg82tQhSfRbThYJc4EypAf4P
7PEg0eYp1/sF2PUc3rBfLH+O/J8qpb/Z+YoLaJSBv+yyIqxVbDh+lIO5Yx/7GGF/
rDUVXalVeHdK0ksc7+9CjUq3KPesN49Ie1n/a/XtOp4sUf9lhRoSwga8GVrImGGu
Gl2gaEmArSUc8AARGTroURN2XOEhjNrZwLx59O4vM+wX6Vryl1RazehsWJYZHcKm
JzLhCvfiscubgY6FSt7/ipqsmLau89RAbzcr93hK9zFkobFyrHTUiSM+t5M5CSrf
tR/4q0Nqr/rD2m3YZ+IXSt9dZi9TRIIWPVsUf9gWMPrtl4GxgpiGPi3xqa7HCOkF
HFrBezSkW+OFIhPKP4yQqX1l6k7qBiT84SIgFNq9uY3Sid4n3hNQpQgPjzVGq0Sm
qz9bEvTteO4aKxnthr7GFjuFPnWiCg8YSfvigsVw/OE0IkORU2reYb6UBXNnSeXL
yBTjafaLJTWD8hHPuBEh5VvLYxtbSj63uQUE4Vwk/4zpPUtJGQhIvblJK3c5mCAQ
A0Zaf4pzFFuG6LyYaP6Jfkv4Mn0HwugYHaRzuK0Mjg3MGwkCflc31z/rHGUQRFv1
j+QToMkf3cytjeXuiXPvF7bPd7Co8VMh07DPP3M7YRacVsR40u6PY6fMsmacmBYn
QCFn2BgAFGX1GdchXnXEfeClCxeJrHEKCwMSAZoisAw5HegvVH/TwCRV4seOw1Dr
s2Fc0kYFAuuUuLCVo/19rbM0jFvjiwtzqU56DQEMtQ7vZ6Uu1FKZ7Dt2BM/B79yD
rDpCYPot+3x4p0XdpHU8OwwJq0kav5Q46S/kXxVicfjmOgZZUbsb56Z6sfvG61ib
m0cYw3dOw/kBloijUZxI2uMSaxJnekWWrCRDNAvl//olHjcAIztmyQWQxXq8B7bM
cOTdrk6JHLEGOFISq9b/jP986X8v95GO41y7mc/65OnkiUIhPcCKHcM3GwK7bqn9
Nv9IGMOZO5W8QQXVukackOFUCF9kLwqCjPQdJf+ZWGalK/uKhRwg2KY0xuDWeBx1
ZvdFt9tMdmgfl9xc+spVVxTD+e3vOmd2VwAqiGxWfNdtO8hmGY2fQelBM2dPXOFe
eVWwL2H99KZ2UJrtmoNC+gbvFYbwjF16UwqGtKDt4eXlZ4jUIhTWj/xXgim+AGNx
P3G+CPsOCAmT2tzwS0rIW6Plgm8kjYH4NXcTMjdM0qE+7PVMlHznYEKFYGeZf65t
vdD44N3seld1xyXLsWQ9QgLDX7xADdW+2Qf8zZR80MFWkP5nJQI9CvsKkoOyWjt+
E5UZzvwd2SEmZJNvNSo/p88ChqqguLUgpqcLmfPqPdwpVIuk+4ePlnz7rRmnbWu4
Y1iPaBFWHDhBGCbk+uX2aXfVrCbo7IDpp1JJeFcZcDAArQVXJ3EEi9lHIreiPjBs
4GyKR4OMx8Dlr1xNHU5EySYxawyTtEDd7sjJBXzC9oAhRPhlM7BRRU/fBuIr5qxv
oTGGQDtyZYhpaDzo9aPrRV64xz8VZI+KlOP7Zs0KASlu5AsqZlJguWQ0YCg+scbi
sftY4crPsS0/zHR6wyDucWH03D8GNCZSeXlQ01p9tdtzOHpTJLatdrzzd0FRH3Fv
GIW7cX5CNpIbVd+I6a/s8HTp4KErQpYDxjxTMLLsd/mSGnIq+TdkeV/1UsC25k1O
4MwAjWhb6yd2AtRzr5sbmUjw7o2Tp1ZvcemcIC4MjZNGIPtIyEu+DzVniZemqtK9
1KA/3F/yQIuYAmtYnl+DEvKUeK8TA2yRIFscBJGnYwBTB1LU9J6AfqBpVxGrym+i
VV+rEZIIf33L6yS03Q7IP+c/SohOyVADLXxic9HoGPne4PorPl26U5mmHjQVCPZE
sgdyBG7p7PCY//0QtTT8SGmmrfPB1zxrnXAW+8/GlU8XQyyWGLk9x4sYrdgn8/ZZ
y6E7RxTlZbQAJ8bnhimmOymRk33fCj5KZjeaqgmlE2h0VdcyKYRA6wpsn353Gp3m
bMswRWL6fiiWat9jARzzqMpd1xp9Hp1yskZ5kBFyZTPgptudP6WT1OMyXAxHtfRO
hOP/j8b04dJP7h6L8liTUFV/lhWBFyjfpL7Ef0J0B0UdpQkOTmVC8EqGotdCfZ/h
8/CxueVHZgu4vB5HuneQBByx60OW5ipM8Yz221t6WQBDkn8ITmQoeSsADQ3Pc50H
fYe6DX0SJhOLN2OfnQLfB+zegwcRFJlQnyix80TAvRvDNHquWGK0ca3zVBBf1rse
DQWOVGSBToyj8FlEuW+UTUSs0T9Vw1fws0ZEawwz8H2Wn139EPkwiE8+UU9LWIs7
QqpWFMOiM5u6KLs7YLDyjpg+y1mVQvNPLQ714qIDMSxdBzbyYL2o+2zWhwORRfOe
ypU3iswbVRsbA5SFR1PPxiXRXNstDyxcnvAOPnMZaoWcsVOmBpCn1D0BPrWS+wjM
7RCkQSMOZKnqktU+ybR7Z8aNWPy9iQxKllOWvP9K/2DTL75MzI81WWatdPgy1tGi
DAmIUfO+XESPyuwHw5BiZTUie6/ssEtbphx2OdHSJuHbUIJugvojWPgs3eJTxA+N
jorIqhy+yYn8TAGbtumiaP9dLAsqY4xJzhnv8QeD5in5ATVJELI1cMosdVIxlMGc
WwAW6mLyJ9Ccd5SEZjfw9NgBOEGdQrAypJpO2fMJI6/vxq5WQDeXUq36vkZDGJ0X
Vn7sxQN3wBAnNHN/aIw7rZiowIz9ux0+gwagMMp8saLhQE+gDD7iiZ5sZGgJ7U7a
us7OdMSFB4ZrrAmpcrmPSVlhxthZV+gSIVxsMGvB7G8HSdoYep1BRCp8NaPccSe/
ydPycGKLZ8Hs0kvfqINm54Id9S32xn7874BZHdZEoWmAJxVBHnsQkjog/S67OzyF
wxdne91Y3oUGpUZYZWQYkoOMK1mYHaHPL+tfb52ce4uyvE9esc7f4EYcGcm12dYR
nTNrI/48cm40ClZ4m0Su0AVLqwMSq1ZDO6C40DG/5yb4OPX3TOnUAIcn904zM2Hw
xMu8ewul/ZotDslNCXT2Uz/yYWx1IKH/r4LHPE3AarMBXqKvP+gXCvtFdpF4dkb8
WKR3Hy0OKDhOrbf8XxSdKW8SmFVbhPs4+PgiDs6N7eS2qPn6lOyaA5pNdQv69YaZ
Urm9b33HJSXAMxGRkKde3y+o7igRpJQy8y76WiQdPBYplZamZNtPKfVq0eVb/tOs
KPVGs61yIIqNy1WUknIEZlLE9m5guBUnnrKHSE3EDIUvSsZZUN6agd97xsifvlWc
A5m1RR9PWEAN8CMQqJgJ/UBwl0sUpEBGAU2LzKjlgULoNQrrp+iGjN6WWdCKZAc+
bpEFaPou+BCYkeAm/I7t7LgKnkGkNZkTU1Pfy3HA+YJqTNL0mFRXNaQMlwMAh6l8
OAvaVu3HIgtQcA+a+3JFAC0MMzxglyliJpS2R5wv/4FRux7tk2ZuaGi8c9xIZGkV
nbEq0gK8+V79KkGGvRQaQe+gfYDhx3RieUeOvQT5iKj9AdfJmJu6aT3Pd3iQVlBt
ms+rn3k9qRTwr2BdqpygM4b/2Z4vhhZ5EclhLqMEQEeh0NqTaoUeNUTNhkZ8sOqZ
86Y2blbFpFYU8RRuiKDzE9Vnnlh+l7lP+v9XE47kVhezwqqHxrNMQzz9ZQ05X5zh
c9lOufeMed3M6tgE8KHGjmPBbpdw9HCdUwqrD//7gthj6gPwhY5emELoQ3WanUgC
4Xlhfn3DwteclEtpSPi0cCf7L9BRMEEEXQ8l5pKVMyRAVcqzwsxg5KmNVAf4teuV
rT3wXBuDNwdoVJynJteBwwt5BKLS4lgUglmT2AXajpXu6XrJSxDdP4qnY7Tw/490
ZW/T+URuNx6nyRbiQs8DzAcPtzcFH85MwxZuAkJzkgOD1Vg8HK8utGVPlpejrkAN
EeFPDoPqxQ6h/VYzuX1BsFF3yMvjSDmVlJAXtGevJvfJTgT00rrLnTej5LAzw+cC
T1m+5nMeaUymgNLNptPP8UI1OW/+Ve+LK0rxZZPS3oQgNhyubfhX3fOHzUMLdexw
j4+Kxdv0EPWX5fO4OyR/VQxWB9M+0M0EFBmuptkbqsd71SeO1pfpSp87IzJXmjwA
06XZZ2gvzTB+X99VZ9iJat+0iqHY5RVQYPQo4LG2w1zDyKow1jNCUP+ePzaUaG3a
iXTqAvkdA+mZ8SXCoA55O/ykISwxFJwQgiyiJxzjJyLdltF/k9D29Ufzd/mE71HT
IO88HUBuHaApJyECFtyx8yxwdyj2yGKrvemNnqo+8OuPN62AGyKXHiBYzH8QgbqM
Ew9csBCUmxFUyYXFARN3sHzbUuYpaTAxQb4MHoxJL+QMOkZ5KJL9mLYFRpDDlks1
I4ePvvuHMgJaDI8+FfaGyjfI/53cv6yR9hy5FuJUrA/vPurQnUMlOtr7S60D6AUN
iVfbV9Q3Z84qXXQ1L7tR7wp62j+ZGLx0ja7Wiq+u6fWmBhNVkGyF0Yin2uulGEpM
3HHIfymnq0FYhgbHV4MKHqY0LkzA8Y6OvJo07z5cr44xYldFgsUiJEpqUeQTbuhq
lh3xsmcAQwytQWBVBjbWVh92577DOvYV8AeUsgwwsVmD6hINJYh+ZcFA9wYmwHo5
lN7uyRbmk3476S2uGyLnujBiIYt+zLusJAGutO4tkHzr2rYCcMaizBzAsysYRxvS
LADNRH7WZi+dWZC8nuVBYzLvs7CH6TrkYpaH0zFiTpbUjKOfSbQDeyS27PFZZZ4n
lNJOTgezgWU+vuYHIW7hCulsDvJOj2LilnZjasfvLO+axxA3xagVkSk5Sg/xj7It
bjP9fkf3OxCwywUWUwVl6Y+lai5+/4g29eQkG7EjlVBc2QvRNkD0shDn4Q6riHmq
bDZ9TDnvmWEkQvqVi8H3t6xfxXQYQROg9ZA336Qi/9GTMxpMlSAIDV4mYaQOv4T7
K5fbE9C+JkeDYFjwmP/9R7zlPX00I+P7rUoLOb1ezpREvAgR1hHU3LlMcG8BRoCR
/5xVd7aOiF/Da4inIrO9sRybX4x6d+jsDRScL6zZZhITiXWGLpfqwGa8m0XUzwFa
0q12WaAMw+5MIfsjDn7HtFfj7KOKPv6hu5zCNOcitw+X+cszE/vsFzVkJNnwvm/7
hTNLmax4LSI0tbKimdUXD61PcMQhU/AO8R8axLGEr8j2p07S7R2myzOvdgW3OoMi
qWlLfxR67sc7kPrjXqwZeUrdK6jZPlOCEJCoGFKVY9ueWJfwTDrRnmVVEADeDQXD
3bUzD3+5VMZqiTYVp891Anmyu+pCYY4f/jIVJhrxnr5e4FaAHeZ4tZT2WLM3VYzZ
pdLiov/S+fxtpwFTyGhX4CtreZN3DnH/fQBoye4frW5+PXarucdqYNLnDcKOzurS
FM49UhZOtfed7AtNnMCKQH5KMZ0dtG/ahEKjj/AO3X9BNgnHfRatA3wqwRhRVZsM
gX/7qkG84uyxuMa7UwN8in1+x6EXig82TI+GTZ7EJzLnW9q66kCxkvmgNB5q5lej
FiXYrYx3Xrw4JUCymng/5oQgYDVl8ZiCeQvK/1uykzseNQqUOd7BFzumvLC9Iqer
11GoCp39TQ4tGcaVF+3tZJFmaUacg4pqwZ6uSsoLY4TSGVUNdIyRFlQZ4qZZGGn8
7sXuz6YdGu9xxXALttXHSakQQ4KZFnwnJBCI0n19uDiodOVNn+rrP21LFUUZfNpz
FNCzE8VH18qehmglNgSwpEAEW3jz2FuMzuqZ/r0AYBw5dXAq1B21aXz/L3JrUfPr
FsnFV+s1gZ1MCPenqu50b2Ow298ZVxTIoeXIkPRC7o2oLwwf5Cmx0DWOrlt9MDZb
py0VfoMNd7nj3RZMRRFy7KZGY3/6OorgUE2bwWp1UBmnOTDM1m0gSVYHpiWVnFSi
hxNks0NbIUtUyz1yuZKE9jSGd7J989NUeWouydUlk1XSilNfJ1iMuM9x0314klT1
pT7y3fY0pKqDgIUSwoNTSKN7dRQHKVruKTxDLWWnt/nAysZWl/VdnQEPenTqdnHn
3rV8kArAPi0G1/TCOA2vKbcXVTP2m0riFSJfQaCxWYee1gbIl4y3SoneTQIfKNw9
grrYjtX7G6y3EIvaaXwiw00UBOJMZTXJM3ikwtv5Vosa9q9NTIYLw8oX6kpCUYZm
ruC8iYKMfcOHcAYRhu1bkfwLBLH/jtiibqUzqIKOLlIm0SYtIkkeq32EyH5RxaFo
7yelotj0Bk+5r/K+jqrHRXLYHRqXiaNAEFopVwVQe4nJnXNZwGix93Pr77QbUYD+
LOgBB/nmdn1QUFqVcMTUT5LMXClvGbcrM7Da5IUZkGWP4Bb4FDKCzbwMjQYa/Q/j
K2Cfvewpz4SJRJWWONM1Uzt7HhjFEGH2c2ecBfffDx+Etx7EIVBPO3tHuRNaV4do
t8UsZs7cUjwiCwrCSFtfUSsQskoNmsqULRmTEz+fJai+JgsgPSUSOVWteBcYDWqr
YR/cGxUIVam+AL8hrqfm4MMQ3MPYocUlKYt/3Nv18N5ec1yZwXLUvnRfQuTiL3AB
lNL4LRxqg91tKi+5WJdQvqgCfp5h+5dkZcfQhXooFsp5G13ZPqnTRdns+LJa5ETO
sgdz8pL3vF+CxEpbpigNkU6qqxR6CdumX8Tb3zbq/SnPJmsWJi8uPWZCPfUQzfin
VvaLxQ2IxVkgvSl6z22DmS08hH0q/+PTyB6Z/qcsL5K2UqZYxUiAs0RKGssmWPHW
BJDLzuwNT0Dt7mF8QGsNHkuTYU47SxPsGEjXshAwkKbp4YMzTm6UlLPxsR5dKwuy
aRVcq24ppM7vsRli7TeFv6ee2a6l5Exc1Y9jYNoKtWfS6gaxhggZjGvKM0z1wc5Y
MO5V3jNKF0UgFodbHdSBO1KSk3NqWjDpKkLon1Eqeijyp4pjsYWi4fwDuYucDr3R
NWAeVn0lK/eOpTdHl3BD48knJjrTblYbUDUNcsPtBx6vlv4B9RAeOjr/avgrrrlI
WkvqYewuAMuqf7MOOqqAvX0AZ00dm+H7nlp8w3c9/aJofH98AZ+22zJRgu67uG1U
XI3KaNnFU0a8BYnKlQaaxG/9aTR5isfBUvs5sgSOvbKh/WCpWrO0nU8V1BXxk5/p
CEcIhGRRuyKi4oi6QpTi6F7uDiTQ4VUtQJWi+44ycT5wASZcu/5bynNSB2yXU+Y0
JO+kz7wqxt16U3Bkevgiqa8mBii6e+Xw4i1XE1QZHpQNZYX75jzTZ+IDjU2cqT7/
WPpnAcBHbZzp2sr+AMfILlPLNIf+z44nb5rz6mYv68va5AYBnzgXNKNRE5M2omTS
p2Ry+rM+o9vcTSrYY8ABJ+6AyQkWiO2p9D0Waw/k+TIADoG8OLpcQw+vymkrWHUl
Wa8PFyMdEEfkfTfe3T86EkkEIXXkjfzM6nmhhclha2X0oMzBF2xy5pk8SJL6QpZm
AJ1yNUUIvmmM1SaPhwPcno4Safiu7ZbANen3gLc0ed/Z2UztmausKR9HxUdiOEpN
UxDCVrXotWMXVW/wHIf9KafDXMlM5OULw2QBadCbi3JRbtBqzRMW1tN3O/8hNXN9
KPnyy1XorgQXEM+FfamqCivY5Qfy1cfzYCu8SW8jQXD9Vi+pGkqXuAHtbTGiMNXc
sPqZ6LGqdhwSo9Qghh1B+d3Nu5he/fSk/A3tGCOwLMEAbzLIWpG0me5KOpx7E5E3
lsEzOgxJThk8XekbY7maReJMp+7nZx6mUv8uzg0IUKxV5d8ecU97M6oX6pdEjrIM
q3AkDOlsnK7YAOqkil8h2CJywrcCPxPPXVEd69lvlDL2KMlahpxSecizVFNw/O3G
Ju+JWzqm8nSg2aOv5AyoCIvZW2k2pspTmVJUc9c1i5PNllCdq3WymqjVLxOkdevk
KSOibRB5s36pHrrF6UBLE46SL1vdes255FC5ssg3k166Vd1aSlrnR3sB45ua3HgS
Is0Pa1UdsQbUIqkSwWIxZSxeyop+Z5ySBvETVAwPHGuzhxuW9WkRe3KMDVELHe97
fn3Jp6IPpRKvd3F1jyvLZQBpyd22qnXKJhBLTQBvjiF1ULbXhzMI4GSdzVtBAaZy
L+l1+uIeDAGcOP/vHxggUD6JalWxP2DqfjkGmC3Ha+h1kz3f+HxBQx6hUo7wkqNu
lPPSVfoYxHWfU6nmy05sMKGbAg5UIrOhCGuf6VJ0Mu9Si9zPmq1N2qSajkMX0eHS
dkQmDVDFlEbdNZVPQrrbZqjzoA6o3E9tt+KylfCl6ZzYahOfTrADV6GC5z0Y6EGm
v6cbiLJ12XRZYnCspkiTz+3IJxz017/SIN2wM0i4g5dJoK3Fe3qKA/cCxPUBhABH
/S6kxSI4heIhHMLyGh3pw2jpCPTSVO+xxnrrejHS3JSh0cJ3SPnAR3koifa2Lie3
4tYXiu+54WRmFib/dvAuWQFWjKlAvXIKykLqYYiVmBZ+rF1/TICpcBZsg5T2KM8d
EAZpowz5fa7f+/HnA+DrbCl9DrYqMOQtLv+PUC8Snr8aA2/sQgyKP9LlGuG+cMu8
NIQQBLtWfJdnABejasOufCaUEI/mUAyvhpnHI1EGLNEpi1JOmQXG9tEqA46RMRgy
LJQxtZ33ALwIrFhd7fnYq7Ej4n7dt56pXASB1k6e6dcGZq4A3LFlcLkV6P3V02G2
azYU915vAaNcJqhEoiGReRUw2PZMv5xaEnVZtJZ9+uXpBRb+ZpHTbKlkxHwKwpnX
c2lb6g4Ak0uLhNw4vk14BERStMW3lChvq3Btw3UC2XA1JPuwRujRuQcG7ln1vbxs
HwOoV72uzL9CYk5dL7tMwv0yf0YK+AMQ0YkSArK4uUAGj5kem0F0XWTfybE6Fw1W
mw1adjVvU9PybMW+VSphHIIudg/4RPhtwfjtshoar19mtiJFqA3jTkjxAlJHOE12
PC8pRT+xQxoeENGLXT/mMmFe0356/EZM6l+x+z4/lSoV/LzKB1qtHtx2AVFIzT8a
SKDfRdYtWxveM1kLt0lqpsHPphMKV7ukzulXG6/Nn0y0NzecnK5rwCiKalkcQjaJ
sMaMK8RHdLvPCGzr7vLPivgo9SozTBmklEgeevrVKlt3uQUOLHLXA51wtM1I2qUa
ChDQ10uGZgYTCilQqirdKv6XC2xN1hFZPF6Iwfcm+o26iyZxCdFBlYIMnb3apuOP
v3PzykIwaVp6ErHiWobbUp/Ol/yqiZzYpsbUFrIVBAOlAnzjjie+2awicTdoyEI6
LRYW7JE6Xx2ZvNpbN7NwQKOyVrF8V+r2WQfJUnfziSyWnryqKlp/9v4vphQrhFmJ
rBlrVak3G5Nzh/UoMw+yCeY43bv8gUK2JhnhS8AZ0gISVFbJvbydZ89RzFDiydK2
M1Q0+9AnlxDDMwOFDcnIUaQZ3ifOCXkBuhxbwBIP8PRWSxm7qRqiNcsoMCW0kNbr
7ZUXuh8tGMSEuLTLR/kLtjtxu29XAhaR0zQxibBQ0DK+7gUZqPs+/7fDjACelSoX
tO2b7JuudyhFQExoivTqyEjGhcdjRpyXKk4OaX2V3EIxQx2duC9BWwvmuGvxvx4k
RKHwHcmI+e5Z6nRzkSRaZlg45VhGhr7KAFXjhV0PaptpTh9M7XBHYzcK6fxD9PNw
w67da2psFtx2scwIQj/itLT5WBBZv8BQAsPrSwon/YOqQ1+XAzLWkMRJlBH2wtiT
ZuWUbLydCUfvUSQmvfRQwTFjIq0p8BD57ARE8ytea1liToTi/269LRfoM8WjKihk
VLI+djOB9mRHimH5dLUCZgfQoJTZBJREFPXDkgasi3WTUckwRrz8uhcamX3+wS0A
VvGsgBuIQfUAm5VSupxmR9SwLqq/KD+3Ipx/70jD8RFDIo/h32maapmTNqUm+/sh
0rjMa1NUyURbnUPMLpIPcKM1hMXrZW/gMqPCJGEk4WfN84OunoRAKRkein4nfbUz
DBoQvUH/eAjuNmwDfHo0wZYp1TY6X04vXiKEOdBFeF1PR0WPjt/0GQkjHPe1RhnX
cXLCmbK5vzY9ppFlb5H56/7QlNjQZY6zQ/dOHkPUsGrDVF102GVoPyjVUlTzsAC2
6OYHY1Us3xrU37/Ee0Qtqs0ZsTbqGNFpjC8ncOKQ0aVuQ5rGrjhAiez1m7zsNuHx
uoZ8tuz4adMeTyHzzpSWMvKwg9pX6+0dXZ4olPKWznc+6fOo4I4P+tD/w1uGcV4i
crA9KvLXL5z3p2s9rQXV+FAGFUEIYIYWMOr7kKDEfLTKS1+R5BzxqkiO525Hy/TY
/ttLVt93fq/dQpe740ZNOoWTtX4Yd0S35MNYR789JBDw2KrfCgUdtuCpf+aeDGPl
qHeidEh0MoRNMf+B8BM9ayEGh/UUj0fR9V5VNdnfmfECbRM6bH4p58NViGlSTHDb
bOsyCSi+74vBZmcPKDSiOn7Hk4g5gJO6yV6KzkfkK5GcCr7U9JnDJ0pJJHzs9Wc9
EyGxSOYIbwXDsZTs8A/bGzkrfFfLS10EHjGmXZhdgdGRqipHdXI2vZn8sI0Pb/pZ
Z0kvPZmMfuZ9/fzoYfx2UtC/krqvhLOCUMbXLrvqlAuEcWRtbj5CQKmvfB8qLc1E
GJZco1O++weF1L+T8/9eSB6sWPA63XRcd+aqfaVgKKXCEoO1xPooB4K1Fnc8EJFu
ahWg9ujzxmQV2CK7q4vSnbmvkb/sxlr+pGAJ1hatXN2aEGP6pM5zSnK9AFG8oq+n
3uHeSauAzbCMh2on3Ol3n8SO/ULdIk/wU1WlLlb0hCEg33/vDzk8+lxH9nFIehyQ
ToAWZgEpm8QbE7oni6FRz9//j1HnzSXLpkBtkeZYuae3S+IKGxXlF8qu10aOacFw
f8toR544oAIIGmt5eUlbGZZ+N0DY5Y+/KLs6HXOkXZpGH0NwccNpRVP/ZgOSIEQl
sWW2ubEn/88echPKnA1jwN/rE+fWq3E6kb9y/RDFFjOWMgblnpuVgBwwIzPsYrCM
X691RxuRZXXIG0fQmINRxp/UwTJokQWMC5hK4XBmERLdu4SDXJ6VtP4FhXLJP7/+
2/E5/OdVjsJ5I/qV2lntvcZizzKyDekAQ7dYDbPmO6+UwH237rABlAITL5J5Otc5
cdPBUkxReFSxgpjwQv1FR7niI5LL9AQ4qzuH6iI33b/rXGuziHeQnwoiZ/1p7HBi
hyibEOiBlEltmaUHN6jX7MlVtV/vQFJa+WpyB4wjAz9fJKinXzoUul/3uRI7cFKb
TsKOSuApoR+THpTY+aWsznuqX1vs0yB7+A6gdSczXVimoDFbtUKS4tLqiBMYAxYk
ux45K8JkA2x5HpQpbxJXTl9YXTq0MX+6AhHb7OuHf0Lr4m28Azcn/6o0i+3AENIb
2o880Md37LEyJqaKEK4F1WoJxPKyrCPxcgvys102ggD6Ii6ZhM93rVlJJiRW8Efi
63Le2IeGosSF7ap5W/GM4wrNQ0f0WdEyneLCWF8xhDcS3GZVT6qFHgo62G4BlhcJ
STebBR14scS8/4ItyT9mG2pGmJKbiT8ExIgWUiz5cAAO7LJA5Y2ErXwAtjRdAx+N
OEfE4owzaM8hH0nPjP/FhF68IKCstrwlrhdGAzS/FnSYb6kyqMcQ0/U3wM9otabb
j1HvAdOoCiaHtRxkwLdGn068r+BEVKThnv66JY0JcjDXzgR3q4r0/qcz5aVyk4EI
nI7heEn0Yfitgc6UD4maXo8BAOtN3B4MLPFqAyo3gvGtyyr0rSemsHRFFUSsPQev
151bRf91O2Yxif0u6QAf/tkHiwDZ1Fd5NX+hViSnQZAkdo4gDxHDGro/EV/A9QNm
80OKRgtzOAc+4jBfLXbKBs0vfPGaTWEqSqFO7a/9hg4rRK3a7WTty38oZxtZ+EWM
xc9yNstRt1Rc1HAA7y0q5/fGqBvezAf1qABUb8UbRYdQbuDj9K7s1YTOWqIfvuhW
A6DtrJr9iBqTA1oMVr+qj5ApzHE57Flaif6RxYwpJ7s3umk48HyBqa6xvjtEmp/z
lRJqUTTvpW1LkY+MHZfz1k3haD4KDpEOVtNXrFR0bK+ENutI1ESWTJpikxgpNObe
moypIRbyBVxvV8BKgMty5VHgtttz03mWkAV9rm0/EtEmq89Ojbjvr9eCrdlx9tbY
W9t9Vb+58vNTJxdhAbZSP5rfhoIPz12AiS7YkCrdjuLu9zGaX7I7BQqJn2PfejqN
IuL2wD9/DMvBWibVwEklMyj9lAuVr1YKPo9sWAQ0OFrSqUdh5LAzg4LNMAHyZj+w
tByXbWPQueTB7g/CYtbldsF7oR1q+G8Si1uGMReUyMKb0FIQYemj08W/SMk4fUcW
lzRRq1coPy8pmZiEWlQHQmqUMtcX0Zt3YPhhJodz4M3On5FFTJHwjBJeYd9QzMI2
Mc1goWRTvS6wx9+kTZVZqfCfW1pfYZC5neZivGfTIf3Trv4aV1Fwx1a7lMXapIfr
8yc1yvQkxMy0VrD/ISheT0xx+haTZTCWxRjcORpGVH324W3usnbC7P2FSAMNEIrB
XtrotEPEdPJdLSqmVjwqb597yJzdzqshIzRf/ivq/ohq5elOxDBc3nbN/gWVLhG4
34btTD7pJ70ii035lmO06PMY+BoZSEUYJySZ+PjGBiraz7wP9JhOHs0N3PpNnGfp
eL1Nobelyl6e/461K1f+FrEgTMibyOP6ohnc4G5Ou0fis8liC20ngh2ZpNarEooY
HH6pGZPnXzFMSMwE9LZpYRrTMQjpeAJPBzCnWEFXtnieJfAwN1IiXNjOHxYg12+F
1AvbYqrf8AcHyWY+l9F/KdmgzHUekk21Q+rblWQHx+eNA0/ifUPX5mmyRudaDHz4
QgZeQY33nptGUA8zJaf3aXI18Alr3OvMFdPds6KzqUpYcVSIvNgPzAYABepTmWcc
yiQ1jr5/bQTlOZGBp/BUtoGqiCqatfhfRaxo4T3lwJ6lOOBXMG3DDZUTulb1eybR
WjsFjQKdEBzrZYSvxPXWgeyp7fjYnR6iLXc29xkcK9nCSxtnCV6TT/SnM33moRj0
fd2cC3TbYIDY7w9OduU5gu/sLqUr4NEwOwL7glHZ+q+QUrBF40TtY3OmLolnGewE
rUBfpwBMDu96+RtjFE9GJQDs3OLnKIDGGNrSDCzmXoLonEy7lswU0R3omUtYaCOP
CL6g88cuEe0n/4xm+baXj2aAEvBQmUjAUZEiC6tVsexhwKfVCkTY0ViJCb53EkbY
GHv63AJspnDmHQIuGBNkMMOdfFU5wWVtFGEYsxy3Ygedph3xdO3eaTpR1pL77T19
xs/0gZnyrELYJP9n/RzF4mvSyUu0WZTc1uj1CFUW/fqNGzLFXMbLcmWYtUVcKxwp
ynChrnehuIFh7O7QvxG5diolegCAUwxTkePtVWkcMiObugaq8TjaVv6sgcOhIf1z
eftQrHiSMu5FwneqqMfGzAwNSaCb1nZMmjD/cl4js5Vt3kmuNegjES5Zy6lMJRwr
uYwBY2vy4kwucBDxOa6UtWWzXyUToRg5FGl89u2St2lwbhpz2mAaIyFEm0Z9Cdqd
VUsERL/aPxA4dGGjIpOu5F3JFi/KqlKqyDuIgP0tkigmqV+gCGXWYAQp3UU8d+0d
wf/RyKjfGWZhuSUBkcI6w0bA56QDxrmkM1POApIlvZXzCjUl+jPDPZwjCe6basLP
xzbG8LAxULmg55Cau/+XAe3gVgq948voujxIPKCP2SxsN4ZY+RrKDCqKp3zj4Nnb
0mLeJ7/bEeUhqVf+UzMpPcWxhuyRWc/lyxD3N/5Ov86+T0bVK31tM5XbLVC7NXgL
mp39qU+Bs1n/qSA436YmbQqv/+71Aab6wkCVnDE12kQlXSx4BcDUGVg0PChic4je
0v0Yuphx+BNw2bV25HCR8wbb1TQY9gHB1EcOrYf86IyOUEu4OxPm/oyOZGmqdDjF
c3SODEqVDtHvdjbv+4HNHLZ0GdLd6wZZK1v3fM39/JsLf2b4XWcXXO+oO8UiqkJG
UAFLMbANWocgVZ2t9atisb26GoCnZImlTiu5GvkAs6l5ROe9sDAUdDgr9UxksdX0
9Ff4UVLIaJBD4yZ5P93Ww5L8R+lPgeK4oAAWJBdFf0X7tFdKyHmMSWZQZd/cSWXH
iAQ6jjPg8g8xIytKeX+Yu7kOcCUO5bvZ3RmkqxnWYq4s+9+vpjKX8AOseHxMa7KG
fnO4zfmA6rOIwTbhmKEWYjaqX5NewNPyqD/VWEF9whBhh1j9R/88wCqif5tO9qWT
59lLP0TIajucml6K7nP3XF+iOfyHPpljnRA/iDu8ssVP2xQzU2avOp6bvfAYBK9D
DqkX3qg6RvZUKWI7KAj1YFLjG+y2MaA3AHfHjKsqPSkhlh9hoycblEnMQAx31bqF
NzH81+6CMuRvRdhMD7Y9H/WPpm0rUWVsVbawcQUV9JEX4zzCCaooFCRA2Zq6NfkI
LXsnQhewA9vt/StX0SslN07PyOXXC9Nkc4LDmbXySNkk3WApMwNleCdhYomelyNX
eej75/2p5XCH6LwLx7K1CYkK5sUbnwfWa8mrH2oZRdahmzRPbizI3bRZln7Sdzqg
C1NRhNkPN09ze7hrm2ju/RS8XDIop5q7yUytoy/3uSrFdY1NXmcTTgximdy/Zbgk
2xmQDWmWDbkdC9yULp/GTHYq6+tvAi7p74MltYZT0UdTY5FMFn0qehON5pKxFUag
+ho/NdTGLcCBU6XNhRJZdfaECyvMUeuHZVe34rdQfFO96+tY5rqL3KLuKmjlld3Z
dICOCiQ3T2SN3LYGqim7vg3VTndNWzhqVkd1SlsV2n+/6ASixQk7BxASyB7tdVFl
Go3BRZSMR0XW/2AlpjvEsP/l1wScFcyNOj8JFnBdq9ax6Xam4jlGb1H/rvap7IXI
BmviuDBHowqOZAKh5Vbk5QsyYsm1NtXtDcpcYpHVKaVftdJ+nTJUMtPa+1XeIqzf
pOSRc/oTFodrEV+iMweRZGcuDQdLS+8soIzkZ+jjRFaXQ6UeJO5nw8WRRvzPayK+
S9pKNsR3UiqhM7MiqV2RnX/8ofy+RJ7VsXOhCBfLiKOXTGlP8wU6ZIybnj3usu+V
6rYusFSwEekN8mkZToyXLpy/GCNWenZmCXtw5z5UojVgughHDdGkTZEA65y+4EeU
qEGgwUGZs6cn11TXh8MTct+DTRHz2N3VSs7AbGy9x2R8WgeimJ6hhMl0qudS5dge
1YLTHVDGz9ZwbDFMcUht/HdSVn/Q63uNwyd+N34wCpPn0lZvxtNdIXkUolCu89dS
t6S5kpyuxj65YihA4jdc02Yli5CPLWslz5xrjdfUxCv4gegc2Lj5s/gPBQzt8S3N
02d8/vq+B/yquKlLW1/gUusGY+eL2NYolcCpm2uboKmSVzbspsGFEemGHLLx+ICw
0t2TVfq4vbklFciHTeZwQCkoQUrbTkiP4Km8Sghb0F7/mRjzaIs98w4xBF6jVdTX
daRCV8xKaJn4zrffyuX59HnVHs428TOIoqo3aOFThwMqDLNBMxsdRT3WGMLsZv6X
t/bhxkJfn79/xDbfMLc/5E16wd4QFgyk4LRNzAGDaA5rZIW0KVlUTUhIXicj8lVH
A6kopu+XsabL4bmfIZV74qBf7BO//RpZ5qVurdGA6/jfuB6vPzWVojfDn/p/HI5w
MeuFYkEfl5crjdbzus0jdMufDv/rPilcltXVIlKl2UhVkAiZco7Q4VXJy+gKtDup
z17pCno7kKP0pBdoT537urzAhwuEaPYSQKY5LpzYAKz37tGEzoeondRq5rh2ysUE
lM1wpkWph2eLAZcpBm+zoaZBvXhc3aeqQ5po5P7rHycpNkPuHpkceMtP+0CJXbR8
zD2J4R2sOANMJARmOY41xCryN1bomU4+shhK+QI0eCWBA48Suy75NbF6kpNoSK7Z
mFehorWacTdbzTrd7R7zb6Q3cNhIvX4EiWaK2SVnglUOG/uVUAixgqKcUa41JGur
ZF1LJVhQbqN4JQITbRDwqfKIwCgQP8+Wxfhbo/XmYlUlpO9bjEtgOLiuuZ7vGnRL
oJbHWuVnwlnAhgp13ZJ7c0wh8NN+/B3PVLkhqtXw+1+saKhS17Pkc/RPRTQblyj7
YudumsIcZ1ob9bNW2Ec6gW3o/AVRVV4wZ3MKjArThokGgLCW7wU90oJyyBU2GQmu
uUlQbu/2FmWJQy72zpk/iFr5vWx4l9ZnRubZmfpX3EhcHkhyZ2HFWOptixO4dR6M
UwkRjcrh1TLDNsUX4+YV7qRvHIxoPPaqRRI5T/VZgcxDT/eT5FkCq1rLuiWOEzl4
xDC4YbiTtiR+C+Nug0O7Mvd5JlDRdRRWMfaqepfhlpb0Ejtv99Nxc3eaA5Lkatn9
+rtOlQ9fvCtH6QMZRUT06fJ+oxkRN9hUn9klJqWi0kM/lmvkNBioxI7N0YtPmtkE
QWR3Fn6OexDVi9u/h897UD7+00bItkXh84rL6QKQRBgCg/EyWM09zwpEfe0R6Tqk
2R9tHRgURZvBNBgTx6zxwTuxob3sOkYaGApSAOxAdW62egBMOc2LUrhYD1urXP9Y
you9iKGiJpi3sNPz+4gMiHhUwPaPfLRD991zzB2fZS7r1EaiFDOOAsaG5aSy9IHN
RINFN2KZ3P38Ls3UVraNqhCzwXHqW2i9MCoAVOXFDOpbv+1mVcmXHf1gKSAQIYF7
zXjrQcrPDY6iaJbAlQz1O4RcSzYMIottTrc5UIJKCjFVvLq/NqqBYG3Ev9LYhqnJ
4mgRCCNRSbxCzeUvrW8n1zkBPLg22L0NrXXLynmZmUwnr8LMNPnhA+Jm6fHDP86H
W4Rh5iBlE+0TEp5oGX5/nceIXNSV5gMYZB7GWlbbCH1s4Js97iJ9DycnoTQjhcLY
W7uq2ZpDoR/PCNq8UzJKA54bLyRAU15sxOe3ZazpPZTqYpxXv7XplS0PmvBydUZ8
yUi30euX2Wi8vzI2jjUDLMzPjKMfj5MlEL7BTgYfZbDHOE+1CX4xJx8dPtyFn+8S
43t2lbgOF+9kE+C3BnvkSB6aCqZmA2Piq7a6VsJkKInP+mogwePJLy5eD/wRtnI8
wcM60bvclpP92Xb2KF9HUZS5BfcTcOhnD6jsuPbMZC6unXolY1P2u6+Y9DIYQHzj
QnqKQfV2Ma1Q4PZptRGztLXPuY3ts8ohknw0GOqSgyMkUTAR3dtRENiyLv/57axH
tK0Uxk+aXjqiZagS031y5VJrB3H/EcTIktmTQi/OwRnbkZ8COKn5IrYdL+5eUeZu
KnOPiCtm67HKat/sxxd2OX5Lcshj4YuaW2ADMvuD84FZxYuzR34XU2mQhXDfRksE
OFr8m+pKmqzE1ULpr4+vVhkPt9MPAB6U+bI/vXGkekihElbrt0Vh9FYBJpG6w6X9
yn0SuYQReb2gyrscaWazw5OKM3+/otBJcW5dgNxUKHfSB68GM6mK6v4qAKeMKGQr
l3/GxPkkQJkpvRunEjFm5RmBA6qW0YSbRXMBR3kdw9YYyPoXhs/44Rsu0VWsr+PE
prxex1hTcC9tKhH7gMJr0qRN5gC+lkG5ynNAIM7WX9h6+R+M/PqFwnaq5bMzP4Es
wZa5ApkyMULgr4ZQM1LYI7hcPA79lQUjJ0JDTp2qTXe3LTPheYFvRJkf5+1vaPAA
An8scBNmbF/75LTjlsF2Gl9lkmhD+rc3bMZseksHEnTjexcG15tesDALB1t19YNv
SUPl48H1pHZrEOmvrx22ZwQNYU8UeHaEwn6gMkHWei/WqbKbcBe0ax0c4xm+4Qv2
4Co7bBt2Y6r9r7Q+lP3mazs7j5RJl947OsBwB5VV6DDXES9Uoh2OY+/wCc7C6Thi
OyXHd8gHwUm3YLx9cdCTDGtdtpS9dFsqJM+ZQ1C1Xg4dtOaGKxoIpPxVc63WKqk0
CHzBkIXQeYSbjDjx5UDxgmSaFE8lAjWajYFJQd9nu/HePtG8B47qVT3pupZWcKvf
3n7+rx/yD5GBsQylQYls+MVwq4RZe1goxavNYkWbW1eyi49TKIIQvvXHgz0s71RI
K5zGjUXraoxZmBIGQ00vMDVAedmeldqJXVxBXfOFuTv/44is99vcodB/ZdUx3WzX
MOvzuGk8ta2PvUnkM/MgRzbmVgvkj2iyv9alQBr3+eEHoNiATXcBr741qtARmqsh
DZLBlVeV3+nFMDVLLo7B31FQrTNKuIk1pjzRJ2U3LNyQFIkxnRnfa8o7dzgp8/VF
LRP/OdOvivHE0fc0UD6Cib9LV8yU3/czDJwxRBX6jCSwUIHgikaLw26rga2Kvazi
xoGMRLcss+9+a+Du5yiQGvP1XOOX3ucv9SalbQfPJKMFONJTCWXJ62JzqiCan0r8
0MBw3nJ7Blt3xEnf8qyVksnoqUox+MYr2f7oniPOlfZfTKnUxcwdtNh889g1E7Qk
/oH+r5aiZZ3or0WgQ/quaMVIE81oUDw+TyA45FPW/etDtlSp15rYS2ZDwwj2DRJC
yHV8XZWzTtT4hpzdNzJRWpv6ESVs/1qV1AMBhUPVoE1rvsfHAYimJeR+x4hWCQMD
DzHeEUUorhrvU5kWsaEtnKzP+DyGBDuh7+y53v/+znna/3mqZ12buatThmeNlEkD
tMeIoejtpx9oT7LaiAI4WFoqA+NJPUAaerVS8jEUFqNG6hkhQfDRNJBFIyU9/n+x
MQRUC9v1CqrWCDL3s5oK4niMGmkNvIBfl7tISp1F7cjM1LxV9oU7luqRdhUrTM70
8rD2R6ySD48V8CNCpDV9B789touDRw3GkSU40vCjk1B5Q+z49/YJ6xUVFgBvAb8p
SScMa2ASs72P98mSR2XbBpoSIBY9psVld5tV2sxHvI/mkpjsP9bAs6pmU7cNFHe3
BlBf4Aj4j3JsS5lFcrTASt7b2tewft/w/dWM2nWFpbyj7AasIusdBm8uf6wBTY1+
mNjEgstet2HcIyli71+bDsF5Gn0dk3TuVL9fpSf3/FpQjmsyzW2ODLbZnnG9KUjw
TUexrV7fDaaqDm6efB8mCNrhRjbp7EBn+f6/7AXNzNrpw86CtPq8jA7xz260pl5G
16r1ppARm26yl5oPT/mtJocsiB+5in9eaAbw8CL7msIrUu7qeMPaauqiaOcGnXWp
AkAYdDj7VCpLAMdycSQVd4SoJRHx34HcibG1rRUeYtO8t+NnorDcB/bzccVQRsWc
Hy+8w3iAZJxmhY+gTCLaJF0+LqaWzjMpjT9ctdg7pYvFdpLTOt4ONP7j5EkMn+2J
sXtsnUC4g5zTGWeXbE7wUkF/yb5ElM91VSGhp0TBtbB5gTdQIXdYEHUfOMfrFKAB
WMtwnuguC3P7ejmF9cTiheFZ0/MqbT3qczUk+POwy/Pe0Zk9dFqpp4jma0cuZCk4
BFFUq00HJJ6sW83pDQKaivCNs6f5IDDIe0xjwEu+S+Ic0lPjp1bLnLXftGpyC3J4
Frj2dtnSwY6UKl32Sy2XOY2yTCuEhewp0bHWIUvLhReQwDvNGHqGQiC5Pn28ZTIA
LKLDxrqGlev1R2cR40X7NZq22rbuDjpKqxmPIK14LD+NBKtVo5A3OhOVZiT9mV16
1bUFS7Q6W+7AT5IardssNDQdeBeaPqIbbJrvnik4zMhWc+30rb9qvSfNpDdeeB2m
rwn+Kk4yNRUNlJUxY6IlBMPtzdA/GJ10UoZDS8Y5so6W5EixDQhI8Lx7M7++dVOI
6C2glRO4jXcQoq4pdRT9muNKd7Em4vWBmyGuHDAM8ZvNAEFtnOOCQ1Iv76TmUKyC
GFr8jqlEACzzxS+v6/29JLw6IFyEbFt1IlcLL2/1kd2xzh/eY3qtvx4jdNaMEh4Z
tKcTDevtsfqJ5e5d09cJ4LeAUYS7NJjWF24Ewkvmw7ojI2K4IV6Hkjgzouh3Y1IH
Neb036aqtzFmur6z85R+xYmq7/Yzsv2Fl4KlWxSAKZkVPXyHy3HVHmncTY8tslA4
+NLifI1zFtHKq9ZlmtuKxy9jg9dXEqBiFlV2vi3A4d3yAgOkZHZpmfU0FbNn8ij3
CPcCaoigv+Hceofzb3RNVdjTsjlhNj1BI197xz9IlcwUVU7S0PvnZ1FSTFueHfZi
InO7hhnHkupDh9ob59RpTIONkOT/dG1dBQzoyKhbg5NuJwH1Ax2hZssxI805or/5
QUSpMC7ejATxehlls4dQeAHXj3CDPmU7L/FnOiTn/g5j3n0v9mIQa+gxqEPwLrb/
u9cYI4D2yGQrssCkb0vx2obEeiqyISY6gt2J+Kt3YDVBaKLPC8eeLGkmuBQiYj7W
RMeRDY7+qqrb91EKfOVC9ko9k3uVe6zGf0iySmPzuEDKsMdjii2NQ5XTj3wdFJoC
KfzmHSCSdn1aa8DS1MYwexWKXUhem/zP05MWM54WPgEZU2J99qKTczCg80+ObmUv
DsSoHV5UclVNOM4mES39j6GUaYEJMZyfskc+ZK2D1zwJ5r1FItNHr6nsxk2HXDZ+
K0DgegSWN5K0HqhnoQicOJ+ArufBW0yfUNPGOxHzqWatUSRPjZNLDWOBj0GjbSVi
f5JBAQPKVw7yr8cl5gqU7aW3Ozgep97dErMJ/xJybeAaBu68HjqZ40dqk6PPtQQa
nBFlx1pCtw2ufCOIVQ+5utonBrLtehEO/5l8xPEJ9GNtqjU6MAeaRFhvJpK9Q0cC
Eqvf5QbSJxe5+2rhKUvukeMVA/qs7gOewa8UVNaIDV55ngHKooKGca87Swisbgqc
Rdfin/6/A3xT1WAycmKWSi77EhWVHDXiw/LKrlKu60fKdzDnT+uFECygsozalcp6
jHxAh/Pbe7WhY5/75DjbWQ5eISsPggcqiS3uPmvJWKkjbkFR5/udY6QbtsJKcpfz
7vkF0Zwf2US+/WSuP7rdRP8jhDlIzmIK7FEunkjINt6H0LXM41nzQw7TTR84E+VE
vh/d5aZsOfEC5UklNAiz1qRahXD6zpaPwwlPIZN1JUPJkjchLzUXkLSSAv84KfG/
RvfO3ztG9cusQVnUKLtLlcMJfjy/MofMlDvzdjHuNt5ApA8S8LL51h8eY17Yd44Y
b6Y0e4D6CD7MSKLJ2n3HjdggQkU0wlHvm5iYwcM64IeLappgsR6JmYJEyKKs13xw
VrYSFiAewMbKp+35T5maW7PL+Xe/npp0qNE6gSoTYb93aRhrC1F9hVyPHx9Jbk57
VV6Wxoz9p+XGXzGfZlLBMOTlVtrB76lnjqXh4R/w+9W8AwPqwVGGOC37amla+fxB
W66hYo5G16TPTwuKydYWZwgI0lae2b11sDK8Lh8RxUQXXiRrHQpJ3VlSoQl4bUwk
endD1Enf5wiKJg2NRYMvy40lxwW7fRCkXVudio9tU+IsFNCwQY57Pfr2nnVKu71N
gyqXo3LnqAC9s+c2FUJSE2SWeOnVlTEp3sgX3XKe7VzPXd7eYBzvrrJ3TY0M8M+L
GKNl7jnUyRSh3IrTV13ilbaa5VYiFJgelV4/RZ4gQY7ZOgnduKMaqtmE3rnEG9GL
lRtTtkuiTXm3TIk+CVh4lQMsxz0QxuiDZPPFKW6htM9dyrnKtmYVvLep3J0RrrXc
F5hUQJNO69AJzjTX6joGvfVOUzyro/BLIG9S+EX2FXaGDbOOruqjR5xPuVgHiCbm
LmjzDxqgOeoXCpLNFSeZmFjtLKADe0gPMleJBedjW395zA/+Qc2rsQh6o6jHAaRE
PyD5y7ObmjFN1FiBIbDuGd1Nl12GAQmGD5UAaUUy5UCVgPgNj6q8WtEbTxrpmVMb
m4wE7udhzNILxNNPptKlv8Vj/o5zXcxckPrt8YiOD4AyuM4/Z3U6lTWhHrIPoi+I
JkEuRp5Sz97KJu9Fo7MGuE+mugEAwq5X1Z8yXuZACYOyfAmvA+RVN2aNU64djxyR
qOSh0Jlw97rbqfZqbsJCtssfmrz7whckWf6syumx7Kyar/Vp5BjXLTa/i4VxaAR0
knRIF2mJ48KX71UWTFyTrK7+kvTs7+TPGWt/9rjUnksUh+Wyi3SjkxkKW0GUE49x
czyrQyfjyPnBOd5C26HL3DV3JN6y772SUX/ViM4omzosDlXopRTbupq82hsCIyku
GEDeEcsEnEL7TAdccHFTDqlvmj9/Po/+w08IvVrvWMxWYHqZ654hiqVdVi9xnhve
8rxLI1i6u/nc32iQ4jrbhIrPCrVP3JLhx9PWEsAa3EMmi5N0K+gki6R1R+7fUj7G
5ahGq9aH54cex24dvhgusTN1QNWbshoLw+LWh3vbdpHmMaT7IqncOQ4DrFgu4MJ+
4Z+UFNOVPBBbnmlzCWJy9uSZPPL6ygVivQrQE5ExrqkZun4pXXwSuIwCFXngjHYD
wE6g4qgbDOPClE7fDpweCWKUs4avxijpT6Dd4AGWbfjW/Cc66YLs+/hbWmI3oh4p
VUNPyqTtK8fMP7FN3YiZDY+3yauTqh66s/PELQky5QW6U0gNjQz1lRVRRKX3L1ur
3rKWeNQR+b5epVSmfom87kleyEi3RaUfohGARc0HdMgKKlZ0bg70ReX01I+ErabM
WRs6Yy/08JGbC/KHLpg6x+5MG6AcxR7yOojvo+p+FQEbrtJfbFEc4h//8YB8uzHQ
pzd1ew5ocFVoX9TIGPkpWobq16z7BXpVOYw0KjpLAx0Bfkg8vwsDnL0ReM0w6gnt
FwqXn0ioUD7Wg2tHvbaOwIm/7moq4G8LD2ZYI2j7NtPXOkT7reEOeKSuwonn+XlO
0rpLlhWuQb9/30UZbVKTn0J/Yb8uTQ/IqQ7soNAgX4M+lc4TRu65r/q7Q62yTWyP
9MHQxpS8WDxzCeXDFsQdibYVr+YeS37OKNDlDmzhNVy7vmDUWZOBNGAX+wwiZmLq
YzLD17q2ljnYwCsHxcjLyd/DFxncNHhKgAT9atkmMT8pUcvroUyMtDlZUuKeDcgr
i3n5VgS+AM2t2dRAwKAqr4FMDqGJnd7hfzB13PUyaAP+MDYyVQPYjgeWzrH4fgjw
JYLa4nkEDY9JzsB10ibM2NsWKBL4z84k3MGDUHfzbB/gQufxNF6Q2xeGfcm9gWGw
+227nmPoZq3RjpPyoiKlPsoyygyuM4/kioVksyuZ8y1kZK87eeOtaxjdwkb8hM17
Fa3xrqwZ2jynHB79IQlJt69AY8i9JDx+wu6mJfN2+IQFT8tU7w1ImWYwASyKl+Ll
akRVWZToxHk/CXJRk7GMTMxYhiI1wRutBbSzY77mYqyn2HTUB4f0zhhOPWpaDkc8
kW4QjJUqN0W+OWAXvIswAree6vXDuZbs6AZ72xccg0mnoZCe2HHwNDeAXZEDL3hS
zMVcVKFvXm4j/ZtZozhoNNgBJB3lsGWg20ZcQltmm+D1bB4hfNT22073cCcfSLSI
7AByb/ZTz8TmdQOP2RhOdQaAWuGcNBsu6EXkksAA9LyJFP0rCrb5pEZzVVD+KINk
Bh9Hi5wveQllxPcTA4F9cLk5lzEJkuA9IZEuR0vhP1iDolla/KRZOXeqMedE/R4T
RbRQAu3PVVminjXE/ff5CK2hm3hl3Bq8zdwy3t2rJw7qydMjH2VUeFlO7WeYKVzP
DUzP2AH9gPirC1shbRmKlQQY74CWPU9XCL/o1Fk5rLZ5hy3HKV11CuQTwC0rcEHt
uxIH7cJvamYkbs/usIKdJNHPJg/ob3pOMYAfjcW9gQVeZx3ZXvaOAsnKoPBG8dgk
Erh8jTOVWLmaT6h1kbAH2Oj8iWnF0Hne4Is7QkQJ8TLGJO4Sv86I4f9b8bjxJv1n
jmx9N6bT4JSC5dG8c9+0M08ciBaor/ar0eHSKLkR3HRTlZEvwrXhn58jKv5ZEugx
I6rDEqxtb5KsED9x5bd4Y4hLxmLkUxB37eKkhr2vlaXPHREBUc4DtDOuaVLWwGED
q+UBNN5rpgODULNWaai8O8O0O88VaV7k4u3BH3NNYYY+vELAmym/vPB5QR+fy5Uk
4yjffiGnHWJil/Hy14oV/5sE5RpD9r6nkjs8sRSGPiGCf4xc0jMaOedhsUVnT6An
/huOI1a7IHE7frlZD3vuB8waC6NplVussbv8tgu9krrwEmCIzAL/ElkbeUDqBKzL
qmoEbvErJitXkRmXhjepMc5moAiPygMcIhx+E1hQagRNAdzTpTPIbN+5FMdocsBH
G18x3pk+GIq6vu2aE/egYZUwvLrDvYjCbpt4Pa8XH06e+xt2qh4h2BEHgKfL7DRJ
b7nWOm0y3KU0JihrQfU9oQZ1rEJjqY8kTEZyGOFVL2WVFOYaGbzSF+lo2ROoepMn
m4lTE/6iYlGfANH2ZEBuxWYIP7b2krffaWAqkR8pGP2f18+EUCy3hWmCeNmnd1RQ
BOs9k53xuj4wwA+ZDfquJNvzlbtPE/pBPVUbAqlE1oUzT58yOrkylWNCaZ4rSuS7
RGJsfH7vzUinOhDnVgaWtSU+nyLi6VL24DAkDBciPZe3+PsqBJcPLytkIz0YMKtd
mPqAfTfb7YELBEOqRNYfa6jFRiaRywybaPUQRun6yqUQ5Xuh68RaF3l9awtSF+IC
pm65mnggr2rg0VTbmPUch5qDzo9coobD4E2CthpoY/QHljI5PrjdfHMjJCr95Q7y
yfoVwh8wFdUh6BsCl/o8J+88QsV7SaAkZx/KWW5w4zOtb+Zq1bVcC8ftn3k2HS/s
Op59ej6XcBBHU98t9QqE4/i9QHeIQwSoxveL4QeXDvgzWvYsFx+b9hyBxRAgXr5q
Yn5F3S8s276O3ofu/bcIBCSvPfJmOLg66WDWtTQAdqAqDYLvkhTzM+HcIa5VxOpu
uGsv+iMtq2uA2lyBtX/uQI4aGO3NS9jgJtCgItjT56uVldDy376vfK7IkDNuc+lw
s+a7hn4kUcgjWWr0dZJW/YXNi2jPaZervny9MRfYWsGErYi9p4aQyL8k/qH8vgyN
Ms0cm1+R6fMg9bUHy8tEbueLN2WalDNxt4zAjRKb0niKpwXZhB9bkrUUabW3cBXQ
psGFw/ZHQAGzrO/vrrHjW1v4MYQB3eui3q4t0d5G9udvYf5OVqo0B6JdAlRghfoc
JC43M2ef5zyFGhkv8NI3wrgoxTs5nyotem7AhKWlzyf2ld9j5ykVLvLdCHsGVo/C
Cvmvm6Fbb0o0hvvVFtlacOifpNaG+AgeACZEo0MSZK+BLP/70gJcreFU+GJyphZV
qq5k/dLXf4nVcPbt+zIo+wYEb2u7kP/LmKBArRLf+oFUpreCJUTdiN6tUSanBFNX
i7dQltNSoiw8ZljPrFc/FYnTPWfnHiGD4me3Icn7MupojYXpZMTbROFKtzPXrOBt
kPjdJvHHrFJj1eRo+y2kug32w7JoWm9NVDsxUaRqkIQHLZZNMmk6Z67jCzSa7wZn
gJyQJ6feXVjjUhIUvl8PRi5feGkkIJswLFuhX04vPCZtXNlwBUdtUCKrvCoWuF51
QQg16IyUnqFJ0iQgXz6S1e9BN8am7ls0gzpN22UY6m8/gq6l5cTJDUaPKe367jsk
upCI9/ED7iNe9XAi/+Y1HQ92qtnt6w+2/HfrX0pn5nQ2velFo/r/Wl6cPGuW2k4W
bVNY4K/H3gzhrVkI5P6rNOOBW5VTkVFVYej1hu2ENl2y2zBKMnOMHHtqUZskcHbz
8+VLwo6lZ46/1SvE4lQAKqPQqRiXt4GskEoSPvUlUbGsv9be4SSCHvFEPA4JBWFq
B5n01iOOFDnV67mE3vRlmavsoox7NdJDEhV6xmv720VhwLib3iB/aYiD1oe4DEMH
9E7JF6NPT6VcM7IrCn9870LgpISWjjL3Y0RS8jPPMCqS6R4HWvl7CNHJ6XB+IS4A
e28HoyuTDnX+J8KpF9wE+KhIwuGfN8pBKiBC8VH0U157iC9PxNaYw6Nt+LGVFJPH
r3OzVE4QE74TJbkaXqU6RdMwgnbWJ97tUAtmmBBiBP73wSeBxfjxku2VeFMpft+g
rAYjhY5BCrnZces3GnLPJNVlu7lNioAXmjh3nQ80o9agaqbWkYajXRzVjXa67OP9
tXMKaLZVbylMxYcDwTa3OkFi4W5TbIjVYW3onEUvTOtcjS5ZEKERDXLzJssFP2Xj
ex7TU6Xlw5opk0Ht5mrA7DZzceRGWo1kDGVR2s5G1Jj3A4HOpuQFSSPyYSvBS2wO
imv5OO0UNOXOdMxBWSN5gLhFlywDbRCdUucI/NajUpENVvtfZIEmgyullY29hmRN
TCFxYDn4ocPkPKKRB4+JpvEd0ls+e42tCJQEVmPjoQNzugkby1jNM1MdJsOwWhPt
7oounyIuQS8FItXWYO3yIs295tF63yB70yKjYvfrVBSrI834BFcXrUHvJneGwYxz
3BCDS8JMsloJZnhpGGQsIYhzDU6iHaupDczkDDhB5Mkfb/4Q7BnDFSj1tnu7KIxd
ltgkkp+U8UNeMeQu/iqBoAgmaNO0FB/ujK+IMSGu8doaC2Qm/p1VUUBxW68HMl/m
ayqvxobWqMCFfKLSbraBt0uoCZ3hZs+Ym19hvt7pSD9Xjflmuv0Wl/U0T7uoBYWe
jiQCgQ2sF+0GwZlrQlstKkW5iIVhLWY95dQ3MwKBeQ4OwlLMupdEHQvxBjyPSWOq
s9uLJIG2evREWnk1ppPPX1tWv/AlRAdn/68HMGvkkxhOcbgavAECj3ziKCVHidRR
xqlZG5ON9/faIFfbgXFPep4MDY8lRlJXzDxeVDGnFBJWtND51NKDOkw5p34ecEMB
USoxa0L96m4ZDMiz5tvhtCg0fQDodJzLhrn8sMWZtvPjuvRq/VqP/u0cfyt1xL/H
uvm8r8xRe8YsgTpcEVd6VnGkX5Qvtu35w8T+KZWw+N/tndccg6M9t/ixcXSXJrV7
GFMW8K0XZzrQuRM4pih5iwnhWuo2EbwmP8MIwcq6WuMyuVoflel/gkRYFvGYrQqi
T+a6ZtrnZwSwPbAoYgSTgfdp6DwEkzVX1V7B+l1BkUa+UR8YYle9D2z8bsNzlhiu
5PNBlgl55BQQrZNL01+Yz/pjJkWoZ00i6LmQs8R4uR9Nv51su4q/jwkT1id9Fd0I
8wa4873BDRN62iR59OwDI4iir5X8y1uAh9KOvWhsLGPomeQvElqvLBMqj6QRMGpK
bWKIX9bPBkbO68Bz54ZBnke7pIY4Wb6iQAwwt7S0ynEiiznTCVZFFBb1XxiGUO8Z
An6YWII8FvUWNTmLuhRgh32g5X6Xj7Ytdt3SqEzOrm/86kSxvreUT+M8UlkZ+389
cX0G19AxZ9aO0/e611HJ4XGPIDUSymhJrwnUCdarjHc3zz2apXvQsNrzD+yQ7nxR
NWAGWUt/9D2onYxY6JHQdXEFIs1h+jAwT9Wg/Ym/NigaJSAhnErzS5uupfuQ4zxP
hFHlDnw2g20fG7yl+Uj7g8hg57db5JwReZjwsxDK98Ch8YOKkVSyQaMyP6Zrbpta
dAASanq+Khn/nCnJqs6G4RpgZR+QArI4HcWew3dxn2+DQJYeJAI/2KEIhx94z+YO
li3/mnVoS+f63C/ytBQFZxeXB3/cQ65aA7eHVRCs5wCGBtYX0UrW44RNhCyCTp++
yXDvXbixpx6b07IQlCbeP5UF8jwohK+cALXwu0je7uVUbX5y7pPJGkhpLlqL7O4X
PdctMSdQRf2+gITzwSEbBE4t//TVfDTENWfo9jh89SniNO8rb09GKNaarWGVCF/T
LymM58/TlijhdsS/8u1GvBcsnYynFKAryP0qmiDCEQgucViAEZKUIiwoWZHl2h3S
CvwdGrlax0lRZkCkbZxZcw+gPFoSmmQEL262NDtN9YCqi/lr2MbnYVEY6FBHaHMT
4GhwPA4U9odhEu303IOKK16kXovRvBn3+9rmRRN2AWHXsQx/m1L3OPmUQHBdp600
+8KTh9biYEcae2ug4xWz9GT6AxbaD0Pl76bAOnKc7ogQpejj2+ZMEeMt4u/mdho5
oNUCh/9nREFCL3SOHrW0UY6adUB8N9x20nvJkqZ5DiWycrSX06xuhvf+r5ZknFXO
EPNBxsDpUnXu4EVnQghZGWGfR+9Nz2s9r/GbFZnTJ75H3ulEAOtFEKUtUTtjmKIy
4qMgABR2zVeSrgeTswQqsHbmUvtpoMLhZxWv8GR+RokDGhnISP4P7eOESG8YoTo+
96UwRCqfDUC60bD/n0DjkaPyPg7gu1thkmpbrgOy7++VtqQVqQeNqpHMEf2swll9
lXDo2FIhr96E9FXtn6FXzbNn6zlhRjud/rUFjl2A3lN+LiQoteu3tb43IdV3Bmrb
5jNM0PMcpJcWjiQErrxbU4v3WVZHFLtHji51ZrVBDeOiDLcPWu44jR5TNz+wNjUx
6CeKPdiLKvDJN4E2BFI+K76C5SCcNB56JvHzsR5eCD02XNZWFg5Yr7Sx/eoY3MuX
79QEKDb+Lj6760SFSgieAsIrnSUOctgCMyyeA+kYhxmJ5bkwmLz2Gu/bzpwac29n
1kawV4i3XzNh9It675jdOr6HAQoV68pzJbouGtMucMtNwWVCiRi2RxY1vpKWuM57
nGfO87Q11MvHR4e2LTt8tC2Li7QPtNRIpf7BL4D3onmgtBdID2vbeBR+/USoyKlF
yD1143jb63v2zP5p4F802zfPDX8Tsmumw17rugViYcN9aFMdGTv7EOK0OcxH6b5a
gJ7BuOAq/rbCUw5D2WpY7bUk0UP6nt5nbeQfxP7k5JHu1ryUcUBCCmQHexCwGk0H
vN4fztjLh5D4Alk7NojxEmlrywfGW3VJSydGiQ3OMkwuh99alf503hgZv2SUDMWw
6UXSz1fsscPBBv68/xYOxX/44O4mJYGRVOHKdUsw7euwBJCI1o9LuUwdrvMO5huO
B8r0BXuGP7MTvXb3UpV8ZzcTZ6E2orwSY9IrmvPRPxTQTwnebOBauOvwOWsHSTF4
1q4Mw1MD5cG+162XlR284Fgfbw5C09rwO9FGimQFOi2iznkc6Kyd/z1GgEqIpOsN
0Jh79x+6owu9l6H8X7hIqdYHpj6fqXBosYxWC7XuYvqVLtsmESWByuCOUgIiTXDz
xeqoFfXJCo+rZJOqcO7jVbqRQcIwn38mJE3/r+xZJrx8DZftcM9lUTleHXA1quZT
ELUonCPJH0ihUFdhUyGyDiBaZEw1mEGBkipxi4/jlo9ZRTKnlkfUrdpm9qdPSc0t
6VxkBjB+whHFeXnSKpbIzLrsOfOMKfje8/uCrlB/AQml4oUPnUwgUfTgNkkJwYxS
DFQYEQgGiMZiFT0Wg6SEjMGmNj77gPIDQQn13+rcxXqnvBHOMdn3foqv8DgvfHiE
9E8LeB308+x2J3R3YAFsOUeez8gcfBL3WnnHriMuuhl7iCRMuaGdpCS5Jbie7hA6
3Cx83Rc1CeKBI32je744KysKeHJxOU8T0lFWt8guab1cFrO3FIT34ENn55q310Z0
adCaT+TmZI4tfoo5+k+u5ce1NAA66wAN6DQqtyKK65aDlGXK10iprQCW4UXap2Vh
9ChUaLfRdNGCPpMl7hMzOo3xI2J4T9+TczbsARfJyuRRDh1aCGJAKHAYoMAu1E38
VoIEDehWE5g1lEGJw6Sfg9bWO0/DfSeS4PciDcKiBkAYDzMHMq8+C2A5uAtrgtVf
WGWWBLEOxyPEksA2BEbcVtnOyivVQXcGTL4++rDrSQIw7l7sP3/3oRm1BOQWBJjY
HuZiudDgxQRtMbeZlW9/rIiVIJ8RHKF8Hd8ltl10cT+2OWxQ+6h6pEpmesCzCmVR
Z4sKQoyUDffmgX51Un15+eUMnqPRUiv7mANY4rl7egMgUPy511ikU0pOddZtOnnB
XBUumHsABkbhMnuEPfa5yEwv6a6hGy4jknQeJaGVG6slsEG49MfDcOWSwAl+7Wug
J0/Ftz/XVpaJZ/aWfRxdUSccShxxu6Pf8K9n3g1071aWAADby6ORIGVi2nMGDvHh
7dARDC6w15S3hgtZ8AQwxqZsFCDVvxXzunorkoHlB6oeE97nYJQHNYwiCiBHAER1
fB7CQvw8W3ex7in0GsHOT7yniZ14e0KBZMABkg9trIeAob75aV4TsNey4g0LMYTk
Rlj95svSm8yfx7RkEacUbdI+90txyExU1lHsJXUK5VmcEjZqZMbJxiR7dVV712Rj
LCk4S5eRWmhU9aPY2DFg3o+bK67qh8jSuP41du/AdLw9dNkEoeHRJOUbIT8pJMnd
GoACZE1Ki4wug5ic2YVt0caqJX8E63Uh81EhW7oc4UkeIGFtrvXf59rHimoVFCcE
wcdgY2MnrXsFvca/Q3UhcPiudLvG42B8lcux1RAUk9ED2J1tTfjgeZFpghjTHV0v
9SctYz0uob27W8jOyV2d1nlKx+lliEKbuCdq1RJPzaHJK9rfZfx62ukqH4jblMma
XOd62EvPJ2TWHsl3IzsGE+0SZ3TGeWLJp7ogzoiahZhHY3xD33TjyTBPwIdQIBRU
KOQ6siobqObLu9/Ghkdp5AEIWJC1Gp1uUnQMYowEj/jNIFuRGyxTGVknzk1VZkYx
cgQjDXNpVxymR80brRSohVlAbTIXyhlFt6PgwSv/tApihLntZm1HNoF+j7IPFhjQ
NSw7pdDSHimvjy1QmgfMe+jJVv4A5kdK9kj9KEaoF29qpItulkceHCXSoxVxjzTY
+gWoZYGGd/aQL9zty43kpBeU5q9H8Oldtgd+K17z/u7BraT95xCxW1bdrqfXcd9H
uO/9toGf6jZIucSJc3UMiNbKVSGkbO51s+/dbELvDCHP+Zq4QaDwNwaWhxWkcsuf
olYr5QNkGGt+c/muN+X025Z62rLJjaI1c00kWstbkNeOwmny/f5SZDATB9P8LPCJ
FrkKmtOyCjPSI13xG+DU57drkodHZm2pqSKJLwOlkT9tANpzxV4R4pJgPncykZtw
qAldzi0QhFZ/EGNQUcuIakijjEt/Wz/H18/3jyvbyGCjKFKKcoYRyGeUaoPKt4r1
qgKMhh6ILQgobJ9BFDf0OMnv9ZIsQaKYTSGJmfFHn7UlSaa3MRUZ3X0VRi7J4jRU
5+WI0+hqNHAcIn1Vnrgv3ky9a8k+B2iu+weIdkhkKGzpQ5qmJMWmlEodP2nRHsl2
sGhXRXRAI6n1GJOKK55RTEWovficEeJAgDIt3w+LAs0SDBpZO66GpdXUO29/+EoF
gXEOJesO9Okann+JrhuXO+y4ARFuCfWawbbdjDmj0UZUDf2KXdTFm+w8ftV2kC5L
8Fri7CVDlOcKsvUwUuBrx0qKNCNKMobuWmTuiiafh/ETHFzS2ghW47T7J77r+zUh
9BZ5WuCmGBCeu1c6ztEcbHoeRabKwCYjYEseMs2BrTGtHCif8YO/Fl4w86HrnNPG
kySIBN5dh1XBI1enWwFIBApycQRHIt1KNNMn66KjzJ1ywxtO6I4tWgJvStw21Q6U
qUCZQVfGnSBCkN/4PvqPKp3sztOckdr7ogfTcX1iasexHQfILguDTRdk686nQl4q
8PJv4XS73mEYJdzcjQl5DI9hrJUht2YDSQ9DmJA1Xx6n0Giv2XZXdXyKrtQ8PhP3
BhL1odIx3sXkAppYmjXquj7/XG4kml2q6eFM4ebZzBwTJbNgTR1akEQnWZjW+5pj
T2gotoUuehOcJrNMChaJbMfKDDAoY9qMCIb2sQQaPZsCELd6z5fI9tRhikEYcgG7
8YD4mf6+bVQAkRY/oxlHN0PEOlr9oenIkzpUAqYNeWk455jNLhvQNkOBLPBgsbZJ
hLxPUtjusGXZ+sjXzAOAkIt5wLktIqdaFvd+aaNpA+E6rLe3+QMFMiZAvwCrWZzI
YFyVmEvFhuTFSHg54YGtsaExhRXVPl0OFmHbxCOYV/nl4n2NHA9hFDCZ1BEShywN
EtplDRmw6ARDKCD1dA2VG3gZkUbtxCbKCs1hMZ9Bu3CL5oUIqfWYzuGbv0tgw+BK
MCEzQkM3R5bzoIZSXk/8lyFY5tqfpebh0wMEfn7KmV/ZXHwapHhIeUYQFLw6vJ+2
tXh1j/eGywON4tPby68PFqUCYNN0jleS0vlBzK9KzlYGKexHkP+NYHvEzGdIKaUj
6Xij4AXL/WlYXxM+IXsENNi1zyHFRQWI+YOh72iA8HIOCv71rWxEhE/7LNJfFIVb
b/95yHWycJCVg7uDKVBkWoBkySBkYZayDya1iN/1K+fCu/avnpwHUlFvdauITmLw
lBSDZNPdgrblgBCqcx713DkCriOlHmDUk7yIlcT9J73EQ1R0phg6ksPyLLRrEU0w
AdXVLgfhts6inULAxtnaHeOPRABz7m8iaYDsNUmueuco4srbp9YMFvQ7gZ3mb/3G
1dwACld5Qv8XYpXzocqTD4aDL+Qybi7nMlq0Vw/n6txh7H/fNqm1bDFrLtDG/kVo
pZ4o2sQCcx+sjWS0pgXgSWkhriDjhwdy6kGUcifPR9O2KBVxZ2uDGtNRwGOvcUlW
r2bumJ0niWeLKErZ9u+MbIOyq/nrL8WjvDksk9Idne3gxXDLwAkY7csAsiROw5Fr
uR9LVtokcIPX2OlxlH8duwLr0RMG3Kh2XlJqFKEcAEFS6TY5B47f8I+sfdqIlZ9O
Hn19EkqA87SF1b2aSHWIKXpti+AglpmIa+xKKVO5WSZE026IgIHBglNTCqvsGfHU
Tg2PVN8ZIEwQGbZhsOCd2N3r7LKRidZQLG0x2oi1ePVn4iCrzii8WHWwpOU00Wdr
3wie/tl0dO5/GiSgJAnyd5fXFxU8KDzInqjk8cSH2fh2F2yijvox03mrQAvJc7P8
+KfxLERbu4MkWMNqj0vjFKQrdGA6/LqsvjbqrpisGFu4AnnG4HHGFr2WFT9wkhFZ
ECCuWRntEfTAtZ797kkalqxvbQNw8tjphHkgWQpzNj4DRlCnHHmrCSBxtu9Icz9C
DncuFeMSMY2VNsrrMkSMPgKK/SwlxEUAHMjSzKfizY/VlTa0516T5ffsxG+v089R
SzWWokMHZ4vzj0iCu+pvTDZJBWOh5fd/5W1bAsNEi8sQQ3BONWy17fcSHeMvCfzB
3iK1sRo5f1Vem23idszzPdn8TB/GuC0VbA9ZC4KNQBk+QP17n8LYvCvEAwusYRy5
upFHkvBcyVd7YOIIQqQVA3TcZpZ16VoSbHAjJqSXnNZHl/5/xamNk/YfHkGBoCqv
a55lVBDiDN8vunz+Aso2j5fKOMXYYNS+DKCZD5pPPY7xt86Q8UViEC4IMxi2YP65
CGeEswf3GcTSsCDVl1g9LpuL7A2tb8ME6ohY58MrcHUU6VYCQnhCM7NP5Zh1l70q
kMV4QBohuldk1MHznZa1+SbJp160tPEwScfZIftICY8t0F12eE6wpQbTGL5TO9gK
NqQSyMcbzh9lKUpiU+YHZMu8V1ZnK8u0isxANSHn7+NT7IYReuDIyK+iMq9RtoCe
o2Ae7MXkr5KkcvwYRV5u5PfskSpb0K3dUseiEZNwi11mDodaOO7pbrTBLzUa21qu
l2zJ0N3BQCRY6OhOFvy+jfo1eRTqfcgfN/LExD7uZtO+BusFkoDgqPf0U0Trjljq
uHcxibhLVcbE+CQc6GFVG0hcbuqAWa4xYD7kb5Dmq3Je0W/j/soRKC1LBCwpVjvv
CZaHlr+s94qKRmvxUEV9sfALo6hP8qfLHgq/IIIkqGgSNTWcYOF994AfPNYL1gsT
IJfzWm23Mro5sCi5E4MwM0x6CpNZ5XvI9SPzXcgFPlJU2viKIUTXJrgE2MrgaTkU
2goHRf6P6x1nYAZcoWXPv1Cwfk08uJC+AnefYCA+6UuVcBWSKDGo77I7VS8WCnzl
l3S/7q35pIeWRytNpfa3EMyjyjCRJ0yY9ctv/YpYVaODPk5yYIW7OZDFBDdB13ZL
bz3DxhXz7aYzG7Chhw7OxOfOcUTeBZD325TAZe2lJe6wKdUKYnLtYBjnPebwfEKE
zeBAnyfoNIUveigKc5mwAs7UkEXkKPa4XzMn1oHTal4vXN2vu3wPN/BPTaxTgZKx
yxDc+EfKhpAj5Fsh0JpF97TR+cY2e2KkySkDCRTyzcGjx8HLVVpf5ZHcoxlRHNgK
idUKKAIfXcfo1ESQbENOSUdM/kOM88AG3YvTVyRHzrMQoJZBFrBK2eCtrIIaYgZf
hgjmTd4z1/JDYWHUFo4jFarKE3EnQyXc2OV+wFAHo3nWxRlUQpV27JlTvz5u3vX/
08LCJJNpjVvw2S0AMqnsJ1BdvC66uE5TSBoj8nag6qoDrx//QdD3G8t45+BzCq9k
qR44PkkDeqw1RaFE/SJz98i7z9pthG7VIHM0yom/007EmI3agdc6TCiCdUsAV5h3
xRxTAJ2XoWyRNYusMW6CXdTn/FB7gSvvy7o7OprNevXuytSfstLJGiF1Gfvsuuie
hTxjhqYffjiOpQJEUqFUdNxHJ3Wvli1XvlXXQxyBR5OK28j4m0AL0DFhm7pPVGhU
IkaiuqGqDK+KGqLZXMQ747kNItKbPNx1h4RXLgGIBYOpUa1FiyKHSAnLbp2JPh/A
yG64eyWNhMQyoJFS02HwXN2HcohJXfKmZYszd4BY7ZRy1JjYNSlkmiOk3e+wXXpX
Db7jMhmBnnh/LgBlqS4KRDDSAjlmNUwSXegbn7Cpmr952iW05FOfAOs9MM098759
qBYgFpGNJh2M+yG/eKd0AN5Nei3zDLfCiGm0ZKIWObndNNbwVYmEUrabqVs88nta
2vJmgIwnQOIlAw/8Zd1Y7b3xa4EwQRYijwrkod1vDz4tdedajBmYWcLheQ3CBx+K
+v23gv4La76yjweHctQ/JVZFp9InUIEKobR76L/uXY6DOkhMzwQKU7OvsI5JOdVm
QRv4rSGuWgyXKY4MGVFRl3ENPlVkx3JxYfUyDBO5iyNrPkhWWHbCxVbf+tGF7J8l
TK7hY00J3LnjhzRcVWI4kcAR4fNwJsdF1ZThLSodo1Eo0agzfA/zQmz9DEF2k3Ur
KTFWI2zag0uC8IHwurhT40Hh23c1qu52SHMlbY06/GFB9xQKHg9AwBZPN1N4Rl/V
hxdUlM+EvCi4LD5QEq+CxZKWmsSsP9hsI2QFVIqeGfFV+sMoh/NuCmLeG2zyhLRZ
xkwTOD9ME4MFtsYcmyKOTG/oySWf/cPW4yia13E1I0pHRcc1BimLnK5H+sRTsTu/
UQdcZVeejaBurezx4OuqoS7a9rKvyOJgsLm8qXXENdiREulPtK2DeUspMS5YdR7b
5KV7e1DhlKmbnYJ22SwgMRH9jdgBJkRdL6VmdS9bEfS3/PaXoFwvI21YaeK1o4ug
2Wap0zNxCQEHrItDGpEJvXlyBcBEqdWNnsorGBkK0VfBS71JkXHPw/ZRDOQ8VGlU
gbW0ElXuYfxOgFqbweffL3CtpOnsiqXeIG5T+6APowaF/usbwP5ygn7GMWrGtv6T
RnytscxiAMVQfJiC6YBxECohQ0Layd3xYdsvGDSyXLVITn4e6UamA9reIsr4XPk8
JnEm4Px/LqdJ4czh7WIhC0EaWss+x9ciVGUBRU8xl79yQeZhMENfFYN1hcrE82ro
a3dc+C9Iby7cECju1p1N8p324jhgEBcCxFMXMDA4msVHHQFnE8TkjyVs3lXOfwMm
Au3cuRBoCh2N2nmJJHpAauuBc4Ef+dx0xQmIeomEmcaYRoXCs7UqsFppEk/qlxkZ
I1mv4SAeqHHdOt9lV0Qlyv1fZCl4BMDzBCAStdUviEiVohieFpRslygfOWMNV/Dg
crJcLooRJASaJcXaBqQOKapamoAabD8B7EOzcBKVt5tsvzJ02mpVkIFPVB8zeIyJ
WfZbsgZ9M1+iW+K3N2W7raALFsdXq0TVr8qixNeN1wZefFZaxTngKgCWzsQs//zr
reHHQ8zY+5V+HMSnvsJ0owax1BP/ODNZig9veUVzWHmny4z95EqFdw0GiITPZP9C
saMlqYNF4ZaGwl6RcO3J+eUmLr7qZpMHhuViYNGZiTz/QwY12duZ7XDtecbfnCY3
+eT3lSPtdBFmD9zP0ihz4pF3T+Kz8pbohMXO/uaH/e5Ae4Q2ABXBQVAncejB7APl
p4OxzThPbT4OVCxKvE612ixuoZG9WrzBfbVOO8J3BVggrtsgugCH662K6nbbPfF+
C3ibNa4qVkVgCWA1+OC4NJgkQbGHUKY5O5IW4Io2WyklWnWMTkCjwqoCceoTcSd4
2rMFV4iYkdMdbZ9lEJnCpPfVIkJ8/I9FGfr69lLNZmpUzZWOjQKA45seEOrFo+Q9
63HoQK5HuZrRonMWu+JPmkaepX74+woLfcjkU6vo34OmKAZ5x9p0YnXWnXcq+gdH
uQbYf9zTnRuL/72OtCsEHtlc5LoCIVs44secsKqKF4s92DeJ214L04cMiaTVp7Ri
3piDa7bil49kJ5mXjy7Nzq/QxdZ6HOhDemGrkbvvZap5rBvTR1mDvK2ORXywaJ7l
DioffA8u0T106YMzaLyMhSQtYYmfZ14g8Ag2trmFGKxdu2N5h9pYoOmhFwf13/cS
5Fq/VI+7sQNNtFrz0VLuygvNxSe2Z1r6J8DmyDq8OBeZQJLL0nV15bvoMX1coYrV
DQ1wiMeFICsIu8zsHe/8zT+FcG1P7/p5gUQ32jHimtc6PdZh2wxspPf9t4HQZJgG
IP96bU3xN1/ieirExyxXMFC2H3srgp0be3TJnRxbyO70EqgPtG2G2ZyFfouRwBe8
vlj19/u35BC5nBhqyzqn57rr7L0I4bDON3jM7Dtyq9vJ3nVNV8BNPmNKr7CepKjQ
CI+LBTWW2KNtUL7yLRlCw04BM4H8dPJqCEUSICbOWSzbGYcjbxiK4QxnKYTdNNuh
dRclFXrxKmo0DF6IRPyjCdlVgtG5TvKRzHIJ1FB/C/UTKz4nSh6nAfeBWBGtvvhg
oJ/DQ3ikY1nR1EcU1F7f7JZjfJr++ui7D4g9wLUDDOCkJU1a6UyVEmwtDte/skVz
oS5vD8aFeYYuY+psVWjGO3EqyJL1qDhxWboTrDKaGA0ahhmbASSGU19KMi3DbI3v
7ND+Od0ZNJzjEtCe5T1nAnMUrBePkvGCEI2wL0t4pWitVYBrBB4FiKHAMzaU3U41
bD/ws8dvbhzUQTNHj97YpIWUYQK7IUK/8ENtI1zy1lmodIbdVentrZDuwDaxFYrN
pq8yVYugjghbjuRre3CpHuNrFOKQc0OShoPojFsXTOtLWCG77VKTJoBnB9bM4fOE
0GPOk19XxJTn4Dce+AilWMmrFy4opr1BNGJcMl27M6QGUQ0AJH4R8xT0YPnlsa3w
hWr1+h4l9ojL4opgTrwgT/94BmFRRnJB+WBggT49xbXxUY4lEB/8KCNR2OD2qvkG
f+BYsG5wKBlFett1AenX7PcHbm+RuDQEo8635qeplf66nqlXO5/hZQx07GQmwh/2
FybNvPGjSxDyMmt8yYtlCkSw7RsisMz8/KkVc7n6mJtXF/vV0FKegJI4E3EAbg60
V8Ulu7BzhcprEw/LdZ6dtR2LXAzKS4E1q23wGQCAm76bleCcRDdcvmy96gxYiJOt
mljOK0WjEYwoxLotvIdyKa2hUbZYyyCtivUBuVBSFA9vyGwHMBID6QUhuBW9Igt3
3RxKJYk9JnAPZXIg705k1iQ2ImsGoTOqACl4m82a3poYeqmgelusAS10jeoT0mAg
UM6KUvWd/sO3ad6J3WxlFHyBmK2IQr2amM0/zTuA0OEiViAAx/EUNMQa+hOR509J
m1+vPJTIxOhEe0kyd21BS7w8b6Zji5OEBoLDjT5+9+5q6aqz3V5dND3g9vuEDKX+
8O+K8zoi+pSfuyu+rIuAknIVJlBbGdNWA6gilH/Gtan3LsrcTqJntx9BQfmwMCFo
iH7625/HNaVSlz6F5zJXKWdBtVwG6/gwMzPnuePyJcjikb0AeZk/PYXL0hfvuzPh
kw22F9repRl++/0E/CxmowK9FKvhkTwIGvto4PInP/0G/qROFE3lPcz4KaKejs9j
O74oeeIud48xkxbn2ecuxen0I9wFlWiwnTa/SoWojYffFnPlumaM1ENPLxcstvd6
u5MsRWTq6RErEyO35dCJnpqXCEcZkp7GsCvhK6A8vo8dnWU0ax0AeTTqMX/ExdlC
OeEBt6FM0ccDV982G+5yjLlPedxH4MNJjGIYD3KO7dVYnX7f0BmFTyYR96F7CSCR
vrrbcldEnACI7fHx/Ca8f5tgbeqjMQcrWct7vAwZFQ+Le0LXDB8VnGGUoHuPTF9x
PJBoeUNd9cjw9YcHBhk/Ed+ERb+4iOJdSlBLQUrTD4nSukauZ7CuC6y5UnqbXdrD
vBWubbF4ctE01ZKli9pfSYhEYG4Ur4dN9VOq93zae4v0l+HS7JmXLIAyFaglCSFy
GIC6QRXpTrncfcr2nC+dOVadVNrubfyJnHXV/aURgs2dQ+dKpLYOcVngfB06H/2i
KGcqVJ2bqJTfqCasN/Dnwg+LBws70DTjkeZD8gJHmujlDHC1TxaI52mi84zQxst/
WmKyxvtQvDLQ81PgXNaNgYPw2UZKEa9z7Zbf/IPYtQ+H04rekU6muBsyBchZ6xTP
2oHHXosofKRdsKuqSYkZYbOJpg6tD8785RiJi3CtYZy0d+M7Tzp98GELbCC+iGIC
K7/2znC462Jfe8kMdSLQ2LhfpB5L/PaFE8l2tARxrTJHadbhlh22RDGd4O4ZZgax
WJWL/pH4Bdk5cLH+KAusp+XhdX4uYWMwjyoRZTAGdn5Mc7qOqoWfksGMOHKztr0b
wrFMcCfCAoBQPBoeViOn/PXD69iZ8Ak6lcDC9BPmD/sVexeJowHhAW1NYXBx4z2i
wq+nGgIB3Vj1DMwYAG/ZrB6AnbhekpaDoVFU1/TXUOPbkz+En+bwqvL97rzF1Pv4
p5zQXrpeFXs2IdJ1+pbQM5Wa3kmSnnL6M/OxQhi3mvZmGrUb2ThMW1DvWgOeREnS
x3CNucFRb+676Zmk3U57zSJ2Pm+em6oyMnB4icLUX02pf7TAXudJ5H+sr6FXAWEb
jjtv1ey3BZ86pRfEbxLkZTSF+EEOtBg0Wm2JL7G7ukyKYsTqr7+dLcWzQr9ujss0
dgcOEW1GMEpzcEaW7p59BdFICr1PAyBwHSqvfdbF7aS+atZn1qQNIlGPUkFLhHm4
mpYHRQwr/HPhWU8RyB5+HH+zMNDKytb+FzXA6va8BE9EWSbFhcEgySnW/KyWGSF4
s5fiNkObBQorrV5QnN81M/sCv1S8lu/fVUlAi6tNk1Gv9z9Svgd1FwreOqizahwi
1cYu9DnOEMTtdDfP4fkgHUionUQ8MmgxwMmvYpshmFwM6PH9XUeaE6V+sEyueg4I
mEjq7LWFJDa9YVpu6wpdGBBmV3k+uD4KfuuDnAU84AM3CmWKCr4vFceb6tYPZ10b
qeiSGGvV42ltVyBK2jVFTa2SKsg5qV2LhA2CU5TWTfoouWMuHbXVfRxI3oxQaHUd
nCJ3+xkT09ER7WPFwZWAOB87pyHBJ+6DpxGrwKePzUWs/p5vHyQcUPMhkZQN3tDA
Jetjd3eo1BxV3v1/u0EZ73nFCLZhgDA79hsxgLPuYEtcav3hTMCzBi2ciOmF/Tha
/KWE6wCU54LyH/kiHev5rYvVJzAnShxid48GP65hFhqMJKD0KtTHULQUnlaT20IX
NHJn5yddNtwU96mPC1REKd/M0mYx0R77xN57H5HuQH3fWpZvVWdVuMG4Jn5eWO0P
68+0Y53dlevGEJ7Hrkd3uBzV3d2a4pkQWm1W+szJjhbMhtjaOPrUywRjEu4Fbxyq
YlfQJgIFYxvcXySYwa+BW+EaMi/lILruCdiWCZoGii47QpcfJhC5BZ+zi7oexnoH
RGG4t9k+7jTOmPneOQxpwySppWBh8BfluOBkFcecNZsKmtNLtdREA+o3NcmEm/d2
gGLlF5aaSSVuVJPy0pcOcXsdaSje/X8XhuSvJLbxBjMujwhjNK5oigQa+mSO3Kio
Co1EfrGxWcnwmma34h77Bj2aKVbIY6vDVuDqKdfxQoZA6ccb86adPFTHfArK7KNv
njcMqUbuhvRsfoM8kilDq8/HQFrIcHydMOXQ5seJI2TypkjqVZHKIxr9ry9E/lmA
+Q0+UND/tz1Ak8ypp0JghXKamvdUUNhcrrmNWw50cYZYSoi5eEdI1O15fIfmeAdG
QgF9IXEYhFoPKF/FG+mVkohCVWXanXdMVELwBUgR6TuQhMWldPJLcIURekg0yFfH
ekhCIVKFEEr3XESo/XK4polOLdJ/wfLOquKiu0ifMvEmgU11tddzC/TAMu9XgV8B
KGZvlxnaMH+3H206ivv7H5RtAyTgY3DtQgqz7A/8kzVAiC63KaH6k8kQ6Ll76Ytz
zhwU67lD9TLqnyqvQPQBTVsh39JD2/o2IKveE6OqjNwFcYeaEo45d9SnJ43l65Ya
+EabAVzYus/thCgJn4RfxXAA3gDUnB9wgzefOEaDBY1G2x3AKWushljhaDefOgRF
EWv9zT636udnWwMnZzCX6SfFqiVVKyS3SqMxg1X1XlVN2qyAhS61g+nIlrr3+pA4
whv9bNsI7Y6bF0UJtiBDJ84JfAXeOEFeJ/p6dVGSoI1SDdfAICTYR921LZ6ek/if
Ag35Fleh5YDmDAee/qPBW6BrY1Pq6G/Je+tcQEXvnsvb+aVPY67XYv/dXC30fJAH
ZPBsh2G+BvloPPRfv4rq9Hut/O4QfYLFZo1e7SrDO+1w+WRyuuUMOdrmNnbWCDI6
A4vUXqYARFqPDxyIj4mSAwSuEtspu6KOwSsKwruwApf0ha/0iZSD71c7zrz9cgTn
nGNHDl0A6Rb7iohjy8XSPhSKfBDMIuCjUhCJ356BU7BaLlsppMWFzNnyXHjegp3z
pd+wnIpSUTbsHaJKKxL5eGAO+xmLIXCKv8K0XTv8TxIm3vsPpADkYWy2XiTbk2N3
NHKA/kER8GOC2F0z275LZ8Jth6t4Byz8y/1iNCz4rX46wthJOm7ZoloX2denyQQS
mhKGhex11lwhiUY3qdGI8PdkfsRT774gk1KBx5eA6YBm4JgWNioeQ7yCusw36rIY
Z/tH5McrGGkMXZTKabkiMoycyWmaeNB1auZgPgSpcCYUxBuYS9BYfCbWiUPybtg6
v7+7YMsHIkkNa4JGLeG1d8VyCvLDDh75TAKq3pvfbk4f4vTSd7ItwvbS58CQHJqp
3ytitMmbEb9XNLR8l4/eq9uFoomLnX90ddjyhPTtic0iTc/f8XRR6gKioxQGyv29
KyXjeTYqM4uh0prVcwkx6J/wZWALoZ3q73JzOKZy8iRhqjEzuyom08x3gB5H6POr
5LCgfCIpkH9RMReozFJVWRbhddzaHh/3JztswnEfji1D1vLkOPXXMouIc7sDhKII
3fCX1SqNkv29erflUyjmMyF4XN/7aq525iMqA9HiNKbtU6AzLmrKlzIp/BDnWjb/
hEX/CWylFFvMcGQxKPSNM7wyQFqyyf4oXKR+U86iArOn+XCst/HIoS+hq1ZwHwEe
2I0LVdRTehFP+iVA9KSj4vM4IiFIZq+HnziBynHc/vMWVpe7FEHI+Y+UOHXaSa3q
pddCcUyJEZb8C8wlfWomxaNoYiNcgrBsirjGgrdSoxJTvlcM0l9SDOw4nxVZnha1
z4wcH/M/LNBiwMIDpOmV2zdRbCNpOt4xFx2v7tyReV6dgT9n8/K3RTXleZ+EyxVv
2qudAWw6p5wC+aCRaB8UOcTPg497qGAqZLfk9VEnrlBg72ut5dLAY/lHSkxPSmL5
JNnEsRkNROy36sttn/sopAb6xTyEjF01aas5b5RNKcyHjr2BirgBfy4ZmvN+foxg
QJ2h874pboNQZ8geEgiMeNaG3tg/JPa3NO5v6ze6lOr4vUKXti8MDo2gzFf7EkC7
idQJkSwqEWofPQ6gkO5SKqOACJLTZo4qixj/v88EMyU535oZnRMIN2QmRKmrZnQQ
lBcjS79UA1WYoSxPVuW02fGki12QWvLrKetZMeleKBw3jBCxkcLwutM8OwO/aNC0
rPl+o2w8gSO10jmjpPj+B5PVtzDNgK4aPfT+oLVCzak5zZoUKBeeNIIgNAAP49MR
mzHTdRBvzBk9HNY2C7pfvPchKKqAQG3aNYbkbA5dg55t6FaAWxGSHk7RuIiMttYC
zVqUSVcnvYLJSIPOFpcnHfCth/tKK7L4Ur9dm9OtlagRtAxRescpAz1sgFRUBYDp
+Yg1B1DSe/TOKkCs450Dey1Qo1nk6mRowZV9J89g5CCItnIpgJqFwdp08IOEsah2
5/ywo/rcMBdo9JS0ZwDodikEBT6HVIzxnbiwCIT4YwdLCen9e0F1UtZ5x3C4VcvW
ExQjeeT3zbk1vJBz+6d+RBsSTy0mnv09nBBlQMLcRIoTqLwhdFo+Cn8GsLo0AqK0
cPD02Cy0B/L3IAmjmTh6EWOuN9UUIFFoOeUhgnpHWgGmJtQIFXCeatgWNHL1ZFTH
eor8vyerBHkTppjvMa1eNzj7Nb69tTqmwlpXWGquhKPP/Ot+vjd3Z08BC5oy1Vcl
g/3/PJpm7S0mMHWZ5byiotzNXh9/RQ0AEQSb/L6Dt1jn/TZXtqacUW1fdL4V1azr
PJEzAWer6TQ0m3hWyOXPoTbVVEn/OLGOJGzVCVnJ6xpoQWz7GJwSoeXPijPVKi/b
6by1VRHsLUl3UHRHcjirSM23f5YFzT/2+GFMU/5/xhZlpoQ7nL2zggQ4R14BCNcM
Sqoql2LZMRgMDPvix4JL/BOVjXqvsqAtiNeY86iWMIewYS6VtF6OqAOeWp4chdBW
lWwi1HnVcPvOn/pfVPyEP7qehECZXZgrmmG4JkOBeNJlXvarf1suAr28vVjcsLi7
IEXvuhuPqeJnSUmIzOTEYjXVWbyguJy0px2LG7LToN8WxsAjIApAmOirU3Ic68Xn
OL+x9kA4uxkb/wR3cKkama/3jLuHMLGZCJCnVTMwxfxD+5mqpNfGz6UVdMFr1I6s
WJvb2sSe9kDLlfD3nlPjs4/hAX0ex9/6DmI+aN8clVBhYR7OptsVtrr1ZBR1cveg
qtEzstFPf9NSXSVSp7e8Y03kgN+0dF2JVrhLRjV6e4qlByNhuKPoz/e0C3OmQTvM
RirwBtu9pW7vat7+caA1d+27TX6CoPkWMrMjyyDgTsJ0hjSPXfp/jv5i+41WHFSB
vqXYaUtplaXwn8EEcmDDcRiYOm/0IphymX3TNU79dD6NDANc8rK3BnhkY8KK4CfY
7RuswGAMcSvgeg9juAQwq7926v8ErKzXK54FJm9lEZajoTYzpfSKfD7zf5LHhxzw
a9vgiUb97uRrWRuhzJZbThTUkqHFO3rgYMB179dbhJIvXZqgbsVmkJzWe5hQc+X7
octXy791WUv5Iag6Inuzhh/etg7Orz2J5JuldDs2btr56TvLPMJ8TFvO9+EDg2Le
nI4C0DkupwX1IEf1pY3deH7Ttc4U7mxoTSgndb+AtwCZheuu8Ffto3rINFOa6lfP
N/R5LPlwsvUYZiqwsad0djHJ6NHtLwUtyDm7hcSMWn0y69jz/kNnhjh8nTOceEP9
xu0j1mwGLNgJ70MTXkrQSRwoopwKcnSx71vdUFwU5zFS+ugJ/O+NYJOQHqR9Fpjb
9lgJJIs9QQ0atrcH3b9RtDPqJXvi2x+EHJQHMRRNbN01UZYecRHhUlGhC9Eqy2k3
n/CbPb87TP1elQD1HVUGumQZYxAYPRHpzge7imdxE6Y/G/ImZm8V74ICWb+zKSCs
v2yzw+uCdJB08xiDuw7/z6M0FWj0gMIOz4icFjJW2OTqE3hRv/M3b1LToU64ZlgU
natce7KUhB8Y+L12Fs5kXTJWm4BqUiBlSdf/D2JbyV6yO3aVjrQcd5o31reZKvx/
wbHEi2n7c1IBw1gA/OaUaTiiDs9PYD4dKV4p+eJsOzK/jPCtYjs5eCmCE/YAJj3G
3slWo4wi2jc+dNLSM3Cqvt3EyJmu814lYV7erAza/6y8973feTjSFXxMLHb/oFaA
UD5OpxHG3TtwrEg+C0uLI2ykijTVSGkyb+BAKpjaKPnW/z92Tr2mE2YvGPPMmsYi
s8tpOQWkeOQx5xtM6HGBQ0ArA2oWoT2xdfnfo8TJrYD0aHS7xCukSTYMXM0zaU5f
iTkhsaCuKYPSH8JgOsxCZLT8VRPIVt7Gd7aK5/K8ODuu+DUYGKV4zCmUa/WoO+e7
eiCkhJVudYO/FiP2nq6PQdW0OET0S7umyKQa7l5CjWr1xcEtMbzY6Y53QI6OLE6X
dXF8rI1QA0ZF2o0ife44g1hI2JvB5TzXAsGEJbjstuqjcCERpjzVHtkB0VuGs5Ay
M27sCnJoBv3LEG9hqBMkwA/j5xG9mn0L2QncrFcKZAalej2c2GKOeGTzFCXCFlVL
+VJcns+06218c3rdIx/sn+NUChsiJeLyCYW/+GuDr7jOC0KTlX23E5YVQFn0i4H5
IDAl5BYfAN49Nw+c58drQqLXut/pFzLtCDqFaaEL/mOceGJkeSfK8rvHDTatxATI
wihfVTsq5wZ115qO5cacInjPAwXE/LGYtorixwgir8KTsV63MFQNr39v6F0wVxpL
WJ2W1ltL/uPaTc5FBNGaZoYk5lhr9KYFidT7RqQZIM6dE3XLfh+wLuvBahlQ5rI8
ORaXzAB/dTtg/wJANYeDCQGaPjPgxzzGYaMitJfdNoV87eozp7l5iEUQod5loylI
jeWNW32WKIuYgOV1ey97wjtpDZIgVTU69yZAzN1km325UmP3Cg+9Hpfuf/0Qw1Oa
fnWECFRV7KXlKn2FCHdUHURrtKZCzHPTLRVirPh443xAxOFFTruMeLQSRXfGY6XI
NnBIZyeUgzkylmR3kPWOLkvBwNpCBI5brnY6QWLmJt7e6AKPKDh+1TrIHZFRkKHj
iFx0oZm+UGkr7sohUVbAq8G/HGMbRfqWoxDMOi2j+1z0cyngokZY7sCSUAXtJpy8
lgxv+3+KOACx8rqGcc4LUy+gc1Ov1MEEEUHvnXW0R121TPQCLQNVClzEXy++ShIE
K8NxDAckYldnZcTQjxvU0SDvFSHwIOQ5F2E5pKq+Z66avtje1Ww+8ldZbmQcBhnD
lzIurRJ7xvBqQRNgelaIC53I6FAEjX3I1+ybC3gqUs96jrP3FYd74o886dfA/IPv
NE/Pxu87Y+5xItY58fXGJzMx5cUX7PzWL2CeBsNciRe0E6dGtQab0imtd9RdM7HJ
YKjYD4dnVt7hmQtUql3fO81FvD8wyUIRprbQ83OIw5G4CndB15Pcp89ddhq2sW8d
+5yBaUUCbgazOQApX+mFreN01yEymAAetsV6D4l9wj0qQDqWTbvNFCpWlCZiIhkJ
XSN04PQyLTjKUj1Fl8d5U9sLZsM9+9I4nwS5BPMYMl0ctmnRWKkVWlURlnEPbHov
aP83mUppYda1yGmdDd5yCZAfQI2LbUUfFZolxjVSjTmQZjVl6uuicMMV7Xrd7Wr1
tW83trGkSygRBFZFASHEpLoJWaZGa+GHT+RmHfcWhpYnjYMUS8uespaJYaX7YSfB
D2mfxNZTdMTDAVwTHwdLWDIAc82tCCICNPrY8hCdATQKQq4JmOEin8tcBPea3/vH
mnm/8jQHV6akUPavruHduOIARgocs2DNC4HiIVSrS+gN6z9ckenO5GJl7oS3nWc+
4vbAEUNiOZLWkMB78QYkNq7E2jXi6NVvP8WS8W3R7Kfam+g5G6KF6mXCUx+m4J5Q
mi8AjbbwX7U3w/b0DKk0athxRVSIBb6544qB+sNRoWkWlA4WtBFovNstwVQMT3PI
w0SeA3Ry824NnsNEctjUYi531Rn5AGXeMYT479GlDN6MrZHVaNWHJ93SYAR1RPlq
hipbtBHS+nKWpue9rZL+LFEmNR3VWJRDD/+6fj2ZBaqUuXbVMyfFBy/8QdEkH0Dj
wyFi7JWx49NPULS1ASC+8FHRRXv13nAekN9mkzDGawcbJKeI4d/mPaPCspplRYSR
Hnzw6840LS34qPJDNyOVCkH7S9AmfGGpMVm9v2y3poiLf+ZhJrBz+Io+gz0ohBBM
BnYxZ4tTqmUV3jN+HZW4W+a0qeTzaLUZcL7W88VODvymlBjlqeSxYUbSbTm9qWD2
R1APvmRum6klo9HyK/oKrM0l3KIXS5jtiPAncGeTK9KeubbDJMx7AKI8sJOIkqoq
fc3KuwO4uKSgAnTeDERfgSedeLkzQyH2tAgyEyDjYDlv7ge1NQNw284u3VwleTSn
5cLd9aN7vavz+bzwgWIVE30hSyfo+FF/XuYe3k/+wYVeKE+Wq/LCj+c0WTKsmmR4
2UP7YF6jDB6GY6p5v33waoviZphfe4pStFfc7QZF6ZZb5JHN7IKMipxZwK1LNbKj
EkzwrXX5XXMpx0ZQSUWL2eXaFwYrwosh5/8x/oISgCo2K1fVXt1T4efE3augORUK
27YYha5KO4PsSw/hHhmhXftshy2dYMV/hEtL95daEH7dApSNl3/8ivI/xUhKpfbp
6lgtTa9ob5BO0SZ5/UWS/zgqrUv5O+m7sQKwqF1wRuMMn3GRaSm3JM+Q8bf7V+Z4
RK5JXLvjUwf59r9CAh2L9GoP3/3KsQQD4UX5J/zZbROXsCO32jInIf0/UlcDyMqC
bNIMLSBHRoVKuf6OpNI6WQKhDVqJ/pjUsGcI1VS19A21pdykGfFtaNrSudU7dSKw
4rqZNW7UyQpA0mhelTQ4UmpcIT0ZNgyqdxKBWws+VZ0/QGpkQC4TUW62QPZ2DrES
WGu7vDksLqpqQA/5dhxDvivYxIoAMY5GbphQ4/EEoe5AQTQ5T6fpp5OptUEQklnM
5yK96XPNm4dzAs53YTDG4CSkz0slMQmsPq2Fp8GDnmLn+7atfNtWMRgLmtDkLYup
NwSflmwDoGKydnylOlOsvhFf9kcjnKArcRKsSS2GsDOLK+8BGlH5dQPfEPSyIaCN
6Yc0kTfg+yLa7WcCn01AtKTLeCQ3QiMAowhIqZ/+L3tgzPUjph4EUcdycflcpM4n
4OPBw6cTPc3rxhLpVfU7kv2DXQPYZbjtePBLTs3ATHpLC8eyzb4IZwDQwgkQdrEV
0aIJTvWsFaYZ1XuUwwHg7YFEvpjJndbnA9DeSL2lracB9GkSsCFD0dXOmaQvELGB
IlbKhTHYH7qd4fOYOOLq/0kUH7xF7ShaCAsC02+FzAIMBjhrOf9KK2zQrsrppFO6
NVVQUh1vJbEyP/kTyOcGsEmGu3Kd26B/httioyGoykhgsxNIrFrpPJleFp8J3GHY
O9XFBBIho81a+b6ZqjEIiGiDMf8aiiwb2NEG33ThSfikglr60QLuTWWNlsYSXn0L
UT+vhj2jhoOwOxcD3Gg3I0CLf8bduUiw4j8rX06XuEucBPBZIfXrkI0axpwrZc1o
OrLDnxRjKAkQFBIyirHvuldP9ZQej2SopCCrP96K9XbYjg96zNqlEXbBEnw7vtcR
Ag6CT0Kz+CWxzTleSx2D/mfwC+uyWAd43h09+XpCWpdg8pECyC+/Qd8+EEHTuOz+
CD9cADxzOfIZhtlA6t1yPcm7DfsRQ2/uJIlzZzQi+JoexWnc1g6ZzA1foOkfHZUk
CVOIIg4yoCddS+tCZmG4/sqjUHh85Z611aAyQ/78cbGkHeD9krCoukq9y/aeTges
6SblG92q8vzkiFHUR1nY5wmYPdPr1R9o8k3mROLasJZxCLmW1yTaLeqfaxjKrZgR
JbaMehNvJsgsTuqpdS5e/kFdJUK7tJ6RYMqBohg+aldg7crS3kEGtcOCpwQEeBWN
UJKw3bdlu0UI8HKDzIuqVhN8B1mHaiKHRURPVvZeuei8i947dBvielFrc2ahtytd
ZmfaqyxkGF7rvyoxExKqQetE6Xlsw5Jt2YfZAV1Tuvfn+blxEo5NbylBX6Sx27bb
oVhFGbwc5kjqGvv/DV13zowfBLnyWeVxF79BGA1y0SpapTQsTWura50w1vEdCcnO
WqAATgkEU3KG9epfrf9GiNaNJm3/rj0vG4MyvSDYUy1pWt5Q6NkUFAToQ/6gEWI1
oN4g53YdTHRVZ97UUoQ8Bnlder/wU959+xe4nEidZTVZVe0dQdovw/Uspz2MTC+A
9JF9mSo9vhZ6RrHWQpkEEhPrCZb9k13kZM8GwLebNc9MMbPHr/grgoBenZjrqcl7
H+pAXBxJwnYNut5lBp2VEAKUQINTSkC26tGCD3MduoGQOvKOo/yDucD4+M2gA4Zz
jHTmuabJeAWYzUc/3mCMz1vrH3JOb9RrNAReRHmkiJLSQIXxPmQdqfTdbdbyEooN
ffbBrMBEG9Bjfni/V8pCPsgWy1/tS/uloViAueNxaa6Yh937WOVZCYGhzQZBvjl7
/7TqBKxU71hgLLUL65wSiXhi2GUNeV83/eUkPQ7MPzeHZITZ6/FWjlrYmEUMMYXk
SCYZBECC2s5XnQma2YjaEKwfCPfOeHeZIB4tquxwNDa/py6Im+wf5jUA9OZcJHJQ
82jAKb1VCGNNSSSs0ITfCIAttbu81FAmJkHqgx+0HwhbZYPPWxFBavB2k0Y9TxOx
HTj2ALSW7uK3eLlAsEO+UR5fYtlrrv6fNLMUR+AgiFzOvBkPfY+GEhMilVNRhABq
PmaJ8sloic5aQbkioWQ4rK1Y5CQ97BK7KXoIfljvsjF6+YNzdgb/8v8tF/iMSqZf
JXgg0i+fXpviblI4BH0FzFQtTm9KivOMzkUz1mW58/ooXxwX+X1/UzaHLIpfwYdJ
I+sSrRuKDR58VR8z4GYBRcspUfckwP3g6P0NhFSPvq+uVHKXU4m3MYP6Jjx+AbAf
IQjIjYLOQTpB89vLq2g1D/Ujm1WXOqYwndrsBYLs2ljipV4WIDKIGkgqsCaLN4oA
6ETNjmo9dSOoKIJj6H+i/HU1tN+NeAcfYV4Yca/Jj1zz4ietfV7ChnTNYPxZxdcX
+3k2PZx6uyPhq0N4GtE1dyPpiY1iqvFhs3jK7wNqlznLup94jJrVUPNmf6LruqqB
eUSPh60wLhS7TcG1mW4FaOP3Ggtgp/9ufNP6gDo3zraCWgU+cdMqOTaKEhYty7RM
lOoSwC1eKpLg/eT7xIVCnKnvG6PsH+JLH1NBlzRp9nYcUtU0wC8v/BvyDeBR0Bem
eB+dPnyM5jqpN9yI6ouJEzDwQoMTo0wJRD7i8GX1H4Klw6RQJ+pum86s7q3xQa6L
OReuaGqC/zr6iYz65+GRmMVqeLxtvC6PIpjWDVFgmXTU2LlKlEqSZYNWu5jeTDiV
lh2AnmZEzeab5OpdQWQy1Wi3L7yI2Z4oVrzJ06ETAwyHY2INSMAxtusoIFesQjSK
ffOX7zZ9wdtNiPBe1o36+soRL8C1w7/XzeFjemjnOtGUmWOjtjfzLiXvjZUx1v/6
kMxvf9T4i6jKzKGpVegqmbPOGrcWLJIIqrQIJnZkt/FhqtvbyfLLe6qE8Q/kBiI0
CT0YxI0fXGAPwTtUX7yHKVh9ZegBEs2TJm6c7L7Yf6B7nQbxvzDrUOZRwAtZTCVS
VjhljKszqXvVZJO3HuPw5qfF8RQP2jk+2PcSdEOXpCbGJby2qkEenTqc0gha2Hxj
fYsaxcYLFFFYWRgoYvQgXQ57iq2+qNVU2/n2aUy9Yp2xzmaCq0iTRSM4b2xUOiIg
FSll+JyOCqS5NE9CF0PyZFOUuM1BymerX2gzIty9Jcq2sR8+TEuauA/SET78jF0w
Uz9xId2uvB8+3DQkOdRrq1POIUJWVma9dp5qpnr1zxDpU9LsqXaIanXf01hbcebS
zoKjQiH6ZZzYsgdc1imw5ydwEP+pCbe5XK7JN9+OqcpJttZeZyatbFbQ6A2Papay
Y0sy1XcYPs3iAtwB2adHDORrAvPqvFY6+UZxf0MQQVeFsghB7i0A4hFwfMh6NINK
54yu8jgVYkE7wIp9G+86WAZJP1sHGkb6U6Sr08nAG4ZRbq1wwEOlnyfqFEnXThsN
Z+UCIjckiiLhV3AE2U1KInZqyqJdCcnJgBZ8lO6vKj5LbRijmxcPTVcbNv2nkBxp
DbWmXP0aP0/Bovp6xuJw0UwMSRp72QQZfgXhKGoe7nQC1VXEVbhuHLTg5UmQn37R
eaFrYmd7BIVTR4fZwRRqsDMWHt/8jfnx7gZlfOTywNYqvE5qyukH2h/+CKwolJe1
SdHtpPUMfqqZJz2lQDTMFDGCmumWieGG9pfokGUOGcPgEUkDLK8n6m4DBRznDUxq
N7WnFeHEsnJc8C6/ioJJJEGiJJHUa9Y6PMV6gz+MOAJ6urfO1TjyKgUHumTFp2y6
zWh896pLSI8EBX4N54+rspm/YXm1UNPNkuPq37lDUNUnsL1sOCpVNzUkK3o6GSHf
BZ88crusbizuDhEIG+h3f/ZNPgt1UyeY7DWmOvpoPYSnWftywPZvGGgTqz95QYPA
qwC9ywFoO6GBHFvOjkWijAWnr/ZplGRxDmfip0xtnykjDU+eG6aJH7St8mrpUIxQ
H0I2ggL9siyBTRnthqEFeECDlz0udZk/QHdHhNBxNgPW6EtIuckoPKb0SF94DSyw
OiOO5Cqc/+XCpoHBpJ/AOpECJRJSYFzPMnMqYk7pkeY9CTRW18BzmF38UZ3JGcz1
RSRahJA94N4IhjiDjv3zuG35uYsav/49FkMMI94YnJtID0xXJRtUH+Y+h8vEETFX
IwORxrFg1wTEfq6ODsvPXXIkQ8tU/LbBXst977HlZPtynCWDVRpQhAReT6zTJb5G
qB9l1l/LUu7IN1Icgu+KMDkpqa97GbTJq8bcVNi9rwru+UrqtIGNQXbtG2ICw4Q8
Glrce2GEudY4eOe6WINstG9oURLMGqMPkL5M/Egk8gGewRLegQZYrEu0G27e3MnC
jSzKg6QKMFPLJ5PemYoMmhpis4SP7mCW62XiBVpObkIxcVwxew6xZ5CZb0w2E7bk
kJhaM/NEYWFYOU1HIN1qdrxUookRzop0eNYdkt/5h8CYdIIJbgGSUFZycjRlwm/o
YLrf/JYkx0OzKFCwSVFk0S7lT7hXgivEXRucJDcvKkZMd3VnSlYZC2MTveaDTzza
35f8bN/isv0KROtLKkS+IVHqdMeaSWegv5QQxORHC/d2vEqDO/OUAYJ+ENXrjMKt
d8a2sxkkZmKRqWcuGg9cH/QeqS9M1uDV9k86kqFdQjiM5xmYwLQguAkaLGkuurgi
WneVjQyeH7a49pgejxs2LRmP/jfnAgpBPfIIRbKvdULmewP8EuAYfiCbm/1+aYa0
XMLJZV4N83YYMewO2NbRMNIfru9KIl3JP1ne58eLuqqeR6bjEZFksjWBFjqdoG6w
sLJH07cUVaQcTAiOcjGRRGY8gjFZQO0QN5unKnBNyI/vPLO4y5UiYN4qWMX4EQ/d
XDxV/iq7qRWDSMe1Sgr+QF9oml4G0fAi4fWVPXkM270kS7o/UUeq3R+V/uoDhXTt
Jh8pgKLIpCKynW0DtPPodsVQwC5FIXbdtscTQi6jlmEkwg7CGZaSMRvqT16n+3fV
JMVBzJHxfOuDl5UiChmaPP17ZXHGtRu4btiZpmg30Tii/9VDqZSW3+87N0CIZ+0H
ZhwlnEonFXAMaoB0ggGoKU4vJI/ztFqCX0thPpJM5kVQuGXKLilCTIBAyAWlJ24W
7WuGdoN8Tkvw4H9e+eZJ+jTFg/k6zXDduC8j/q2DowxPlJuFuZsRoCCd9xskI56s
yXeI6G2p0aloO3txyEDlByitczKyEATiXCbYrg+butRlMulSMsRAEu5HFfeq/+d6
fp7uQlF+Yz2deBU93AM4NCECYNnUmC6/hddXJnDAFs4eQwG4T3QNbLSrR8wdoZsc
Jt0LH7yVwjuTuBzXV92qy/HIJNHYu4AtzuCP7gMOyl0wERGea17VZrIEpwNM7gBA
bwv40+80SD4vM8mr8eG2rWNN3eruKKy43B5cH1fAA2deE/KwFa/XOuvhyLrR+R4O
nzNbVJqC6gW7NF5GyjUVqMqpHN7O8hP3mQJzLrFEQb+5Hcpp/BZpGAZaadSuUMtk
5vfAm+20eLcdVGCSnUSxldwlUkY45W/7xRJAqyGTcqKend0ow0lgQuMt2Icv4wE0
1o5QwGkTuBakAqscUuhZ4QDO6kNMlG/dAER91SaItIu4Yy22FP+U/YG5DTamJfcn
0nLb0Br0oxoTtplQithxdSEB6J9JLGBkoFViWkAwcHiYlE1Po/CEv3nXCKbqGs/R
GlCEVTBpkfW7ntnBgAfzFhqT0H8+RZM1Y/iPo/RZLC5e5AugkzEFsb6tbf4B4oPZ
bIYvFSo48R5hQruQ7CvPZLhUyaFPLoeHURXsHYpBgWzPb+V+B8yleOCuVsAO0RYA
B6aAgOoS+zz3FCvxZN+yNWIsoF4yumOG8GOR52W86ZcBhkucLdcsyPndM0WWLu9y
tmHJiSSwilsUaWd5j6kVNcxZq2gqLfGAYYdpt2DiWmtwGv68aukCyXQ+ltTQeSbs
mGityElVzoKUkWp1EsbQ0rytm+X08mvFxVi2fm+DY+0d/2r8QJxuf5KPbZ3G8Tn3
xBPY8vyCw8TiwXhFcrCy1HP7X1z1LzVHE4N6SMlm47Mr8edsQnTLtRBsHPdU2nHE
l1u26mqhTUIFt5p4BQ/TG1SivuLdd0FCevbe/wzvYe6BkB1YPUh85ODw+L4EkhPo
r07L34XwLUBE1lwstUqfyU/BjhlKl3DBrmWz10NouHB63ZUunZdlekXfWw4CA2hP
sDrzsslpC2IJWeD/PRnfcF23SNni+HFXTvCFZNqVjOiqDjl2O5paY7nyQ0f2K0wU
/8Cnpj4VqamBWyOzXib192WZ+FyWZFg7brgRp6d1ZU0yPyf7i6el3QGMsQ/W0PJW
9iaLhRY9fDwA8ZqJlkQeOZWx5o16XOz8Gipk4C/5BPsU6VMI/SfthUszyy5kdN9n
SihkFb2zUzEd5yMM9tinQlJJ68XYGxYuxuyuh2JaEoFm3NL9MbNsHVZRR7TlCuQ4
aZ7hdeH0VxkpyJFLLpd5hekxF6w8ThnfdwSiX/9H2nwCS0A7ZLP3ZfYOvDfUIyGm
9Rkryx6rVSSRy/Uw8t9UpbhvxVbCdfy0sGzOAdyEUH76u4Ohb68ki9jD2kaRIP9C
Np44YDSabmJjcmQ/NbQxCFbV4h7SLxdP+Pm0TqujEbOBQUynP52JUPBiwf1ElE8w
Q6rQ3aI9E+CC+XtPD6Vg+2AAOwIasgwbCtpE0d+lxohDRkLdEmkxg6bR3mcJ0d7J
TI9iReGKnAyhdXQl9gtcS/W1mIYAeB7HRT/4cYKP15uzmtKA8+807u1MV/BkFgje
jG7yoe02swLV302yH/nc+CiiLsfUC96NaJ31eVG7ksOZZXRuCB6kivAiaFqOmJF/
f20bfmZsQW3+b6lIQl5/kmH7UNwkxEyGirgKn6+NAcFF6vUQ4lZlLRU84AZqM9Te
1Xpw4wITKBeQJDQsDfNJpHgf6fmH4LQ6HnMvDAaVbpPEVXExXuuYcEwGWLUZY3RX
If0tbU9nvYmfWFOBpayoRfGz/imkEFbSOwg22IxxbX839Boro+DbsE/F1cc0YeEd
YyRyUHr3sWc9q82B3scs2RUxmUzjTe4FBPTkhGK2Jghbsj7pkpbJujZJkCq0ZJR3
34RWhRgKSxLDWt1zPUZ9J8MBEK3ezF1PwH9ylk+FQz2gI7zLj1cxWpTgFi502Gfj
qAkz3PZ/jP5jGGzINqxWnL5ObY7zcLWx7z3d+2UdfXESWGV+vcM09HuuF8BclvWh
MJXBAaGgsHLzADA8D4whYTvZorNvonePc1Sv4n6yt8sTukzi2/sqvJGhkSZO5aMV
FfOnuARcF3l8tOWXSwKGsZEUKP1+zvznrmipWBiTYUfjkLAC00Pau3hkjuZyY3AR
k96Vht+pzkMvrHqbTSTX4GwsC7OATj+vH2IrfNX10DNQxLkoHywqI2M8ksujBzlM
xI1L8gPA5xGzZXG/zqT5v49I9da8YQXouxR//c+V4pP1iAwot6NunvPMMBM9BnHM
B92OOPTxVvtJjctn4c0xFU8cMt0/K/gMPNuQLMDtGdrsEssNWi9EscDkX8OoIS3m
Zy2DD6uG7Ccfxr+nMCGkSAm0867Z2Dv+nzgYS6MScmLaZeKNrDWaaHjxMgw66GoH
S6M3lapQV3pYydSUvBNc72q68+Dro9uGLCtyXRcP7dY/ddsWd8VPIFFGdi5f+A9T
3DZdUQf4RfXU4t0VTrmZ5AVK9IH9+phI/wQ6xGPe/6V5yvnqUYHVfxjwCwnl+H6k
DbPEqjLDaUlMClU873aVMtABJH3Mxl5rqJHYMkF4S6kNsy6kkOuwbnyUKbwBhH7O
RwhbR4Q4ZQhoM0/Fr0zjpOsx70I1TqbDbFpzcui+WLR+0JrPtJkjZNdz1QevZciH
Z2SoOA2LHUvFXo9UtoB8yM7Xv6SOeRHtUh4BgFldY5YI+iINwEPrQE8YLEnEEBbk
gHUAnzR6nb1KopFdtG+/bWgvvmavW4m/JLsw62ugWTpJ1wZbLI6mgLn0/70oKBAt
Mir7+ZWEJNz6r8QTPnCjNsxW+yxh/t3//8heS4VdpH8Qk6PL8hGhbXY6k0c0pu5O
OKz6F0/+vZOV6An+VUJK2CU1VXzmp2QQ3L/rSiiZinbZLNrzzTUsbi6zjZpvIe3+
lvOEaGu9DbD1gfGYwPStfdalk9pnvHXSzBadqKBItWwlkoMz0D5R8J+Thhe5N2qR
nwJ2x9KV8pFJ3CeA5HDpj7WZ46/S9QtRD4LV2VpS6CXHeiC4BTnVyivhh2llenKC
owlpqBHumVuP0uslIXecU9ZHrCLONJ2SMBIvdnU+k6fbfUpPFW+xRIXkDO3BKgd3
AHIPYizeYXCwO9SiCF8S2IKoHJ3TP1E8cmaeshu9PL9MlhZC0lQn0wV84uadIvd0
BvPGEntrw7o3JUwyXCTfbC4bb+Reacg8A6zXhhoJiIG2u/iFN6IVMbkIETmRoLc/
hNKrrobAmhX135XTk+i27/Mu5FWIngtMs5L9RhIYYPYd7DZBwbsFEiexYn/tRWa9
mOHDj8ZJr6uMFE+MMm6b/rAU+GQdwAcgfJDxdwtWLrNnkzVTx6A1DgeTmc+pyLLB
HpExR9TufL/0GJ+LNH42XymZGdig614b5iLRMOf/+Y8p8h7Ihg+v+Ch9oIg9L72+
ZnyXMIYZ4kt/M2WVx+tFF5AZBQV9saUzCSjnyWI+BuCImLwq1g+8ONF8vIoHwAye
1rJI1s3UpFljdJZ/sXvs60qAs+H4vMGRrdU5lGzKK/h2VMFDfXH+CSOMeIbK1Nzy
KFI3fRaNQDghsumK4HEyC4bxd8LBN2VUrPhmUG/LNL8MOoTR6CI5O2F1NgDQSwbW
0JocNdK3gGweCN7snNqpheF4IxRoT4ayll8hY/Bkjv8dbXSqAVh4KlyWXKrx2tKE
rFmTX2QlEAlMkAqpS0HGQv3JLT7LAwer/1MwqKrjD4iN8+qDjbEJso2A8Gf8L5tN
LV09qqHkiLrWIuf+PcKwbMx6ZlL0wQ9HMGnLfB32iKLutG1DCRZG1nzbKjiIn7xh
P6moZwjm8quxsjZaIWkQsyTmTjO8m7knUOk2AxmYSo2d0JDGM8/PFIseu3Ds+ECE
O3arV5ogx756IIOj+rbwVusR0IQEu/1ZzPaU28JMyo0/PBx+yaKzsa/0i/pDoBkt
mrZvw6M6T/GeK9tE3pDFrgeTg3jfnUv4q/UobdjpsF6yMqeDXbujDSHSJiQluBqU
oUCmzs7lNCADs2ccCGc4rRdlstRobGcdKiHOmA8kfteJ9OMzeSp+mBAc53VdX4pI
zIfL1sMlnzNcFLvHc69frMHamYkw9FN0HGk3KY91MVUmlBY5ImLxldTV/JMwlgpB
zuozvFrZwY3K2qM3zrqleLnluysYDDBZdnqNWlsZPvC9Hnu1MrPUjTN7Jenhl2sM
ALb8veM6BO2nYiX9i+VzbnhLoegnHZX82XHx3lVrB2TkbV0PVGVMSXBleIb8pZvX
OeIIvR5x/wocsYuTIL76yG6MBdf5Cc9UYq+Zb4CmEs7srLh1qiAVpRA6l9XM4FVK
ZlWiet622QcdE8e13ghvx9Iin7ySQqXJ1RwW1VT1xPnwEQ86BywH3ES1wQTYsnFE
M7MtftZNd4bmwcsbt/G0VnWB+btfiS3XdCi0W4CHkdLBVFewk7PPuPGYLUzsfNAp
bLgHitAaiSoEIluu3IR97LKnptO1TmTMSUlD/79WYCmajfdOv0AbWbT0nLx0+/gz
fnXkYeUoUj76mZHKGc5pcOAsM7z+14vAcJVdM0Q1XFBSfOaQ6DI6vvNShpsyeXSY
k5vIj6h6wrpPxt5EUWwOZdDsQQkqYFueguIdkI7qFV0TiBn3yCpN5fNAC/igFX9z
KrnwIRSXUL7vJJHWgS5BdEcxH5M3NsvzcxLnSVSu2XzgOPDIMx51CNuPVL5SU2YX
FN4dGET5udUmiMiJ+TlASJ0+b3xDSq3TsjR8eQnMPrJEwixgPJvcejG2mPMaltZh
LxpvkfnbyFiFuoBMWi9aktnv3eR/fu1PVbendD3ustCtcc6mCTkkuvNFK83WTvUb
G5E/xzpssYLAopzyEq4USFMYOdSIyzWUnV/cTlEzUQ+BfsqfIhmCIFbsDVrnCF2I
HPFJDCmgdWA7Ap9ma0/oVvwghK5dqZ+3jBC5LS+Xm6VobKTyHNah2Fosy24rebWX
/RXtEWMiZ1Lrk/wTTA9n63ZFMmpMjNUfMeC8z80DuzGxEPFQSZO98uO4SfAdD3ZO
S9FWoVdDCeuuhuGBz3jKOU0d3ZrdS7ScK6tOTBRnMaZhEobCU1L8zBsp5AAlR/q4
KVgKa6MEVRIsI8DlrkjMw+SZ+JpULWBOlGtNAEe/mwEFLyLd8JAwQGLJsmQda/mg
W7kfu0SkK1VJr5yPvs6QQsyFzWbaXDgSbkn4LzOnghRVLfZ6oUWBOvJJoUef5vWN
VhtVaFyy6cu1Pz/R/9yns0zjxE+fWFRa14UMDTGxhkz1rctJL9Uq/fxVqdWNoLsW
9k2RUdESChKdCu4W6bLBUG6AvK5AZd12scgBZfWj7JgVqHBZUuUd7L3TWMs8xZF/
GLNmxOZTx4VVTgGH5UpAs8wK7m/qQoG9kiM3l5rewldAdW/xBpVyMv0G1/5/vxLE
/Dd5PkfUV6xnsB6kYvlieyfKdXw3j3Af1z3S62QVhm3mv/euPsu4apzKTmIIW4d0
ygc5uq60Ujikqmra7LCgPSpoyA+SzvRdyKOq0WQeUU4xkxIkeVMDwaoGsVTup9PA
fpMSsnNDApTMQ97Lmd4NY2/KpaJu3aglEDROt3ZsR9ohiD/zSru6FY/1q4ffjLQF
ddVwaG0XkH+tYvmLbXFUXxDUjTC/z/w/sEWdjjZfHygJxt9ZK5IezkxXm1Gj+Eep
eEIWEc6Tvw2z/QBR/bxAxix9o4rcFfyclNE9IoRfZO0+WqcC1dYexp2+LJULsN2d
PxiKLKWOybKRBsJaF1ju+gzGg7ZhchLkGD/n2UukQlSP9SEstQfUyR6wHznmCRSy
SO4m63GJ8pdA7X/Lby90b9e+v7trTMDAZagHZ2ZxEIUgdIQTeuhrIJWJ2FCZtVzP
eGqv1db5/PdtBnj1qocZw4jwOYfyaCGGF/FWNmljjSd3V9L8wXRUVjne1k4UChPJ
Nj8ZpOWeNJBL0wOjGe4hMJsQLGSGQWDv2htTeOLd6zvmxFKdTuO53n7ecFUhrwPC
+Vn2eH/SufE4GSLJ9MYQk/yW+ZP6Dlz4tmFSBm5y+Lx/PyOGduJkaGUn2Y4NWyMO
KvcXS52n6kOqjrQ2sHhCsPFX2Xvan3S3ooIREWo5WhdE0QsQM88mBNRzXxXF8co5
EBJ9ZAdieAsM+M3UL6aGz3VbfWVBZ3/Sb/xsvu2WieHTAawTKVAzxi84t4aMcGvj
HYifZPSWXz3Rtlwvxdn7E7e9T3175T7vIDgFCT81lCG97NWjTTv0ptPirPtjHaDg
DFeXgjPz6A2DemKbuDI7uDcQ1Xm7rUUoP/3j1c90sVagQ5ZLBoCkCU/dtls3b1jr
AGp51Qk4H8XmxU54bgBoH7TvC+UabAgE8Y0xRjgZiU9LhvIFbDFHustQ4rc8d4RI
IzsDwL/Z1VOn/5jAB5cJYPEJ7efTAk+fm5aTRDPSr8XohcrfVXoRRiz5/DJP1lvC
Sf4Ay78uj3B0BB+LJXkkhKqDhnWYhIHGnH5pZXTnsd/p7dWAVBGJ/qVP2NvzyAMh
vgScIyndUi+OoaN9Bf8sW/PO1gY1of8Y53Hf1Ro45tFdHPs/lyt8qA4XI4xM8ngp
IVN8wkB7AZ6fIDYGZCJRMgX9YQB+lehYDe+YY/34JceYAt/TV5yym26TT2bBd6NZ
9FynnLVMXC5EJ0mmRvd8+vW1acm9WqTxD5omMZ0P43aakQYn7UAynbKh8Zc8tFW8
JT+pSGGIxLnpVzovUqc+oPte35bnkFPfZuLBIJZfAH9Lh5Eja5FsBGnsz4LbTbbP
L3zH1OisZM7O3DMy1+qxZ/Whm9329odIeKGBk02FrjFE0O3m+JZOjKoCFid7vUpv
Fe9hsPegQ5LftSoUhkdFOsbMRzR6lXw/t3iRv/c820FArJ2T86mNGfUggGqA/V0G
yMO1n15amSRER+AGI/nScIa4W56YpAYcBTcYOSlLH7yvd/h4s7dO0o1P2BAVL/AV
9mtuDfX5FgCgHKvZB09dYNf+5ownKoEbC2tJiIlX0NkzCUURiOcOOAa4I/6VmMkP
GbzdfH148Lh0ouLrSG+ITfBnPnFkQHdHfdjKZ48NmU+9aQD/MoqXnLAAXipAlG3W
Lc0cx+B9PAgwrdAKGnTuP7Rapu9qc31qRuhk9Ui4HtnZd5PrcUe5Mgcifva37EcI
FBks83KeSfHUTUnmDPbzqWp53hhNy6p8udECCEiTT6JzQukEsOBm8eQInDc0qq5W
WopyMJND0BcbJgGyLTVkAkNbh1jzLR8Nl80lOH+wyA8IRzCULtX74jtqRZgfSwKd
A0Ou7UPyIJcxmgBz3QbZUwH2eaPcarrA3ZE6ZhJVfHj+FnULg0CLnqQi0LgVJ6Qo
704MuxJcRJwX1Gp6o3uS42+Q2672F6ldGq4wcf2Yh8E7JOvUOXWOvQqCmkmC4LaI
g2B51oauOfWlty7HbVEeCYJ4Cjm81OkaATUklABo7p203mXmQYGVLT1ySHKs85WW
04IGGJsWTnKwbkbLFdw7rFcJR0fAWDuyM/6KosneefTjC4N7LlKfIXhwqPSjeB79
snoQxNkYV5KB5LrX9bRBaEeroG9qGnKh8LN/PvRsBXiuhv/rHtyx6ER0UG2PavQD
mS2tXDlN72WJyGfS99o3IBazzUkiXsUUaVDfR9G1Uy4zkLahKrw7YxiEgx8ORs42
eW4VFnZaSjL/lGG7ctVMkepo/zURwnsfjjeKlYJ7I9qIlX9gQsSBRhzPZftoHa3j
u6sKhX4VfNFQISBmEFxUQtG+6TX1YS3D+xDYG1DTssVl0glgbEP8BkYjtOLz7IlC
KpwY7xsNnjFRG3wCYg5g0pkKW/CwTab/eISOAj98Kcvcc9eP2StT4mVL0teLv9Y8
W2xvS1X+h8zbk0dVzn6ZGM+FgBe4RNQ3wbKKgx4Sgl0+ubK52Xb3zWuOwI3bVHi9
sZW4xc+e7iNeo+6KSPyBIEyvu1ttYXLekbj/DsIOe8WyuJCiAwbFIakvAmWZT3Yj
O2V318sKvG16GvltybnLC0igDEzP5FiPmhjEaRJgmRjnD6eCzIW3PFIorLq/RsFE
SCcvif/pN7gcG0E3jdPOnR46iTaD2WrGr4BUpyxdlvJuIXp3Qei0jQXVSyBNfw/G
EwKvssPycb6qWwFB5BTEkWfniC3PcWm6s6HGZdccoR6jxFtuGZrpw0sn2W4FhQny
NFjEKVeBCJmvTqOHzjyg6nyLOsk200GkGHS/849BitZHSzH6bBcpOtSj+mbCz+hF
bpHkxLB3d19SWR04tysVZS8egSXRuHN0FaSTvYhW7VjaZZ5uapHPzqmqGLpiVLXs
Fju5OdjwbEgaMgWCbQAW2wvkKDePbYHV/KeRAuGFBBgnlpfS00rn5OKEFT/4iLJD
k6DtOp676LXyjxAN6apLQ1aMN/wRgxUhwIt7hWQ0tnDDoVl9tJE0DmOa+rTHi3PA
fIm4g+cKweDhj7IvktdNZuC3mCGtgHUNVlacEYzMg4yeGk3dPlyh8e/7KpR/C0Jt
Jj46kJGxR2QrUEDloAzcvqXmNWZFb2ebw93UHxQMIzGewFML6iWGkk3OZasHuphB
LO3b5sHYdacLqmnVJTvg4hZWTdZaZQJXArZPPqnnuDPPSdsAeKCBPBn6kNYBWosK
thV19rp3+vZH83WNjh2Il+Gxww74rOctlk4D0+aLA0UMcn1rn1cxLQ9DcuPApDyx
Kmkr6PuA11s0XxWerH51B7rNJ9vspU9nAloSK6/jZ1HpHSoO4bsPQRf8IgPXAg5V
EjzyZHiUo36YDP7SfXXvY3SSSqs7QCl4jM6KdWAsEZKN8A+nkFA2/v4rvhpShd+4
H8N5mxu3H+ahKKCI7bSbVv8SdxizxPx3B5gOB1DSbPeFH2WzsB2osK0xfLDTr2nN
wh2+XLIueYTxS5NimfwxwGi7fG97NCr/rxKUqOnX24CupeBSRuQ/NU6XEe2Ljqrg
5KwLRCV3Z6OIZwJQraYcz19N+bpSim87gqtzeKHRIjYIoeEh7tJCiHCeLDdLWdbt
EGnXbYlh5b0a2gPeyetH4Ir+KRdUCEUc/doiwhkfVXRN0IpsP12mYPM67O8M2YG2
9u3Yjn1qSFmkP70gAacir0n57Jn5Go9V7YxFp/y8y5K8CEGrF/1Lp8FS6cZlzY6P
bgK2rrRJgGzJjPtsKzIJg9hDrda+uFLXlt6YIE06bE11CWxph9G3UeaT4PwKVmUE
L87bkVMgh49H9mK1+6UilewGYoE8Nw7YvZkNaLvUSM1nAf0+LzdOjTLf0fJXPHUN
4ujkXbcKX1pwokEa1H9xuj+e0P/9sH1RgOwYkUJEfyOoI4l3ml23lCSucFOErVqf
4SXceB0rE9iyGy1Ffv8In74ZOsUmBrODiyzOrvmB19GxCCA34kkuDYR0ahMy0bDP
71bAh71wtzcIpBOSBbK3WtQpL9elHKNA0YaWYOfKbFT8A850LQvjbViVZiOuEQOy
N0m1q3AkxoyDxuLwq3jUGQS2pYElxPbu8GbOWj0ur3UjQpAkfQvVG2T70cfGQ8aa
HjotVcs2g9VrwKOreGL1/h6IGpLZL0KBpVAk+xtDpMAHnm906xVIzsnEZuB0URLB
6JfIKJGbxi/J1EYGeZn2ARFWJV7BaOaBKyzwcG6FHElxEzLtOIv2J9c4PE6FLM3F
ChpHIX1g7yIcxvq2DwzBYwUDlR4SB6oHhSoN6z/D83tr+b3LxTJwoDTljBi3s6TR
tcf4gz47oiWkEDfITv7U+1qpaSiIkxVuprhTE7c9EikSrgdI8BsjUutNPsfRV4Xl
SswZuwG4gVmxOgb7w/w0PrqqLMlRJNmAyxe0a+VjSxZWx9wvxAQjyLE4EKL2RMHg
PAkxI7QWi+fNfFWiO/Vc1Jg1Dv9hUIseoVZEUHOLpNnrBwVTQ/zgE15oOjKbC51N
kdjCFQ5tuZg/F5fpCr8hX05Tpxrf3XNhiaYcw6mhu/e5xr4TTgWT5dttoDiWMfBe
zCa9mG4l67MpvFQEnDH4LfRkyIfO/15XgPDdk7WMHjRUYaBpkvVyRh/FODbLm/Gd
ttjX6UAH4vjngHYCqSJ/7cXrY4RXVw9gixZemjJi8q1cOT5pfGWWWng7nySG/+Ht
+vHFrmJAhHRZoiLdj/BBoIDYfBpZvXIbL7Bd78xziSgNI7HWbOuyNdIbI5cYUdw8
AdGbAdPAA4coOwSsbUUSvyJiKKZa9JD972Nh71EIrtZtQUdmvTOhd8DADbTei7Fh
ltevTxNt1jRnhfy4ncFcA2NyOpbS24JKKtyz7ilJujHKlRSFP1l8wzTE7pCW8/RD
18zisl5p4Q45KhZU/5Nwb9ZTXPAyVITOntp3ILC6JEZbnrxR62j9hC3R0iPavEDI
WTUk63olYXJ4amH2QjTZX+VfyYLhI54hWJEXV91rX3TVOXr9eCDkR9dPH38Uno/1
5CU3/KOl6Q2lmrNzkhzvU8j/0sWucmUgxlm4txJlyCUy1x1xuLs3/AQnb42HsNHz
+HToRcLBN6lPWCq/Wk4fQObTo/3EmG5VIJGDLQ6kIVzOQo887YPoOStW8HkFZmcc
m+d+iUr4QRk9o2meWIfDjdeu3Zb40PN+D0KBEkvo30M6kQv0lH8MS91G4v6UsXEu
mJdn4dyYH20yxIcItrONLNoARhB0HApew+45+I2cEVoN1CGWOrqig+Y/tAELWT+m
vVBWHYRcO7/LzPCJoFuE4J9NZ80L7jQA49wUKH4yh4tqUgO7tx3bkhNwwajYBqEr
yUZ7Xbb7tEVCeq0b7Xa52XD2KotDwH5w8OhUczXLyORbjRqftedmpm2YRB/ze24Z
L2XJee7yuI84qWvCGQkOsXpD8GfmzxWMYK1T0H2UyD5kH4Uq3lIus+/n7pqycfmS
ui+U0Df9htLLlaMpGXlWBsjif0olgyti73YWp5ahjWrodFFiCslX7+RaMnoOdfnc
CkdSSEXQAY6JPFI6ZQEN6YLX8l75ts2Kht8f6Vmr7+x0xXzWigcibQtMYIL45g7z
Mn6W4O8NV820ebkKaBhremo06M/W+vhRoC/HTKgowb+laBo+fMKK7bQXHimv/FEG
k2Uk0y8QaOIXZgvtl6CDI7ZOJlboZa4yc8S+WNPzNvi/aIxUClMDKF9mBhNIgcqw
4LPRXRZtIan8CpB7JFzI9SLUFe6p0WZ501iBa8u+pLFFadrU35McfVYm6WB7iz61
jgh8ptNtGjPxl9G/lYD2dQ7tyidVJ9Ygv+c85Zpmv80viM1QqafavgEG+LNpT99X
t0WlmPfyrLa65uByHiZS+z/WsGRKIvBASTAQExv1BDd15zpQmb6K9zbOKEFCt2HK
Zwvwm3HW5J3hrUGixFGOZP0NG8cdaeS+pLgnbr/x2o+4xh9Gt8RDNON+Am1F4VB/
pJ4GhV9ml0Sn+dn+ekrjMPBRPUYDrVonXOfRGr0Sbk5DdJ7iHbts5wWUftKW3WxU
l02fS5zEzjcfn/5zDHHXG9xFkYvWXV+0Quav7hbY249vrYUjxUkdmW4oRwiWPQo9
7I2udc+Qno9ruxcqx/pkSr5VkOFQjLLg3UOAn0EfnBq7V+/q6vjEVTseAEtanUe2
2FGd2tsmVS4NqOKP1S0tDaTNw7CS+970KuYaKEDASQ/gQBGk2a04N0zZII8x2nQA
fnzjd4Qmuijo2HVVckpUbNzRO52+EN7tWrOhVqM/d2VGgzv7uvXkSOqh9jGhl+8L
9zeO/ZJyh4jtbdqR6UKpAIjxqgBcQSj6gl4o2UtNYqRZ0h2vMHmbVP9qsPRJJWGU
mlg4BALRiz2/bKkc7kj5+wuvl92ngovTSdkVt1PLiA/3xhVnHe4bdF/ii4pRYK2m
Xf+DoDLN766+cnkh7BD+R8HOhTPbnGEpYLU5MIwxlRjMqwrMAPrK6A5DkwonSvj3
6lOEDG7rkrGLt54KbftYVQ9hlU3sRKzg1948ymoqo7nz2POsM5H9qKQxIplnM6x+
Ui5hGtHQ2dTsX20no9VljPzQO4XPmTMArPThbNN+/WGwLWhzlUEobOin+o2DrkXA
d1wBPpZ/jA9xFoaXBXZdR5qnbthuBkPF4ypSqZMsDwyAotDIsqXge4IUsfAIKwCL
Wke3ioi6QoAjnupiMBCSBWhyK74+1rKsfthsoTaD1O2C0mwywpaJJqeeyApsV+vT
3VG1XNpDYGHJgVDlmf3FP0Or+pcVYB1odyt8xzjlYXOj7wLaVlzxW0x7CnegAW9O
Iv3uKbsmVwvs1HcRtYx7tgRbiHjRkKsVc/JydoQPUHa3WLpliE8dyxNK9GL9THll
biAWKNRQpoGzDWHth5bke9Onc/gkAlhYaZxlsn3pybjGxeU+cfDWqicrzJQ/CHCY
ba69a1e9VcfsHEeaV24RzG3/SkpHo7ddMb7mNG3BfUOG/pgYih+fzf0zi6D3/47Q
vV8hXis/AFn0nmFrVLjy9kbmyc9X+4lYyzLzVb6jZS9HuVmKJ/BpkA1qbCBV0FxY
GF4f1qm3FdehA+Se8feGvKypVyBjVEXO08o1WsOImMIFDs7K6BdbHtzqFykeKDIE
2rKyJ9MOeodNaX7dhS/6vQQCv/+IBq1b4v3fkiBSJsblTRrIRx/eDJ+TeBu7jFtp
z87N89J255GOk5KzLuAI7ZSG5oOE1ZSoWqjxK6+VKVEqc48ezRGNTA+T13m1+LzK
Zfg+qBtnfVcqlMRluzDWwRosBbv06gjsWq2BKYRq3H+UhGAAMgELw79XG7JbUzLk
DmHMzm7Pn9oQrf05PmLFnW2ewWuBbx/tV2N9iZqnAiE3NLmWuYWC06INdMdJhNNz
AtwwroFmSWXxtZPYr2n79eIvgcirS7L8dX/1lp+bwW5He5a1A9gitTpJGxJ4yYX/
28BE8ZQ89I9KQL75aCB1i4qjIGo8PkdbXth8aALQlrJe4MQulJTGDgGfAHgNM2Ux
usiKftSKnFkaRz/N3+zE7RO2JyoHVZCHIwISkUG0/h0EndneVnLOZjtx/TXETBJX
BLycLresx0bI2R0CRcJdRo5qt1eMgIxi4EeohkIKl86QpRFgAbbTDJ/i6YPhg7Fy
viSiRzFKiQG4rSbX4E64QF7fiS2OaSAQ5704IkOuydYWf2ERG+o6/FaU2IkpdOtN
Man9tOy5f6S6ehkj897OgTnzcTuhQtTax3agGQZu21qgh1VkzqCJrj/um36QgC5w
NqyxGB+OIVqAtGhE/DRfi2GOKlavMlCxu+BI8mqIT2F3Zjvf7YuKeafdvtlnKtsH
nv7/ldK/6tf1EXsx95hlGJttFRL0XV6jEzB8ox0WC6GgSU3O/GRZnwRuRNyi6lBz
DWAELyONn1cW5zgId97kgED7ZjQyGycd89eF5C7ZYm7encZyhkxS6w3asux/isgY
t+cphXP06CJVubZXmkhc3iuIUVNBsz/edhzsnQuZnqXIGUrxbBADOJ8ZiLwCTA5F
p438TdJ8r4lSYa4LfEOJ/LiK4MJ2tRDgkgLLGL3SZLzVp/IF4m1Ha01EK+roh9Sq
5zU883PX5FUNvF/zYZEbsG9qGWdLCey+xvnHyIXOmL4a2Te+vkAabvU8DbG2dwC8
WdB41BINJa54++iFi0kxPjf6R5EBb+gpuMYXAeDn7NbtR/l9Po8j+zNrFUqqT3/o
nbMDKvygZM5DiEov1Hnf2GqKbZfIAImMZ17k8TG3O9oCOlmSvLTbIHgrxjNEzDY/
4qMfM+cEmCPIHqInXpwPKOGKd7bdGCCXUw7APgGU/FR99eJ0Gsw5VSEJrui+g3i0
4IPW3h8DWh0wugtk/hVsDft3oT1rOj+ujhTHMqHYP2T/QrwBhMKZJYvlDLUzxvuV
m/OVRDkNybvLP291MFBXEt8xBPU70+lrnimlhIRDdod8rUXeqt5DoPvVpMoIBxGh
tgKsQ01sEgcuvpI/9pdhnzSQwHK85ztVs8XgXNO8o+mWugjyXLN5AloUaT1bUiQ2
eelzrHKg1NZ6Ce7jjds//TYCSclyWr6yR+rmijuPvJ9ytl8Y8/6jPiyAMhY7dDAV
9DtyQAMKCJMvdpAYtk6gwQiUWMJb87sxguwnmAv0BKS3RjUvrjUc4iDTo0VaL0Cb
1aMbCoXDRKG+g8Y0Tuaawg9Xl4h85Sj4lkVl5By8BuIXQ99BqUG9VXlFJWnjUULS
VIxtun/iOVIHZ4RY4Z9Rn8bQwB407MX/Qc8iBLv6qx2+GitcFSwY39OEoS46miuD
s2kpR4uu1Kr+eMFYDU+sTSc3DkcNrmJd26SkXGqavlAK7B364pEY1gOMH/QSpLXf
dQWziFpSeX7HrZRoD13G2jutD+zs6V2jVjlIlBWqAJpiBp9c/tPT+gPc9FjlrzBr
aA1GaoeuGpcygiy+1t29VNM7dK5X7u0yyvVFGHsjnYf+Eruqt0GKDu7zNv+YHf8O
oeO3JKM+Vy6DWOadxVNcScee9eLpB7ZtCEgFKLdeCFExmN3W3j652hCFUqaKvH5N
BIIibkRorTBokoTVxPDDbVk40dNviwLbco2aODP+lGYO05b+TNrVA+CCJamhSLFA
kStWB5nv8hu3gmslgH2xbqHG10MyFY9/7Cq5p9wQ68DjdITqKkRhCTIK3U92VoDU
A5BrsWYv1V1N42V0r2XR0OpNBGCgDTjMBsUIiSVAnQ754Ty+9s+RIsAoywoQ03XM
xv1W9FrcvUozgzP5JYsz93KkgDa79ULuR3qoMmGx3zBrmUnbxEFIwq+G1v0Fqrzy
IDv66OLdqjFtcsQ1K/mhaNjxKv/r8FJRuvyame3NQ4olbGzjfADlD9K93WvbIvHd
D5pAEqzsgJutkiqKttasealX+8ZXxwq6KO9OZ1MpQVsLd+H4X1nebMlzCsK+8gLJ
EiLxTOp/D3YX/PaaEmR75v+binjhM0H2ZCs92Q9FzABe/C3xgOq9m4GEkyt5vViB
UCR9Wn3I8KvMurxD9BXEBR8LVLT/B647kR0i+h7lXyIPGwLZEBVE0x4XlOaw4IRx
n8g3k8dQQ7dG0Vc+4rXUB3NpgLa5sLCTkNYZRadGR5dnuNrtlUJ28248Ox2TqeEE
zZdJTvPLAbyBFx0qphltqLeBLxhFh5wD7zQqC2+q6Y24UqOFazdYjXsuR92ilZvX
f0kFcCK4uYeAfveKkqpfEv+4O0r2qKPj1SkipcWlbYR1S50T4qeVJLHI2jtwtFCh
5f5yCD4r+7WuNz9KH6qfqLYHksvDf+eNiH9AiTITY8qRh67LXamVVTZCGnfRGk5Q
+YmPsAinPe/FZ1zlAZcNT9lVXF1lVNe2FQ/paOm7DoolgNAdWEgCwwgMuD5gmtWU
VWUuPxRS0KI4O3HhgSFroL4UCfvPkLes6f9XFFIjmeR3fNGkI7sj3MbySVEDcEsa
/ixnTb5ITQPFfAmewcoVLF2LzsA8k7+SiWWZCTDEY0IbOn1XQuuWKkstJCyAXgWW
Ly7LaOWJ4O+FabruZJ8Qw0GH0m444OUlkW583aeWZkEHEmx2gyGnr0nNMFBC4XX2
HmULh8+HnM2ZywipvHJy6/+c8/C6luIVKmadS+kQoELesw7uLAZe44BQqTq46HBD
EpvQ6h/jNh5so2YenqEHbDYHddcAvdfg3hPUX4N0FKkMWzGcEyWz/gxSy0W3CeOm
nI16FRFKI9RN8IIEruGuzf6Lef0VE6IvdUeuTJK7kZOypfwZPddoaPaRn1bEljAL
VFEXmYjsH9NJQ+UMFjEbGXXTqi6WaGNVX+aULScLE6gIBJ698bTwOqvLVkJwPn+6
BMxuP43yvUWt83Q6+nM8PZDWZV7ao2jw5+xFEvBYGtiyG7XVcfnZNCQFUIpo6zKk
W/ABNWv6BMPqKmGMCjQi/qouXCPjQJf9q8IctoX59IOKIZ8ZwyqupvBdte5KZNbK
BVfTM3W1M5jNDvrhXutI9ja34Nfby/Qmx+YwlkGpjmKEWHRFD0AEgdjWUu+9K+iK
7oAhpBsd8r+ptDv3dGcsaH/Xk2P/OP9Ir478malI9oV0Q5WD8wxosf/Y4C5DnhG+
BALGGefwBLePNfyFIKXgCrSc3sT3ZTZjkIwj1dq2o8FHrS1gnTetsgWhI7cq6U3s
BbpRpfgFv495J1oL8h1YzFO8ljYKh1iMKh6ARcCbSDLh9pV6ydmrrCybAasjqUHY
yD/emelnP44DxOiZl+6XrVRPzOJxkHoe6nqsRVlGrhqKYb81k9iBjYNIPX3KyHpw
hB3DQufYseQST/nfgekPrtgzLE5K6b+d8qFuGnJZ9LFjXhvy5dHSJcoyDWZ+PZiz
X9t9qRPfWK1eGpFtQ2u0SJS8g4rEYCd+vRE0G1aDff0Qn8k7PWpqO3+CgVg53ggP
Yfvp6tvmz34RLfPPqgd3Ko5LhcrDiBOGZtNtkunFurVeMmNqd9YGiwp92NTgK0p0
2Zme/TDYbl5DV/WM3KSvQ6d2n6ZyqKzdPtohv9sYN9Clg04rGewwEwsQ0OhKcPtG
drmW05E0DGObkz1Totn+7t7ChUWz3L4orvOavLWMAfAbQhsg+u151mO5B/IcZAc4
F3R7d67n80S9+6jomRJ+qP1Oh4CZi/mKDtL8FcgPTpQC9VxKbXQopOWInYt9ZjSV
ol0sSvrzrRYyMHi4kqNpTmQ6JrtroiZ3xOKl8ydRf/Ob5K2Zs6CPwrCyvCXDOCT3
UYr3iMrITNNrgFL3stJXTUHQVK1v6pai5dBic3GYGyu3mVZULKrlq2e3doNWTP3Y
0ciDFRWeZWLAUBo7jKNhA9Ov+GEu7gL4Ak1+IA2OQtjojEjxPcYXrGj84HCQ3evz
sn6Bn7GRO7p8+TxXCSfgCd6Igd2HOFZMSU89hkWdtcCyH69ACr6GDRtHN0uR3qdI
/h8oo/b7YROXN/EDK7+6UyMF8j1DtBLC1NTox/nb6FE6sTUWU+OIR6pzSKaq2wqD
d8OBBKjOmFvTI9OQ+mU14ueOR5tXQZjkH6hk/rVty9DnKq3LiSx/5oOrldoROuyQ
6VOcijq5q2hj07qMl8PVlRhf3qKEPtewmpGkq9r4lpdMsm6Bo4ZscUIeUwjaJV87
7LGu6w6R7AP8Dp1jhxz+DYUN3o/ZS5EoiuU6m6UQ5x6bEqXXVdvnUk/wgL0jTeZL
sp7TkR/GYsH6CoGS44GxgXQzHI7dMJo+TPJTY/8r5E1sDKxBQHyG8sFvNFs24pfI
ddkUtp5Czc2SalsW5bcycJlBnq9icjdOgCX9evtfZE5bCRJiI/AzY97p/nM8pkI1
l6nMTi1W2c92aZINObFdcimPDqYPBr7G6avDiheuq5SGYG9xTqOv1BLUFJC/gOLE
tWBpX+8+YfudMHXek61W5UbQth079AK2wN1RNpWN0AvScPMjs5IW4pDITNkQ+S6X
pgHX5MBOVViOONlDmEpOT1bJeT/uQSkGzWzDq9R0shq98SpXiV9ax5pcFGpI6VPz
JTIZiTZ4XaRVTHbstfiT0jv8ZIxTSBihVg7BN/fZ2Aw7V5nSLwJE+09IgUpuTRa0
EIDhsYjMKVGbi2FAeZnIjnqJWeOVWqWo3xYPgvNZ51j6cB55rZ691yyLA26iiC+B
j3cNLdwPPfOtrsfwdQvllQNAAOjmnoklRpAImGVqwoGn2p/EQQ6U+Oa1Lcbm6oTD
opSjzdYltWWo3lPpAjb4UhwYToqfJ6dCTTzNeDTMzGQkq15QIwzjuCzGezOBCZU1
L7OGZSRRRUWwe5o3VtLAofRhN/mAG3c/3WTDbowxMxxXdi2cwVVRPyEMG6HNWqAV
ClCiQwnZ/UJ8JSR/riZfYqIJ9kYe+SjKfhKjdNRqmYhC6cuIHuJpMdY27N7a74jN
LAEcVX/MTVX2Tg2pac5feBD8cK1GGTz4PnDogQ5Hyu00ZcqvYwJfbab2oW0wepwv
MF+KaJyE0VMCzptWkAOM+1YjO3yzXEMJTi5M2hRIrEEqAjS2VCuUbhTsh9OncSm/
eOkOCEzV8cNET4khZ/oMrSWYixZ9kE03Y9yBmZPHKyWPQIiB9qh6vW/PYuDyPF7o
FjPz2INoYz85957UtxDh5CNp+n0Bva3LNqcqHQsYr5vkllrmfAEScsmboODo+GMl
TY6SjSNYIzh1KSNNKEFJw0VCQHDVuytYPfhi5DhF5q4Y93SpP/och1F37cPTJwHV
JBi8zlG89YW4/M14G4sJs82MguWuVVhCRKMkvAujvPUBCeTGUtfC6xJn6DfZs+6f
clMj0H5vM8+2YY6FHuPZhqolMWBajNxee6LcPKRgz4HOwYBNmJylsyjvQLGKrWYU
NzY9OauUt0Zg+sB0UvpDh72DVol05XrIiWHRcXe4HOzZROjNbJEOSX4vW2duT0I5
5aVfm2NwyJxug3uYBBaEJaE052mr/IwrvXQoSkjIGMvzWrWNB/+nDSUX+yCZQPsx
gqAXswBEtnObrhFxdFsSR8y5xD5kTWs8M+8ffjZwd1KqGiSDQa7oNciHAKOYEN/0
ATb38seM/gtSv6yshDZttZPv4j31GK9NH2yk0won+8YDOIvp/Jf9Utp6G3bsysd9
aPYHkNEJzC1FutfL5UNcxBtIvcg5tXyyHlqYWfS2A5RBr5VRkRrZ0dczNoIYvJTw
ycHkuVb0Kiic+VG20xEdLV1kyAAFBnDJnpMSBp/JCVXj/eFZvAsR/aw6j/Nw4XQ5
oQcdJrlIP6zoSPGsWwRjwShzkkV5NMyJrRDaZ/0A66fhxwfbS1DD4Vd2wzoTkXsb
yTQzxkx5mbp/h5o08KdMF4sTmMd7+5i4lIp+Ox4dt13Wy4VBQGqDW88kSvWTci8f
7/L7diAFKO2A5ecZuEdjcpPmA/NIl7R16faCB+pd5h2l3GIOO2pQoy6bLoMi22QK
JcJwFkRaH5axTS5s9n3xBomoBizwIWMxgE8Hnsk0wFCe4S6B4xBPY3MltuKNN2kY
XIZknJzR3eMcskPZD4h32lBVQpZ5K1606li56ChJ66FV0JIQZ8DeLBy+ca9MRvLA
8E0Ytc8MtmuM+Tq6hQDlY4dP0d9yPSiHV8FTUY4freh8rrnxpynXOKIq+ufybKAi
4h3iO/MsoOfawHPZOHSjIAAlSNzMSwQz0YLv1hmin3Xb0hxoEJPdaG56VeZZk7w8
yyUtuJFitTeUbEwHmT/uq1OKoxpFL0X1qHx4bnnEflOSOYOp6ovZT6a9okjCsWke
zN5XXV4H10EESzzm1mhvqmizCELIis6I0Z2Bt3rd9xEe+rjfBPDNlGret7yxGDa0
Y7K83/4CBPUMLj75C2SH6LImrbvqbKd+pmd//69ND8LK1ahA1pS+V00KpVh6f+VS
64n79Pe934Zh00epaeiytUKfdCQ6pGzok8BvaVmDBT2KPi4Hn+c928vDOUgXCYf4
i8YMn3JNI96mWo/PZgveauVFGjn1GHsj2odwmWAZb085E2od17FD3uZ7BzpYwG1t
Rm28esRCYIbNE862s8ZSUbI/FBxpECoN3MTvSm9QoRbzO5EseYVQ45qTkvuHTqip
VwZPNUG3tiWVqvWIyvVA0anB5xbAY3H62pZXYnodl0AkHguFZNpZg190/88EnbbX
UqRZdsIETk2UA+XWDKQOXRzTMwVqX2bcN92xvY2hTQ3Uvl1re4P4vRFd3bHlJpsU
e2ilFeGVC3Sh97uXXXF5qaG2h5K7ssZC8Gtxsd6pE1re09sA1DsXJib9qDOwXZ51
5jpiyN7WiYNarUPBDiJ2vSk7Hm/ktSGMS4x2mYw895Nrcbtz1z0Bpx6Z6j8qoM6s
BMdO8mDFuMt/9i13xrV8MShMcuTkB2eVb9uf1jRVVMWp41EixRBs99IfVnZusidC
dhjTPlgwVq8n/timCVBecTmyozwwN2WJ6Y6Zi2kVv/Q+R1aPtEvqxYXGkMnkXLHw
BUzHEUwIZVneCQeukXaVve+KOdQRugrB1TYz2ZL7Fgd9LwrJj66DIYdmYye1z+59
rp80xaUSFa0nLCX/UttkmYLYA/XanDcqRKxqRjBLAWVXbD/c5wxl24vaX8LdQx6o
mpMRuWzTHY2Bog96oz+4RHXmYTBRi75bVDpy8yULHpi+liPnW3FGipiT3xpZh6iZ
pBllQVyakvtf/m0T4Chr2yVhQk80NsBJ6wST7whr42hcMGmodYcpOuB6r0BsXP6q
Um0iO1cGky/wS0e9bU6BPH3NkNSeh10uorh6tq+qpBp/mg9hw9iJzrhR1UCf/g1l
CWY1oykZ8EGaiEmEWwQG4CWm/rqWa9L8eytgj4Mw6sVHKNybE7U36TZwL11/IdeJ
U+81ajwxS6oVX6Yd2SjvJokU5+zE50FPqi3zJUiamet3nMGXzaq6l+Hgwa0rCJx5
LVND1WlPDv0xARYounMWy6HOijY8ZzG+grOVYBxq3G0UfOq3lFyGHZ6dHj6UQ7N+
gTXyM+lNg19eczeSIUFTyDgpGTd1cxZ3Fozxf66lWVUXkAOPKgX0v4OPHWBctVcA
PuKKECVb15EC6oyrtAf88OeNEexew7OWDwcj6zs6akbfBIfo23fgt8Aj3er05cWg
Z6s1S6JT8JUv2LrTRWFFklXdqOsoFtoFpmFs0oiW3yVYYfuEJZxY0xQzr++xiTAB
z72X6OmBK5VECZGriIKJfwWVozViaJEVo2HXJbtxlGpHI4ZNkzPLEmRYfJGkarp9
BOuRvd/xL5rTI1J+2y5aRwOvbWv+D+8xCMy2L3b/6xu7MCr+OgbqN+i7igZ2lAF1
tHuB1n+r5MRSp2izZxsILWaXStdF6XEK8PuR1kbEXy94LvaGNfb1laPOGQQn6MJH
qVb+evocQzRBvxUMhCMTsxorDPPSrGZx1WF8lyxjcGJ1PnpL6rRJ86M6+O9e0FvQ
qFXiYDt0L9J9dKTL2Ek7txcRSHryOMjWNpk5RY05tMYNGDAtXPcxJhjzFBbci+sE
7VLJnqM1bLTM6mrBUlxPqgLfokw3MWRasrAFGe08sVA9dSL9d2y6N7kS6MUYZZyh
kkFWFJ35n8XiUla1d2ExJGeJHHEMvVaI6Ymgn0deIm5/t3wMxrywfRmPXLxKrcUf
n6u0kH0SYiEKj9EHIEeZXIdUcOg1+N7eGpzoljZFQssvZo2P2elyCx0AHY80UHTi
Hz/Yr/nLTtjfRBpX9xptpR/W0D42cZAUlXx07oi8TRkzGU519aomEZTmWiWa0wSu
yBu4fdh+7gpGYubgBIg2i7yqJ3WIaIEgnzAED55JkMicT9RYzd22o0x30Jm00oKr
RYYfvQLJgCdTFzJeNea57+j++sfjobpjWTSg1Z1s7Ms2Y9Xza3jnN/RbzVI+Uypr
WaSMQIZ6oOGtq10xpUd9R91MmdURHEOBzRcElWCOE4suW5Ty+ZEM4HaigbLDIlbd
Kv5tZqaA6FSyWt3kDF9RmGqjHiB8CvGlSD47OxWHfUH+PhQC2nm6aTMQvCDPWxLl
b+2Uwb3P2RbsLdX8XK98QyLkmN0M1ywK7VDcpoALjqVF7WkHXqagvY9O3QKWOgd/
FInJ58HF1CDJ83+3GX4kUCqxr6Qwby1cN02h044z8d/0nPYFrNoitoGRtbldFIIA
PaMXBFz/ez83VOaX9KufIBxir9xnYni1yAUzjHfNPN1zRNM4CGH8mhZZOrOhIuxt
0KOHONUDzhx4O3SPMk0LXBKXNA8fiQZYauRolB/TpbF0xR5vFDSIL8INJeT2///V
dH6KX1UqIyN0wyhsC8+WjsqymrCTbj2mbuDO+0KpkCt9uGeI7CzjfyDaSe1wYXLD
jsKGywWnDGEP+bIrZOcgEpdGSXYcL+/v/D7ph8mhdONrL0VLTWrsDCVfdc7Amgtx
ymgq3QT9wX9YosSvyFXb1HI2DABNaINSMChloQUWaNJ8DFMPsN2OrUUcJx8TB3xu
RtA5quGb6PPnebjUj/r+MpK+hQbnRK2OhsqR8Nv5hYkeHmmS1rYFvOpG4j3yIjpa
UK3ZfeUFRAR/LTdk7K2eh5dbJOKi4ruFS1BtC5tcCb70OaSbDvrfR8rCwq05kbDn
KiX4NPwdK68TxqsnfC3ZL+J0ojf0OOIbBj3xS03mb5xprYXjH/wEBNscpedHSjGz
qBmlQsedOFA4QiCWIUGdgeMbmd2jxaId4f29qC4tSLQ68ZDxgJCyRL2aDmVI1eas
GtuXp1X2arfyzmpWdNrXQ5mR9RZjyTECQmuGG+lyjlud/rADg9tzfLmnnqhi2Q1w
fBm+/Yp32rRQj37VHqe+W9nTttbmH9V2+cZzsE7EYFCErRRCfxODa8TZoXaeuCeH
SGNZHGq8CzRMkBnURahHflbKvQzfdTNPjDOTGwG4XgsCQEsE4n66Nwqvb8XVkMl4
+uDN5VLkjQ1YyLahupLVj7IwdTzGAinU+RnCAX/Ay8CbHoLvO2LK/W873y1kKimr
8L5c0tPHO+prhb6zDSj2CsbHKoTNm0fGm3hyw8bak60VO5EnJYV3/Nu1kTrHankT
+Lv+UP4rx3Wx0qcqsgkvaZrSB1FrzqPZN4r8U9RyJ7eG74+pPFN94B0gBjL1YpSe
OoOYUxfQZLUHo8b8v+EDjFMNFfz6dHUqL1KYXTQimW9PSOEN59KcOtESiT323s0x
Gm/fcgmoMIxX2thxU5ldVBAO8aM9iICriWhnTjCHkhI/BuPFyk4/hSqitLQkJQb+
AbbMCC7c8Ia+gdCXCg4LtSQVNxVppFoOx7MsDWwu2eZp2a+ObRbgJtOG7YuN5YXo
Q4kszpwfXHjLS6w8ekfh/r71R5iodVBlKUKEuAySMUFjNwgzsrzQo2k3kJQDRIiy
Cd2GDkCXk5BHr877UBgfJYZJCIz3J8xHhI6z/QhYAKZDR1eoDF8tZx6vn+I8C2V0
8ii5Jxb3MZECP6fDCoLboXoY+kejhGAXizTzLKL/XXnVIVyIlah0AjryHnvUe3I/
EfxW+j2PDVJbUXcGXJHRlKYfmv9ECBjWXqm4QOHWGU3X5v985kBAgMmKxa963uqx
BxoB5eSLCjkxvSWkCbkZnAU6WfdD2cDoXeqwyUADHKlxrJc1cebCtCihpxkSP4q4
7SUcRGPLhMrEIWl+U/pyuV46xoJag9Q5DSSyMT9h+PaJr1D0MYTk1nflFL4DUMH9
xo1m7c7CgsNIcRLsdeC3Y/uCZVZ//qBVRQ+ZH13gTYVnwkgxySFuWlfV1swq9JHN
cFO+zjnizhOS3gC53au7hRJ9WdG8kVxLJ+Vv2SQtaegtAgTmcLlHpzTUm3JeYlvw
HvSE6ZzEuR1xp95GaX0NkcNN8Kqg8c0y+HCCbCVpB2zzqDhWLTsi2jhxKveaOlqZ
7N/jAhX3fcP1sP8LPN7h7CjhohmY3bnKFtMwav09agveNPpDcOXqU0yjo3k/jCDq
1KTE6F55/U8YlfTAddCSQAPhzkCAwYRKIl1oNpHopCS2wp5TD3BLxFdtzaFNXSR5
K+wUutghxGDpX+MlhS7st+1s8gG+1g/TFjZkx8jW20h9TsQFBDfIXC44tw9pmFRy
/+OwP65ubksMmYTQ0dNaAUW6N1KZAIg9FjNDiaGODv/ae62GWCVmRdfvrfwTcFHa
FUS0ICUBvPb6Q9+NWO4Fa0tRvhpjoe81cOmYi512IIEg1Se/PN7EVd+ynXgTc2kT
X1WxL64T/Hbrx69xEror028YRm32Se12m6oLlOrB8KTrAv8uultUe/dufOZHvrlS
cS6B82rFSPeZy3C4kvnKE96cPWJ49cYdOqc1Vidu5nHo1/1R/4wd4zzBVWJOoHNY
DscMT97o3j+bpteDEojr7vGBBK8N08EWeJIwBaKqDJlIPf1w/ctZmfxL8FHaWWbR
ZT1UVtL0yvbB2sRZE4VRnFAYotCGXOrWqvSLV7EI5T5NDaYX8XZtsTk1+pwED/dj
IQATFuvrKzCfu6ZAa0vd9ony0vqfhAwaPk2RxafkmJsciUY3xhju7mzD4B/r3jkK
NVN7OfmpB14c2ff/JwFD0jcQplG31T2xkpiCKI/9a3hb0izmmOGZqV6FNYv7e8Jz
b7rBTSxMBqtnVUoCJm5Z8LrUCe1oTxtsZJIREVGw5/8IfwaeTwivz/388wcXPUiQ
oB3l8JSqG+Mzm+HyuHW6DgQMjh/zRTNn8sdDeDzpMrJHz8QtjvxNzTYLXHsk7dD2
tMU4hZVsr772tny7CcJFE/CVl2bohGnAmWPIqfiTk/cfBlbP73XEFDuFbeDpJanH
+ju+bef3aYIhwnIqYw2hpqfSf7WkWqI893BykXEWNJ2BP3XW83X5lUOCx+9gG6fD
ogInsMGQa5Xl55VQVFhqHy7a3pbU1ouDHtKKdbAaELSJC345Z8nvKVcZjj4L3dWe
NqlcMaIpPHj9AU5PWd69haSfVegopPlVHpZPsOksLyl2W3l6mwcMafvl8mll3zYb
7o+M2S/AbUBjXtqkVmv0dDYiuZjW/ocKkEAvBL9PNe9ABdsD891Z78nQzGMV+MQb
PnfLgwqoxa4kEzBOVLgZtfUxHy67cING6Le8jgeduYSnqIgCoaMKTHpvlHxYXUZW
Xwm+gQOMWBhTROHfZed3foWJaB7WGGk8itPFRUPV7Zb0IaV7dFMvnkeLUR7flh+m
OdVFOR65QiFj0PC0mUOOhMpF8Sexg1nBPUg9n9aeq5LjOmZa1yXpM9mJNTkCgv6Y
xvLCk42nXL1jVrc4TabprZ8ZBrpkMvl0m4cPscxnyrvBMcLPzDk8G4vjPNCyqpk/
NJi2DKo1wS3IUVtyUAUbAK0b7vkh8TPKaHRub49/4bBkRyPXzDkziy84m8MOQl6m
1LDdGXNq6ya390ovER208FJFMlfSyTaohO5PuU/JXv25lr6abp6G/iIuWKaojSMe
JNsrq0RwtXYcgCk+ywrMXFSYBw9eur+ndlw6j7q5e/m52MEVCpI4XWHE8Vf5tATA
Gv3wodHTjQA1hhoFdLUudkUPwy5xGkGvz6H6VcFDF+gdODzTG6layOi/Aby5ylRy
y6oR8iPWZoSFLsCKFkoKidBB+fPKw3bphFyPzhEMHFOkMN6NBgdb1kGNJ+FwtWiA
oyjtGNjIf6q6JjUz83X3G03Rc77EEubRplaCTVqqw85V5Oaop/khbFWZXmCPHyjs
MN2/CCzbZgalB+XFGYUZlnqa0KrA6ZOmgYm1Yzn4CGYi07n53J98CxhtgJ89dC+L
q+NlnTRYty3YjXAvNGQeEEKFghLShUouDl6ctJC04GNcS/1IgeypKOfq4FHfCsIM
XLFKZDBhnngwioYsw1rRyXT0tmfuScl9LP993ai78cKmQQK6uW4movfHL2zs05ge
UZm1VOLd3UNflkdw99XE75Z1t9ryHRrxqkRiYY4ypgK4UKYfihoBC2OrFVgusMpj
QrKW1/s8iM8kcVQB1OSNZGMbj1+lUofi2eYqczKuIQ9/crhmB+wWf5c0JwZqN428
PGKnYjWqLBDZs/3otf+JNHS/UY1Q+3tl9pETTXFXzBvAacgoUxz3RFJrfOAF8esX
MOZld+cddWA2223OZw+pd8rE9vEm8u8WZeToiZsw1L4kKPRTVoIUyzFRkguIYHQQ
LWkXlKqvq8xqEaNBA4vvHYpjsq1+XkLBgu9YguQ4wmKBVCWG9oJxqQMafJrxGQSS
DknrdvACVL7qGhllHuqZkqOEoBSlhjCvdDtpLBgYw5zH4h/a2l4SRj/JT4vfrN6Y
D6EhsthHhFNYjhqZcQzmw10kDbbJjZDer0IVDb6tcaAXOgVFTozcS7jJ6tXqp+uS
E6JzvAUs1ARZ2riErzUfpBJkgylc7EUktHxwYwIqd0o0U1LjrMwHHmtUWYqF665d
BuSNxpp9eBvLiSS/UqiVLKEcnnJertUSjAvWdtxZJIt1pL1NZBs+CPwG47EVkB/I
h4KJDGw0JkC0FsGn8mgCgeoNcLsjiK5qf4SYg280Zdn3WKqwLaz0JvNzz1FbxgGD
ZLUHYRGfDdj75dg65Oqu9wFkap1SE9iz3Z+HF0cRDs0YUDP5zyTXr17AvZLvCACr
gWZHut7LTFMis/Ywl1vF/Dgw+VfUUKFcm/ywGNA0XfpdMDoatNrxKhswV72RQkfJ
4y5GqpQmKGEyPeUEw9FfkjEtMDDvHuithxnmU1Y/zcr3/oruYRGSvHXArVwT+V/0
CGMngmTZSLZnurxWyvvMFTFi7dhbp8QKkcTCPNC9x6gP4W52NbuXYvHk3yKlpUmI
rfmhWBIF5w6FOsXUIRl6hl+4SFOHK/5i3r2PsMi9DL/IyNLnWtdWP1xQMUAzATPy
V0Uprp3ar21dLNH8jo3NwcE/p60jBBTUTxBi8t32aDVZehjK4EhEKJPF7l628TmC
pn/dOG+lUJkOCiEN1G61cEwPTKJMTwwE6trYEc8FFoXng7AGRm0xz4XsjHmz5wSD
q+yH17vcU7mgm9YdUhbB2dG95rEYaENAd+f8/VQJuWT9tMOBgTNNw290vY3wzzUd
xlDz66VWd6BTcMjoMFKoIoWHfOGxbyz61iLDz8PcRP/gkBQqojsxGdWhtC4R0mcw
YM0sw5DUuW0fijZ5+RTIT3A7ey8EC308mwwCKhQztTJlf2bsljNQasXGyFkr8E3a
RYsFLMD9S6xr4Mbw6LquSV73FELAi7T2KEa7C3LWTZa/HF683N9pytG1rSkcIFwt
lGurKjYfBSn2vMgWTZlcpltexaDCr7yqTAT6bv5Xy//DiV2XsfK+uIdmhRp7VcGj
SHyCM2oiPJnB5gbC5YnW8aGRvU6k4OrLT6M6ryxBvUCCJlbZ71V0bgOSQxzuoxzc
U4qZZsRK7yGw3/oNOiAdyvFrq5HTmogk3dWbGR4/HRQql2d8pGOEfzDZ90phajPI
J61O3INwwRRCX6Ui3zc7cBHgq9kFQ9n8OSMuWHF7aURe/N4tWUz92mH9ulkRigxK
cS2K3M5f5tGboTPf3esfa/rIHcbp6aEoQJ73NKNg6oi33mMKen9zg8sQoYUv8PEq
874bl8HXqAe0rO+Wo+Y5fLY1XCF4BLic/lbvsIf0rhifnRA4wKgbXO9XFlE6FNwe
7GSpk6OL++QAT+gmDAkCsDs2BBnpIiaV+vgGo838hY4Aqx0CbPkLzGdZ99uZJGW5
2pKoBm/3W5Q4RPuWn1st69G1k69T6SnjyVfl41QzGrZfkHJnnWxDXVPXUbisDQwR
DYYErsUJedm3ykuk73RILCG+AfU4NWeghCgnDKktUCtSCnv18OwgIpfH0CwR7j9o
kJ8hSnxgs+vXSDNLL5gM5GQhOYt6y4bcW1yqE+G8KEPphgx4pm1xVkk1akwQbVFv
iamDgWT3BSkbHT9Il26E8zBwEgOZBkMmYViwgP/9CWDi8XfR/D+ugojaebv238np
j1UBnmxYSKloWGPxFkMdOvzPkIV3uOgead3ee849STgQb2IchGRYLqlbmsrbdzFo
1aMZgUL2fa+WCjeSmpas5ET8R3HA8njJTEaXSHsT2Qu9bzYuFkeD/U2qoWVVqvDi
JaZo6kwt963nWkgDnTzmfBc27CtWHeo5LhZOp8DMNnVp2j4Y/YGg05pMhCnS8d1g
Je9ywYI02zO3sLSgFXiIDHKMwKblq9xE/DuNjSGaIxWLfSV6G0Pk0xA3M5vgpKqU
NZYQ9TZMBqr6cwxX4Psew0sHD/uG7mQDcJ07ypdqTXTTbLNYZchRY7EBWgWg1JR1
v3QCRruG3frEm1L4xnsoyFdMuHfZJPY1gGlyAIo5ioMNbXeQ62wq38pbmLJpPKAc
Uqg5H9FAw2cSjGq3G/qhBJGT4o2/l1JzQKDTAtxX4nARq6xsCVEPcIO2wnrkppb5
2nhWTcIOBjsb3Q8FzFV5dbMibml/SJXvVT0z1lrPdMlfVgLWh4nUBS7qDnMd994e
/gtbfndC31955o/prtElBdPw4wcKLsDcYdpSTTz+ZqbcpgHb+LUjAp77sS5rtu/Y
VFokf6mLTjA8JJG8LVMt6itK9UB6qRvBw+mujz9vikhka6f69dR0eCFWc7nOjZyZ
r/VXQtqCs0ZyMWzhroBuUCcN/nnv4kfUpsi4WX3qlHg0B3TyhDrrmTa2qb3Y0hLv
N6GEUL+t7nBuW67ROT2+lqLHsBhxEdhUC9ThjqmzMbBr2lvFeHGwqmXB19p8KYDM
QFko/W0pc8rYJXpdn3tm7/ssno+izjN2yXlcY5IwGuk807n0+qJBl47ZPQi22/+7
vSzafLUm9YcAUUItpxRKk+raKcijyo/u/csImGdJB5fgMeoVSLjE2E3iYoqPb3EL
8TrofMTI+c9V3gdzlxtmrCSCa1MMsunC1nv7qHE3qIwLimEFejAnkEJxBtj2xiFx
e/szS1REz0sE/bleEG95BQXb3xIUwobPTkYnBtgHvwmeROgMkBIK/CYPBhx6cAin
uv6m57jTYCyq/4G3pJhomt26z9UQ4cxJbCASP+QduNZDhefMa5ONAylld4iSAC8e
2iwD+BNFhPlaK2bb/aA6/HMnPInx0cq6R+AFI4cfVwJeVjvUjgfucEjjbc+j+NBm
c/LY7jTOyIntjva7eoligu5oDLq6+Xpv/8k85aSiceM+2tjexpZSYTxr3UgNq4yN
W1FTbik02VjV/bukIw4UncxkZbAzSNDdqoAtGki59zl8DdoKXd1H+wAXQ8Suln9D
+6MHvMDvXC/2S+m5A4ya3Jn21wN1C8x3DouoSi0Kybu2UWFj44Jxxx8v6/zGrutE
X2UorGLUlOOoIA1FPDa2wraOr8iEXPinJhTm1lHSPR2u6e4dMf3yWZG+EuvSYvsZ
bPuDGBYnIzWNWy1fWnLo2a91WPHsS2SLVBTdbNoJ3RjMTvaATjeBwDkk3D4GMiMu
QLKr1KbywAl5/x3VLoBF4pxaY8Lv6/BcuymILv4qH7hjRdzRfIlbQpdFzEDD2NCR
ND8Yk/jpO8UFcGhuVLiFx2gH7wwK9eVFkPDY9CWi0eJd+TokXjA7QfmoRFDaLjhF
mwt0UCRL6XUvs56wvO6sw2q8SFJ8kE6DYiiWFcTEN9SdVg6vZawo9EU+fGdWfxCC
mE8Ji99C8fcFHKTfY4i6ITK7Qiw1rjlZOCntR9RVihp7jLw8JHKaFBrHKfF/qevR
GwUiKHLq9zzi64lvI6H+lr1M6RQM8vgToqYAea+LgXL7p+BCpAU3BjGkxx07nveG
UBzCOFEVotvegnNDY3RTZyVT5vzQLZFp6rufWDfd8LTU++wK3uji/bWV/aUSyH38
TsjbY+7XcFF+OrbyAkwqBRp99ffyzEp+5qBwRGlI+mkDzS/Sz+hYHufuS5Zs5YY3
w7tBUcswwZirHE1wXuKBPH6BE0uaf34PbB+f+YIkNDudO/41ljRR91GEudhfAtcX
DU0RtavZ0fNL78xPPDy5eBbzta2mF7R/kdw3YHBCWH9OHqgpAJiB8Zh+pxaup4A+
EW2XGd/B49uBmxDqZj1WrcPGU7iD7diDP5xW8vRZwFJIQMUdlTJKXWQjkvwG7QnZ
pxkRE4EriX1RneeQv5uCGZpMcGn8vwsUOMw+LREbTWxjJQiJ/awPYKQ6ZV5AUtkj
0BoJLEv36dIBg4Z5zZkkaUFUfQJ2O5Qf6Dzc75zDwEmYR79gjqK9HIg7OpTrV+kc
VuF7NBh6J3NZizKxJrX8Et2V8SVrXyDA/g6Ls9ETPeCR4grTLSqciTrmi0sKRHAz
zAzGoh8ljftKV+cnRezqiuy0QCxwNuLzwBg5jTFOY39xydKyzh1T8fteRYQaJuIy
yE2ZLHUK2iEgmxmFosKRJUttv83ZISXPHCnaOAv18ggWHNBoQum0r7z/z1kKVVun
zSnpgxHAt1miXv5FYDqrmVwy1EbqwoLvB30UajYZ3JLRGC3BItdUduBh+d26wytF
SsMEw1mmle7sUgoZazm9+IhMe+Erh7+ur4ahMNno0NccnLNooj2aZrf7Gm/uODFS
PJ5QOYtp/+gfSSEZUCp2qV9SoVNpuOs/lbtEu2bAT7FvgvJfvUjuSY+mnWdOweTu
lf6M+KN94HaRMbbXbxxmsv5dGmjJwFb8SAALs3wcsw2NKt6puWLDFjdcZYl2Wjaw
RX5tgC2ipp3TUKl6FV/YYkKuPyE51S/Tm4ipFtYDaU8KE4ZfOGAhNWiyT9J/1M4n
Vwtp4WN5X7wc+NqKh8my8WQZLFzsC3UtA6J1IVWI0Qr3SbeWtuto9fw+jm809KQi
EDK7YsPToUKyQeelTWXA8FBFDRGfkN40mEpxAqjzOmL9rGmOxbfuRYzxpXt1zBkh
5CHnfG23OCyCR5prZT+tQRwQSmVbAlAMs3HtSS0YOl6VNbqXcyHGjA5gzmBm2CjE
hFzNtfAzZRtIUkEYoxXohB7KxEe88QLWCbreG7kUxywMwBinswY0TlWxlbI23SDp
6SmdnS4x88ddKY7pu3pWJiWrUTgXRibx9DlD+bD3iqoCUEL19XqClarelt/crMHg
U1rO3QCh9tB9D96Hl8ye2onwv7rjLXmC0hDnwjyu5XR0oXtQykh5MuGJPTNkAI1u
Nlh4gwpiEy0l5IUipAH3JRa7NSyAvmVhSIingegzzM/vU9MXyAqVyhIG9LDNxQF6
czqXvrPQ3A1GpEJRaBms8q35Lxcm1agQLBHdOXXLilBck1WoBSRAoG5M+7SsVRX3
dVBmn2Lb72vPlem1RVuKmPgdrq35getMUlt9SJW7xvQylPgXDvUg4puGq/cMS3nC
mZbbBDMB+hLv+tSMQvszPchhS/9HhdSWtOBAlXnKDviTVJkZIB/BrKcqqqLLDBbQ
zbaL/vY6DimhW4aMLPSb2xdmjJ+TwBWe6RFkfg3zaE5SbKWR4sB0lw2B8lHt+Cec
Orspwd7QMjkspztKNx+0b0uhluQ29QwTxpK5j5RCtIIo/p5YaqwtqVGpDfh1Nudz
q8CelHHtbW/ySIwwu2rctizb7f3uDHb/8ZU5YbShXAGdlj8qDSVXbRKdJ2aNZY6K
XHeEMNTgUcm3YTNHZrgznfNIoI1VL3vxDoCYvsnjmt3LmE6LojxKrgU5fRXtzLGb
TshjPDTRPj7r6pSvCB6Gl9ApJdKeZ9J9ut0teObxHNJbbuvFkljJJJNc8YKFdLon
q2AP4HLAcRFPuAAja9uy9tNWv59v1i2IeQBu6GUDvj/F7+8gpJdf9oNyV+5NcJ6l
ETQ+wARYO06xC5Jn5knZY6HljbXciH/feeh+5vOfbykGaTQ0LS5BJnbQbHmVYIm2
Zqnl51de8+XIdmAMP4by8eVJlYKEa3LQUlZU8OmnvyCftFWF8FgT0s2b+F9l3GiF
/jNSnmv38w2X3A777qX5kPKjI5wnjHknEqek1elXK95LVioyugyouB3zMMWXTlcX
HXROAopIKHHPaEOk0fyUrWAqVbbNPXyu0TmI8oxMnQ0hPVB1vBxOpT33Ra0JCbBY
aFaIki2rxb+MYOp0xyAh83QNN2PZWlF/Kk8wly947Jsxcbk5dWf5bKK0s1d8W6bC
rOIvImMaO/cBrAvqm132N4QxvDOlxDcYCqYBBKllN65f9BlP8CYBX1O5Zj8payfK
IhrOSKBwGCtfIzdAtgZT4qzlSSjZEz0GjrT4Akz7qls1v5yjAob2KK4uXldSuAgE
rq/Xn7mZpaIJGDmzjb3Rqmee9fO07KvDWvKdHYqxjwISWj/wrfsJAc82Aju0/nEs
0Y77lUvdJ8o0gt2im2jBIPqMcnRKMkQ3f4YZMFzWiYE9YVJUZxEYfG35wppWDraN
6+/oDfi7qIJoAFQEnziG3xhJFDarqbuLGBTEVjBKTwxNqQzQZbIS7gUuxdhodJZd
6HdndWpJa/ZGvwH8u3jcnKhA5QPovlAP9aDovBzpQlhKf0CymdGu4BRgaupVLtz5
Zx+xUyIg3X+CY4c6lhqojxZhKMZ66YcV+7dlr9E6oOEljAsuVk/5ATSPBzLZwsuo
yarVdge79ghOmNqqUOSdtdbEnbjR3072DaOUcXXQGM+SmyN7yPkLseljtr14EhUQ
X0rDcURkk1TIsCPyGjqOYYVlLnjyhJPPyRhdXmAkFH/ohmhI3CIvaN5CPZIwqSem
N5HRv4P4W/bzobEVsoEmLGPJ7BazQrHnH77iiJ1S+R3pa4uVTsNKZvwpiZ47aGyn
b3i81p3USBKwNMShKH8a9DVrwV6dW2Ez8yS5TyoyMdcR4DHjGZ2ZN0eDpcRqqtKk
QJbGQlEtwLoyIVWfpeY6ZiiZuY/DhJy31eYpOduZxVaj/u4XurnWA1WariD1jCEp
K406SO4B71MhAGt/iiP21/H/ide5VrGx1VWZzEABx40N99zmqrozsd1/6edpYsjY
Jk3vTDadApax6GUIQyn9ODe1rhCWE9gnSYH7J7XP5hTzGDsfzug5gPHAiZPR6CD+
epY5ffdxD9pC67E1EACn4R06VgXEIeu6CQXMQpCrnx6iS+Cu1vbGhMmQ2uXrcU7a
AgazVHIngOwJdUKj2XZ7/b04Y5bfNtEPZhLK4RNQPW98EOkC5rjDs3hhTFhPvLy3
7oIfbmcZv2ZymSdMa/Ahr47x6sl3S5rpwR0vSiyt4sCdQ43vpb57Ojqcyl5oArqF
mKX5t2wermhwTwEfMlelt8gjG96v/BzhjLBivmbP1fEiOAkqFe5zVjZKM48h31JO
Oovj5B3XpTayDLDaxe23Hd5sVnocsiqBGwMcfrcflNeeVqg8jyiy/zjXwLx/BQU+
w6j2nKhnYZUHdeJQDyyvlqv9FEzCxqScRG29xwqUQMMUh/emr66YdMQER8JWO2do
yieCjLtWSPoZS2gm/nO14NZ2L9qYfK7/CoAcJUxuIta2K7HNQS77UWfRbmpyyJJY
c9wio74x3YYWf9cp2PFjjQbkRR3C9UGnrTiFpSKz3dxIIRSHNgq7f6OxXQbbuO1r
wZwxGtfDFT6cvRBpJWQjISF1VuvZGCMGc6BFrKfYVPpTWSukYPyQdygOSD562LF+
9s/4W05FCAjHVpU5zzhfpI7K4yN6+Rojanq5QCn2RHZrlep/IFIBMMUF7+gi3Hhs
OGt0jCh3SmZcxopOTaPGUXF6F+ToSCZDI6mo976toiCxwmsfnKvy0iW3W7PN1+aR
5n9vVJp/dwOyPQO2VSIm/aVROreQxiPeYkLvu3Fa3TCSE/e/4alkKnCyvZTqNw3V
hgWzkiaPflWzzCY8fl1FYXCcPNtHNym4IveO3PHOLP/ycxoeDxqU08X3p1dYJnNJ
bB3B/2rFvgR0CxV9acNoS2w1SPhqVEJesvW+jZsdGy55Nx51haOu3qUCQ3Bmlw0G
IM2In5NUQlfQ/Hc/81SRtfjRV+n1427VvsAXcJJGaHxTFtwNa2rOc7TeWARu0NVe
C0u75lsMuN5jth39FQ14vyqhrK2X66l9REDewQeMfyPvpxQC3N4CxS7lv6c7zeJv
oewRHJ2y/21krZ/mNVQjfax7bw78oZDgTySSTmzFMSnyMsTphLicTqQ2SCRioHjR
mVIDuOcq/F2fu4/4zJzMuqVw25ZsfFNeNREVvlsb1zenDB25xt0PHJcUwS0kKLS2
uufQAfzClueiK2y7gWfXyvqmhl0JZyiXsbI7Ah2fAxp+8MJDN0rAHD2U7dsMWzER
fCfNGTiZ9lBrOK78c1MhffSBOGMwcHyr0rd32N/rg2X/+bsqO8bDjJ+kfJYpw3SE
7SVDjurd02PYozlT6u0Go5pmBVZdkdEd6QA3mQC+jNvC1uG0iiubTo1sEQ399qu6
it0VZlAMufujutqvo7GaBFEGls2g6u7TYklEHTFYJWG4VbTzwB6bWbTHNrs/MUZA
rHq3buVZoh5fKmHWqeam5yhpCW7KNp3u/3FBTVtZcsb/UYzRxXvMti8PNtpJ1+fX
h2C45ZXDBqt25UQ0aXE1OSb3eu4lJ7V0fCxFVFzY+bQw91+nWQ93JXJ3CLO6uRwc
0ztFfc64pgGQFgXIR+f50Uprt20jTQzxG6cZoOD94q/ddDOnmXLoqxdiLeNkHSjK
7/ATzIs+on0vgc96/kHalZ1tpaUBH5lyIr2MRvBMioqbAH/+wjW/5tGkGFBTbf0Z
ubXI9R9IH6bkPJ9o6SS8yZjGLHJj/TPprFTZp0/YBIVo4ihZBXdHkGdBoOigU/TU
nTRTEbs3tZpQc6cqooId6T5v+h31fQ9QOJGrJhUzbCzjKr8S9hTvfl8j6+GRbExP
UjzMzQe4qkI3S5IfBuIv0XUXCp4uA9Cnve/Pufzx29WkGvswKGEP37iUyn+c6cyM
dxJxJKeMi0RxseuCsXcQOHndTePkRbuYtfH39gbohBAUB86LawqKH8179yaiPHkn
b2bYOvXfD0cJQnjZBryVgOGd5DqX9BBRw6f62xhGWIInrPFvgcDXr3ekdZjxi9JU
yt5tbXJzVVEFgEMs5B2qfgtmU/GBaT0l8q67ED9O6EHnz6Oh+oTcrUnRPBr4aoQp
qEVN1Q7tXak7/8JX5msNP1LoNE62mwQPkCUeIneDgXEi6CMaBwYKM3ZPGrIMnaBv
u94LsesF96m177NlCInoHhcSR4VDoDzGLitCKwAEjVwxDGpmMXUGnz9VaMEELMFb
upwffqCtTb/uioObXknFWO/qKMwYBFLW9WIEWQ+qx6cwv6ZGROxEYTYn5sSJwreW
ZHg1ObfJhhVWXBThF2BbjNNnirtXkvdBuKQT895wZpRaFCBDRjGkvLdTQJW971hC
x1Ts8GBRA18szG8OYIpmBvNpeVhUXLOutO5etNvkaL3IGomkwpPzAExgv16YL7Xj
m8CAZWt72D8kxLOPDnRsQelHmk/XRboGL4Zh1Ekp+KU3NgZDqLDUPPbTh/4vy2+o
Dc3pTHsbIYQ6BkHJPqn5EZEXMJsu90D3qz/BDqpdz21Ubu3SNd5hPCRNm4GJAGAe
Y4zBZbL/lm0uvGzVTs6R/pcYqwrnzJemTvRY8Mof5FUoRUjqyDrHAsju+0AqPzec
LAUmc9bsA+Gx8KbtpZDRN+g6Fq+yYLk1Am2eeB0/6WnSNeEIHSI4i1iQnCCImcto
TnprYXtHBOBCSSTYQhHrZfGdSg+zkGWoiEio+ZKF58F4RssNuMj8uCLLgHRNssMY
DgQD7ozHc9KTWeh/JYJhzeaO2Cl0azJkJ+AAdSYwE8IAojYd14OGoF/xZcy4NZOa
ZHHUC4+kCysKYOpE6sk8C9VeV+PE+KPsb6Zlwd//sRTiQhZdh8iNdPaPDsju2yhU
JTjHX8MGx6MLaozS8mXbt1AmN1CV16A93McXNM389nwd3HCUChnks31d5ti5dWrg
j/TkC0o02Ie4/qnlvWpSbih6Uqpvh1ncc9LVpDZEO8od7eZjJ2j0BEZRaVahz9Lk
QYyI5tL0sz0SidyRofOjooDywl2Y5jggjubkctrhl+zNBWcmrQ4W0cvj4iGbJiCZ
EyfG3wLvLLn+KxzNQA2pi8+AQfR3osgDvlmj2ICZr9aKp25GZ8hpDer4lwNRDSMC
RV3RW5JPKm4IXPrUYKlyw857OY76R2NH/8MyWLh3pKSP7HjmJDrBGuvwmdWDaUN7
yCNm0FpBJj42Jxi+RW1OlZ7xNyTh8dllh0RslWDxvuQfbsKLoORex0EEnCnTl4Dx
8sx+5fdPgrVFLefj/G0MXtPsGWWGLnGmeDUG6JEa6ZzNt+dEGK6ACFdf6cKDiugx
HN9D2+Gf0CsSnhrizFGfTg8ob+XzW1OXBV12IzZaMP6lNlgymvtjAP9oDVjS4xAt
9VX7u9C9SBV83DaJkh1McnPcfNdvjXdLwlIDeT0Iv0E2hyjV0uhJNnz7341jLTdb
8VwvxDtBnuY9WFeIprNAstiWt7jc5I7vaeMsvH5vI604t1pG1CgIy5xjcs80TXAQ
ZDhkavvIRarMbUtmuKK1iDKCPFmwzKjJj/HAg4VeExq8BA3HzAcPjigAmVoUMwIe
t0AMmrNjcaC+mjSVn0+877VXr5mF9sWE3vaygHF3LlK7SUWK4XDfItwWvr56N11X
lEIYyJm9HmmHOcVFquGVyVgw7xb6O59o/rjw0VppQnwkza62340VdeprwN7YRD7U
RDvw7i1eiswH5Imu8iHSTON7k60LzMoi6SjAwOcrlflvMCQ2V6isAWrXGiBXMP33
5s/wkZGuF/5QJbdxDwLlXj0fdOITnnQyir+ETYYJ2HJPZH3b8YlQZH9Yeor5aWnD
x/Ky3SJ30Kld8PyEerSFWiI4dEFyCFkDQlVFvZtruMkR7TWwzeWPcd2ksnGD6p7r
yRaQ7tC4w7vZSqsDnN0GcDwY/q8WzO3yJ1PxvPdM019bAhdpBMrquKA/enyCdPmE
UEfmmiU6JuCW6OetwhLnYZCkdJERp5fM7AzfRMtdYaAbRZUrcdMEBlLFkDyHsc39
ZErXvb9Cgui0EhkdcjYaSJhEYuoD6jEPjXRbcWv6w+PunQnUmWeiUWgiw3MppFor
IKdg40tMLR8ZmMCDhgAOwbYMZCOFCHWefTPsGLJDX/w2rRNWLkTee2meRpGgzrRX
urpRK47rMJxVaCk9TypVz8GDib3SfNbPcUmus5R/WUTdQyiTy+rSJsTcroeoYnuF
eSoyDZ79ON1AHN7IqPWnAKQj/nVfcTm4PPYHBiuUUrX8gAQmozFBipK/8delkUw9
dlIG2q865SmZJbvu4gEQFSS1kx2CGtfytsq9c3jjnwL0IJPYXAde3F9v6KpLCCMj
CF0GhcAXFNzmqfUaaRAVg2cZIihzr4VjixldFhEC+wGJ3CHybowDgWMXbFri8UTO
ccdxNKoBYyXoFtkijZO/ZP/eMFyWUBD59XEykvA7KpLjGRdH1gslB8kOKG3RsFlX
2eHOa04uzzSCoC9Od5h0ChpL6yHmgCGYPvYjFib+3A+CGo854xNo56I/fZZNOQli
uHIlBhWF2PClt3nrN4aR2dApbyZHDcvgOIeF5LJREFRCMwCJAueijbW3Czo/khRi
EmYlFS6yrWOAQf/e+fpF5XnD/UcaS4UyAgx/aNZ/HqMcxOJ2o1qbPvhjJ20QRhOc
cYuoFlQvQoxPAfaaTHlsqg7HPVWTUoVuyYTCLNwcTDBqX0p7vK8x/rtOpCI2cqFx
T3hd/0b3tOD9SFjvT2cc60eLZ2apiMc5B1POAvaeaosj0xcKvAw3bJ1zyjfkk7x9
TSnIRsXc28BoEvWVVeR6b8W10GGKudeRY51zTSOLyJ3O4+DKa87sfnaw/QO72Kt0
ex/CzwwmbUriOKiM7gIymF7lZbvDNzokU2Um+QgctouJ3SUKc3LLbc5vXFXoScQq
uFpEkgCgfEZF5oM0bdkYbFINs2pCdgEIJ1rlDC330ctxfq8IHinj5n8LBCGis37W
ps0s8MFmTZ5cjGdxN39CFukjAoMUqYMy/AUs4mg6leKWCmkytmb5tI+qB5iK2NVV
wJsQ4ZBvofuD/el9BPgtkgwu/asOe/3tPGXu0c7FMsij/mAkyK6AekewJqif9swC
9dbsR19Z6hUMH8xX9bk5KSZPVHdYKd7I6qmHH+GEc9aalMLJ3L9cxYDs+TlJaVNl
k4VsGynXQD8y5+7bl5xpUdKmmsYNXAje5X9oshPRKZDsoQFTKbsBT4dSUXxnZTnx
enD8X8cSaSvG9gEc3ceETgyplkM0g2fG95W6R37w+JeqLMJal5BAn6scPhYJEaMV
WjNF3YzPSnUYvTCyZ5cyK72BNf+Sk4ureCs1wZ2lZ0qRAzOGfbJUMKdeUqzYd7hv
wuCiTJuF/ETJ+RCioV4G2w0WQIcpk+VE+RXwa7iE3VUij4QF0zLVLTTfmG0ZtXvA
ukqmH4oD9MEau0vgKu1pNZPYA+m3ZOwvOhTRqbpC9nLCe+5k1e9bt59mBXwHp3aa
IuozpHceTww8FeBr3MC+/cAXhZk6mn/jUv2+siBsa8OAOrs2lM+YSwExBjWbR9bK
+a1dwwrndj9f0cOCB47u72SIdZU3VzwB2m+E87piTzbrExDHsISn8E9ufvICMq99
SYX58yv0aVBaJmgUT/1725q9+yoN68U68EUvg5Us2gMu/hUSoRG093z5ICVvMseD
6I+V/TujIk7qfNFhykuYmH99yaC/wdS10kQUo0hM9K8jllzm6rHmM2Ad839RPoQP
sEo40/XgJTNcyxWDsHhtmolDr31yDaG37Yshj28FDRBLLzrjxv0CKIpns9nornEg
LVxk68fUe+CfnDh6+mURDHmDq9JbXsOjCD0R6ht46wBimCqC3w/AKK4KHXO7EIsS
4dg+CTThwv8mh/+LRKM3dMKr4ukPcmJsf2JNq+bFut3dMETr1R4yZ7gSQ9/8c6CH
/GczG06oJ5hpBErPognwfqWX2mxHhJL4l9f+TmQe9cSNHB1LQdDiO51gMCwctQat
hz3GFgxV3RVib0393ERM4lvUFYCFT2ErGng7OnJWVo+IRtYsBpjrc+9zkqk8+7/w
GfjYAIFTyHOsi6ExZlFLxBhya7uw/Gj+s2i1iEtWtpPQ/7Xc1RZ7EsqrlnXTZn+J
OALpyQwFBxOUjh/0ounnhlNP6agJisQ9xLb+mxMcQ6L+x2Rd76ly6rB8erlDfJ+P
hwBuzHM63k4Dknwbew4HKcRmo7eUrJOg4Yw53KxUFyiUIMO71Lo30s3fowBHA+lV
NdNDakYLrA8yu/ZvcwF71wBz6l7nFZA6oc1/33rkQD8bJ42CEXDklsK8pHQbzF89
ElqGZkhpTa4dJg9mc3wUxxJtCpaGWAWWyGE2rW6ds2wq88YctZv92/eXbgVgGonR
/jgNrmPbxzJy9PCwynORnqjIkpwzvFfLOnQVTBtQSqYRULOD+pU+de2lUwurHBxh
xxzU/I9kpqZizke+dX0EQvT5glbuHud4dQ5l/Qxzvcy4ZuH3rKPJehZySt2jgxuP
kd/hYt9QCc3RybC4kDri8hED9mo1O6gI5liaQbKqVr3yIbxUyZyflaYi133lD48X
jhPSlWXw6Ey+9CVMOZuRO1YtW+NDUmT5GhWtOYYGjgQFXKL5vRJAK3u26ssU5tN3
aj2f4rZ8uGbddbIVpzKFeo4oYfzD+olzsPpi6M5rrp5My/09EmZnVz8klKxbPkfu
onsW71FOVHhRBQdNfyCpsO9GDFeCkK6n/IDAPm0oQN+67QiUwnhYB+ZEM+hI4GcP
APXxjLq+FdvR07/tpYrhw5zY+6fwfiWukggRmS1r4h+tw+wvTzb2l6CNhOP9ahf/
hc5Q+T5mi9FDUuq3av/JXeCMrt26zTbEL1jWEkGI+BxCILl0RoejVMge+WWcQcR7
xTy5jgXNtW8N9Hpr9ZMePEsKaP8DCPD14ekarYTduIujdmNF6yJH/YmEkeLCvAp4
nulvqQBoHVkgYQqYNyQ6kHN1D8g7S7Kge7dN5gZZ+ka1PNC4X3mxkcYMa9GNb6U4
uwFLQ9wKdztaFSKDrRkIsmMCYAZuWcWqCBf1QG8yUHZeaNZcxTAWt+LP5cxKdkaY
V1YthQMUcXGugu7vYFT8w4QNUUMQNaMDdDEszn5Jc3TOTLE6TKHqy6C8HCOsK9w4
Hqnp0Pgnvn7Kit3vGkDBNTTtwmadBcwYC8rV4m8PV/MJQ6v9ygTf0HKkxPYDzA03
CNVW2v0r2Y8i2ngznBj49LRHaFEhGdpJVClwaThlbU1A1+lOud4Gggs7Jo74vzPc
Kk9GrVlHL724fM5Pa7Ax3NDyhJcDaHFnyJ6rAPH6v5GGHdj5BpQ6bkPDM/C6uEjl
JQzMTCoZedZttdbyzFE7wrVIkd3qqBVI5ZdQgrR92Ozczx9ndjZe7eisPJ9ZXLXu
VkTyMKuLnTpE0MFmYBlxusJ9rlW21vyCwCBdPvGUP8Ukp0pGbJEtyztPVWilK0Yu
HsJMnpZSAjJg/MfT6OAGp25qSyI95+o5lYfHwRDWrMZiNz1IboELya10c5VJST6w
FrQvwRX0m1NjOD36G7TV/9Xkms9LeGk9Ypc+b7Kql4F/lUcl+pM4wwMgGhSsx2dw
ve73sz67xAm9wCTe9DMKro8uUETbPE7adkELxuWs4C0fwlYvVheHdacTkg7xu4j+
WVC/N6k686UmmQpkTlW++ebxB0GMF+lN1i53evdUhZvD/t3fhvheqid/Pn2IUn5x
ahbOwe5sX3mWgVb757O8gaEtyc3dmSk3KRDiakWBkLnBdVTTgG5/jxF0Wuh0LfQ7
MCxgXTxiwKctGv3D4AUeSURJMJ2TTT2Q8ygRimcvGct3nzasarJAdocJ9xRfUgUt
zgflF1mY7wdvRpTqZ0OnHWqtEtpqI44I4/oZxl10QZ6Hr3NqgHht+eTNcxaSRC3H
Yp8G9c43ECSScHNXAUbSjLtMmDfv9XJzcomvlF1KrLI8fxzkgFI+NRWwRKRO4Sw6
A3MWDDPh3NmNSo5GVFpjVeduTGHOiijoSodHWYzPajwPEgp0ml0GYZftEyaSxPmm
39hkKMI2jzTrqZ3GTk2BCpNe127q3i+Jrx6GJORWqg2LX/m/IvF03teJ7Btv+kTV
kzhT50ITJzlID8MLKMt0imibRMxVgUK6XyElxgS3hczl0/84IuiQJYgSLoT1PmSi
n0iPKiSt9WWopno2NbXpi9wjkyTRk78xG8fzFUvHcUZ+HEoifPIIz3LqTRacXDVd
AZ+Em2Vrk9ahrc2Z/g2bDHNHrH8f5CtWM7SVgpYZajGI5orhEDHkBEoccwwJHDO8
1aghwyYueTfVe9nmHpLy9oCRxMuj0UAPp9/+AFOWoKO1L6S2aeGTwAXOG4EFONv6
Bvjof7sXVzKPSoPjSpIjPq0Ao704+xQm0Rx+8GWBCOUjJlbQWDkNPza2CkVB2+Uk
G3CPy+1E3On9aIYLx27hoSYr+fDNFhgdHUXb0vZTn7TfhIwttt9BjzdsW2UQbT4u
cMCmrVlrs/5RRIDI8BnmZAMqiSQpdFURc7o189Zb2h/16WbtN6JqRc7eT5CWkLlS
d88oTLePb9kVaUu1JyfP3OqpzZoUbyKz/R/1up1FaJz3IJzWMypfEN+M2VPjyt5b
HdaIZdfLaNQlv0KR5vgMaBRjRiRHT0W/Z85pAKGl37rKmkyW5pobMkGPNxSyVVBm
hWFnxzSeRvoPBWXSL6tPYbobhkTsBq+UX88KXYKU88QCslWeBHI+BuTHuALgpJF4
vEBSrUQpJagXIVgE6LCYKCdu7mDQgcc9+uI7WhzYAon/9Tjuhgcet+0Pn2Ey2q7M
pkNFEq7o3e9PRa4dq9pqk4cq0buSbkln6SG92HH3AHx9Px0IOh5b4RLf7SGDEYLl
GpTVvJAwLN6JSCwIq4/2+sI4MStYA3Cm+ARjadkGCG8tHGxJuDIStgMx7kwmZJYU
nJIWNd/PYx2hZ2CVEpXnPfcNMnW0dpnuxWUoJtIFsvUDDylLxbVGbU6E/OYUMF3H
D99QCHVFM7LWN1X2uu6hzXoWx+gVPzWt8KPWqlIbxBOvkwy8K3BazdsVxsgjU6SE
5QDutFtCGKZ7yVPfO0zAANYohPvd0EC7ISHjPoOssTShedWbf0aSL1unGRxboGYl
sU3gX6ttVSFEJK61C1dqb4AJpCxDBzloJQKm0U0EmX0hvuzUrdbYJ6NDCfx/OBaQ
YXAd0YRwDJsz+aSPBS+liQ0O4WpoFuPDDZk+Z+dK9s6qXyATPEgIBVblxW9a7FJN
AakbDI9KpCQ7ioG8yt+C7oTI5idhrgb5L9Cygqb0e8e/IU7wLb5wmNHE8xlujWKC
+fvkONaURsFHs+FhvIJqI4D5MkxiZkx6hNomhyUj8n1InIqxGhI9tarm/TgW4rB5
0ydavMBKjVwEahCN9Wdhcy8QoARkbq2Qczu5oVmPuBwylmbcppHOZCvcL8JU6ts6
meh8JeXG/Yc/T+5DLpBLI/rOTNNS/vO0prw/LDPjzumiWeo00kZyKcuwSNoXYwlb
YVkYe3xLabEonL7EmihsytA/LBBdVMjkayPU4iVriZ/Pn1wOWe/nuX1DmJBY6viu
iNdczvJkNLj2H3u32lOTFJAYclPodRAcdl2C3oc3pPRYjNAajEC62NyckfmMwwDN
a0LfHSkEmYPjSipIeVz0/t6zYrDItpUZ1bqZc9VfsXwZXhMw3rWRtl7ijLTr+Liq
24yILGtaJt9THIePLvYw+UA9lFFk7oWQYq4yoMGmY9UoYNJDdTHsZK0KaMjtXNiN
na630tdgUdJ9VnqAPk4sqG6kndK04Rc1jMKnjVrw9VDB6yJgn8N9jk4CzPOgXV4y
AMG+YboAsw3w54HWas4VxCgeCF/FfFf+6JFBv71oThDp6HaNgnf09veFm53tDWME
/TTYpxh0A8gZXcgaoAe4w7fG2MoOpz4U9rea09CWgtP5ocxdA5yxXjU+BBltq991
0tfMW316sO/j+dibF1fIxhB6yYtACXWmvQOBOdRrr3w7V9/7fQWMhN3ZxN6CRHNk
H/tBOYN68tzSgwyxRziST2raYn/9TIXtqgMwGohzTgJ5umM+IptxwXErCoFcfRD8
XobxEG9Sqv7dTLhFNncCfSZZZG4O+hzclyaHwf7Va5cng8V7hkVDyhtU10/Ue9pc
xmqx5y1z6gKJuwxeqEYIESeW4WEokOT9C4mJeRHG5RVOPMOwhregJGUAn+jX3Iu4
sOVEHeCoo4a6VMBNbjQwWiW/Zq+A8+Fipa622yxfq4fVAYfgc+YqSLWNsAGMyeHT
zHQHPNXuidL1ZPaDmxU4nalkYfXvHu32nDPRnkjqEWvUBELWu6sxT/kSexBu3JO4
iPSkonj6W/IY7CA4Y4yENa59O4Z+unnNM56umdMrCe1thq6+Ks2BI90C6zqWaMhm
g4S1CFoaZuvc/0L81niLcQtOOKmZOpe6mmxn3CuAc7RUBkIsHhvSRbuzIvoZzTma
4xQjW1X79I/tisYUz5GPJt2KksTEjsMgghxd2zqe7WxySU0xWM98xiiY2vJTETlq
r9GvLe6y418b2eZDXMDgG3ie4SwC+Ct1W2uvk7dIQKT1yKAa2zkWAiST+M9klN8L
1vBK4k0XVYDDDWybvOEbIlBEuRl58nQR1ZUA2GD/4Qukr2xU0JZEI3Qh1o+msE9F
TQzt2fwhNkT40Z2UN56Tu4bELepsjXytr7HWHjUOLE9kifdVe9YbQcXtOK+WyD6A
822DCi8AlFzm7KDhdwf8Sr8m8X/lc9xOgZ6kIC3tsL+HzwLnhd/MXDA1Fi50XUTZ
Q5zxQ0jdEeN4l8YitmopnrLJSIcNE9l5dRdd6tqt1EEP2lO1PG0CWzmj3FwDPkBk
VB6N+blwunbfeHFggsfXMLTyFoCeqc9rbxSHvzPsmA4moGEWyGOnLtjbuBusuqYj
+I+jbu6XYvlyF4X+/SF6CTCOSRwICHCzGWqrVtKroXk2jLrjT6GURyjLHppj+Uhc
i8t951pm0/zLfHvexj2mspbsZFBp9RGmfQ1tuHo1jNDvhqFepy8HiQYjdrwAnbX0
2agcNujqKr6jNX9OPas4VIix0V4LRuabloY1lPOLiVVgVC2AnoWM05+XijBIgJ4X
UENhBeeWJ0L9CcweY7CuJfsi1r1i7b+CO5Pg9uh9jGUkRHuQJrjns/GMbAZ0rXiD
e3FRvj1cvZhMMqUaHJGWY1SLRru1sKI2QiQsi6Wr5A1DG1c5l247L+TuzwuFBaMN
jtfSc/BkP3JV7FlOUdqRFwJa7H6G707Mx4gkI7GZtw7wX1OTH7cql7T3yShnZ0Il
lzciBKMBuCNfhtKB8YuCC5P70hQojMsQAhXnb0dlMqTMilvcOWf9WxvhV6yy1R5K
TR2oby5d5mkg0OdzDo4/1Ja0r0U8xfI8viLqEdVZO4535eUucnzofsCNSIHar1Ee
cHidRGT5lWeIb+BRklDtX9sGOoU83zHB61cV52f7CoiL1z/sx9hIkIJpONsj06Nl
Jd8A6PhfFSuGk59iLTaqHXrxGiZ3YzEyY4LjXP4Q1ClAs+h5W2rWKNxwd+bz9ERs
7oh9Gv/IYnojlZl0tctyUzZrA2YlZKb3DuZJ2wTewIG7ecHhCxdPaN66i8AdhQGx
QmjfOP4QuoUnz2HiSF57/t/6ukMvRL/PZSrxKUqjgM4x5AChIE77otKJPIkc3+PD
zQRJ40FbEoCz9mozzR9y1RGh4pTaR7L4XjCAgcFBv5WZwdqYdDLLBGxwIyoHGtO5
LKifMMVQR11ncR3LNic6r9MfLxmFHMpYbWAmejuhvBwxRmI9lC4ZEkxZsmE0+XFU
Eje4A7k03rv8ESwuWJqlKc1jFQXInHk6JuLfppisdYPBdgYOEILa6ptG/3vkKV/e
KRkg5AZ4ua069MhwW9iren3tL6YBZQJm8PzQjqIh54NqowpTfKsmDlTKxJLXibHm
XlCvZY3jLaraOgloK3xB9iWEYp3OgtE3z4DpwIsAq9yB/nTQGd+TNo7D87WDpM1u
x6xEov2XJySat0AEoV6Hx8AjXPGW9nWccG6nN1YTto8jLf6JO7D5tOgPTWQppQps
6JA+XGGNM8oNZmW8fS1bMVyEsCalG4Ox7R525T8qahwPNeKXEkIkN/NTV44V6xNC
zk6i6yw5YxgsOP41kAV6hXrnUy1XdClmMWNn3YvzXDMF431h7pCeYeKY32UqLra/
Vy79ezWAueCNn+FAn3qU/R2Vz1ahbSM4Usy5FsoLEiWIk2hl5UjdXdk7br5K1C/Y
DKIthcHOGNAh3g5Q8TfILrTNVHzO7uxltBrLyRkkb/lICkf8S8G1kJ1p0HYb5B+W
SrX4gUsLwVVi86UrWNyts1vNyBcggpen+5fnj13AHlGADNpwVN6plV7weFPQ34nf
o6ofiT00PBi5YNqveZKegPX7GZNYAVd6bUwtXC5J4DUODWup+Q13R9MT2jMO35b+
66wQR/5sL+ZmUUjVAwpdWmoFdGsyimOrgYrmjv0dVsrlS89e6cvagagCHuj4zT8X
ZglCRBSS7VcCnyDczSACFYH4fEBFf3v8/4aTBYHQn9NgP1/96PkxlJIlTCZVSY0S
GurfOrBAYdYnLoczBMT3s/St6NsoIAtncWSp2wN79xca+bU0U9TRACRlSS+J4Mrg
KDN3WAOKae9mLXuz2XFZz5h3vi/hz7UiRiIeVdOU01VfdyfZrvMyIa/rneyR8fIs
WuWVl5uz7Y+a4bj4nEVWTw38SZVjI+EqU/Dc2Mpmb2UApie8LNBjVnbzRb4BHwWB
emkM6Th8MH3uaUKmKxDeaxO57jQuAa3nl8zq8Ry/eketFdJfCWewWK8DVdFcPo6h
XZ2sEREE2RO0f0om+bRKk/aDiI5nuSFXvduBKfE4L2nf+OJduHw6Y1Ops6hzbL86
nk9sLRX61D2YZ7iS2xzfjGWwX9ao7WdWAJYCnB5p03Yh65MB9+r00xxvWnX9dIpp
rhkAvjTT0ThKFFvn2TIce5yWMktmGHdQTJN8ZyK5oqvXyJN5OorQ0HUvn2/+wmLx
A9rX8k3hQOOjqu3L9eEYoLkzWLXDYxKYsFcF3yOUANf7/6k5e8zIx1mviOj/4fdC
JPSvOJUO+oQrx02UTZyA/ovTA79fXtZdKnLzj1DXGXSHJj9pQjLNlnBQZ2SHd/Bf
CJUZ1JDo5WpDu2g4+cVG75J2kKSj9rK/3SK/TSfe03BqJC6sWjdzmuRV23p7Qny/
onv+T96ivC7/eC8Us/a0UuIeJFJ0OEBP3qamfxoXq2EoFuIF4rRcW5tAJCJKukT8
NsoosZcJSNV73FFEfvdhNXdVpDjFELe8wMH5yYwhVfBQkByFzpRDR8ozSiAQwDas
IrUf0WU3SZKFW1Xwv4Ff1D20sAs6wGhdplTQ967h6Dk/DtSIDyj3WVCDhW+jbFDY
cCuCcLoXgSVshv4wXy4uTt9HCqnGRwfWE33EQew1Z1BASB4+MzwU7Jrouiug4r4n
+kBP2i90h+0G4LvmauTx91pwYVlH0eB0mPRHYwQfi/wflmNxWilMmBRfOzKH/AAq
mx5Z0tjGTKlHw03kfqQMjW9rHwdH3MZfdIu+qWPkNi1LThIjqLqTyXYa3arxUTbO
vbMmrvc3dsJyB2Dxfbbac3RUFcZvLlQDt2Xn1/zX6Bj6BfeYZF1xHxGcrhxcxym6
M5FBwzBKxTic0I/g/LeBG7ZCulUHWmuotHqydQraZefBg66MSnmh1JCbpW1EoPNr
eum3/mgGOgYgX/XDqPeW7WpHnuGWPxLgOZy/Dp4piMGeRW6Ed/56FhIHO14iDNZM
BeZT76FYwEWvBAVgtka/DQZDAJLEqAQndpWTLbKSqjbKFDN/YY8buoOVzw2z9W8n
4Zu+CHevy4XSlWwNcybCX1BOzCxMWIaUyTq1QGYQ4xgFHKUdgM9U6NXJHV8XElOy
q2Wk85l2nCoj5hMHfuh5XW+MR7EiVQ2dKD/XMXprEt+hqDwP7I/cWHzSjTgDYqBP
6ATHKn4hYs3kHimYFMJm+FJkENDDUlzRfVKZm7TGdjCrrqgfv8vgYGYh1DOfqmUK
oPTfONHFg4XxCUvRBzWej2VyQ2Z2mHif7aO1kBf5EJxerMNttgFWII6R1pmS1lLb
qk87E3VJshnw0eVakMz9sSOSHOIbAgd3r0qB+t0O/DzFMhYhhAy4Um8njxQPbw1l
74gYFni5r1/aoGOX8PjjnWscRBCIH8z5qVX6prkRryhEcesPxbSoAnqf1VKKLfHL
pwgVp9xe4XY/EI7OjfQL0siW/BL3u7/9Bcs7QB4YaVBDYwWg+IrGKMya99K9ADxl
OyLPu1mUfjGh7kRqAQFHLy8BdD5JRGFz8BrlSlJ6cIqqJGY2qLQ3iGqNwQcbzhl9
QBfkupmh+tow2uI+/jlldA4Ih3Z9W2vYOG5J5x/qH5I77L5KwS0rrnkQ4Clj6GbI
PezgqIZ1Eq8xLCJVssBTSYNHmpsqDZmj6FQy4HZB5gR9j4qp0pa6NNqsxPsPCNao
DggvcTOhvFMrQjgfT42HmxYCCIRmqkYvH5A44EoXLkjfhXXDNe+qWS7jVPWdY5CC
9pS3EQUITMDAmC0AHlotSHtYFqBGLIkyJF9stmy+484mtubdAt+2bimLF5K2RvVV
TXxD8s9xs8PWJFccfejC0HAgt0OSaNLYxzET0gxvo5Wp8r/cvjZev2QWCrZq1mWT
C+hFB3AreMjPJ9wyNbemkwbXXBZqALZZbGHzm6EVL6c0nNJKJ+lji5wToQ0FZ3TN
iWhGVRllfFuPoAA1yjDoBuDwzxmXJedTI/MDFan5nAXCItftq263rOwP6A9SUgQM
DwiNNxaBvI7/6PtKkQmrubpmyV0KIjaxJH9gfBINv9A0gdnq+mfdOEzvrUWOZF07
MUp1EJRPzAWl+fX6DnGfEBLD7cazaHZOUoIMTa8L7Ou6gn28sVgSQi/EkyAMQq5f
TvvzpwB+cQ1MJ8pd+L8zI0Y1BGCwJTsNcPwn2rSbA6TyhB7KuKmM0lgC6k8ifD7L
I1iPMtxhm/Gcgk/IpmToHjj2+IvSbBWD3kqUd9Bg3ODQHo8yckdSXzQiQmbNLlL8
MBOEc/jK1lHOor1I/hS0sKDaWZHdYCk5UYn6+YQYAXNN7w3XbLb4YAZRoR7DfLBk
SUYL71gUTaDSV0VbeOZpZ13gZhCVT8TP3Kg1zCh0Z6KNqjnlA3ZAt/V3xfmyPCuo
TX4PsFp8+7dkzjk8W8txbpo/+h4WV/IqEyPIpGDjwa1o0HwOmpeKeCFufxK40K2p
fGYmdao6dKVnzKxV0pI6A7tFO3zj35BccAWBn4tmND5u7pDMMILZNXkusnTbnu7g
CErCQ4aRP2kV5m0/c5MIQZY/xRWERmqoxP7WWnnK9h0lXxufBeyYc8bU6ZW6zGNy
dO/EUJhGBTO/B8Rc/OnO6EiT70yKFYMnVAAq2SbaalH018+K3ejubvfDZJPL9Dy4
Fb6j/PH3sStBACYrRjPTgu5gUwXBeHJFwPBYy8JYW8aRV4tAvnQo/fswE6lHU5mM
vyIBRzxjhntGEXvMEJgQ6WVLQKC7wYO0HHNKOkG8xbytNZ+5pbgaL9xqardguaoM
zaBo8YSeBiOPl1u6QdxWi7luEJFNYNThOKZdfj1VhWd1zAchsZVDxYmv5gthBJrf
hWcLrYj4wgLXzorEiucLgGmBMYXXzE4E3ucTI/OFk9w3u7lSk59bO64jm9xV3GUV
60y9yhesRJCxAgS0YvLJ43e+CsaU61DGk0vRD8hznPqtoz7LVX3lQuMc5ZGkA+NN
2Wp/v4Me07H7mZwX+LOl7IQXQ8AWlLuu6d+zxWdqltecdtBhg4RKt0NKdOOkYEsD
r+LZ0k+MWlSInIhvCH2D2mDYaSP2w5Ie7iIRZiUhrab/bZNifeSohK1uGyL9KUml
t7G3jAd1gPNiTQSlE0oSoA7KJrW6Qkdet2vrqb2R2xvI92SUWJPwx/3KHgHSzlSU
xr+LBdvYGX0ec3tWIlR5w1E3R8rldi6QO2arpjKrcCnLb65+ayuvUpoiNfezyCUk
OIKD8Gq7ePuwGACXKzL+sixygm+ajzKLIWHZOK4sYzNDjGbQKSUMjoVSHg+q2RCQ
kififEJPfMzjrNQLqk5SS4I95LqCxTOKRrhSwSvWNhcn8XorjbRm344VbU1u1M+O
2m+InXJys5eZwf0nxY2H37m3xsDVpmw96rAG/yefMdr8eT0LcJ8Xkt3TlSWK+ydb
rcz1DUs7aSyy9nd/oVPE5JUsA6762s77SI8mRA/QcG8KrFNWJoUXtIMC0irlRvbZ
fYvfNxN/UIlDcchEpxA0mpwPzSKBdNciK5nUwSzSHZ7vBbheBkzNxC93ER3aAafs
KGJvId4CydK3iOMRl6VqgDC52NLE4XWJTZ+k4N6PDHi6lJ6zt1p3jQneOF0Ka0Nv
pQyTX2DpXoQVQRpNBR6cUTSWrO47WAe/Ud6CY9tSGvBKGkE/T+MtVZTaAknAyFMP
MwAgKdJdOtDJTmHptSpbwRMYOB3GXmQfZLuPR67bgKkj81dyDPgfiUO/sx94aNb3
+lUQV3VXLDz1FI5RpIDvW1dJCI30gviEn98DdoiuADx8CMz5c21nFQt7utKDGMqq
uj42QL6pD6qBT1kXhQD04akLAE1uWEQTfAMw8gzDROET2a5y0H/mPphML3D+0FJ7
kxlz+mIV+0Bz/T2R54L2lfvZV/BXQAhBwlNt95PdgZaVW2QF9lfPiQ0rGHFtZGiV
sK5sEtk688/EnCBu4qWREPk3oJGOCYmSSwcVPX8nAw1Qx5/FZxtbhKpE5pf+XH/E
W4uUNqXmgUe5uXJ48/aeah3ofqLHteO2wSpsJ8LLHsG3JAXUnjn0FwaCL/VnY8G2
8ITYvhU6jkePgeATmd8mzXuQ4Bv5o2axb2UsdReswexsXRpH64sHuE1ocabmWx1H
plMotZgHvwH8refyjQTTo2R+22TAQhOGmuVnFnPTaHGxsm5WNsakuBQLBzswLCx+
xx7fGVFpGOlFEDBdIBjRcLjI6HiHKSdh9KtSO2f92PW1R5rNbM8AtjTMen1w9ltq
o9tsEU9pG5pD7WFnYHb1Hp5wxuf1IWTdDNIYe64HYeJ6GV9Xoswhky+Y9ixOfTXn
yW0I1wGFEgkyXrJbm2pgLo7Y2Rz6h9SZfr181qs38VGC/pG7UPT78/5Y0PFIwjMs
3OCVnHMAORyikUaSMjATSZpRdB3ajFga21H9ODWiAIcDvn53TGon6OPvlnYdLFRc
gVBclzyW0OE6OGqduSI1RxyW4HDFxzrG3tffahzYmu09ChIjAY4C0QdzhGveDBla
3kBHhRj8XaOi4M8UywPjUCV4ebkBHaqi7kTF2l5650/NhcA6InvNPjMpk/mQNLl6
eGbs6Gd5kFZ3gphOO/qmlaH7hd1YpzhV59NX0FrI1tIy6Bc86zSLDQidFet172DC
KgWHal7qBALoeTFil8UfeRyRNGRYPHL8+6qjK5YRtg7jfDd9tl0wxgW7V7XV/aG9
wf/oUV9iMucmC4D9G3nUxG1j/vVgHoEhpN6cZflHwB0KTBMVP6jENjOv8IdYWgjo
euIFXifLd7JiRTDx7irac54ZmAyCnIGWFohJOgx2p7WgLQF9DXrkexZxLqiOL0lg
Sdvso4ivbMNdP+ihB3iva+pnVEutiwpWnRVEIHBcETda9dO50Y2k4JXnMuaxTH6S
LkZTx8XYmIHz3oSAWrHa8PR8hExhOY4Hs6uLt8+blQkz6KuInnncrpt6i69LUNN/
Gs/aTk7cAmCcJHnGu+CTVzIwjNWz87qqBxazKY6bot/4e9o26wcSBZKImuNg36sL
ztjaYvRpkI45zx31HcNjq2caVHPgP0VGshV5u/F0H4sPGfxVY4r4KA2KlW3BhSSa
tPVKnYXqJiU2KDJbKF4inPaOfU2wVN/Ijs97oMmMfmR2kgUZ0hYcCSwYarZCFQzw
V128kG/r4y45iNSywAFmo/bvzVH/8zG+D3mSTGeo+tfDM8Y4dDz8H9dya4N/H9uH
ev/faF8mSKFQPy2ycvpPip8ZW/fcFAtq0GFB8Tl2/roEK2KKbWTPg8d/RQzKKElV
8H2c7ZWJToEyiFr9z5Xdnx4HiPKT3j++uWYp9rd8LUNdVbq/Urxqc/Xt60CHwj5N
KlGlgUoNCabB2VYsDRN69nWM0z0+oaWgBPNo2/6G3hSO2tFgOMpEPDkHhgH1f3Tu
iW84BHMVhlfKVo+an/FqYJ2UA3sK68iHa7ZUxUEfYfWq59Lgtx/AxlQhUt5r5cK7
tgxd1/a8eMUthYSlLpt/WM0WLUwKeNSwpRXpnYH2CY/zUBH6xGAhEuz0i1T95MDc
3mNghqKDvXJqtIb0rKbKbdxiibPvcflJC7JLmzeIpBKsitS/VQ9JP9ohLJjOQPb5
RniJbu78hlGyCl+5DxQFBLUU1DlskYHdkgZVTUVFghGt+Rt82A0we4jAfXJXtUKK
u3v7kMFdOWL/HBpu2iObhF9wXpWdr7E2sBnVkh3PLOwMx/i+IVs8TbBav8jx/VCd
BVrobYy4k/BMj5XiACHq2on00YPfCoqJP9FANekHJyOdqeLxkjZkhr3UxpK27kqU
H/defDPsCqsIC293fM6U3BIt2bU0GCVw/H1uji8ApY1wXFUJyVjFPUhcB+JVXv7G
2YDnzDL8Kc9ws6AGHyjx3cwPsJQ98qfEOMHQFNlXOafXT3PKeKHE+q3YoOYM8gph
29a0ZXM91QkrEwsrc52DdHOiUoXduK2erAF7S1bm70ABYsO2Z7uN3rQq9u8/y95n
u9WTXagPYSXr02CCEKgkxQ1BCFm0i/WXXROD0qC8mGxqlyKrlp8haAb+N9wVjeM1
w7XFNOInfYJBYFIXd7OpRa8ajVxki8ys06tz3e6vkHhJtARDA+EW23OYDHEnIG/4
VtbuEkyS2PKQ+llgo9dSb5Z83ROWrDn3jWWvZWxvUS/68j0PgwkxpV+d9sFRhNoE
hBrDji0waYzYBZd4tBePucBpXMnkv0dsUJtOZZL6PxQxP5k+BbXBvsDI+seRBxFB
yZ7MmVQQtMKAbxuAzyBWDZRe6MiGlrDntwOvR/VW0y01iYzUncMvAHJVyoZF5dm/
VyUccKJDxllxfo+bPD9/8zzHfjT+rV60F0RvFqwSpy7PIZJ9KknZIniVLF4y19RG
0/BE8w2Lny0L0EeL3YgSG2/YSQ5bl4UDniPD1TfoCIL0OrAhDsYjFI4F0kAtfj58
oryIoVd2MN/6SUi0f9SLytjZuFNO4dITnTR9PUHT0BImRf5vIjakouu4k9akot9w
/0hLOHV0zj2RKgROhYnExFLidE52jOTh5tWarjfN2msLne1fyqscIKbi888fYiQW
URjK4USjlb6DJq+ueeWFqqxKn65e0DLIJdBep+tZGptKpmEy5PGQISuJjQUffi1Y
45dV3HYgfs4X7TvCTAipNq9/7HiSo6/pkAkxEvqLRBzveN4/HdS6e0ku/Y0fLLnO
X67rI9m/tC+Br9oSrceD7WfrWUHM6e7XmX6UQ5+0mdaoWDTpUx854IuSzyRGVQD7
ANoSt7pNPH9OPXTUpA4R/D1uDM4fVhujwLEvZpxyWBb+uAFeYrNWqOGUZRfe0Wwx
JHh+UA6MaG6NJj57qoWBPnlCT8FdcZwnUxr8UBcmK01QpzAV9XsoGYFfkqgGinxO
QVXfphwy5DAWM5Q62bb63bOdFsYj1AqcMpJSHRZWVcs7PGVnlzNPXQubRvNXEcgG
X+t9mUCa2L0nED3R26Ny3i6Jyv+2GKjlxtDGlD+E/NhDvI0tGeuAtekJWo/68joc
kOceqBZBY14UV8chwnEgd1dJIaWUTWNZS4cHMhhWuR909Nx9Tvs9xUZ41NGl28ab
seQ1fEDtFx0U13u7XYoijy9uKySP3k/fGa7peRPucikdv2P1LfTprdkZpYy3tRxR
IB6oVhlKAPyVSDO4YHo16LRXyA2qM4OhG1OA6OryKFoqsDQTPIuJxdU8sGT8R207
f4V+quc7qRDcWiNidLCUWn+nj/xZgfGt1eQAp3wJANt3rkEGqN1toGCJtwvIpHAf
dS+jqrvgM9O9MPDk+D1Fd8UX4ywHd3jKaT2KG2HwmMfodJbH4jd640X78lchRUsm
KFe9uVmUpyAae5ovFgmGLpm9n8CcQFkD6985Ppf1fruQsXUQWKU8geKXXvnfcU8f
1ZTSPAgzSPVDHpGtZvC7opvB4iJkZ2VUqMaq85JnCGKnqboBJz+cj6YaAMwW+b+B
AAGT1UMP/cWMMVjjW3Oq1S5SvMIhrEWVVfQHbWsgVEGDm0Iqd7KrCtLj6E1RUToh
Z2KRGZN9TlLWKne7+waAmd3Hnb62K4EIQlp1eg7rEx4uJZCn8jRUM6zX6oDSln+P
+57gf6FQJYLUldqbMOm1x8MeI5pUBzoGEOrH+8u4yWVeiTsEqDqYw7qmpzwcUOrV
SktOootbVoAlpycFyxYDJIpQtYLOW37WXk2ruQSLm1VFhHJQ2IT0B8XN/umAzDd/
pEZPe3GD8YU9QAjp++1VgzQIuV2Xh81vh2JLDKvewP5I7nmSNorwfmPUaBBBU7dG
EAWy4k1KBTqJp2pfko7lVWoZMOyiFw/t0aHOhEJP4Z6UVJkuUbUNXtYxNyPIut/X
8WGwU/iKIwZWeSKx+AwJmOsOyv0qKV7awa+IUWNdA9kjBGyArGbbTp22GOXQmQL4
MHLJ95tumUFeaIeYtte5ioxbkUpy4dzWL6ztPvXkqQyxVdLtak48gpTGnHObe086
yZqsrZx4WEevb6q/hJA9vE3ViTTVxyg6OZGPFmravdPQ1ZlZtEoMAs/EsRp/OJr2
taiE3KxM8PDx52Lo8tTtOUa8PEX3dR82FXU9tM3NfHQcADPU8pz4OKAV6+v9PQKG
CAPQrnusV8sqv1PYAR1BYqqiSBOJQVdeF6wWOFRL2IukMYZOYq+JNcO3MtJYvOr1
p8dzSMWCNiFEFTVVY/Vz00bJ5lEYFubE5AqTRhQ1rr1yCIirZfqIRXaWZqWjtnv/
CYE0hnmMhUKIMt4tNk0gos+qLyUNf7M8Pa6Co3LfRfifEmz9r+qKEtmii43RLP3m
8+80flA4oo/BjeewLQfuQFApaVHMEl0swZpPGmnbPab0VqLknhiOBePBNBlCQwxy
DcWX7YMmVkcdj7m5vMD2mhhzsT8mRPF11MxlTz4kvJrsP37SyAPEtZoyX6weYQ1n
OBhw2YhGApdKn0F7V16UTuMWc7C5KfbODetx0f/C+k1FSk/4oAvsWmNP0E2+AA0H
UWii32RyiMPCLTnVBVOFKKOjEct7fTa1t+MpAOonLH1EW4xN2s+dsNJrERWnzys1
QgGHMA+CkIz1vlO1Y7R82GHuUVAEN7D0V1XLphSrxIUvS/cmoLHVLWQtEDX5wTT1
gDtIyafFIqvOaC7RbNNTW2ptVVhuFvJfKkmjr0HGBskVGIoinJHXtUo4swFNcSDN
Xbyk6gm54gQpZ2IYENEIeIZqlvkJlsoZOWl0GBBWY3+fzuJlxCfAPTRuLTutcvdy
eYsmvXfrHDBXIkwNKhqcIbJY2zgrWqASDdZ73J/NX7x66P4WvSFBRnKmVsTucq2D
ZKBCnydyXusZH4fmpaixpKRls1YcuQtd9DCpG4oJ3wVddGc69z7RvBMqgL25NumM
YOL+lsoGT0FJffe+eTobJDiBTO1+cbvPHaKKSFeGB0UPYG6AgHSAqmT/ETRkfwKU
xSWGSkEQTjYdgVxuoMCwdiQEVgd64xi+iLBbevTp5s8yqP+EAXV6IaBrXn6+s2TP
aaWypJJ2uTm38SZti1kaLU58qDYyaJdoTKYzvQe+5Eev9toGgqj8R/S2hIJMzwwE
mGc8FxvP91BJ13Pmk5jQY4tvala2Yb/nR879NQwmB8SOyhByfSStpHRu8Gk/GQsM
hxSN1gwYYc/WGbEfwbuNQ8qBfEQLzr4JeMQHs77Qy6FXcqzSQX7pqEJzOrVBQxxx
3hmhlMTzkH3EUbqeyoCyrHbRNj9BYn1yxCBWuAgkXV4HLljBfD/cxgPCPiztCv2i
487VLNbj5RiCseXNlBy3e6rR0NglDdNdmueqAn4Mc4RcsAu1F++KUOe9t1J3LF98
f0EFnYRuMu58Co0h4NY76lPMvMHctnvVG3ERvGCfoRcPEj1mxlX1tsLdBNiBhl7O
iyASDagzPFR18a+u/CGWdfDRNTK3jvAEQlGmqHGWiLD+ba3d8ogI9xtsd2DzqOlR
zUA5lzbbuq1cvKBXIvLlq/LYK1MMeX07KSJnfd2iRfmrN8nepN/YyICLi/l3jdGX
GGPYR/QzErZhpvIPmh/g5gkDAgeHgKB6Viv/4ASSJWdqjfBR5Yo/UPGj/otNI1kR
XWB+I2pS2q8H3SLwfDs5VuRNNNxwKptlSEdfZF6Xwig1WW7CCFBFd8PYzgkg6r32
YyAX+WOFf9Nwq+oZPNoxGdtojtXL1oQI9M3nwDe2Kpun971y71AOJD4eraXgH1J/
RXMLM5wVr9B3cdD+76isI0X8uvqwcMxrcyGHqOZ+p2QvSB+MBprmvs1xM0Ck/uN6
KSb8p+GEC1+MeFTRVU04iY7+1ITYudimVg01ESi8WOV3LBzkOY5u4EzEhkq9ENl0
/ukoha4oD/hqZ6CuhjP83bsevKayn+544VyLWFsxbIioaHTDw+LRPCy7aMyH9B9E
3+R0MTrm2WDZ2b/EWe1g8axyvve5VUL9Xu/LUqmiZykDoIuK22V2a/WWa+JrHj8e
8At8xVkYTKDGo0Eptmy5r80nAYFvcmuHQfhc9fmUF1wV/hHrm4epbhfy2LZTW0Tl
3ahYVCKNUzp5srAWlWczmknJRs85zfni5ifI+WrqRLyAeeGE/4F5pQszq0XJEqbY
Us9MmoUY03NzIPfN3TdaiIsRjrzU/LLhWje4Y1N29WxOeELOKMPEORZPYyNk2MO4
nMCfDbxGnzSDLY8BpZYrDFOW4/R2X2As53Hn8tlDFlDRQuavHZB+vBOiBa5pDM4r
xCjeehXCceLmzjE7M73LEjbfpRj18eIf5WAdx0gvumBs+qPAUkbGpInOggPsy/JV
+XMjdg+0tjsLwRtqiWSUVUWTXaeDCBix0aIrFqyt96Q5Bu5HpFbBz005XgDfZ2Qr
T3t+fXKrvmrzDT3irgeb5Om1zyct7r5Vv0tJXBSYJdOts6qUjJtZRIEWAjaLa2B1
i5dxqwM7kP/g2Gsn/uj3sd7Y2NLWIdJbHvQYwGGnJTairnAYFL70noeIZHzNOVLl
vYisHQYWLRH/RUlV6YdVsILEyfoBg/f6Jv4JYgN+zwfSLRgZEY7hwM5/RUcAAnnP
nxQSafhQCPsQCNAm+wBik/e6rbch8rbtjtoa8+UUzu/+q8CbhO+eYMbPCMYVhh9R
/ir4LeFw/SjJtDBiLefVUai1/Ow2n9pqyo5fxSlUL3oiQ/WfPQhDX8Y4nTZAKlAW
JxWZh2voMYFNoi19X4TJqKWTv0JgAcDCyPOtyL+kA046X6OouEg51nZAlM9l/mRn
2rkYi6Zn/dMbu2xh5GejkisL98FA1URwaoJ3nHYPYIFzcDisTgyZgPcpxjC2wqiX
Ho0ENCbBetn3t7/LjiSj+2g3SZ4Nr5meEoHayKUfRwkbvKqCOADB+iQ3OmwAJuav
XU2fdhtmsrECvzZiWY2Ouufnk9oZIDjSnVR05QA7Z71YnQqjLKiSUf2Nmymd0rFy
DZv5HdXL+DRj2cVQ3jVlkd/IAzLlTPzBX2d917YrX7arVcEreO+WMYfv0r5/Xoq9
4EW9dtfMOhxhN6GVaDZKhAVSdKSc60Lv+xDzpmnbcV2IyhI4IiVrB2zCODp7n4Hn
49ehFc5d2PUCTm4xX2FgmDWec6V3LPrqqs0eCxwm4g6Zxj8YA3+cM2s37GlTyCiC
zRxpiStF/kgj4CP3mPx7Wx+Wm6MJEnwx7lo2d4BrDMGxcOkYwiGhnbd3SnXrkN1M
fnw6fEwKYW97QdUxcTYpuKxzE0uEsHLaIJgwfb0LiiMKMvskoNdXCZ4KJqAzXjN8
ZuU6xFnpD31/w3Ca0tDAYHoL5hAWYKbegCDWLb7HpEBwl4KPluj7Y9yi9anEx5cO
4zH5mDNB1+Q4dkiOYk1dEAOjfSCbt0mXlrdf9ofH+kbSuaZI9AfvpBhVqbN/YC0J
EeQLkXJ0gbJjbwSVGCcbal7h0PHV1rVw4VOflwV3Q6/SjxqUyhCaUxfgiPe73Sq3
VCRC+Cz5jIqv3iM4mIcY133Xuo3FZc2xXepS28dB/bQxe+A0qVkY3W2/pHOderv7
Tumig4kckqMk8zwtX+Pwx/XFJywz+/J9Tcj4KjtkbU1cC2gxP8eBG8SoFXwXcmM+
6++ZikNXNLEF9Inblu4ZlkOl3F14vPleuIA9c9x/wz28LH4sKmM6mhR46ZabC+u4
rEE8dMlK62bKV/HUx1P5z/nzLWGcyxj5Pcgl1/CjQJi0rYSzQ7Mj+hoSUsp1KVwS
sm5lFRfU+NsMNOiQ1EAmljyr2mLyv8oKzsW7/6ocf24wEuJKLAYdo33L5Lvlh13h
1ZkSDJ9j/BjvYDkNSgfzYiA6UZy2oPj3tB9fw6B7JvHMNDqVQFoQfZYPXYg+OYv5
ATJ3xzWngCFoxfWl9A9txwmOp0u8tlvGmB3mMYLBuNG7voROF/rurG7TBNvxv0Ul
Um2WeE0fqH7Zqm7U6z2KS1wehm+mYa8XrWOtzz7AFTSivqzGJ0hSTfd8wvrARPrv
suEDK5mWiM4DwiGreFSrgKaGmeioeiBQgM+bzg0zCgARBs1qV/VghOEvjX1/EZ+c
eEXXWgxNJKr1Xx1rxed6ql6tF886ss9YkjxCyNu0Gbtzh7ZNiK2Mv+95s930hvnw
HgD5UxQjPukLQARfAEWuO/Ha1AEBc6u/UAWdgVJkL1uw2PdxSEKuYemWzBAK2ifE
nwplOzvj0GiL98Nm5iYKYdrOuWqMhR7RR9N9ogMHaeDvnxWqHq+6WYoxZ0RsPQDg
EoRwNZCCJSzD6t+WpEM5yWBCc83lLHMK4IzzdqFX/7fnqdpFaPu4bc3QztnA+QAr
hWCMUfOSAlewdJqQklngCSvLagkKuL81i7OK4HF7PjamyarcKjHRp/chGBzNZJmv
y+STjEKSdJqBJjrCuHcDpESzAa+N4goTdMxPrHE+ky8GUzDfIF04bLi7jPtliQb9
KTa1urImFTywY8bjOari/0lE4wTJGgajO0fG3eJ+jgLnJz5EDB3l5CUM97e4VksF
cAyMpQ1GtnxbEljz5FOBC6mayS4JBKgqHm7QcE33MFIE9PAQtNajtZl/qPK67+IS
xvr6PbrBHJ8Lf+0rWmIul852MPrLqQ98zDW9610n539fUiplbbkgT+vSw0LWFkN8
pD3nuYeUocu9OYfrGqgCnMoWF/4riwbVKb+Qptke4RE2OiadW1U8hxrC2BR3iNMB
2NvCS2rz9fqj6hshLTukxX7/wflUl8fdyocu0/jFN3tNA7rFD6dlYTiSPtDW2/JX
vcmcWhf9WVo/HKB1Lrgg132bY1ylPhVTzg5EVo/Y+pdZcqmIfkQ3C7b9x9XNru2h
JvyV0PHkL4NEkbx08DqJinNvVE9FXRnXaQ4NgaQlGRikTXoRlJSsHjWraem516fl
xSzy5JYuJwezkTMPlJIsgSsm625RqcGnr7ZbsMYACkObtOpTJg6QFcUHAw95Kai0
zoekVZ+MD7Ts850I4YTZ7JK30iF0lK3rS+OenTAZaTqZx9B3mqGFGLWgd1rAHES7
R8YSCeTei9a4cLhDiOk0euN0lnmFzJ+SzelusZVgeCfW/g531L06kEPHzh05dAZk
VWkmbzTbvHs2DS0H1NLOfHvMNigXLyHsCAKq4Ff65o5TvOMT4vmcNWsbjkBEtEqf
lAzKVLDFxjz1kHnJY1VveAtie9TFuMO2MUlmtU3GGU9VJpIfzCuYWio8ABsLmv6P
H/mvaDYclQOUktLmQ9srOTSuuuUzbeN+zSxR5Y+JaW3fsOvZCw+Q6S/oVAWejG0I
kYckirMVy1vhRgSGobSbfIz86bj0EhveG3porzR/iwign2RaVotZgi9Q/ptJw9ew
p8j0xNtZPMyl+HcimVsWD4kQ7/z2QRCSo/AzckOkjqhA14HdMZORnxwZ1n/3qv6u
Jw+Epsa6wU/fWHxA7/Wmk6lJVRqQ0DblLpeyY9JGGEQwIU8sGwcDsBwkCMPBCX6W
Fr6ntFefRMwYa8GLXYmYafMT6NWjUHYnCldRKgN6F5G01UeZJAnbpHqgzd2uGg+x
eBNZI5o7drArla9sWiOSdCvAdi/7LVyZeZbTFGDxy9Tuom/TV9ORZ99duGGL82T2
xhxHkeb2S8pC2RSRt0XN5i++uW65PzUw2v3g+TsNmxIsebFTKNBoZL2GLxFpggma
eXdzB9ydoSMYgn1mExe3VYnuRBD70RuV54UjYUa61qBAVWtRSCUGglEwreViEvtg
ycMELqZwkmDL0g+KiJHErwh7WEpLLLqOFlh7bxO8Q/dXzLDTAilwUDqEAB/txUJQ
Ac4/F+QDKJdj+ClCuTeAaoWxotx/69W38FSo54LFioT8d7qCp/D8R1Mox/0/CipO
IljpaJ3bS9uHJ0OGBwHVjuzbu3wK+9vtz8ynEQ5ADAYY0M+7I1CD/f6qA42z0w6h
xJuAuMX5j98JE1SOo86mkamCLlPF41hA4vUyPGq6SKYwyAUFG3NuVtJmvdmRdfOz
l6SnYW5E37a5zD6g6Vmo5DkGMWEd1WbyAdaOhqf2CgOGqtPfhVef4OO2ytT3mQT6
AtYA5dVg762w+xocCEMcq9U6bvATadmYsACzZm7LJHo8CcROklnYhn+ACskHimnr
wxKZC2ph4T0gnFhq7eC6uFG3Ml9haLBc8PZv0lYljxJLKWeem7FQxKq64/J8imLK
Pl/0VE/3jYjEiP1tc4opbbmuc8zd+x6o+4Hj+lMY58hUDnJLfrxe3my23spnT/U2
ZoEW8geF5BAjI5erV+vUF95kO+mfJ9UpyhIGCeT8aKkGUSJlvRGc+j6+jj9fQ+n3
V8MiNEQ4HJ7JFdaChqIg0ltQ9I7Y6g6y4sTRluYEZL5silboSxMykxCU7bKKpAGG
jZpZOgfrjcAoK1Hw1fryvO8i6YtUJrvb9KnCjagRZNlhFoM5I+JQdl8JSfzPlzS5
mhmFphICGaBAV3scBm/Dot6wETxEfubHcmRG3SdFn8eNzDzjwLrjN22AVSK6UNh0
2A/TBEaKExEAZtYnJPdV25hrry4f7mhEyhnVJIRrJRkS1aCyl/RL3PMxE8qQpW06
6ABwF4V7DJ6ver2t5YBztmTyYuPDuwy+jM5H2QCaU9cUZ8ekbSIfvHVCHoJoJyYG
kYgtjgsanJ6G3YPcK8QN3aeIfpm9+qCSUTHfKBZ46E+QwLBfuvoODuS4ISp0+Xpj
NUt8okfETR4tt68tu9YIT4npLcoan8BM60+IJhYLbfAmp0MAtf1Bt1HBOrz3XV/P
LqQaqD2zbNkRkn/H/HdSSBAb3A+kyOyipOSwgwszJrFdqcbC3BQgZ7yNghMzpGzp
uHrtjZ4WfllfqIStfqQXGnchIL3BCdVRmK/XhFDWZe6vr+lVfyFprNcnBXuP2a5z
1Uvtqo/eorqFEUEg48Lr3J/1UQiwrKJ2om2Gs3Z8YKQ5FME51r1CXQSoDYfYeDoJ
nhkIT+5Otgl1EXklMSZn1R6TPixSrrZNji7RjbZZ+1FHw5v0pc8s/aO/CmYRlFYY
Ox083cbIx55NzWdtcYci3pdtgl23V0Cq0miLKfPTuuE78TkDdkW8PnNTYzKWuV7Q
TtpNWu/5V30JAogI9UpNmuhlyf/yB1ND18+4vCu3d81KyGNVgyS5DYDebpZXoskm
p+udGPmXb21aUwqi+ynMgQna0/CokSYXvnUC9ycAAu946aLt0eNlK2xeMBiIXZOz
WpEJzo7pj2SBRL559csFw9xy4b19qLKyvx9ZoUb+ZGqU2B/y6FjOB8TLPE/Ugb6B
GggGkGT6Qke5LNWRe8PLEHaSeS2/R89NOBk8RG0Kxxor/5+LVeekOhh9I13rqDZb
pisgg5g9QgBefqzrG6Kip5KCKbre8AW2F9ckptGlcYc2ZzQV/h6lxCWv9ePzyu6A
I+Epu4YUGKWw5OdDVqFaYgyWfCkFHnYfEX9IROIYjcE0eE8gxpjSgeinovqP3U24
n945/26ydtlr1nujJc/cyAIOxXchG+N46xi01kZc71i1WsZu9LOuo9yOun93mntR
W+r8ixcLX+C2Td16LnKDAiENNeFFGIdaYvqNDVIOPhw5wNLj/4T7plRvoFv8nyEb
zd847XhL+aVVjuanpub/fMQ/QQCKhlf8R2M5WDtZiTqI9vvNHMG+EYoKImUqdkOs
zMu+PSMNyS3nw1TMDz3kepEeTOOw/Yi8uFf2dJuA0XtYEzIHy+Af9oQInLfOpA33
Go5juj8HBQ4n5U3neoPgDKUoip+UfA5Vo98GFLkcTGpeyKLRJM8pfBvXcyJ4j7WZ
uVrZ6+mTvI2XCOEBCxnEXSPIjAt5NepPd6Uwuz58Wd+JpeGPIxKGa9rGwZ2pG0tK
dQ6iAj73MH16gG1U9IWKa3dP+XbPldpW+VWxy9HNbqr1KUMYtmXdJaedvpemcOq5
KeQOlceQrzGQgHhbyPOvL1/YhDEUdFj3f57PcryAlC2diaKS005IduDf4Cu4fkeU
r8lsvwedalXyTDStvr5N+bsCfI9d4BcmUjr0lF6lHL5QMBX76CQlArj63ANY6zQi
cAGfRc0Bj+zuhJnnOOgalHhfDmRcaLRJiS6RWSpvnN0qqXsRx902U7QJhmnr5JPE
GIkqwSLSxv3HmMIhzKSt6NIYhsM4yN+V8alH8qMkRtWT9DyMf9lRIsq/y/r/NNxe
265JadMGSFaAYLl4JaeZQd3qqZMIZEcrICVJG/VA2R/WIIUvSusj/0Ap+Gu4wH53
2DhwnSwIZBJzKXCk2ljDnU0elQ6Z3IwVhVrdAXj3ir4Fh18tylDOAby69BVDDfaW
+eaRG/GRLEJnxX8YwITuPWeTIG+aV3KUgwvYnjAyWHB6NgXmgkj+DNZYF8o4fQ/m
dvQQHV/yqjiQXbZsXc/lslv31wWpROl7au4D4aUpGKVevLDPOkzMD9NzBIv32e+t
qR+pApymiEuE/pKTcxfAHbcoxKS4YStxdiA6MPdRF3o/6xgS3aBWIgHV0Y2f2IIv
zZ6UU0e8N5UN6oTtFMfcuOWRm+DMkHcfanbvKb8DAqT6dyo1EPUGGh7MQhWLcIC/
Gkr4Xnr086e5dvMrMb1U8O0WMV6rxUD8ctmtMc93YZNzWOQfzKN9tt5Mvw8bnkNj
dDx2yzdEsH7jkyO9BVYNKpabMLJeDS/IXTHMfbgOYhUUE2JgvAFvOHy6fnPfsmXj
nVl0A/wWxMJmDzyzKX+1Gg0j2/zoLa9fbcIzEEX7VMpNZleB5nTmsVVzr4kgm42W
gCMw+TinG72EHyoIxzTFoFWUhuT9UXtTWCVDgxk7our42ToyUDI0d2DDIa8DCXom
BWg14ujH3aKPOnulGvB2yGZcO20NscfwT13cdmqFUoJzPZx7MktRySyvdNUjF3Mt
9CNP5OxZSb2vX/CeTEmfDAR9JuAndvxDCtWcsTPQ4hECNZ1owWuZPFM40eb0OEJO
ZQ8cAd+dqHKgBNNLMiSGPp0erNyVHRTJWFiiGSrEo2TyZ7bSf+MlC8oSL8FW3yFT
Y6ncIbk3OMt8mS30GTvseMUtzBoa2d+a0A4/aJaYlRoKsGfWZPBHcunHDrqzE1zs
JRpnallI3HJQLRa8dhWpP6jHw7UJdSU1Q9KQEDA9LimJsQFNINyyMsC65CP6E4mG
RDHnVEWogxT1xsxD6+pr5ZnH+saSAqmGDCJlQ9w7aq3OnK1XsQ8iWnpNygPh7xQJ
kHrK/6HQjaELCUdw8rQkBqnvtW9q84llyzm3j4pIfiV/2nC1q0V3YYPqPHj/vrXR
jcdlf87WrxlL8IPhdQYTudfM9Bl+/4KVmvTXP6w5ZzIdgYCaEZ/ZZ1JSWwqnWy4j
6eVj2AwNNb0lE+21EnyESYo+30Etl4NtYmirFBell0m1N00S5iXjhOhRXsbuv7rH
Xr2lqquJVmUZsGPkz0X1p8aej4KbB51Ggk0OcfAGh/e3Q14RzHWm7etsv5qCJ2fY
29FrtZQC8gAPncd7T6wHyk+DNX5UQ3ljy0FHNVPd/PfKq6TqYC88FCVjuBv1aZAH
FWSgoNItBZhl2y69ocNeAM1GQzw5IJ2N1Db8FvqZagJ/tdvIMJAyz4BgxFJU0G0F
L3+UqkO8M1/3Vk2RmgqYS7dEDOAKUbvQMuDS0PR8Idu50q9AdsH9ZMn81nx/uPY5
Pk8yVgOjxEApW4u2m8AiNgQwNqjtPDp+qX5/ZoswfftqEb1ZYAuoJTpeVZX/N1PO
fe3JlXHKmuTuYjZxR/n8ofMGXe2/U2M4/PaH5qL++zHFwufVxZ32J1lOEZgK2M0u
Be4JPm3Ms0ZLDCpEfb+gmy5htQCmXC2t+PbSMXaSuOl3MpLmbnUgka811Q/Wqisp
JY2G+UvCx5vTC0xP1cTF9d4Gqig2RvONw/mBgIhrdstz+BGcKy+gGGnso39s29So
4Zv3twp6PgoqwZN/DpdNxyMeRyAxx6qT1FuNSsOkQV0lXGie14ima04sHmCx8fa8
Fj4qROM/Z17uPUj9gvhDn7lPL9jyVEEsguBuUDcBfuESLvgcCPQ0UHIREmQh8fML
O1feKU+iV4T4f9SJrjZXMGbk7NxN0oKQqjuJRIpfnLAvIYrEzrnXQVGhhbDoJGJ/
J3P5QCQAuNT/TtP17FjAG8/xlaHindP9uvJeceJXHpilflisCdO9clGHT39526Md
5J0O9IXnvIh+TPSbNHBQpOiak21vl62kdya9syhcScRuAOz1FZ0uaR2J5vl9eem7
mKMndNxN86noPoXL4Py7tT/NkhbvQRLTK69qU5hGOla/mEMbtQiGi/TRFmLBp0Wu
xWNSiWz40Qu9eXtyeZvism9O2dL+ao/R9ltyWVvSkV7GxVAZJSUiw8kKums7WBq7
D+bXeI8LQhiA7hJM3pL/N8HCOt8vZqu8bwOMA+4puWBi8HlBPmj1uLY1IY/USoHw
JrKHIB/xOImNzgLs1NLkgLcEP0mM4xsPm8NunaglmJ0aCL1qMNtW2tn5gZntFU+2
jmZ6YJOMAcMfQfwCV8gZVmxEB36yRdXApN1DjH/OZ2C3+pNDg/KktXwdDkK7nv2A
UBWYYgRYgsNsPXXpLq65A1bwUI4X6bhGpKzJiD3ssGRK7WcGtwK5jlf2Jor/9XJM
4SOJd3Z7fT6v+F5QoleTInQpfca7tHthDnOH691avQWqOTPn5A3jJ2hm8dLDKuuX
mNpNB90REJHLdGIg8TbtK9GFXfbdQ9kbkB/FT+5umy2dC54ckN+oUomW6vd3LjT3
ktrjSHicTx1p0TfJuyaBp0lvZ7F1J1B3rmfh5Nmp/eGK6kHFnxUEs4HcXkUKi8Nm
wGsEKCt9PArntrrcnGiNwWgFrUdY2nfqx0rqlD6nQhnrWzY+7xUBjG4wH1VJ3Zhy
y6L/YctMXkQOeMWatIMFS/HGkSIdiNPOOPixg1uREse/aE4AMLCto5gLmtczlmu0
YjDvLu1Ti1ebwVcoGdcQpX+oE9XoWrxjB3Stiqb5Tn5paAr/XiwfaKU8/y3TXj+P
PcQvTBLkPvzWDsJ8OB6e3xrQQLfTNARR0fG853nWNqnZOZGUDq8bvFAHNZKqBz9n
JsLRZGGQ0taZu8wPhanghp513W+MBxBP9JzMyOqI8QixilJFkEh9hhwgVb96H528
lXpjT0Y+ox2+ovuwakQLmgjuo6yks+I736TNHNZa6QtDx+O9h5FNs6aTN2SRJXuk
AT5m1Tk0sw8f+i9Ev8awueyqbDEOfQWr8IzPppjqtyz55rmw6OMM/XFnJ4hCOvOK
7uuQyuPMd+bVLrLa4zQYmsdgeePJRVg2EPA2D+6/v22s7yDw3BZLL8jgTLdbLohC
12nRd8AHGx0L7NWro22Es/83IjPZQ+OPPLaO/uWGJBw0XMSW0p/fY1VuJvdXj2pf
vTOzXNLTsMNw9YVGbZv7wPfU3mSifjCykzo8l9QGEybTXoOLEcdi0byenTMelbiC
BIHwZcouADvDQTmiU1p0Txug5PmuotwBr0pyyG/pefKI9QlKsAF50ttzpFDjOJmn
2M0/ihudnTfUc0GXZO/N/csPkL0Yo4WOY82orksuZwNz/bpbx+nECekZGI7lIvOW
VTSGUxGbXyC2uiAoImgJ1j49bC9rfCpI4pYV6XEd1tVcPwztY2SWphKOn8V/X2cC
yiBnJyTjiOb7vDBEK/WZwiG5cXMaVAw2GyS+EPqCCpZ/EmfSD/rUbBtitaJcvVIl
OPsQiCJFAQYzfpfLnFwYsCoTuUTxt3oKhI9m6gaiQnQULqXkB8MZFycUOWhcYt5t
8dpb8uOF/1Fp1GNlELOcySY8QAPunak/yaui5Xei8szT5B2ADiqxUGVAz1hFCMsV
ZMHSGoDBaaFkqx8Tm4XDImf7hx6QmXrjsjizEawAhdz60ljHLDRNeLA77re6IfT5
G0FRyIsx0Wg93Q1KvQZ7fd9uqEVZKTmGXzcpF/nbM6CrEb11JCMTW4tS/p0ByFKv
Hj/pkvZ6BebdaV4gH82Sj9vba+Ld75/XSrwW6VWg0lrbpOzRUInIrmxosBo9vpk4
bj4+1mhjDfhYll78JSTbq4Q55FFwpqB5YWPPNqCKjLZcim921CqswxYM1Ouqf27F
J+6M/t+Lmhe1UOQFtuBDTbud3/dbrLv6c8D8i0bdw7IjltCIS255sCAXIuw3JLSY
TJJuCynZSFtKSwJDU+8bWlW86+58/XutxSVIpGTu9V/p/liICeJCS9iRqH76WXlv
O1HPkip5NEO18jF1LZ29qTATe5gQc9X4gOaGuaxzqiP7LXrvDU9mfH4oqHWP7OOK
gDXmUlZmlTZkYjgSkWXvK12H5VSnkhXnhL/51bpKdE5GCgguOESJEydqQch5qsQK
XEhIMY+hTfAncQOFRRlvkmatOmiw8kN5ll/x4EGpVHTL+extwpKa/MzNK+jUgtXc
RLKQ728tEe9xHu8oiHSB2q49qA5ly3hhz1amsXSWP93QOEUgIBkJ3hyFFVY3Vb3g
9FYbW9e8YSYA/HDQv8eRLH+T/TY1gsncHx+aihrBKf/wEVbu0KSISLI+LQCG40qF
M3tCi/tQcKu+lmH9YtX3wDU5i3G1kRFfy5gETBvoGNBQEbc9g+d+5wA0rNzx0V/S
LkLLA7ZCkPXBxkOJdeukn0krgr4Ya/2xMGlIMFJKsKSMai40KDwkkd/uaK2WAVKm
7LvNbYHNlo/uOHYCe953eK8KikKAqO+VQeGWDJOYLjfpj36Vrxa1ymOLswDb8sTJ
jOZt/W1H0bjw95FDUv5rwsmdfIa2ABl9HHTYoBsAyhFS7fylzbtrs9l6NUMfmZa9
fXnr5iSnZB2UsQ3+H07ERw/18eha5ow/UgKbDxnBmz5FGXVNGxzZ0nH4iGluBd/U
99c9ZexC3VXvFkmUA1IMuHgMCJXAOTP4eqW7UvI2eSNb13pe9VIV5K+vxWR1wGkO
JWGih4pdl1iEQgVvOfi8FMJRlO/7fO4NsS/5t7PPGhrVZckD5XLol16D6XRO/UwC
BiDWjGnnHJpPlkyepw3eTAoX/5IFT+kYI3C2VcwO+dVPYaEvHc6UQG7EFivFFwcx
ra3rYBag/wnO+ilWqU7urn5tvWrb/RIt5xWmD0FUwVWH9wPHrodVVhXBKZO7bGLz
ea1hYTJTXAovEfdmW9lNYTMm6PeiMFmehyonoekdN1tsQ7oz4Xg2qtyTxpNFG5ip
orsL84Kq8jemgDICOvKzruNsN6DofXtzOV5qfEkr2F2ndvODL8ZkDtWATbBVSWkq
UO8gIOveYx6pjubTYyGw4yjzehxyMzQHw4rDFVCgoONoDd99fCzSeTrXm0XBKaW/
9+ansKI8OnfhtchAJHMen0Onmba3ZxYaZbrNqWAT6z2IDRs3lhXjMFmfX2UkPEnr
8finook0b+yXED5P8nj8fjHbzKlglnso4cehS+gFvlvAP3rVCxNOcz/eTMfJb8RE
kRrdEIGncn7Ry6YqN+6bRMjwPDMmBTBBzWKtnC1BcYrveGwi8lQo6hUER4vJh9Dm
RDGB79O5n1kKOhTeJ3Ewwhj1MdGkTAYMTi95Z3kw24ikRaa/sH1jlAS12uHFF8WD
xnMjW8BANTo8QMdw158vaD1W+SaGZy19KnLghHnQ0eXRTfjphFiC8p5nU4dvQbyU
r0r7spgb5Qfgaq1I8Zn7hMzScEmQmvPFxulZBBFdLoU0Sd8Qq7NY3ijQ7h/w1HgZ
t7kbO/qsBOfqINZclNwUroyg+ulBJk5TLs8+CwVFBl57WWcrI/QEnln68ENCA0nH
/L2ZzqD2OkJwJrLQHaftyDssIYKJVgsVUyaAa4UGnbB2FEYFwlW8iCugETvvPujt
Z0PPHzWjUrnuYLOEgfy8r6zQNUUvapTvQipsQee1nIGMuTBquGacI7Wk8mMaFqwO
mIZ0CFckf0MV6E2FXIO5dTT1otTntfCsKQ2DxN+A2shncwbEQOc7dlLauxuiXH+p
7EqbkzkFcb23bXv13bzK5qSZt1LGuHVF6VtV+S50kxZrb9TgFNgQvEEFtcbNkR1B
Gmt1D2kjYJM//tyudVWk64iekY4vYQV2aLHlMVvtYu46DWm8pcCe6A7P6qIaxgB2
67hzkb8S3MAYW+bqQJ44H5z5eQvsOiAydqrZNft0J1juqgcm41KkqNqKI8atKUQ4
XS0ECqFPhMmEEC6V4ueGqEApc0NMp7q/kxk5OWEw0xkhIZbr4upvmNwmTMiJPKWa
NzLfQDQRxWGkJYS2ASntTPgwq/HvSOe3N/57xD8CUuT2/NVdR8pOYAeFRkeYkSEw
US+Qj88ILS1QKifc0/00TulhL639VlWF9LiOwqXXguW0pfxLUZmoEtEl+EUvO+qQ
H8fvnkK8U7KOOBgZBVYoGs+WyaUyUH+AxkjizLO5ld4LGa+Mkya3AwZD4iji4P98
ZJLrRH27gMbcWcse1TOzWwq1oDLd1FUivNHxXCn5v94bu8OfPrbgb5XOdrpQSiah
3RXtAwI0tq/TgHT4bVbmbXE7HYCweShtRcEWqz3FAeTiL6Q4WWSOpSzQMXfGAfVf
lP3iACZuU7ttE+5J3T/3Nsct5M67qJ5Uo2uRm3SObq8la8m+Su2wJBq12KSEkHbL
TNybAE4eCmpD6XQjhMMxZpbjvKOgDvlN/V240X2oEJCjH8y5ym9LnoH2FAaSp2i6
Hqq6q1jswagYVs69xA1kAW1M4RkH7Gr5WHnBmTVe8/R9lhJTrUzP3Lo7oUcFacK4
hP0/jS/26RLuJzE0OoZzv95tKho29if4YgCxPMg0gjDtl1Pk7a2Crj9X798C/JmF
OakbBcpY61r2XHGDPrEbFBV65YSYqnVJmIgAJecO+5WgV4DlZH6kl7ZaiCR9gsd3
8gzkGJWxsFoVeNiTV1Bs99H8CosiYIyO50LcpotdxZ5z+TldKLCACn576lUD7Vkh
LbwKH2vlpdEUpkGGN6Vcba7D++t9uzq14XXzzgmmiurSRQcckFZmdrQfmB091ej3
Ys3UAUO45dW7HgIuOYT99LTTkHcPeRvW+QFQeergJ028o8TsC3wZoexdtL8icTUk
vJGLBtXKv2l5mWbnhDNRyTa9h9dZ3VyTIrZ0xTJyN4K28Pnz2tVG2qQhk3UYVs8Z
v6HtGrMOiiD/vgHXWx1LEWZHYTudf0kIW62N+JQPSkNOBexuvAxDXLE+/3EeLVwe
FBSCChtvKV+xJ4Y+5oBWIDdvXqAYt3T/XyBUvCArpvcLlNkyW+aZiEspbkgMJwez
hEbNWt0m5KP4dmva+5VKZRfAeA7ZTkVCM5f51fkdetlmbdPbT2j+SXZ5dLKnmejT
2jZIoMq8bjWz2uVaQHMsxFboX0HfirorjJvTRcmKCScPZNZ1vNAqtO+46S6aQ2jm
1bTRGfxkXSo6KnkURi0GydIIzO/92Od87fagVLMkh5DZtkDfEWsUJshCV8RmiE4y
3FS4i95a3OtHzil9HoRlBX5kKlLJrXhgfl+Scn/syzTCebJv8RFrfrEQMH2o0K5N
OClf6LMYRokJ+vt04+13bNKoVK7U6YDCobB4ocSEAfcqZ3DpGU5/SeExNYf/Whz0
o5ECJPgPkPeLr+XXEXsnJcXoPp/S4fFn0OzV+Qtq9FoQKdfyVsnixmEf2uQrdlx8
ao/UIDLaK/ri668qSvaqFytEDxEV1T42r92Z1/h1suHRUOds0kLexswVg+6Xd+Ey
Z6qbE7Rg4CIYjjZQNq6iy9Z0x28R/yKbJMUjrWib+jCVFKiE3DLqrTlQU77pBoOp
1Otr3VuP8Mv5JBwZNYX/BKhBWtvXLdvtg0UmNPOn+8Ts7ZompIuL40lZF3hXMaqq
QOf93dnZ4g0RPZ0yLRhjq3jPmX2aw0LIcR+KO1OSDwo0es06nVIPNdweTF7QYa+B
rd3TCm/iGO3vagYO5CLp8vmLx312bJYTTfxSYqZgLk2vPoEvwS/ZGR01LGYW6fqk
aAyF5MUNYQQd6a4qR+X3HWNcgqUJQ7MSVp5p8sFOeETM3MOuDFNI1ByHQ9KpnRAM
Yvbi5DU4nLa/EOTUqk6sRje8dnP/bolF04JVe7KVjKo8xHgf6Ks/BXmvknuN64c0
b1JvJ+0CRH4fbHTBoKCgmxIYy7PrMwZfTPNAsV+wlo9IRU9Gfd2qU7ivYEeVv4ks
ugPJo4q0gCf47EjKUuCtvP0JgVAHQYLkXFaoqUijrmD+56PSG6BVF+DsNh3t9Aff
tBc0O6IdgRmkkuoeHluuvKA6inzXO+6rz4thjH/AtSIFQdcMpxUx+gOVRz0IH2JQ
TZfH9P/f5S2TzeHp8j4fjerfG8pUAMqkHi6cdb5/nXE3EqisfU/PWcCtqAloTpml
2YhfwdGrDmfPqHyYY6vxcPaE1hUGeG4Ks5SOOOkA5OENNc40fX6jzu0+IWAuQrHg
aivL/YQYiWpaI5WEQt3MEfwkk3AVK7i6UZwZy5eGsYzxiBOt0+eTEEv5YCN+YRsV
y09UZpm4tnWfQegw3Lle/8TyOi470OWJsBZ72c2flSX2f1jGSRK/ls/tRzEsuhtH
aDHdU5pwZDMD+tBK8oeWlBZj7WSkmVbEDUNKOowIMyXgvz0dHjqM59sioQunPj30
9bih4InHJeB6I4FjdLbNTkfIZn/0vXLCnjqHtYoRxVXNqVBJgooD65AlSodpXy6d
sMH9aIuGATEVCFMxZI1uwSnpwWb1TEOy680nqdIExtxloSX1uhJuprVf9qt5Fkpg
2pIrW20i/pkn7qDfwS9fM82gy3rB3oMtGWHVVg7jY6dxHZy/9Zq3Bha30r3Fl8MN
+wI+q/27NQUchMdd0a1wJIHyTxRtzasoODVGPrVSgf3OOIUMPJ/optcTr55obA21
3wRv1l0ddRezeWQfddQfrDwrx5YFod4F4lp0qnZpYUYiCXcpj4NNXw1iSl+dqRIw
FPH3fBMGwHUkU6VtDk9WgVG0+wOfZfPnGrxkA8mNFBIK0N6JBwozYl5c4pbWZgMX
MuuT9JJl/N9rdtIP5dHChbIu5xUkkRTXXcH6bgHVDygZ+uZkXn0eZQhUCH+FumP4
NA22YSxMYN0IO2xENiSrWpdPr2828Yad6cqEBUv0iL+1osoZCQZKuoSaHI98bjc4
VTKlwE4U7VlPoHCVLWKVC6HrTKzU5Yg4vY20TTfy3Wz/2MtLxsvzXMEoQmy/I2uj
dQrv+NX6Pk4U6KR30cSVfWLBtBCvQKGxZZb+rnZ/1rInZocVE4CkCH+mJ0kbrcyH
sL04X+3RdWniMOqIsjMDIlhSW3Kzl4U2vdhoLbwW6eRXE0WhGI2oPLAbDgYhum84
gdzYXjieZSOaEvsmSTfzEjDWYVaa8EYIJnF2e77pcl4be32VDTynONiBCjRZs77n
CXIp8Uucqfi7yjVIq1NDCmAWImUCpq8l88jXwV+YMlSmojm3j2hCssFBqYvYldqO
T5rSIemhzAK6Q7jVJ7zsKzt9/P3lGUP9dWktnAA1ib2LY22hx+HLLJ9FLmCh1s67
9SkEpPUmQ31F2uysySv/tP4qzT2mquTJqWp3dDMCLoykPCl2IsPh5yYXP5No831Z
eEabwdIzFo5XAFoVDGI7Se5GE1zr5tQ/w/FCK9xLMVJCulAn/bI47776m2vqwviD
XMLSsuE6jkg9bPxbTLjBHcMsD2e6FY+m1euAN1t8T0RxFGkPnn38kBgiQ4N2WtsB
iBhsG6uZ9n9enob3HmFqZy7Ict56XKtvdNP2Xb/5PB+/tWOCuJSS83vB8Gwl0kNQ
X/8Uygvm+lnubnegZfFJFs6iURS9ZeHYizHVjSKijkb8egtVVEZMgBF1Mhp5bZSP
JGxnri8IYN9KW+DuEEU7NWtQ/qltQc7TkG95uT83GQdf7G07AwA2uuuCjpxHxgvp
jIJC5Bqq51rHDYPQhUOK+Ty/stdAhqXYpYGSRIoSNfx4OPqyGlnI87syjItdi65U
JkVR9h4v12z/Bhq5cn3a8T46i2tyH0QT/JIcpUbHX45eZbaxlKQ465fKEJn2vved
qF+kVUQTuGVkVS2pZTH+8LT7ol0uakg8JYCCAZrk6p79gr9jvY6Oxp+anLW7YoAc
T9lKdcuzdCZ5Ls1Xpb1cadsYcelE4y+qSADPYJiZw9NdOqGyBq/CqPE5AqFzB/Q3
zFZ1D43+ahzpU8OTIjsRpxIE2juwHY4O3cBclaGrCCA3rY5s6dM3HHGWWnIWpAEz
D5WO+ea71Ir3G0iVQOwo42Gyxb4Ltblyq7b1ZqSksZggZ6q6I1A5x3+tB/yK//vE
bRsH+FfZoyDL9iDfGylBzUBKU1V2NxUWyQ51cWJgEOgkjIXzbGaMdRIYszo6I5AO
8TzYYng21lYbR4Gm4WK12vERhPaY5v8Shwkh/RWArGg51U5LoZsFMRxy82Prgvn5
AeA4dYIl0FWwExoiK57+07tqtxS8ZigRvJluVuvXiq/QpTe844jcaPBjSYxJprJ2
bWJzIjRd2Da3eKSKKg7SpgP3QSSFsXbjPxaoGnO/iOFv4FVA5eruNh6ayH2VnMkn
0fA2y13Ban40cUrTSC6kmN1APBHooLXbk5uo6f02KCueKVS0juYeCH6fjWzZsueb
jEKvZ/dxf7WICqGNjYNzk9IyZGnfOwPVgjuxIuZD1NXQTPTP2di++PMlKlZIOH2J
VMmoi/EaHyXHa/JGJ6WPKA8uAJA1auyE2EMU6Fq+Y5c8VFStjAS203jzv+RPjGzV
5yaeXKwzhWNMRA+BV+lw3XtX0U82gdRtCP0gvDacIeH/izmZ7MLHl1j4oF8NPcZD
bwyFJ51hrYnQNPeJZ0CebR9G86uV0V/zaZgG0MWsa5O3xZVIxMvBtfQhckQBe4ig
nn421GkajgmGVJ1W7QjKI+SKJaQsorJ8A3IgEVt1HVuVTrVrXw0GVpAqi66qvn1s
ln7gJiMU5J4BCFHitixb8s1oomXKtMq3JPc3zAApYXTU+ZOYXOCw5BjMc4rYbMXb
A59F+IBUgmj3KKX/3cRqUpK5U86K+p843CPFQpXD0SrhXiepwCRrLfoJCnM4e02x
oZ4uNfYk5kYGQApGUscSuzvdLX1EFIlmR6x1Y+vv3bG3x5qPva+iYB/MzLrxROf8
jzSQhMFFqtppJmZ60+BZVwUONWbSdSnfkn1PgIEToGZx+6BP+tEdS01MNxe7HnEN
2rF13E4sGNwV4VVwZN0cMlwyv1EJyg5vU21au5DUY4igY2umpN6/x3Wn1OubXW6/
eBaZHiFUaCmxZ2Ri/oBxlFjl2NTZiVGOdsrdyEAiSfEpJG4rsEuIhes8NZGlsZDW
VVbjpdYPy8i9VA8Im1+VD4I1PRbbblh3dsod96BP7tVcaOujCuIELa+9CdphRchA
/SnvyaAZuCaxBZtShr5ck4DzBsQj3lmvc6YRBdkVK19GKc5Xh5mSCqbQQOy6X4QR
nPYTUqI+pWsHKwBT02ieqYdFvPvDPtKV8I0kqLAAu/FK4yvPBw7kii2LPT3u0kW1
rzCTsYFWGkNIgcXqxMCcF7v+ZsatdwC/d/k+InTfmMk9X1s6YIqzxJShuLTBgrqo
LeokaCl9C9gxxngpAjyJ9N71PuDz+C4r3cqrcUiiF+kECZdBj6G/Obr9J13iSnC1
T1Azf3ZxXOQDYyzA8oU3rUIb5f8O9/s598MlYpdY7RCNgE8P28hVZTdsTEZcPEn3
WJ4sRatYOts2at2xe6LGbiqI4jJKozjwu8krvBd2XbXu4icvzCSPuxss6j2I3M+4
NXOLoFXADFPdhM1sotYXxTjq3oP+PM0TSVPE6DfpgJ+AycV5Gfx4v6fceFX2GmV2
HpDwByaCDXYT04nDIoKJyyhSPUJ4t3OYJ+uJ3FdhQ2wxThuilEJYAgOdNWdS8B6v
xbJ3BuJxW5vQhqS9Am5LMORoOGxGM9wkSg3d1Jqm9MrJ53nyiev2NsfnrfS8McTo
fp0xFVg0udoLUW75Skzz8x8G4oI+Vy7y3AkqKudvGYcL8lvk8cuAhHWxdfpaHL0u
/tGuQEnXBr3mrcwEzv5OzSfVSiy1jZpNxJft0bKTK2fnL9QeYaQxtyykTzu8HhbW
SOgvveyDBSMgRQiC35LF4zpmalAbF9c13aEvizgSULLPoDYSHgVT2XZPAaqtI0mw
6gl1KzLq7NxRB+7AoTDO7xtaRooYnhCgFiXhvAT+akMsORAf/12oHaFhnEUc3woo
/QYm0qmHUULHLCb6cS3U4iNm46w1Xy5313b5djCDj66UyO5gmD4UeplR5JKR6tDE
dkT47z/dn56SIhii/16q19A21D/rfFeYYWTil13xa8nAxUgiTSt/agNTIs4UdTVP
KcHtt52XQD2JK+BB+YMmGij2OpiIoHR0UtxPxz92Gbo+XiV+G/kwz6qhPO8ne3a8
S+LXMVGpHSqdGMbfkhb4vaur4GpFENtc/m7d0B+8/D7lgkKQTiRrAF2g1MirIxDT
6Bj8Q/t1yM7aEhOV/s8uCuxJ7Ha6dBIM+eH5fBzS8wR367V5pGeAiBquBusgfcAX
Nja1aXRfXsOfFQOyGcLAgR5sbx5R2gU+37kt+EQbmLK5nzpEOw8XZv3SHWim+tew
AxSMJuHiHJIL4woL04d8sQOynv5QUtzFNV2MdF9QvLnHpwXU6/kw8T7stF4znhmD
c8xWmAvBDoaTb1a1Ai4VU4LXnn+S4tqtxSWV3YQJmDz76QSFkhw1261oaXpvMDIp
kYsQpaEuBFz4gzlsR2GUsKtXOL6hxQcRuqlhDvFwj1dxRyy+Pw0iebDxlueKEdlA
FXvOftVpAL1LUBVvqxjJYfqjMPoQg35Gw/0ybPU+vcD1RhionrzwWmHCFPq+1HUq
0FPbWoFuEJAO3iDn4zTdXG00wDBzZvX83g4z1sxi3FCaz8bGcEKsCZRHYXpu30NY
6itCMz4Cl5pNr8/iebmBpJeQcYE65Eb1m3zafdtzwCEDg6eyJOkMDgQ+Ve3uY620
nh5buo+IC/7GlXXGgmzNnsmEx8X6NIUCiPHK6FyR08eJDWPKDqTIDiUSHzS8LhU+
+NVM4dP8BQnyra9lRbNetOvQqfDFQmJUmx1SYY1/XJu43b/LhLdUQFRz+DZBlyqI
G9xtFYklZHUbP43Sj9slUav0AUxrisEagAZvX9aZ0ibNiV8hUOwnRGUVhxFH5KS0
ZIn61JCGNcsJGCfYV2tkXwyKhZaIAfExm0BrhEPP3a7Jac45Nm3eVGFD0OZyNCdc
DCIOX0mOF425gEOuplLBGbGGnkv9HM+7VVS4L2bnPiBQQUL/A9OxvDJOdhUUAF7d
c5abELXmXkQD+pZA2jzB3zXWuSubpaOpff12mP7Db4QZhE/owCli7oO2jiIjsmzM
litA/QdyTJTHiosHscuieQdrBHkwahRnZzf0aIi1dR98vY3AZSLhkcQAcCM4G10s
diuAH5jP92SGZvhnvKuH1xsNY45beuPbBhTsBqNZLG4gfnpW+4k7CGo2P6AN1i1Q
NRTvyrURkktMuUh/p7eu+ulbwJljtt0jD5hMwTDIfKXpHXM7Ct8A8Znul5wDLPqc
epjZqdwjtA7IF3U9YZqytiYUeLvd9x8dO7JxYKriBphZ44kB8Tca+gZPAEsARi3M
yJsOlkVqm1es4eSS4BBCiqOIYLd9aZ555Ar09gYWo/fiEpnHfpLYPdymTyO14KL3
aIylrOUlbvPdWSNL2J20HUs8wbyo/dnJRfCK+HoOfe1vyiFGoiSylwQWQyT44IjL
XQiS0qo/ZJcAzKpzbMwvC/VN0m5Ur0+NnuJfQQ7ifUE7KRwJDqWtdfpxooYx3lzb
tun9WYdlmGa+2qCz/xNRwYiA+QHLxtwjofZlT68vdzPJ4ScyW5BCtFQXpli7A2hn
63TSTsv4hb7vkxbYb4sARH5PwkvKNswuvq6lfengi8vgtFKcn0YEKp2VXKqqdStp
eQcIV5FcRO08rq6udfIyz7b4txUQJz0Me8j6l9JJf08h/96/0mE3OnbSAYeC7csf
IV/wmSV+K5GFuNxuF9aNOotjC1E5DZUpAsthiQ9G3X4kiHpq6qYiM+BvY2g9hcFl
nxUPD3E+tFjbK6Xm7o4MM8ao0vrsbUQ0GO+rc/r86On7LmDFjjLWXZe2Q+uxcJsD
/CnOVA8quH1qq2Yc2h0lsGMJ8o+fqAYDkyp6hnkG5g9iM2nR0Ejm3+rLuQxR9qre
KEuVX/5eXH8f7IFAFE8+GQFj/L3EvCSTo/SvL1yqAmubJJ0pTbz9aGAkh/NuMAwy
04hilgnZAmQ+NdaF1TvKGdw9gLDhIUhFm7Bb14ZgPCVCQOojmwAuunXVu7oqCKRN
K92mJ1QZ3MXQVBFmji9MgMkgSeUezQ5ODX1qbVHsWLYQi0QbM5iDklHk89klCYZP
uj3mVYHOIikzmJX++brThTVd3tFtwILrEQzms8koPpjsPOl1YPvTudedp2llq22f
N3jBxNqaJFEWAuE+ZbHdGkutHjsewPaTfL6OVEHIraXXu+OO6tbn5Q4mRNFDjJ9/
nuH/+knW7GFDLUcl/SeDhaEW7WWkFDWxblIeOnXCQuTwKmcMZGQ17S7K6f4kmOLz
FnzwfY6kwCHGByfvEcvpgHuvcyJLwhfFaOVQE9kvURtGej9FWaa68yBKaW3nl9pg
WVECbysEYyoA/glNzP2LqhwV95coxIoCzsXoNt5ysZoeFgwweU4s5n/g2Xjdx5ut
jnEcBntrh5e/Mmbso2mGuJxKFsy1lr+shlgOD2Rp9nunmVoszsCtrONElUGKLL11
KdExfnRV+yWsdaJtzOVb0NFprUKrer8/R4S3PGY6EY6wnQ/FK4EYUJtBb2sGocEq
1E/kDxsd96Zo1bYC/Og/9xEI2Uj9AUS1hYUUI64GwGFdLaWwAKhW1OqOyb6fb3il
rFWtdDRcL3hymLMvpiuSsogDpjXScoJ4JkAymCtdofSX6cK0hcTCpAl/OycOLmmR
RjjsfnkNtDrkFniIbtL5uXs73cW3OXAj5gIpjyJ/0OnlENpdrjxUoKpD3F8ssMNG
nczBink2v9v0a175g+y4a2u+IaOs0rnFYTpG/4AQ8rf3Kjipf6xZHd4MyXo1GUPt
RSa0hlnKYiVnwSPmsNIjXAh4K5jaSsEXS0X5p3MXtat/QOWjguniahJ93zudGLdO
ZbLSv1StOUx6U1rhVjlDZeP2+xFMqohB8KyARnGi5J+8aWviweSF66mz68FstmJA
U3XECLkbEh6NJYQJbLYqMcmLFn+e9XN7iXc5J2pxDU0G7Tow1zZjEVXNieosxk3x
t1dbkXcrmmuxCKY18ZwWFgulcXOBpRKo0vjLsKT7I2WWwAThkgIgr8vC3kWJK6WG
Q7LxDI4oZU8jcVsdhgkuZHnrfNC5dGCcpqM6YcKrwPuG/S9nEr4rnctmYjjnTY3x
oPqTKN4doVKeVJDAb7vLEcyYL+EgTmQJGWGq0dpPz+Ga/vRDt2v4/OLHEiOTZi18
7rlQwaBvapQ+7usU47MO22hbLV1yqkENQJcymyJj8zJxvrINPS3hpZpFJvzq6iJ0
0THWi8QI8fTOPf1L5dwPUsgvSEa/AUpX485nWEgGOGh17UFiXi8XrrmzmQG3jAh3
xvtnJEjwTWGrgMymxKY+rdTifnb+P2ZyXX2MGgROeAA7BnA+PeZFq/Ii8c6gEpJH
ptVqJq7W0YjaYe1RJo1kMDginwStIr8SMsr97guwO5YXjiq4OVk7aClaNLFGm5ti
VMJ/8DUef+QPmuxCJhxNsuCXuNGdwm/jb1Uk0OGa6FOiNjHPaTPTkOWdpi8Qexdb
vSskUbsZ8FI0w5Vds52F/zxJ3tj0PyNsZtRdSzlxEcFSKiqgQK7tThLoE1QDRcUW
jaOd7XV2uusoR9SDKGE76xN0VZu/9JxLsdUmu/YPia0qhtmcXr9Zq//xl9BjwGKo
+Kf2KUPpB5zSWq4abgmpY/4MIitRUL0GPWbsY8mOVXaOeQVzZWpItdDxen6iMUBB
05sJrUu8CI/tAu68hkFjn+tiDkFp7mmc9IZbSfNNuVfuA8CILJ97If87EJwton+k
kAi4RD1ynvzmKzPfwTwyNccxCoVNej4IaXLa5uRQQIdO32G0z1cortXnl3u+qkUe
bWmCdjhpO+q0hLzxit59bQgGA/vJBdTMtMtFyDW1pbBpbQ1+4aYummbkIy4cd/Hb
pfsSo5oMEq4AYDVzYphOc3o3GTgyQ3SjVhnVX5zdlxfyn0DEDLjXlp6lIumBfXHh
7jyvgQhmD2gkV/teRanomuIYaZzJdH5SULGUtAYdM5hBtl6Etq3Ogel9ik92EX0B
C3AaoyMyybbNtgI7FxOWc+UBMPXHNmNE193gg6dC7Eofm+EY6gMC4mBRUis85jz9
9aiGGwM5+5ieZkRS+LWsxKc0/JTiuk3A2vgXhTKYDDBNrGJ1zyr1EZyY48K7KMqb
dl1X0BNdxCJkYVk+hXPusvcnFsnNRX83TDFbUzc0cAuK/TIpYkMZiT7NOcIQTApX
43NT9ryUYucPf8yHFMk6U3QG4XA8kcC6K1shve20R3oIb3W8vxEwMFIuz2AGY5AJ
KZPz+2IratEi6yQSSTUTKo+rthqcuXT9oJxPOGkr+rHNl11N0oyyaBbiLLylymb/
ALM4I8bqz0/xZ6NPt0uq0JYlnLfiEL+BxmSiySInbqu65FWOpKEwZYRb3bgh5RiA
JKZ0FLkhoTTZjfuYh7oSbCMBnUJFaxWIR/h575sGpGy+tXRDfWuH5HEyBr01h+Sj
bH8A533EwmO5ekzZE2qUNggW1FQFBzZkMlYJTyDulhhMD7Av5Z+VTd/g8Ncm7aIr
v1sGP9qa0u0pfS024ZWNXBA1TxTy596e8MW4g0rYm49H9sfW0ZX4WrPjWbEiUD7X
z7UPrQW+rtbB4VWIrZ94LZxJemnzPN67kUHp1euW5K6RVcewOlFAawUHRRYUxQq3
WlYAm6WgMDtSgPdYuG1AuvNdbQ4kpM9kTH6WazBQTAqzBliI0HtK/EZR9cCqVUm+
eAcHd/9DK1BnR8aNgbdd5wOF9J8jwy3B/U9mUG2ZtdUeMUsgvTk2+xDsdGXlKphb
St96WKi2xbFIQsyr//1Qq0w78ZOoMiEZyPpBbrQ2NPy4xLv6ReTlUVo7hlHUYfX2
a7mSrdZAfCE4VLJT2aCjzD0XH1FE97vYRgUcA6CzpZwtHY5dA1H5Uo5Qq58t9fVo
Jnh/IbE5vskGIptGt36U08QXwHAORtQWfkJ9NbDZPXArnoebsExzOz3qJR0szn6h
0aCjo2wfvBSQrU8lk6JrPsW0WKUpkCzD+oEeM+WFRDmmTDQoqHa3YnUG+bx6S+b3
852xuotKZtYsAU1oI7iC6/7flf9yfBhyrFlrYbrLXjgt3f1DiQWtJSEm7ho2RxWV
kmn/4EZ1Xi3yawmCziIgnK2ED8WmbypvT8rCq9ymWcmxnYlMI8xxKrWBuneVcB6O
OFUrjvirXXspVIlNygAzFLtmMqv9p1O1AAB7MocP2CfJ2L198bC+seHOAqti5TFL
z5PORu/vLfUXZiUX1/agG7PRlcAemPTbGb82VFd7hVIUHdy1CQPM4xR0VqHsjAJ4
7atwwzwZRPnmSN4Pg2vHOgeBiDl1JrXF3Jg/wcXuo2bmVlyLZMnSVYKqTZGoHQYq
/3zcbB0hmlGG1ZCSvUEumH6uXIsnWOqJTy2zz76Fg/jc77S2FuCx/ViFUjNA1W03
2DgXp1tz+1H4Xc4CqU1E0iDR3PxNQAIFViVyp3Pvumr6QvRr6FqTzdIYq7/UlExb
bpCBpKC4trBU6CI+71D7bjjw8UbBaUghVzZtYSZyx2i0CttkINyuZ1uu3Jli+mQw
SWQuQqkIbBIcnGpWMAvP8lmPP/jczyzLDuhOn9os4Zl2X1MKoFs6rYpB08Ma1S5T
JqR5dbfDsVaWnI9NtOz26tSil3atZcuqJda4YH+4ROd1UkHf1K4zankbnvkIu/Tw
duPgZI2WuKc6sD4ObZZjP0O4qfJkURy3KU893dSWAqunhqVWR0GS0k3JyouNQxMt
p9JGO7SR5VRVY7zWMX6w6sQuwPNEeat5As8feG8QEtKKpWS8hkPgnUkMZ+noKftF
D4vEDvNwQK3pT6Gr3/N3LuCT3UfO0VWC0vmB7v5GW9JzeCVD2PnyEDIysGUOz6Fk
3uSNfveksyBQJvNw1Bdt/tkHtByryg4SM2Kjt8lxWCMzD4I77R51uFZbS7Ovdouz
QOCcs37lYF0IdgjY3JVwSKFB9kd4wZSUdWnHFp5u2dKxIoDNYQ4isUfd9kGIcm0/
DAFr/K3//j89OTLUZ/IqXvjOwcqSLGSL+sobEZzaSRibgC1kVr4aosJEaPAAwuLK
z7mtQzVtolk5ImHnzhqDAI6tf0/qOCSIMEjLU9/yauwQEczQJt8wAgVOFnDtGu2b
s04kiIWCU36HvCALq6Lldh/C/yMaRVxgWla497FGbv+Y4cRy1l+X1Pv6Ag5uk8tF
NGgblVEEpb+D80P+G8D4J4Eon5nTnGQuzGtDCW+oNErXXaaeWWFRS1+KlDmhM6yB
nkhxOwOc2Bi2+dhn2MeNoYmv2xmZbSCfErJvHWCZMtRIUT1+6vRiMYzwhLnYXUzc
sxMs2ixRMjdFub5jhHyJeC4th5Obv3+nPBD7ovf5gbTL//q7ZFP/241gKobJB9ex
aHmDkBHJdJTXY8IvH6OUs6A1rUuyRruFIMpdwsRtyOhVoCDPHED76CcfKd0YPJM9
oa/exugeJ+5ZbhTXbkXbPdj7RTcGeN1qDKmXHiF2yk+1Ab1uNY39yB0JPFW8iPd7
zS+lJj0dVNfs5lhZwKDumHf0hfICSOeeoVLn33R8KJlfxLlZIkNJkaqx6iqs81lq
mjYmtobRyxgsSoIUboChOtuxLITLe5pHSz58mSXCoKnQi/LORd4snH9fKqPCcBr0
B7qKJVwRKUP32MhaJFnr3aZ/XfONVL8hOc8MxllrKHlKVbla34x0kvAL0w66//pr
KOrlKvQ34OrW4hXXbN6KvE9pkZPus1fW4oritnk8nJ6fhNfEgFIIFTp0Ue8pDvgA
SHu9lpJ0skd2PgUOg8BV26ni1jUuNTBZGCuj7dHsBM6lYBV3ebIQ8M2A8YnL15vM
KytUyNdKcKXTBHFM/ailpwSKKsKxrzXgxWgM7EVnib2IYPjoCzyxPgnRjCSFPNnR
hnixL5zeLXRXKlnias0xgl3lc3gxsDpNJMKRpqI6qQTgqh6jZkZbZ5Vh+FQj3anV
nz3HMhuLQGQq9YZqrKKn9xR/Xiq8C/b5+xybcV2yIeRBvvncPfK+X5WyGQeSbYvm
DjXfQN3gmC2liILnqGS6gbOmoCn+eIIpb2BnmObKTGz+7GZZ43q+kfMR8Jbvq508
XE6rfg0sFEySgMIxtdC5ZAywsabodl2ewdWIgNCsKGmx0HLng3jz8UjFtvSRxRWj
QMCBwJjovg4rfw4HuVEh9qpvWEOraV6s0g/X6ihoG7DQRIUdUSOLU0FZmQHOKdPF
fqhcFk4cXZ49PYve2MQDgUfuemXvGvq3N8efrlD6wvMGBy5N0CF5bPPzAMH0LdwV
oVEe06yDg4rRMOOXvF2GIL6URwZxyIF/znAZcS4j0Jw7tYzGIazqs7Dluq4fL2HA
Qk6ZFXiAh/lH3QB+fV0MOS2rbLwA/uGZ+FL7wKi0Hg+AyeymhMElm/EDtBosaUK6
BvIptuRjJWSvG+PKQySevyfro4TzasVX2NUNOTVKDDt8QwPZNVN1JD1RSHJd9TnR
fa4nVsMoG9qdmTSmYqao8neTR+4pCPJOdBbYt5EgWmatwpW1xie/70EPTV+gJzYj
4Kb21cw55GgWsot8k7Cl0F00cKjyTNS7e2+WgY4M6RmI7m4ZnvNahGgjDHCk6NZo
cqdL8V1aE3lKJPKW8mNYqAevYaj9Swwx/4CFWDPn8qjHYhjVLx0gzZZLdilIOI+6
80q1RZyCBx3x78HFVFrlhzRfbOJ9h3swBm4UqsWZ2FU2Qa+uNRoPJz1AGWdAmX1R
LszUPQG4FEJ9C+ICmzP58geWymGAaibBhCmtUHXemz90UsE9QrCAJiivmLbisU/H
x22ACvtO4ZcnU38YaQ6akUsDjhwhuQW6YN0f0cpiLbQk+AD/hwbBr1WvlACKv76P
0tkE18epi9dFI/WTSqPOcAOwX/5MRpkQbDtWu1GCibmpcWMzxKVE2gK9+ry3Z1vp
2xb+2d9y7ocBIHA2zzNvkiS4cIPCwV+zaZuvLtkZVVLl6FmkSqEFmG2OzvMblNIK
EyILvDst0gKTiH7iVgBEamxwQCZ8SoDYELsE9UjZmuaq2JG++2FRV8q3BMQzq6F3
qu4ZjaWHWshqdt7CYC+OYYlvS25tijf1R/ONPLzjMHBqPB0A7gETAgNAajsDeTpy
SwRoMFJigoZZuVq1yixyS4eiwjB5/rI3FKJ4ULGoPMBYiehAd+Rk62uPyJp6JCHa
o2mMh97gvZZ6cgwtBpOjEVAJUHDjnTEEEExpe3EOBybYCSUPTKuJkkT43nVVTwfn
S/rzo2z4TiIIge9RWtkxOBr36VN2nsfEZOy0QbIHth3Gvt6GhvHQOBRvazb5P7+v
g1U/HdAV+FwE3ab6XT857K9u8oL1EhKy+4KMNgY9pNB02kSE4dNXz5vlkb4r2fol
XjEKMB2k0Gtj21W6T6kMsr/JSyMXYnykJZ7EbET8iZgyQ7n91Kz0gvKgNF0XEfaD
lGYIna4uvOqsIY74h3rToe+UD1ja6JrDEH2sFix5iUALCoN+/Sh61tgsTsBswt1V
yys+r1pk+eWXhHERdmq9kUvNuDd6xZXWvr5DZ6FRSJsahGgJy8+KU1X8JqyZTqje
0gkFzrdDQ4sFW8uG3OYDZGIlt0Z6t2FDT2hksXCWMRA5G45VhUgmpms4dK7uq8wy
9GftmbvqR9D4KycZM/rKmLu52CdRVp3ZJGOGdlAYInVEyed+eX5UTCJEfBimNGmy
VTwjEF+NsId1xBdNw3VJ9cp5iyC06kIaKGpYMVohwMeN4ACwXfYRzf7jgt+3NVQx
SbHYyVOariDL9Rg3wGny8H7gF10Zmhev7EaG/G1pzdyCmuHUQgcclpkPCMjdks1v
Zf+Yf3CvR1I8/ua7KC+lPiP+eKimGn/W5+hLOjA3H+k52SzQ0kMl8KxiQuJACBDK
t44ipM8ED+bO/ZTdG+BC4ZMtGJqfJwoK9y/DPzS4E2V4YVx3mi2iu0WdNh9hX9Vb
ZzfzxTahwBC1rtCMpdvg7IMXtnvB49x7HjYBA2bBM0oQRy4lG0aeVChyWz2UMBjy
CVcJYlM5rCI5DNuKk5bBagppMLnPttHZQGU+glWeY590+jAsLXHfj4eHsLTKv0lH
+87XCauOdJKJNmlEjOuhHwIqAASEGd6MdPIVKJwf5Avy9r2K/f09TVElIO8hdU97
DJg4qoORFAbGzwkPRTWRD8GnoS2ulOqouv7oXD5Riv+kNKe9+Ruyfj/ToyastJaj
pqwqmRSqF4i+tsS/GNFIUapZDdIAcI8f0rGYhaFPIfmZZT7kKhhvAfmqHu0phOLj
Gs9E+IFEO9czJvy/inTHx05IWljsuk0Hh5oqoFYFHhtq06CxvX2zk5hk5/lS1Xup
QKzKTDXBmRC/iWFFwhla3keM1aMgjoB3oHf+XuoqmwisyV3+TIedDvQYOPNzPG35
Dwz8mrj6TtSzCfFWFtIyDE8Siby5XRA+tF8FafclHDRbFqeNpQM6q6kdh2uetivx
tgCZY7DDIwPhsP8NwGFyvnDzrZUJnCc0XsfPjWAR4/128/nh+m2pkHqoJEattLdY
8m1056T8Xu9kH8fHftfx2qmje2tIUXVrHdZYyi2G/rBnKcAD+2gB9lvyvPmXtTJF
hyeVmQGyDLyeA9l9+RVII/PlXOci7HtMSL6sLUA2JLxTNvXdB9qWz+9iJBrDKM/p
Q4uhxnpLCFE+1ahBw0VfwWLEeS7DIxD6OFfnAJRZoWos60iJX+zCI4RS+mku1Xkx
NSrXEEhEdh8udh3N58tTrJPjp5d5R2tjp5bHbgcD0sbEB0ORgbnUtPYsr36VhWU0
3siwqKob7I4Yq4Vf8EgXooQioeplfhjhwM2csV/wYWoNckeYkx1hsdPIG2gJWOZD
liwEpmRtn7OjGVCkPJAjpSVz1EvvbZVk/X5qKk1dG+d9dc+8fObaqDl0niLWOWAm
CssvUa2nnbKkjQSQe47CtOvNrEHJvOfos5GDhp8T7Nf5xuCVj35R4/YLeMb1h6Fo
RQhRbHjqJhbZYkQzVnjK3sYpPjQcYWvloEyARR73SwVeARIfTFM1saxkhh1OEhTM
Uz79BX/9yFN+5dsXx7S0qRntA1ZQM1SSeOlCH01/X1svbapWb555wdzKUr42RNMw
2dLdcTgkc+fySJAPRaXioIKPX+4Dj+/I0+99rzf6aARPweaQBQvuubAFWjSPVWcj
vOCAIIQO6nWX0/BBII4pzlyq1FXRuTbcURCLJAJ2x8pk5LQpDqP2F6INAc+SpC7l
+ehU5onC3phWC0k6MRqgrpEwiDbfRZ6+h21LkqKkARrRuFXi2QdwWRjJuWBP3aOg
+cnIvIyjfaO2yqPpBWqnYnv1nAn2hnaWMQUc7xkBPiU9yx18xwNEDAPTBy2qgocF
6fhXYgBVNvdYGFLGfuUuzbYBa24dQzqpTTEm82ejJQOJJhIgLhLUU7N8eughPCpa
RXmh61aMgAKZZKI2b5AV6bl+q+BbYKFlGZi+DKFs9lt2dDKtNIPZUqoJdrhk53By
tzyRL0OiqdOQQut7OMZFlpdk0bTBH5wZSEeQYET0mp+m9g6Q8+jK+efRjjoTN/iF
LL/x4hlC/KXhC3ZlCSBZusVRqk8zgk5ppVlUm767O2R0rsye6NRucavqFGumDz8z
d0VEUaG3UQO8aajWdnJspKyXAEWTjlWyVyL4tN1A73HBwLCEMJJgcwIFvf8YROki
bllh7mHDNHydCvoN7BwrnHtZuFPh5KtZtYTHxkUfi9d+fBS/paK5zIib1yJNXhbG
6SxVvc8LY2smAgoRNYkHLRxNYvOSRJOEuXNBfuPdQ036hjHW8E/owGcY57woB4hA
GG8OnmotcvV1eb5rzU8FtUSofPEFyLW20PNoToa9AOM+oGXAb7er7bk4RGCitE8Q
k1PSA7YVv4vtWSfYEA1/3O+CF3jtlKFdQ4RxJMZk+n5AAd4Sn+8J0Ri9z1gQAy42
QpG2kxXqtrd+moh0EEtPp171UNHUSDZMg2Yvqk4qv44EmHaYFEcD/56juFbGg2G+
Qa7DATzhkK0VhcLB1N3sxNc6Kflv/Qbm1LijFvk28lDxAG+JDf6F36RdihctjK4R
ZTUNa/n0nhDvPzhPV31XoBcLA36qsm0RC7hI53k1agGB6XAv+43nhGAPIGePNPkk
oYANGHcHS0AthRN5ieXZgoF2BNfrjZW7qBN1RjHPjfguO0qnsxb0j5pFxsDZB8uY
SSWi6/Y5Jc36RQw0gT6cwU37h1BPjnj0chjLtbmODtD8WeKlQn3z78XxZrA6KHXf
RfDsZ9SWfJDkfnz1/er5RdrnrVv6fhMjZe2l55YkF7tJIT19kkOkUigUx1RXR+6F
ecPk9NehQOu9MxKj648x43/7HHc+P4BZ2PSij1DpkvEKw05k/OdRmRN3rfahuy+3
eQRdKA6N9Q8W/eTFBhFjie3X8qQfsB76U+T7/XqXE7h5+Yi3REzoHGxOgnKUkob/
B0AsR+xf5BSEqOvpyo0dCrhXB0rKt4f2LvMyCdUoLZpHUsD0iUCRfF07i/IDSjIK
Czm3By8K9MTsrFSlihEJBhL9SOdPHEioTXv6LY41mCj8O/TX94jeGIRpvuJQXElo
FTvdYURXT2cd/Qn4JArz+hLx2poYFlb0+pM9Ai+4ivhFttpnM/CAP0DU69QhJwri
kgUhfytOC5UtyvvvutzNGxRgKByFo21oV/9zylcC7TpOiOFKmtlNFQmECF3XRixq
QH7bvOZcnD4RRkD63dFC8BGSaG7bpY+YPKou0QPogCG6hMjoL/gXdo27HSvhj9md
Aw9oFPHH739XTmDJhKkFxYwr95HKyH5QjBw7MJ5yVi39oiu2d5liVp4Hybcd60Vv
x84uV3NwEg8nMLF33PA0nbuueU7QGqQZ4XKwZ/w1iUdOUlhRzi5d+JqvSycyT5Zb
b+No60PMkUpACXmmJaaCEXtJbY52DkOH87Ckl2BN4QupTl666QO+0O0Sv8Tj50US
0byrcKe+j9WKluUW4p2eskW/kEFAGVcXncINi4JHvxHD++As5i/MpcLWdUmukqW0
dJSLoWAhjrP0ZpwUNEk7fENHj5sSh2LO6oGXLLjQnCz56r5b9Zh4qJp7+P3g91+m
ewReon50bkxRWJsma26m6wxhnhZCiMwpsL1cg+OnLWQibHUo0coFIPDyhHsJ4SHb
YgfBMnm9zoMVU4aNf2YClm4/QwYxuX+8xaQox38PxddA3JzSvldGB5OL/GuihHLR
jl3rj5i2ox90ldQ7MKEp0aFZ5ANtUQLQbImjgDnlpv9N+vahaz07kvHEsEVKnpRL
6g97wVmW0emkelywsRb1Bhtrnaf0ZJaTqkLbjaQq7u3eKzKo5FA0F68CoOhz7PUH
cEQeHtT6yBIYRVeVHBiNPMOWA0s55w0YfGL8GDDVTQ2d9ceIqkAfhW6sWqVwVCW9
xU3CqmQdRR+w1PZ+EJudibAYHa+LozKdW6FPWbTcEBRv2ZkwsjVcZW12iDGg7jA0
t/1RE5zoI4m6lrfjDWZZYBj3n/h2pBpruTsplYBCXjGSJY6k10SEojZVzHWKCoVe
od2um44S/jPNzqlzk5AIe3k7dBC9W2l24qBRNSLfSFxU0QDQET1ue0+hLJUO+Crp
RmmhWrResLQ5KTLNci/L8538YxQCZNSzEmLz1RQWZ2figiNY3Pn/gaWzVMFvqYHX
9D6TYYBOkKip0epexXoFJ2xz6xip9yRVMzVhaWdgJhreF4tPKD9lwiBoURJYlBKb
VM7sLZjhZsMtzfLKiS9LglY68GpWDLDwSoAnrLQPw4Pg33pci5EpS895PkbCw9hq
Vi0BEksKe+ekYcm6eAhQ6dtQsE84/UmEFL9zwMKWs71chWJd50KFRFQ6pSS6WKDa
WPeCWdzF5navd5/fGMqqWZSCbACNcbikzYcktFyLEApEqi/hn0LBPglYsTBdfVn8
GIytsxkyrqxu4r4XKVruX//o8N8+Yt8ra0G49AerEEqr9BVHuyfisUT3iJLZBsfM
Oy7T5pR6UeSfV2dLSQqKdbGuaGGMJphYMmYW7A2/t5nNcVdh1nfuBDG8mmlsnhvG
xiwZXmB9TxhlRdCE6lacXTuVjEOMZFmkvcwQx3RAYNXHrk2J4TCSnJqWMpbgLlov
cOlsnHwxnL/lqLEx2wW/UunXgiOIZXANiMOcOGgvoNGOKMYkednVP2yv1SnVmb/D
kiV+zOLSkzBHF7HVNdI2H5NZc4+SN/O9uBjlPm0sILZKNl3IkXYRfGPmz/iSGXUB
5hnyjWdrpUGtopJTAPSXiYpTpx35nkZqrubLbf6tCEnzgU8jXWQ4ylc4pWjieE/D
Q255VCQGcY/K/2x7aGIvGAPPCKT4VNnLgnqqlxDjXYm6aAWxcqWoPXcW4jdEQrwT
XQKbJGba8bTHEYRYW3TSdsNNHxq0kHtwkfRxU8C691HLcWfGd8BxJhtkACI+u6oG
CM5341gAK3BysnYF72a3PgWWCPP1IKCk2VB17lNOxTbwF+Iv4weusZTHc5Q7Zxm9
VT3UL9L5OvJv5W7csVpHwgBNUgSW3BYM2Mfu/9QW5zX4q3cd5QHJegWCbJSU5ir2
fZ5cSBENyoSdZbb4g868munr1+Fm7sjOrrowLEAhjSnmTVF51vgRyggCfL+hc8GA
ZJYD4L8MjzxhPcztvfzHXv3P45jkNmTLumndvo8Hdi27KjURuKIh8fSSlTviPQNL
G1SuHBFxnmZQl6ANYJYQXjfCnJzZYStReGCTFGBnZQ6FJuY8mfO4EeWFuKeqm7Lz
KyGq5Z0XFq9r+CeCArEi2eoBW+WGuh8j28/s78b0QtqIoVRT+CXsGdU20Tc5JfwQ
VBYL/jpAHSsUTyIAqw9CgrLaVTJ9NAQ3SYNM8h07jawLO8u+nSMNMGsypuylaGv4
A8o9NZGvvNVPK4neT9Dfal4zEQ63+gqQOpI2VBJ7Rg0uMT6ZEltg6dN32jiA33iX
Z2xHDGAUarhcUuWPpVOzL4Yh9DiamakrqMI0P2ME+akh8IaAJQ47qgpuuDZBfj3Y
FiCWOA2iYBJYnCovD15FE2NDcjEzgAxV7Hgniz073Od3j0oFwARU2PFzcNwtppNJ
IvNzQosuCG8hlzUclXpO9xad8TAUwTv52oVcSSwyvYBACkXxFKk0s2fvU0CvuHwu
X9Ej6pO57yjOO23M5D/D/on4U8q6ZJC7bdD8LPhooGBj5oxmipbJANuSd1iijJiS
sd6AD6SCWsXyVHRqAllL+x1egJp9RvEeUDiM7mh8Z5eGb/2R2UzHeDA62d5oHyBF
H3fIUX2rqAfWd0wAn5RqFRhnB5Zs3WERHx2SK3kYgK6FMW2Di5XonbZFOV30LpiG
viFY/G1IItBIoIuyBOblpOvF6e7RwJdHERSe4MV06RJ8Qh6eRPYjiaLW1X7/hc5p
Itl28qhr5UcVNhxost4mx2y/d43AKED6S6I8UO9KKn16f21qBHc2YqWhHCl2/Uta
EaYWyZEN7B9vSU+c2wEgTGDZsNhg/0N1TvaiI0zRrNC7kFNRojhz9mUdyWFVMC4j
v11ugK5XyMct3wdYNfIF+M57mk5RgOllOkaZoHR4CxGCYHnSl/+WylsRvBxGzqmC
UHvOWN+zBXxBhS1GqM12vE2WQ7NX8jtq8WHFl33usYJLJu5zG+iVU8Fujg5wT4XT
BDYQp+SMNortcUfAZNMyCA5+bIrXH6F8NxICd0m+Fj1D027PQ+IgRohGpOJCbw2k
h3IPLSXIxBVY6rxde8ue7D1ziQWiXwnc2H3zEuHII4nes4O5rvSjVDYiRWdDe9YV
W/JnpTNDZqHcMJC/syC46zFtGXNuTN1fzG8ou7t4lz80MM18Z1ZguA4gGxagr9lH
0P+5XvFRSpbYtT5HrAFFJ/aUCxs6yU4E5RsxWh5wlKBgANNecEOXYcSKmnM7H50w
2Ydz2mXfg+k7/7Bc6wOm1HqbpLtPVbOwwbZ8sYCcM2aEKphUvssscvV9EJspBkhO
HSLt0lpnX+oLJ5pQwauhoomR/0xvAgxAGbz3y0kDFHQcLbQiCOBkch3UIv8Fp7Yt
usSBc73KSgY2ziXc3r4wKdUskkHVLZYEN+qB9GtY9BWENnLm+KlLp4QP1XZh2TVF
2fTE9rZJdQoVJf13wd0ViC73vXmnd/HQIqMO/wkvKJQwsAL4Fhj8BAiC6ktl8gaP
nVT457TxOUJE0Q7GU10JCfELN8Fe2qfGReql5si+UmwoYMOn5m8cLbUkm/p4sQ2m
cHKfPaPJXgCzLuikzY2PBRpGyqvbCFMEh/gx5IXirbpETDoCAgEIaUKdQt2MAWOg
tlBNxuvx6KX9UPvpxQCv8wRITaSWhr2h6/yXFgxDWHUz8NB37g/Vf9T4wfFLb+Ok
EcAVAD35sKhddVlgMTLx8yR+t0emKNQuEHBMW7J5ryBtQSQKPNL1hjEQ3QCuMkx2
VkVCOSSsURD67iEr6nu1LWvSM4JfyckfpixcgV9zEn4rAMTsQBu87EIU+QbUc86R
NX37D0oZY3rI9oOcgeT3FZQVXy52TcvYTvES/dU7yQDnMj9JYV3BxGkylY/TcDCk
h4AmaDPdw0C5y+5MLckVyonByf1LMfM07JI3QnLed832VVLtAOzDQLXlZOrTnV8x
Pa0187UhaTfvXrFufEClY0jbzJzMQO4hPW2KPMx3AbZb2VCx0K/shxsm/khLQJCL
KdWoQFril8hsUwR/vxAJGTJk+Jv/Ktc0vnytpt4eUwomPFlj9D+yxU+m6K//+cgt
M8+4LcsPNdbueL70Fi3EsTMQ9yU/BI1VwVKBkOknxMtkR7cBC+dT7dPAsLmInWwD
8lHR55vgb6cS3nWYsg6tNIDK00Ge2+z6mEeuV5sUFnxOiX8nkTkGjJXId11EPrHq
KWXj6Ng4Yoh1tpCEfqLKZWqSILmavrHUstyFsgSQWIP8uI5CeB30zrd/nW7Ui5B2
edjUn6Gg5NF7SbG2bZkbLhk0gpR19x0P2XQ94F0erSd6vbSZ5KO1ptLYJjAcbVvE
/KjkKi0jcSBi8b7MNFawOjLdY3ssZe0q6pq6UfpmtDyW4Swb3wGwX0g/6rT+hEd0
sWzj9jp8dEVIdcETzqTpdozYl1s6zdGFdiY3NjhmzPfHxRcynczreylTQBiTSOyc
tDoe/xLqy1CjzHm68c6RUWqEKnB2bvHkfWhbtwpbqcIy7t9OBF1T0y+U/aO1Gbf5
irYdDhS5in56x6vrfJWORGPPuyU/pqFZmn7NL/MI4trlEhpmdZqvNCv+9dHeNDL+
k4tCnHIe2a4zTpGcD+SRExyLQP7mwho2XEb899bIL6PTA4rHn09yFQ7ZzXuJqRrO
RNmn6fahLZY0FGtwXA3/MZYMTVi/wFwQ0eFXRCd/QkauUXr0zWqEKpqFYyiVuh6i
A7fNdr6gKChe/XylStzL+CGN5u6Woa5yNmvX4AiQUJXGe6amyMjbPt5AbbL0ysbq
iDU0a+LUP8ssx8i+WLHY2u9qMuzEuPsNUeGe1rLLrIYLWfV5CXz4jkgga0vttvsU
Bjm70rng3VOmlamq5vT0u7eWwAPcq0lGAgHf07q0AomKM3IZrlbeeD6yex2TOR5m
lBGKuTCj+2j4/4bKVbNafKO8VF82wFPYLRxejjJ5MyINNDKpsyjoPWMIcqqps2hz
6GKe8eK/TH/jByffrhGuldaKjyquuWhLs/jFlfDyunLv+By7GnFBxgOU/Ph/f/St
1a3oH23EyIvcaWs5WnxEtDudPevOFzps/FDGpg1npF6aEp0k883taMPXVHLRvopW
zvNp67UIziDjZdbIl2suO0Jjgft8hAoS2xMISzs7kErjN2k02mjBtlZ7sr3cWtkN
IlbPfriPKTNWhkS9MFgjFDfA1BG4FvXFhJPMOooNm8ENpryd0KceIxXuWwhKdBWX
JfJi4f1C0mOtEhJ7KwOf7sPAAlJQR4IWbO/U3VopY0TOB6R1hsLxYM5TgblnaQGx
gc2rILZTg0xviANSSh2KB+EWj0d19qGIybIHTlF0QXrIANLjfHzTTTf/7+rXtFGk
5I0q1VSRHR++BKAb98IOnlLdedMOYla9fhiXN7DZd9LOr4ChqUlkNqkCzRFfOWLC
pickZ7wx/YUznhHQDgvACZc5vp3HhcldO57F7VHU+MvfJ7928Tl4KwYkcfaoJBFn
yHZKs5IexurGBjzifEj2bCQHzJLLBvUM8u20gYJkDFZNFhZmw9Tiu3XvBM8wnyE7
x+pljKVWSLXh9mKyZk2xQKyRxYFIIFsI2NOcHyn9R8Lw5T9uFSsY9Yx3QwMkNnn6
i1/2Jn1is1aAcJlbNmW4yw8BpXMESUiLqBHn/ZpxAWDz6ViIBThA7qw1YDM6Sh0j
aGEKx+S7gNkSpwTsKVjNW+RrCF/E/ceihFbAwg4BxdXuOzAULvLgsPygz0lTrN1Z
UUbCj3BT12Om6vIwYPI0HUoer+snB1u3OeCx5LyNG5gO75YteN79JJYYhcpHb5qI
9GeWVRWX5BnK4QnVXTbbi9u9NxobAFey+TutMoAPFe0WvmuOAIqn9oFeCC/t30yw
HdAQfWEAox1tlHZM2K1V9sBsLjbnbVqFmBrXwhGOfJMHBGDY4+gwFZyDr/FSckcO
/lPp9Qs0H9pUxte3/Q9q+a/qHb3PWCsOUyaLloa/rAaEVusrkFm5fqH6P6RkS0mb
WKiiTgIz5j02QKAXQQxGhYsA+QzJVxRT+to59O7u6WX7xR6iQ8sMU2wHPAWBTFRj
o8NI53pzgzRvZ5wWVPTcp3/qLOWSgyV75YDZjQa+iRMyv2tEJMfxGXjAL9VZ42Dz
rz1fDyG7jXX8sK+Yc6Hi7F8bNMgrzoF4SFRtJDkPHSkVRZbvMSOkj6rIxg0uCwZa
nZByWTMRXONDGdnedGrDaJlaio7kSD3HHYEMLXLsBE5zHyz6AXfZYbqTZMPARiJw
ruCsqTZfyHUQ2XPpD5KGSuJP34nXlHZv7yrHM/RPLQOawXXS+y6FkS2f/zQxlumv
6judZ2JgbUbrvZD8BsTPBCOCIXRsTHTC2yKQwoVG7c+rZJa8Ph5WL4wUwHbVTQ34
wSS/x2nq9erNXQdahMmBaoDS68h8UL2MqIwI22erbSuOeqSWgoBc1BgUBHsO+2zG
JJW0OcGNiZ1OxGuqVzjosfnIPvDsHoz3YqxgIED2OATbfhEeFJTbilbo+bhcKmf5
JKBmDFtly5ZdV1QVDOxu74prYB9JqI4L5lHcOtkOwPRoe4xoNs5M5RjuY5Y+agAQ
qXr+DfkEczvwtDHPoC5YC+SdkcA9QefaEuI0ZQLtEoMDt9ZQWy3rh04a16+mYl32
gyRN4Q8wP2PG1x83S9ve7pPKTR5BEwxQVsjuj+6jxHXPaJwuNGYEzV4W8hwjLJSa
mEVrCl/5vzC1/l1njH9+j0m3GpW31SSdWolWaAPWt3ppRSGZ/1FpuP+v1KsldoHc
c+JEDGA92bA4NQXF9b+2q2sMMPcRnTyl0O1QN/hqIf5u2LuGiZnXJ9fzl6/LskZC
fSHQkth0fPjTuXeYV0Y666t4iwjzPbXLW6/FKKHXohYN9rcK9oGPrGqHF1HhncrT
7dZxnqK8GHa0LbwsedD3sRw+daV/KpEZNMhRLzAUK1dpYSehRh5z6j5HVvgwVaY5
Z91RypYjsciDYph5ZSYWuipXElWVY7NDE6LBw6rO/i/LeV3vq0G6o8TfUvOEFjly
sxz1xq+fthRHxmduWkj7RrQkiKBPytq5Aw2wtZCWojxFvRLHPr9ufA5GS2YE7SfR
JCe/Ovgj1aAgSIroS6ZewhI+V+o9ufvCgVMh6qxs2sQUEWslM/OFMhgTbnROXQvO
McWwbJzuEIUAuA5Wds7INLRYE4Y1DqSgtd4Y12Wq5JgK4DZYi+J8Bo5BaMjDndta
xqRdBpGGpCNIoRCNF9aE7aoitmkfedyQRmQEGdAXxlMMMns5zL6uYfHvTrpQ2/E4
BCjfGIEL3/UqDEL8+glZChbDFzUTge/5d7nWK2M0klX/uo6ubTQx+TYJAdanmEOi
cL0j6N6h4NGD6qRN0sCrQRsbOkL0NBcrHzaJNQq1R8PQ0zVYB5YZ56aoi9x1JiIJ
RhVQmEo86wEYEYtSSgtg7pZxv2HjUs1uEPTvhxZ0uQL9ttatKoIR4zb0MK0EPZ0F
PDVsU/vB3decxI5T8WeeHv5KOD7pWKDEe651+FN8vcvf/U2r7jDdnx7xJLqvNuj0
xa7NxSxZQ9c8Rq6EEIOv6cwUq51w7ojewETWWPzfO4RCwDQ+mrQ6LogxsMJE7XEz
ZmT7rOY6SU4V3gRnFldWF8vsp1kQjzHZf26YrcF3SxzGAMZbTjtNU/ncDIVeZMOz
TPLBPNuiwobvyYLa4AqGPk7A2QDi2epgPu6ggYjV4DUj2x5NEvR3k28VOBii4tS8
A9cy1qnV2cORp11PFnNqbsfNHUFYt01T8VAP9QTgK8ry6NSJF9uWvBjgPyjRDjM8
set+Lz/UARymR+GXOQ4jg9AzZ7wUlxzLn3WvdzyxGRyG8myOHqs7JDzsoREWSxIC
6OyerA8im6ZnKsCqCd3kFcP2atA8Yg7eP26V6/vTYjZ3TmV0u9b2SM70c7IhGMZL
2bqK/c8H7yw/XBAom63i+pyKmp/hKLTgegKrmzfyrHTdBUek/SIYD7/ymHJZ9Som
I8fK94SdVini0VOMSsehuvYETb1+/U+17xsUEaHONKYhA+e1eQY5alvVIPhw2S4D
AftxpnuLzUt9n2mKy1ab8w3qj0FUkvKz0MDeIVzxmrsDbJt+owccsMJU6C5L9O/Y
uRxgkMZs5jw5zcS2Jy/p7k/SYu66YIKbE71wEGbeK3B62kKSExmiVg6L1nfyev1I
qYEYliRyDCfqa6deM2FqWozqyvKIM+ZgokQhDPo3K3CIGZsKlrpuVTCuidbauUf8
n0pSbo5LOQkFc6JoygIvLuwv+WthyD1akU8KsiaBiR3A/KCOksYuRXBaFmjYNUEo
nKb021w3Y5FZqhrH1ELrutLlBI3dzWoexscOLmjAUOEVcH7kBPIjEfAXUEgVEkib
TLb2g3x0sOkUEizX8aVn2e3gcPgoCX++heNu3LpI/WW0cbSOimQJquVwSVz4btNU
yTPYlGaxfb4f2hGsZfyKR7/1nXKgT9RgEojMX05MSO1uwgWpw3/rw6zeAIh2cay/
osyl6C+KCjFqmfo4wsQKS3Hx0JbBsfEvRFT60pKfsr+Nqy8JjhZodMreCl+cwJM8
MycZFhHWy7GK3H0DhH+CVADREDmIyWExKbTHtf6Kuz1M3mcZMkebUukua5/8y4Hp
Oo2QV5uVRRFROoeOzhnLyhJrB4tqGjrmOYFxXMIIHIxketjQbNFPqjSZXlSrpR3m
kseB8fi3jnoMAbXdxWxG1PGO5Dt9DPLtNatqqoE+YUDdtoLQxc0ntnsrU426bHSd
sQO2MmgMwFntCNmAOxcLbAVdFxV7zPxhtaFx9eq8gRic38xGUsiL8VwxuYaksO9F
xMmqVU7bTDclA/G/dZUxEt+6YgMFPucYrvvb/F5NXFjDHbiNlGCSINHgoL/4aa8x
oXj6FV+5D3tIci6cQaeBUwH4K2AsVwFuFvL2WNcJXa/1He0YTE2JMubB+2G9BqnU
ZfBHux0pgCM+biM7cioh5vhCAtnBQzhZS5afKDSY78dzGq8VeEPMImnJLx7qBoDp
qxP5OaIuNGOb7P7U8NL2pQ1tYmsLhScYg1XFNET4v3Rj4G75edLcvyzeHwy02q3Q
YoA1ddsi6jhiT28jyjK+Wopqu3YwZK/Gc3yg1qJ7WJFaEuYVUue8Ii8CtC1tDMUD
rJ8XrXMCYAwIAtLAfl2SEWXrqgxcdeQF4Ml+3pu6cMrrSBLbt/++BBL4upGGEp07
s4OugEo9P11qWGVJI+FJVQ2IKtGNLz1l/TXT3y2HHyBVtr+hY09kdN04ChrlEDXt
rOodeyH4uFug2t6mt8YV1y4PFGI+eDGjcC/Ryp9UFczMoYOm4p0ufZl0BxKsITcy
YSQEY/Rd0pSkBd4zmH5OM/FVoV5zTR1v1ct2tyViMnuAp4w7TU/VOnT99j6aWN09
giXyAvH1Xd2mvgGiuOm512HHcff1wX1rWUOiY1u/jqLq9jRyretrg2UUjT6kvIVW
g3LK4lDY5bwCIVwDp56kJF0jemIQzQ8FmInfG5JM7uQ0C6gTwCCR9AetIafzBuFX
SKb2Cvlrc2pMSCVgbs3exb4m6RMBUh+OhIIbrViwNXHc0jm1z9spegF/TQISIXEw
c/1wXaIQep705WopUHHxb6k6Is0le69iTaVEEZ2HVQqZ5SY+S42uZIqTbRpHoghp
iVp1FlFqFzlZBLTK9YYpoN6TbBw5tTOLcb3SLFNgWWS1mp+VW6Fri8LBbzwpqfGg
+6Hv4PmdxTPGe+PCbuE1kvQppi2yYKfN+6Q9J7FnqDAwKyvndKq7Vrl+9d3IOO6W
QmZS4BikcRdxblh/4upM6OplSxwkFuAdvjj94OrYgE3FtoEdVpeMBlY8W7/Qn52p
OBwzStvWzGSoL7x9Sp0D2mwxdZngyqPe3ezbuLQ78oM0v+Fc+MlG+k6TY6TtfNxL
lgN4WQwm4tdJbgdFHDcGcgkEZm9iTWP6rFGt8gbWBfHQj8l0K+vPlV0Wa9MDAUBj
AlY417IE3vfm9/fN70dXXRbzh8p1URjCi6kBr3fZpb7eNywadj0ESc5fZ7/hr8nh
gcLJxvQIiQ+1Rc1/eOdSbmwG47Drxwjz3FFbFhALaIfEE9zlJ8jUbQ48ZaOfQ/Nm
wPJeehqrIw4f96/aHtV+gBcmHN/buTlrOOuOgjJldB3Dq45RjhEAmuCXp881i88A
8Sy6m0x6kbmXZyxsAWzAyIFXRwOSygysmTwKdE+7cJJ34ukIKOB1tyecJJmvrPV+
yR8pkJWYaEy6I7bRomM3B3LPpUIpOg3IGve6jJiQjfq67nxBVPm6KbLXvBhOONL5
xBCQl4Yuxdf9lk6w8sEbbn8D70wCulTxdoBwI9dP4LkvJ3eUTKuHWANxpIHVJHNy
j6ggA3YGrimZ+8hrzPtKrlABGYSYPyjNZFkB4x338kFqqHDJU33PZLihtTcsD3oZ
Ko22raMC3bi61bOf4Jw92US2/GwBF8rThLauK89NU+vkE13gRyUsl9UvJlmXFvNz
OSgO2ZkDM66c9brNYx5gJdo5yOTOCkWPWDpkqgpux4RCxAF+5f6WFh3z9/2j/plB
nYqpcgbjerHfugxtMbvO0ZO5AEUAb3iT9499KuBhiMYJdNq6ccEF9tx6rQ6EAeJ5
aIBe/x5zma2QAVfSe1qw6LsYniPJ/caBUkVj2IwsGZrlewoGlA/5+uCtCzPxOqkG
5pVXChAq6tTt6a3lLmMcLUMTMHs8p+pvrocfkcOK3bQUOhL2MpryX+OfviJauv8A
MvQBTuwwcyhNTjcp/3NyPBe3f/PxEH+wqULKnlmx+9Qpl2URh5MnUSNz1Ygzza9E
1ThILNSA8pKZj31hxA0/JNSZdh5vCCeiH7vRnivwSgzcyA/U7ZvukSbWxwie5SZL
xLDmh+TqtzzXI5LbU33WX+r7IjuDwJZPUP8/89huVJF18fEtw2O6JYfsqjSN7IGE
Rem/gBbOnDaxC6gGW1R5Hr1/Py5JSQxXN6CbnCy0m13s5OMeA/8MEE3L1sPq/j9H
cV2eAr/gdAFfl1iAgY48K8gc2TDUk/rWjjzlwUgDY9vxzRlE4VBNFYyR2lnEMZOB
cG0vMQtqTLw35bIVYMIOixgKbQiA+AxDttcsGXPgrugItWs23DD42NA1Kr9I1sz4
8+NRd2f6tmqn7JdqbP3V/Q4owOLjJwu1qBT756oE9UcoYE8osbF8rfqeozouFhi+
XfY71LxEkBzsf3k6OkzolU6/Ah4+jPqTh20yktEYs9eamG60RJVfEbGN/klvM8KO
usM1CBZ+30wiDK3R3EV6oaBuncmcy+jZ/qYCujDXdySgqKgGPFojzDUZu1eQlkUi
J+GBQot3IHVrXHdEMkxd7P7PQrkjJJgXRFVFjNNUj+iUdfXbDUS3UNjytakyRKAE
ziF7szud9RwWfgT5SGUkUQXxB+/fCbSffkhnaeK0icE49tVRt+SeCfVWwu88usSr
B7cmU6LeytbNDfud252sVOYZTwPWU7e8BWBNaP5HXZl7QqfSyrYsmDnhVdxqAYJk
0Z4AUMbB7R6ybMIj6RF0GJSNQ/7ScvnonzT4nlX6kN4qIllThXP3fhDvI9MYR0EA
VPJ2ch4i+WeP7sgKlg9Imf7R2gaCuI0+o+PORZLra/4DbuYFxdZGLpiR+oY3Rn+4
4eYn5kq7rxoRpggN55qycAhHjzKctKGeOg2ZY+lucbjXaWI/enHGeqSOE/0s4Ox1
2dRXVUIOfJU8UXuwedIMYeVANYc0cS+3A7vDm1aWS1MRleqlq4winJo1n9uB6Jl7
j+bQwtyLK3FjFpVOmaqDcovk3coS9AdB/xP5n2A9bC7OJn/uP8Smf+UeCyWjQF99
PlcoQIkz/CCsIz+2KUg8XvZpUKQqbS5oFjk+xikdFKUgf4tsW+vmPsIrYK+FCf/G
TcAH9MfOJK8dqP+zXdipQhKfA4tEOTtO443gQFX4wwYuTiv4lIZKHkZmQUti687f
9VU6SXZR0fatsfZVe8KgMCGuFiAWqOCfN1FHEw0QOzTF3ZwGv9t7CAYD7Jx/E683
SCDq34JvCIdausqh58CRPLQ13zlXJ7HAE86QKMUmx35BF7d20nxwXgIkT2AI1zU/
WNY6aFT6HCPBOwXmyWA0RR/31917IsMMDLDa70HmMD/oG3ll3ZSSWdy3z2pSZ29Y
4w20Ci5QPPs0F7G/O/4B0YcmR/4HG/1Xw2hwhfHKN6QZd8OXQDZsRbYMOsBMalaN
Hv1jD2kVtA9dom8NPeTxTWEEn6RXf3dE8RCJeFyuTy1BsyxfHZlRHPmQY5UzIcSd
XwVGivIBZD9/fVrFNZSzl9ilaJsDw+Cj1jdQQiRnNu7rkIL/eHR1arVmv6lYkNZa
lr+p6z0m4cBNEynbV1dsI2UcakrOqUxfCX74o3wItO0KDRuaWQHhaw9MNjZ9DCmc
pkctytcjJXB3PqczRavgJjo0ZDWT4ryEwjiAj1uvUv7HyZGDlAQTLIKpsq8hWRIY
OouQriiEdBY2rNubNKjJd1sGgitHi2U6B4NTJX35rrS0ndKzxnNIuQ1W6dM/ec0l
6OTbVSy63Its/HjnfxJw6X1qihltKa4LapS+UgqFLDJnZo5Z+mnJn47AZo5ZK7Tp
SQQaRs+qvVB4EMVjg+P0ZzoRyMT/Ms3oQ9kkeghMIxTQHtlpGKvBOaIuHuQTVWee
TtxDaIuCdACKW+Ek2mlSlSdq+8ovb++RggmlU0QUmxyxQ+59zlNvLMlKqc776Zjs
aJAm+prVqy0a4bbWKoJZ1p8SSBLWfVfwwNkPB3kg8YqvZRwf+GnReuIxMSYl7lvY
1aYQIaRLZuCHOSvRlhU41QrTYfwAq2+x8wAPLZPSrY78DLAKW5eHWXMyQzONlW2d
rrDFjmBi9juyOoZ3j1uX2hLZTILBa2hvLIJ4Z82P5abTrg8jBm/rZugv1N3yvyMy
/7oyudB5zJAtQ6/43v8gvR/mKRRacjCj2EJalLfx3Rg5VPEQX9+wln33a7eSPFXt
k1NgrFd/MFdBoqMgRCYEzIdmRmSqwpwUUhY0gg6aPEsxWGaqM9xzF47p2MIA+bGL
TU8clwdhE+IVkbmcNBJzzF8dtek+HOO+Qe2+z5O2YbTaQ0yiIkk3d9ttj9PXfAEK
hymiK5gN38CiUCZQYZMgibWUYq6GOsWqru2oUMnhSVo+qfanHq5NL1BLTLODXBf9
sMtolkOcLjNlR/b8pmn/VbRi/j3Y/JHYYX73ilxGPtYYEkooD3STrHmC0nb3nh3o
0dX8iBqonT0CCTR/B50LpompFIuX2wy8p34lr0gtexrhAJn8hkZk7UkeoukfdOmC
RMhjlh1P00xAufxnXxbVBgFbn04Xq0iggXopwyBVpYjPPogFIhHWc7JHKak1lyjy
cd7y3fHdL1OVPfeiNBf6yDAaR2Ta6iQ5/M213PZp/6xwOJliT0DSqChUwwd4yRPt
alGnEmhGRm31PugIYiHyfqeyBSkK/jhDwz7/DlOtEVyJwpF1aV1ZzrkW5B9W4CDL
JncClR1jmnc59wHkXS3c2dgc0DcvvnGBPR+Ahc6RjNmDzlp5fJ3PBB6U0vTmYvch
RnoYbGAaS5U6kZ7CTiQV75b64rOx2al6hFwRx2KT0hKbJWgOztpbKQy5p0BjCAmY
QWffcPjermdKlzytkKoHKH9gt4cT2ZL8qJCGhMi/g42gL1aMglUrMKS5J2PdZ4nj
B9n7pxoDC7MqKZrMMG9uzwaBhwbEKNmsFAn49sgWT6+Pp7fhdTbcu7EbAq0s90Sk
BBld++QV8RKxzA4lE6bfb5wZS/mnrI7sW7rszWHAohVUr/iy7nV0H6HOWynQoWDh
RSNbRNRHIBrHxi1X5E+gM4liDZOl5F7p/64766Aa72nBXxESRY9zGl5SPoaKUkqw
siXU5y1y583BQCQ7Z3EPK/dBB+65VkcMP4IzXLCuvAXBnyomxrr1dCrncbQZScLg
IsUBk17O2C2n7wpScLlTY5zOcOG9Lu2XiiFRTfhelfnMswvb/OjxMf0zMglAtNS+
ZfvKDaNy+D+EyEkqETN8e5DsCxGd+wOmC3fGYcWvOrOD5urFjgjY9yV3ckK+0t2b
gRUphEcKr8Zvi0UoGHqV2b3H6q8Uo2ynhm1NtAmaokrmnn0+54DwRKG1zR8DhVSw
PtCYNHCiTBkPL3iKmfWyxyQ2ixYct2FB7qCEFuVkqiLzu1SMPDl2qs+IjYRHQcqB
J0aAmfrInruHH/3QxpLjMz+ql59eqgLWo6HMGkv/iZ70XuUL/pkXqovLus+DLdUJ
aC0tk7I19d4OuSyM2GTxvg6izmQv8PqINGFpKQzHpl46B6of/SbBKWaVx9sMU6AB
Qg0obuJzsCXekhkFH38jvMCMQqE1Zny8FSGoDeATxxybeV0GcF02SthrnTAXrrOG
Hi9ETfEehrKKU7PYSdAAdxs9HbaCwq61tU2l5B4wTsEWxBaxbjorRarroVGQcwTb
rPzaxowLYQmTyhKSji4W4Hm0hzINQoYYfY3xQ4IGnjHWpXMLFmdArg7GOs/TvOxl
IzFQ0DZXg1e7/roOTcNdojK2R9pKBj3IfFawGS0l6DhY78haARWOXiIRoR+8QoFZ
xtvEqRezMmdhWhS9Jx1FHWzWRWO+2bW+zM3oo1MZDNpjq7xKFFsn5yRkomvyBShe
APj2xnE/bDLbB9R6p8/aBXSv/u2bqZ6SEuy4og8AueslgMMQsbYuL8PUfy3Q9VlZ
SDAIJNV+EfjZC7l5eNY802ZfbfBUCHdLzKtpaJlFeJAYlVMtF/DksIkjRnSxV0Zh
GDOSlR2h5abP0xCzkIdrDZwWEpKO/FzJ3J/psjg2RNYlFCyS1ykn/xE2hpuLy/nx
bVpyUQqNiOBTA4yNOvL/NTJGQ3yH8AJpKNiV+M/iYZAo0NFDAezkFIBlb5N1N4Ng
F8qlTbm8pXLpD2FWseDdOGUUzDXf3Jm+X/VQKxeyIYxnWc9u9kgT1txZmhNRB5Pt
ztcBsW9jrl1KM/pOx6mM0FBmb4E0PzQM1lyKvMeGI22gZxNN+VhemXcJ77VKamIe
CVo19QgTi85UFjqTLcPPcw+iBRGgAu3sExDZJKsr6dbZsAW+9Ov586VigwUxtHa9
E2XAvAO4Tzn1MzHevYVuGAalhwgI6nBaqY2WXzGk9xrt4fmChz1tM9y9EW9iNjaE
C1f50QO5TU/Z4yNbKolW6CA2q9+aYLToEI6cM67RVug5ZluDilOXuT+4RVHqnZVO
lmy/HRcmQClMjdDEANfOj1OmHLP6rQ6z0f9T1ewt5vRlPsGa7llr8G/SS4Bo5xIn
Xg7QC2KXB19Ph6EWpPp6zyMrn/E+gOCM0Y/UsMatGJiNv1P+u2w+RF3wCI3zKhGY
BPjMD8ActlwN15a+QWXPIZdxrN6O3YedqaZ7HVvSA2sN/A1sW27roc/3z8G7MeXS
hgSSoXwkRVmciIqwKyHM0QIDU9Apq7d/VqvHPNen1XUaZhEnnQWN3Qeoat8QL6QS
bWjmnJPaB9O4vo+ONg4FlukyYQRbu191fBuQGRzwgXkoK4S/yHwdG4l7y/1239qf
Hox7mOxNlHn/M8Rl8Tt1pGaAPJzsHGuoijRm26RYsO0OUi1t43sEHYuE3qJmFdru
iJOscXxcC4JDplGP1gFnTzlEHaynv9zPSRaYI0rC+G8XKzE1UrKttK2X6nm3TZYD
Sw75z8nh/5kLUL09MMdXqMt5div813bAIoczt6Wdzb3AugKY4TCdj1pCzBQjm6kk
VZZzk3NFKXUHVIwFTNNGcB/4LbbH2BtAEpT+s1Ttp0WHodAXvMDVre1yPGm0orrU
sGuc8P+Bw72FixnZ9DmqGdSOnkWStfakqKZy/X49Ecvu+hO+14ZjkML5wEURvNqQ
V5eCAwi9RhF09QUp6lN5konLIHPFGedPmNDJ0E+bKJod3hIT3NDrC1APS+G3GcsP
SRiGKB9aCedoj6BJlIbP8whvRoLjff9k0CY9wDDEAezqESPLRXJ7QcT4Ta9cmQ+Q
Kds48jxY906Osgq1sfuSEW7vO/ZgJtN0mzqDwL1cKbvx5KgCejnMK5FmForlhd8F
RXAMNFPoh1FPFFL6cb0B7mNfcxkuTlbdnycNsxESC68V9MORTVxy1VqCGyLexUt6
WA/9QGbvQ1pmwjOXymhCTQlFLQTCC/pTnFu6sB7Pnakq6rSPUTm9t545zh1HpU53
I6DK9lb5/xPzQUTiY7dLW8A8MgFXAzAry4fm2xrtM9ZEGYI3UDTpSInkXFA7eFsl
fv22/kv3yekHU4/2ECRiAxBKJrxlBtmM5K5w/Oboa2HNvZKejBPc7Co7qQu3GSEk
+LQxr5yJfUjz9TG7S2zKqDie3Ls1i8fjeNDqdDiO9h8yO1lcoQgyy+LvYwCcPktG
WMWcTCBi+AKTA8yUtZT0KvNV9s2YSrd88fkOkMTknUh3mOufW+LbysV6RimQSu66
GnnUS3xVrOUJNJ0Q40qYd09peOJ59Tgm2kFK6cXvIR8QuZrL9uXkSLpgrjAeF/8y
xNm4qDZnFnrdJUsMtgKV/IaDdHz/CJJkPj5a9MPNoT5jSeAzL9F6NoQ3lW47pafq
j7M7D1AlT6m9KzoYrz6KOoBMQeJ0WjtmUakPaD0GW3lrq187KW97UEZdZyTyvWGF
2kRs9RodWcKXoaAkektf3r5AUZBpF3V/OgBVhfSoILGA4F+0gLXtefLmNjoUpnEK
bjbnakeQVj2IDfn6TBDMzlK/cgLOHZJGWVyw3Qg5xt0lVip4YPb/LZEJfRhovXBi
ij/BZuP/NM+d9lHgJf6PmCw/6bMy3JBO5CrOyFrUm0jiW93w/LXivJm8CoUNiIIp
yjoKnfRFtL/5OvEruHcJ8Gt5i9j9Kh4u6CcBaNRsC57dahnfNBsv2vgYa2gczLME
LuGPH8XNOr7qxZ+Ej0apYOtURuUHqhtXrF+rftVeRROuNfkSwEqc9loUmti5UjW2
yVuv9H58GCVxXfrzCIUr4pU3X1dmtXPDgil4a9rRp3PmWG0L1BD+51kcGlLrxtMv
/t+LJClCsUGgw0YfI4KPu17+7w//ZtMxNCeFCTalCPSQgtcMOA23/9ACyO+HSNPA
rLJrY9vDS0aUmSh2PX0YcYzCZkhRbbHvAdAlPBVe0M6zrE8+MRpquDWJe/VnR+OS
EezTbAxGu4DIzbxFo8MR/olWCm2//JT9MoXbxZEhvhKp1HEikPowvr8cKeXwnQHf
6/A2/tg/rE/j54Aw5FS9xf4qUxyxDUUjWNI5dk/ysXBIvuClIlxC7vWHu8+DvFOj
Tg9PdTZUXaiwcKI8iGneqgXb7cShzKcQ/ZqBLTqrIAo+Yc0rNAodw0JSFw3pkspj
yDF5O++hhb3jh3wUPrEMcwF/c8pIr0+PykBVQ1OTdQn1FAl3ijCSr+V8yo8vbY6+
0v9b31Lylhftk4+63XoIV349FJO4zJAArMQ/f8e9WHQOyR+JqthXpmp1AAGEN05z
CaHJUL4R+hZrf5DNIRsSKVCqJ6oQI8NfZlUZ+HMEHdzue+pE32SsjJcDqnBGBC6e
nS9DXE8eUqnvqQOTeKUlqZyV/yjPIo70B9/Q12quZrFpgtv8WBWbxStmSyvgZ/jx
4IaL6XWdr4aRXhdfOdiV2wYYv20RAHqrDoAGp8Ky3W8hGURzRS2ybYAmHryS6oz4
p9pBnBhhYpi83nah08H4z47BWsCF4U4QSUoXV2gTd1uiHUNUsbeHgBxmouoNpIOb
8RvbzIuworSUfgVNbuPs8vkfgXgXixs4b3e7Q8ArjGjd5/AKGDQdVMN1f/uu8P3a
h1Uwuo4yCSeuZTBFqFpJDKEAmPMaKWjGaU4O8kVRMGeNY5rSzfU9BxszfaVQZxdJ
xqi+Z4t4dKTeJr37gwvkkAHOne7HD9lVlqWpuI7mOBZaiKqSL7oNLfjUnvEptyde
n+06GGbtR2SdgepM82xVQqQtZGcY6XGHDjsdbRlVdLg0l8JCJZ10ekQXnkQMnR+j
iv/CUEdLaBA7DYr3mk+8cHtuDNGznKsrL+r5S+eLPTUIGgkYdf3/+pqg8NsbhtEq
ZCMBaiyRIBJlzNSGq8+B34saLQzOTZ+2bsOjg/lTZg5OBGrUlB6iKQgLQW8KDp2R
N8RVHYtUKdcs5DZqSng15uARaHKIlVthgyTFm5EJREstac05Zcbi4kwvfQV68WR2
KKOrXcsJDcBOQQXadcS5LWE7WzsX57qfu0aAuTy+uObeJWf0oIxRAyGPF1Q+o9Jf
CHcU+saoZYTYtoiz4ahDTPYOPfz9BG0CpWTW5hchVXxsXyw7icXMX5eKV89j5jgi
hmD3NCz0JD0DkZmD/elo4FsdzdaD+MAwzXhPnBh7TsNacUUTUDqUigYkpwxWJ36c
m85WQjCj2x7NvDG98HxCxO2XezaceRuGNC0zRsC+IFLT1R/Z8AU28ABfeSkH7D1j
X+us5YOdQN8tFHPqihbhfOgenBgGcMWdfiywwsVe+zU6XncXfjdHljhJeOT6Wzv/
QRqL6IZ8zKTbDl/l/WcSBpRB+tz+Y8jWAAWPD8P1VcAPcVnHCgHgKBqwnryMu99J
b51xIoCB+dXxx3rBYFUrNRlYMev06Od6ifUBSt3YCpydq/BrD2s/88Jg9di9/DlN
fByYJ597mhZs9UQZI+KcR6RWuYEIsB7cpay8J0sGxwcKsIm+LMR/FlbOIzqig5YG
AqJ4lVgma9i6q3ugp9I2A1yK0bANnXEAKPxTLMdxGTznnEiyezv5dNGNP9Svu6Z9
rlNtjFRA/wIlq0MqSarQnLU6JwpLlaBgScSIiaTU+45dYABZoTiO47HVf/jSMkA5
0eQl0PH/SnWZckD4G+W3PmM6EhpzRLQBNasr/WkaXikaZChSYj6JLjysssXil/SA
s3rH16CsgkeRDr0PXaiRNuva/9grY8D48f9NyRyG7Suq0KJLrkA3fY2X2Fnxtt7B
o2R4sKUpCkNpgXBFXNNzMpS4T2o++LbgF1vuTSWswjSCLiDzqKO7ZdmuRkcWQqbL
kvylawUlUQnyswrky2sb+T+QJOhQV0XO8ZNu++b5qj1UFaUj+I8BDrkmNsnCwtfA
XmpaYdCPbZ7HnytMLCETms4M1s4MkS1KgzbWzKDJYyGi7Lh2g/oqLq1WXsIghFnK
D+WFMWijHOw0261ONzHEb1eYwWOIxW8m0hQlklDtWjzZhPJ9Ag3StufzXXUXpDFD
CZb321Tfu7JMs9fHUC1BsbRlab/G034yW+YI0uul0DuyeoezH7tGBvoS0855BMl4
1ShLBkeLrqUpNDn0bCdH48Sln8spGd5OxYIKMlQ5+WO9aF76MNUZMsw7TnsjflXN
zkdxB+Dl2xm52BgUYQnEwH5bz1iHKrkqaw/ZL8439p/2M14DeLLpJZ83fLuvlXli
mPSD31MOh1N6XAljZtLjflUILcngJBraIG/dnDaLZA6h1rX0DnDMu4zklmEjzdkT
dynpWvtrdMiJzrDhlshvOwyCI0aLg1x3OtGxm3kHDstNtMLg+VPDX9ocuPquIHGQ
VK2CnyiJr3tHwZscCODFp1AlVoYzAyG+qmlnj2N3G622xCsDpbhSTagsKmnKkauY
G1VTKaEl/wHCcwajLINDRMeO1KY34XR1yzZfBoAvY3tdp3HHdPK9CoWedRgTmGT5
Wd78kuSQkUVy3hp1nj8m4R/G6Qlo0DgqxXduKMr1yf8ohucYzDer4aWsZ5vOXrt4
fYu0eDNZN+Up1MZMFj4YFbRdmvnOJ9a0OGgbT1w8YjL1B71k1pg2+AkyQpu4F1Bh
4hsEeqI5Usdu/U+BhbiznfbaM/XnWjcS8LCHhkAq0M8OAh2Bcwf6usuquaijnT6M
ri16zSqoiIVuw7CLnHHaaHuId84vxjkJbHNYD0W50CUZLhWIz2yrI685oxTyuFO0
4GavQIOAyGQD4p9WGQ3gS4pVd0VQ1vXFlShafg9anK7+vpiCW9mM2ldi9M5lAj5Z
4VScYx2L4DooE+mHpCDYELl88Lm5PhRs3ujwJw4JJvkY0pDj7f/kDGIYk8Xv+muj
H8oOLG7yairCutIkkrv+rnjPXGIRNlS2D/a3vZof38NbVFMxXBTFbDPI8hxpMm3b
gq2NKZLfLaYZbIE2EjWh0cEtqw/vSMHTBgWXnl5ZJxpiYh9a3aba+GrxwVNWRgnU
WhTrO6sytGodqDkHKxvtur0/b4RBb9OIzALaKFdy3s0SO4N4nsCpt50nbN3ZRL3j
XLtwo6zbenKVMX38/e9pnLW6CRFVb1R2VjxiMjLV42vzUds/3UKrqyVJHk15DpFw
cOEYtvZOmcDcsg4BNELkfg7teGp0/rm3MW29eLTMMj8I4iQ+t63rUAnSKeqXjU2f
K9WtKCXZY0KNHMXBLCm6SUt1zVGZSGa7DwnaGr3k+sRl9U56hlmy900rFcjvK0Yh
2gyDc3F3c4vRShTxxZdGYCsP+2w/O7GgBFxa8UT0foH5axftnPxWuJDZHIhCV0ou
9UFoCJkRJelkyXyxs3riucxc2JgR1ASt+A/rGPueTxeBnwLHs0MX8M30zKUqE0ZC
Is9Cm2Ql/hXK7AA3/YKZgBq6T0bGuSzJymxPWatE1KcpyOZQRTlMW30owmXcQMxg
L753lRRRMHMupetSvTKcr8j6778KEzvUy9DBruq9lM+Ok+P0DaPw/xMXqCngQgnX
UkSeKHL33tBTKEpgcVazY4hlqCYQEb0vPzpPF+Jf1YKjGs1GNBdyf/BZrMG7ajnw
0a6abIsdul0PAPK5b4VGLtE1cH0G7/XbM72WiONLQe0Xz+ezESrfj39MvzRUP5UF
EGszi7jFnOPY9UEyoWpHFQZoWZ5pk9sY63/iMVp+SY6MretvoMDZlZ9hko14Ot6R
nm3VAtYl/3ftV+hFB9pGhZq0fY1VdREPRvGyzobN1AjQojEz84Oq7jmWbnitvPun
5GUPt3uAU4ZUY4Vo6FwHP/urw11RIRkEGUIw3biKiKbkO4/dqV3h/zfZvlT7bG+y
G6SHlpJXN09/0PqrIxaPRV1uVQ66J2jmfMmZHVrFitUf/ERlHlWE9blO274f5BsO
SCqBvS5RoXALwcYt8Rag+Q1OYXRSYGc+MpKKaau0aUd4r/7Zqu7aNqY3vUW5sMq7
gVBUMO+yQ40nMcIkjjLIaLFpfgqm6sirAaDXX8u3uiLnQaFEaV3gNeU0mHQ/dB/t
XARXbYpqGCYBStXmqmQAWR7SoFMdhTeC+SSfW1p6bWZ0YASDlvuveeJ5fq7StYLT
krGJAdy0W0HiuD/bOjdsdExihv5xCHhlIcxEiUQf3fqxEY6jkfvy7/VHBt0nJ0lS
JxW7ihWCSWCdfnZnuHTR4yiFhfOk/1v2AdsGiNt1ZlPoY68zRQcvk49rfA1OC7pu
Zq8kEV69XOBYDNuGhjFA6qw04lhhCboTy00GWIbYr0DfxN0Q20wGj2TPtOxenAOq
0MrP00xNC6dsG0xOUfZHkhXpgNN+f84q7OPprEduTjCqYlc+WbMuKih4+T6GRArL
uH8yW8Oob2hp8V5Fi92UQ380MpCP7kasdiu9Jl/8OrjeErHprHcld6AmArje5NU/
lnAyUiTpZzzpNyMzzDQrXgFbbyTGBNjrVeFijKaep6g6peEZHZTm701LupH5l9sS
y2nR853gHsjjr6s0PTOP+dLJCfWMFMI+CR4n7tYI4X/5LVBUhwYRucN4cjvPArGv
Gt9I3EYK0q/UJ+riKsUwPgBdrsRcD3/NgVzW4s1OKWje277J6YIXf5aoswH13ocd
qZtvQU/DT7Qo5Ln3MJo08ZUAYdh438iWnj57apoBvJ+8nrUUen8Lozcp8eJm+Qf5
iC7iTwX1cm34MqeywzkyoEhkAJWmqN8bUjUcOV1Gv8EYUkLgn/O5s8sfkFV/8bkS
Ffok6rdWJNvzNoZv8hgb1kroswb6g0il7ajYTB/5u7WL05LmZmWngNl4dlD6lzXK
oq/XgqcrWUYeJ5OMtOigfWpa9+gYpooPSgEc/0P4hm618sDgipXLp6CEcQqG+m/p
Npvu5fbwXlPZ1lBslpd4P2Sqjjf0G0FArCWH7EDSndlRODvdUtOjtE6A5AofD4JC
XirqkOQQciov7hCSCkb3QH7TwEpsp+FDKRnt8hGhVBKWw9aMrFcC4tfy7uAUSIYL
nILTqZSK28mUN2HLr9iRv2F33wKDLWD62QLuXiT1PmJYEktZPRg+cQESzp9B5264
H6KY/211pVAOMsmeaxYHewiIbDRku2J80SpBKHUUH5ZS/eZJmUlmFVfKiCmfrwqD
P7slDKtNI9flHQJLHlYsDRO7sgkXpjyKpM6YE5yIvtusO1n3Gnz2ypr57t/BN956
lrDPcnRZNoHuf1yCEHsnyTvSCmVBdXNs9eZ0XWJEl4ApP1pYO1LVi1e8o+ZfZRmH
vHgxRrpiqW5mf+f3AmUkdjymSt7bQKWs+TPeTuDyIckKkwnNqLCFJwEJc+Dbl5ka
y8zAbB/41A+zjT8NsQYMwInWOgmwx7ziZ3huqM55VhHePcCvfr7JIhaw4nMFEHAy
/AUAo26sWtSf26/tXLmXK+uFBdJcQYm7AnN2poccRTxjwUC4B7scgCEb1ldAQg38
9oMHOY6duiMN+QuJQe6PA//45G+JDbL7Ot4QIVzAsgHaR9m2nH4FSEhjOVkC3sAd
UL5FjHg2EGaRNLHts4y4H2NOPE9VxLtzxfA3IItDFpQrX/Auowa5B2D+YYAX8d3W
90nRvnWYfZYpOTWyxexffaAtpcQbwcVxfXPIyoOdOMV0pttPhWT2DqqFPo8cYhL2
Xk1oi7ij2vJlLeVW/HYtaGrsWG8VZWpqywdqmuRrM2qtTHjfkiimk8BZK7Gn15OE
LuhI/lFn8F5ij3J0ZQNKd/LLlXcR49Tz1Hl4HEzm7VWz+oqz1xpDYXc0D+RRm4NP
+mjE64fEtZbaWqsGSuazq7hUG0W15mpSgMG92s5f01jOqVtj9ma8g7cJKr57ycUH
+jNsxy5AbznOPkO5cU2iA8q2GbNiSsi20eEvX9oRXABDA09Wand9wHQkwbw1iu4W
TKa4Fvlyn0xJgR/Dd/k3cq6cki9sXnYPy7eTAuN0RY2FM6LXWpRme2Rxe4Naarkn
SsxNge0jjfLy87YkboPa5i+vkTDD80GXkTjew1H5ZEIfotZ6in8Cuhwm9/xFfGqS
bSWGi0NjsGuwUZdc7e3HBuTGaa1DV9B5az2xdkMLUk9fUwFQJamHraBktgoo2RsB
qM3Z+qQfeaarpLmVEZGbID4UcFfiNJ3wFWIeaUjHlGc7qKcJssxqlVm2ajZ+p+z0
1iZcT7wyC/CbIo1YoqkV9tozrb+FiTbSxTbq2op8JyccrT5nwkQImtSUzOLhk1b4
PDkSNIKBb0Yc4zsgHTDkuQjdEtBbOa/b7AJ6cKa0WJ1yN0e3NoOzRHauAsr/WuFE
8DDEX6p9hpOogUgB8WEWfbNybKW4hh1iy9/zuYOWQTFrmO3e6RFXxceGgIZUT1Pe
YCirHeSdt2Q6uSUhrOg7vYtG+9te/ho42U2Y2Z3+Im3aEV6Bs/J37Dm0aLvp/5lZ
dpHggBv4/h895BqikyYyRkcXeLz0oAU7M0nb+0G6Phdu8YS18EPUZ28LHpya8m3Q
USGjopWe+cSpYunhFk5TIFV5H471LqattapE0q9icBBXGc2tPQ0i1QHRTYH0Tl9b
LaaCORDKzdtyTs2V8GNgtdmGMX+WqgJNXQnWdj0iNaORqouKlfRFgQR883La2onv
1oa1vEDo94QVihXxbyJiQ9aeIFKeA5iP2FG4WtJtFYZk4S73+z+MiIu9wt8KAJJ5
TWBC98YMStylb8suqKbbEWE4xn+tMCHVgbFjyLZAo2Id7xTOq8D9pJmdcV3uEXoG
O7qwkw/CFTPPRJVcu+PcJMsdVw+WyLww+emq0Ltp18EdLVB7qalm71pmiSWBONuc
hKEFIhPoMNp9MXuD2Sd09L809LqKsets6T7n+GNvUOxSLMSUdKIRDj6qV91VoXyo
Mz7NVwW28JUVMTb9SKW4WkRHG+MCN6D1kTDHWrpz492wHJC/0Dfv2+PD5csLa1zC
ayViPPiMLsfCZr0x0Hgd/D/X9R/1KmTdugRRUbbbYsKg7Nr0/0NlY6vcfJzorWFr
ko9OHPw1T5XncbjyHEiKJVxB2VlZAmFnhQQmbrfF0FMDcXE8cA/jyg+Ei67afqxp
tjMfBUQx17no6OiajVTldOVfOO7Gws5UPku3iINHMN9dO2S3yf9+AkKeSjBFGjmY
zGzfktqklIkVtsm+rXILNorNkppDAwDOueG+bhg7X70s3xos/L+swPKI3rz8fZKD
IEMNWDwYMe67nwme7JtqUfXmLpY9JPNUOPXdDYt76bo8CZimVfrPhDKdgkSgOPwc
pLuNm4dws7WzG2hr09RgGciYXSiF4y3TLtbUk1UHOtHwdftHzuMkVwhZh0C7ZOvO
6k3YauP4wvTRWPNK7IFJaeq11HCmy6NWOPFt87Ijt9gXZyKz6RRQ2VBTucF4Q2U+
01y6K2fhvT2iYansMczREpQ8HeAGZteka2U5IRJ1qg2ui/lW19Cg4sa36JEUCzZT
43z3GWPqhWa1VeDM3ZANGKJjV0AhQsnxVQ86G83oynk2cY4MFaOhlTf3XVsRCY08
+9FY2oknbU8KEloKzxIWxsoJbp8oSDrmnV9oIlXyRH8wZEoGGEEiryTsIhZ0YEMO
eFEqcxW+pt3vIHkhVAcZ3p53y0hYAPoLI3zkspr+3s2FukvEdmL0aXow4Zj7StSv
ZhB8PmWNOMi7kzlohfbtKBUMTGgQGMCbHtgZYgZ9RZ1CDgMS+oWpA/4qp7J+of2B
Lzc6Izt6fKgzIiH13eo6WyPLOwX1y/pR15XDGiM0gw9pDX23zp9yiY6N5ueEg5pE
cDjAq5DK1qVJneH28A4cxO5Q9h/bkuRUzKgOR6Y9ELGLanhBZv3ADix6bXDxiLXt
ZbxP7aaz9PiFqiYRoctqv29wg/Y14k5yTVOsptzBxjCb17FECUpO6acygKbrbOy/
9ZajQnRu7PWTyMVxrcYyihFwd2g+g+ssi1m+SvkMWcQVlf+Q5O+ylyGGG4HXt4Sg
z5yyzle/pz0H8NtGgbwnZh+YJKubjlM2TKdHzmpegdZeOwWx7WbBZEKixqnjwqHl
OiDrD6UL/rVrrC1m8xuXsp80jPuDzxbjPKBrVG/up0sDQIe0ICAn5PmmcVANwKas
/MxtGxGC2Prc1ZRL3e194OPp76qyCV+IIbSWdIr34195ldMr9r0x3Bx9zkzXlukT
uy16e5zKkGw5OLRgXekCDx3HzL8egatXLDYP8JDowJa04wDvH+Vz7rR+fuRpliJ4
ZKSwJB62iSZDv/AQNLvkGIoIguFluwJ0w6nsFEs+qNlzfg9j/RZ8kxFNcD+Urmuq
B4GSxyRnbu3adQkFX0zNMXbh5owexhp7Mln+g5l3RIGP8WnnFTa5IKDPMX9VLbYd
LCdJCWQrw4uwMLn9OHDnO/fCSL8aPAZLVbSBVGSo/iyC3IrvJ2gE/RBwNOerRhs+
KX1uZhbUTvJhJE5Q9tQBP6i13Hy+Z6R3l3gWjZzNlmGH56whLXFfdC3lBlZi7c0x
nW1mHQrGSqWPAEAgXBxAiMNGjeCZvyGAorYC/FyHBmx41gzFTpO0ZLSVU7xG6K3i
CZ913nHnmCKBvD9mjKWr5IgvYtkOyBSOu9JAu9Em9u1yDdzfN9W2KpaF7oOkuX2m
XubVXmYx5965PswOisVCYtFGBCQygBbCZaMxpxn5tjrOKDq8OguGtGRBx0N0iYHT
S2ooCG83+AAy6vGVYXpODGdv8/sscADmF/g7Dd53Rk02dYmyxLCM4leVMsvK5N6k
LHFSG+QpynF1pr5Wh206YFbOdTTuC/lg0R0ReIRki07qmKBZaCbXDt6jeHBH1sNT
H7d7KvtJ3iUdevMa13xkENYIZbS2GzuYoEi4VPoFbJmwMz5vAViNRMhKWeIhlIcn
0wR3x3bSSFggciNQITe6neL0q2PBmCa6nTYBO+HVdj3B/urSwBdyPdb45wICc6Ja
9xYv/OSzx7OyOcej5Ytlo0M2wgkTE5Hk4yOplD2URx95GF9OLVU+mIQ+FAkAyp/B
87VdqX9IeNfbVWD2HFsYeheL+pDqEwBXVgjPzIAh+AVMWNdIG4gkJ8B9AxI8j2yZ
BnitY2r6DhfHW3Nm3OgfbJQ5rLtJHrm5j7oJ2J08X79v5bHgC6Bk3V+3isFJ0ROM
nheOg8PrwGOhP3QLJQ3OFNL4WegGFYetRoNPaXi1kuITVZ9L3sJLno3rzugeTxLs
hy+aiNDG/QtknRIgDMG/w83WZ4NdiXyLoHFQbPViGIwdD1bR/EGbqCFHI1DsWWMy
faquhoRoTPhxbcd2RpQvpOPvhfYSr7kGWHyi/O0uAaehlnrusQW9pnNyB3zP0bhZ
T1xqodzp26U9NKyFZLVV3XZ5odV+Ur6rFnn6k3HFviGxzKnxH7lFkhcULS3GFYpN
j7KqKrdP+g7O+SHTFrvMQX1sX3R1akH21G/LsVe84sjCXLyfpzOjGg1THnxFsuk9
ouz8Ogq72ITqyivY0Uo6ILx0LO34C1Lz+wHdCLUxo0XtVpXDjtDaOt2/NO/mtPQv
J5xbSk02bKKgIOrCDL4FvzO2Dksg116+xipJqWwrODeMo3LDy3rZOqzs2TLQTUkO
my6jQ3kmRjWPhOUXb2lg9mBsMfvkUFgdCA8ah00IjJW17G2yYfkeB1vAjTkeQLjY
n3dxletS/7iddogGiu/79O+4ZWEa51mAhMMdx1V6EoWBc9sf7206eWSJxcxGXCMZ
kj4dhH86nElka+6oJfIQIN/6skIXUoCve5k7s1VA/kFAFgbg4xrhiklEPHnysKkY
HczHA6NRo7+tsP4ZEjE3dLwd9rKsxWlbcvV7GpFht1X+9EROurGa7h+2wJ+r2xJn
1ynKj4uZM6OcRyXpviC8SCjAAcbV4Vg6DlTa230thVOQnRWFuKzjfL7EAIRx/PpX
xHcASiuYRu9Hjv6HXlCxXQeONbIcXp38JiDn4OIYBa//YPtU5fJiBKdGLHBmWUaD
m29I8ho6sVbHadFrXNclZbQeGOP7hg7YyuyYQHj65vM1iAxarLpKHrUBQ5K8xWjw
WbvK6G3L979YIEui96SygKbHV/olbJWVpFqp052d9EZ4HMdjjHMir8zi4D/AoWNV
mFj6epdmfh8dEVZOPJLw2T8trlQCs4/yLawTMpLXXNNiQVmLbmns96AMhuJ4rOpZ
CDZjlfF+cLu8Oa/kVtMWkbX8qnxzJkO960cjMQEo/ut4Rad8xHav4Ul6Ewi5Pb/e
jhByd6/EPnwe/iGZoZt2aNdjCsvy8NRX7sJ0pMFwT5QnWq/IaS/LvIxVKFuxBvIa
eIroHzCh5oxXq1ogRky2TuKCNrh79A2nn7Fj4u0YQ22OR7HwaSnXguYGs5wcR2ii
iYiWGmz5GTNp7uyQgWYKfajwGU6r8gIkSa9nsRwahYN1bbzpn4ORrBa6sZRQa55F
K9n5//AU9vAWms3bY0wmEnZgHekWQ/2uQfZW8DrIV699VQWvHt7YXRM2wUsJsdx1
M4hjf6rS5u/++KJUG5kYVJ4s6NECdjb0PeiQ8mlWdZTJ2NXqQiOAaOu9PfuEeqbA
q8QajB00ZC7itDkfZiHXCHAW7q5YcQHSXSBz1e3JelYLG9iAnL6RDJHfnOHKH+s0
tF3hYbGWxZnqxJ/tN/o913TN3Ew3UTY+qw0n+Ddg55Md2gnZpr0jGpNr1reZfOT6
iIvKxG7ak35csyAd/H53bnp5hPajVORaC8/JkSrR6B8hQ9ENuyW1yiYJlMNy3Ob1
Za5ihV50/lEf/h2b8nWOd1IoFYJamaIWF69Vt7ZLHQx2BkOkCuZoAtG6Dw8ykBYN
LOB8ONZn6UOMK1pDJ//QYtFDjVk6mzbJdaVzPyaP0AmZ0HcaZLy2RNjkthEMdO3P
TlxR4w1K2BYROE16ccH0pdKCnTSk9klJtuQzxmUlw3za6s7HW2K2JepoNYonEp2L
Rmr7/Eef3QfMszZX5dalVzc2XEYHd/403zZbyE8AUkHh9ZIhoLYsv4KdpKPg/ch8
clmRLmap1UKlglP4QFSr7NexYtw5H9sfN9MfjZD7KWKTTllJCB/2c1QYmpfvgCIw
Psu+G7FzHXxitjM0MxcONpea0aBYyYY4aKuB6BmjOhk=
`pragma protect end_protected
