// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:56 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kK9dCLdKq8PKySotOC9t0iwfR8fJslTQhCYfL2IDk44ebOJrQjCCXRWUNtIKIAxv
aYWN4j5fBnjaSEddIpqHYEDJWCo+W+jB3lwpSC1+0xWopJGV/9yLTPPHdYR5BSyx
gRlXpFwH6WADsO1YRgRpELlHV3sXCgp5E3L1LMflMjQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8608)
76/09GFew6eoT82pT0l4UR0lnd0Rnt8TZHikM652A1pIdeyN+wpYHkzlzeGvsSgJ
7IN5rMXIEp+D0zKWznNCBBXzHTEaQ/DP7Y++vtcUVSe3yI1hAmmVmv5VHJ8omjSI
Kef9hNaEL6UyKNTbB2Y6K+fQD/RltJ16OVPf22u+26Z7WQspXDE7S77gmGtn/oHh
1I7+r9bfv+xAJ/vPftw3ir0x6MBW2OnhQKhuEsJmP3muW3Po8x+C2gFGzrpPHKbi
k1G6njlbBqdArQJDRKhXyGY5JeVYoa82q4DB/6N4uQn8DEq+F3Dpgn4ufb/4EcqD
YxOLcsKBQtYj2B3FNMGj6oNFwVsCQyJxP80z/iha5VG3++ptPZ4TrKOfHVOIsuSC
stDu04z7Tu1Ba0DNhhI1T1/StHQpLg3bfUoEC3Elmnf3qm+2QDPAMHLuHf8siMdo
41eqmSE6ZB3NIEpbX8VBqU/rm/L4zCO+/pKS3iwHLqVKs08lQQUrrSL/vKof8YEh
Abozc3IWpVkjp5mzfd/AQTKv9k2Lppwu4AHy1myCDOaOQPI3q4bGwzssfLbA/ngS
Mmg6BVciZXsJSu8+oLLkErQtRs1XFx3NuduDM4+NHb15noievW6bRYryJpbfA3hL
ydvKb72uRw7FwQ26TETXbyxX7zcxVGhnyC8gO9jebO2GEHbq58TF/KlQ7mwzpFKK
ojzIlNqolQCSwxAqJ13FcKyeyBA2DJDRp7fjqWccXA5V2mtUOyXKWzGpXhvth4WS
3iVaeSyPWRl1B0UTwAYl24H0wn1+nQpqjmBK7FeS9IfuFSg4SfVaOKtnicpyIsLN
fZc0szAY7aYzEHywc1LB6lZr+k1uUoYQbzGFFjpad4ZVjsmu+cwCwMir5J6LXMLL
WMAgfElIM6Zz8UpqGPYs2Fna5LsENobTrGR/dqJtK55KJnQdvAFI1aOX+UQrk71Q
mVv+uY+G+irP8VJa8lV8s25zXUf4EHFa0kfFl+ElXOA44OitBu73CnLTTctLfiT9
3ZsB7dve1zeeHKCtqMkUSJA6U1LYqz5a4x7cf+Azb7VvDlLPVx201yH6QxBk0yJq
nEj/qKOx2xKsG/mPOW0e14fNr7FXtlgCBUnqKdPe5TpCKVNo6jNgPAX4g6lvKNZG
zFY0SBqgcyfCAdv9MyJickwhn38BitZse1mQ60r/csqeb1Q/3Q3E/Y+m4yUfJuMa
WO+/X3VHP49oSKy+DjkxXpRwlwTSXND/fdi13MgoHaBtwlEZ919y/kySGoWkzRn0
Phec1JQ4GRv1ZOTTJFQdIH8nLlabMFmQFlVGl37Ih3RtwUqo0j606NYipvzBUmE6
Hmi7ZXteDiYeS3PxIfFRRq//Trh0wu05U6AlpNDm0aPkGv9qe3/L+1e5J7nzZjud
bcAQks4UfUGTts0Gp6R+XsSa8Xpb5pu7obah+vF+lW+djsCvcb8fafm/3u4trqfU
3H017yNJ+UIiqaEMaQEzVofIXTxaaX+E6sj853SlC6zf5+2yeJ51PSrgaCYNpzuw
ImaRPxuWZA+0mMr4wH5mtz6FEriqAyJixX3DBmFw+iS5E4yik9cxF7XzOooMp6RE
u6PdQdiHoRR9wowOUImcJhtSUaK12RcjkFa+b34KZgp454+gpPw3sx9uDtw3O51z
OXNJCu0qiMelhucVbndDWTTNHFONw0NEpHDVzJ6n7AaKDwaDibpDUmarK8eh75/5
1rb4icpT7EzAjBOzwHMQA4j4K0sMcJMkp8alRFKhEQlc7L/EwG13CeUM2Zrbu4rA
MXBp9PAT/oLZffbMKC8DxOAkGjLndTgIOGvTPhYvi/vb2DwRHvCkXaVnswCMQsjZ
Vdk2fuiydRRHTa1oEJ7uLOE5Zehwog1PMF5OWfOamK5YKiW1N4oAq//rZulQ/rQ5
UYTqScVQGW4Oh5qE92CR7QshZSQv7UuWremnwZRPq/vuZ06yJdbGDK5SjlNLayMw
3Fexet0vi9rv5UqrvAzR7C0MevasqxxUPSsztEj2iZfgEqY4CbqEUSOf3Eu0U6JL
ib/Ea2M566Gx9WWwb7KrGJ8LpPdSFkaSuOICot7fuGthMHjRpwqGT8O4C+HM3a/j
iJdjVS7pGaLa7O9/HOfgUJyZdickkOsUT51O+Y132WcVXDkrU2x0M0HunfzxBM9S
5Kiv/DgpiMKj5VQ4mH8ELJ3HNm/whHXWONfLw0X/5hsKm62nKi1vBmM6E3AW3s/u
apQ6CIkKbM13iB7V/UC2fH5AZRFrpQ0AfDbvnA/zsKFkWHYi8zZOmFd8fOitcJjg
ivpOKvNXGMy217WSBH2SRayRKGsIa/cr6Fr+toXJPqtpSt5WJ7LvffeCGbLHGvfw
bbKa+qREJr5JrNzzGuatlq8n5XXqnu2UvajxI1ca4NM4KqkRIMztG6APi7TaRjkB
JIOOz39FLsn/kwu58/Mg1d8f9kv+SFbSgz7yvmaKGs/bCwsL76CEFcUK01cep9+R
7I4SnlI9TZWErW/Zaq2eSdMx9kK8rhd+srL1EhCOT1iRumi2C6cvizI4NcjOQ87i
geaYNArt1SLd1/3nXYYlzExIJ1c45dg4l/+TWExLrOJqGgtZsxB3weAsUL/a4K75
VQykkh97TFqgn0C8QHBXXiPXSG6CsmHJm4qfs9CHuf+wqhqL1Yn6jHSulmu2I2VP
/WmS2Ow/luuCoqC0N0RthjHUbs1lonRcRf7vFvTEhVtbJ56XORS4OrsM9H00LkSQ
S8ANgZzx28FRPtF2jPHIkru/HPWMLSq+vgy4h9c/VfIJslWA1OXLrWuRNcZNcWQk
3t2St49bHcFHPdo7XLmUukUAu3tCi+i6MH5w6pzVj/Tq543wjecH3poPpJ7rGUku
ph0yqAumz8gAc0INPK2ChDBYjTywo1u2EaHVEKZci06QanLpljpoIGV9b16sQgy6
FhEsmJ+jY9n1VtTFvfN8ouJmJxu5cqdiS7+inpfxgY3v1t987rBWXltN85HBqGxL
w1GDDc3pXUugXXcfHGnKO2HUCqmCaQarVTrq77vrNJW/RBqEeMhcQxVS7PgSJksc
VBFbfAd89aRs6bQ7SINlUd/wzCoZqdpThST2Vblox2gd/CyXJoddnYYVE/3DCqRT
4wrkRccLmBDzfNz1qm/90+GBcRntHnSw9y48YrpxGrC+P1PlAPdNoV2myIUmFVTA
2XPXrldo4K7FTvLZw0K6olYHS4ZTJfmC20Fjl/AJCi8Q1At+qiapWVW2mKvF+O88
I68BLNG/K+TKX+CZ7FS293fsSXaVYzlR1tzgOXoYYg/VBUvju/wzN327w2rvapda
PBCxYZpV7apITAMRIgynhlXNXeVdAhp1v4vmyWa9zDPSzldu5oMzBlC2frReerSH
I+IOJQYl4XB08j/HwimGJMazg3pNwqVmQG0TpJVH4Xqmt8YS7D3E6GTkXoHxnzIv
AOONLeNXoMlcQB0bVi0ITIXZQQSyrz8j3hAeWWsuMyUdUR/+xR1mKAiwhmkpxuon
lZtv22MdumXnE4+PgcPbnppYFS4vGfTy+j0vUBH8pH+Ez1ShkNaGmWb2IS5Ouri0
wlLSr+vdYX7CeNDko16pDvP02sviWV9iCcZ2nwhEk5qZilFG3HvhCqANBI3xzY3S
S0EjBJAZUfB58kXp2Q9csTaFVTB0vzk6XqYfHov76UGO8DNpTHZ15vcNa6R9c8bm
vwZFsO8x5PKN79X9TAy/m1dNODH2Y/ALROzJrccWLqVyLO/lhivvHOcLQwltUnoo
Wy+65ECmRH3I7Yjyx5tojWLvFbofvaAoNqFRy/F6QOmCwrMd5kq8gyjep/i0O/p8
inCw24eNNs2IXCz1gEW8EmU3y5mj4WFrPozebyyXKTBkev1YqrC0deFlc9F9QmkE
DiiKxsDB03PqXbGRf7SUbLrySI1Dis+zuCcl22Lkr1FXYx3Ec/rNlFN3qdjioyrT
dYw53OvOimcOrPrJsQxy4AwIxSSSSRZ5BxAog9o/xK460YCpsCDWcJHnYukQcUGF
LJ/0UmkXO3xwGvaFI4Jei1Q4T9QRfbvL65G76Jy2yuGy5MYJj0y0SibliC+mKnfn
gWlFeXj8rzJuRh+6BnBOxinb8jTLli6IOA3ywBmpBiLhaUyyBhHY+m7aFola/jDi
DbJuwniCVmUx0ZyyxzeGvpnBB+EMqGsVZvz4I0tfydutWOsdaFYsvvLOIL2rad+p
lXS/ugkatr3N4zifeiFLkL+3PVbVSIpa1E6ZW4e8zrxFTY/jNNKK1r81dRqEpnPv
D7KKjaZc0Eo9nbHPpg3a3465Dg1FvOv7/ehcjp8GL+29GnYaFUfIeStiu3bYHy0+
Dc5I3VcfKVlQBu6M/J/cPqPUjJIJPmIhkMH0QaKx5QJ2McrOWTxJw7Rdy7pXjHY6
JRSEl9PSlYDH485x5SH9gbKiV515E+nLVDbBL1KJSvoEKIbZIzGCy56cJTkP3YFh
9kRCpMYH37EVvL6nWw0Wbfl/YOa4zRYy1+YeJ5DaS4CnJ/IWvX1dKVWyh3yyVIdg
BBrRCBoG6pwVm7JEqnpvZmattAokwt9q4oTmkqxqjnd6Viq98OL/HXsDrIRpVMrB
ZiBmEj+kWnYYD1Il8QaZ8miYfnB5yt8F68Jw/ZcHUZV7+7OVKqMFE0GR2mq8XgjU
nSzFzKK6n8RbNqLcP/e07iXJ4/oY/Uozk8RvxxDQuxIPOT+eZBd02vtelYg3RIA4
quu/Ga6/XcvsWCDPcVFWNApIrIWaP9BupRZ1TbQ8neEtBQdzSV9aZN4nKi7uH5lj
7N4AMCj54C0VGMWnTlsl0frDdJkI5QPsT6UvtvdkLULwpfojWDZcSBD65S9tCmx+
g1I8vfkqvVGHdWkDVr103hxCElHUnnKGmHU9egM5banGEYu0+yV6i7uoHnZtFS+w
HDPEXfhn8qBB+Rl9RVEpQkjExMxueYC9xy4q7WuMLkDzPkXmb1q5Xh79Bxzr2NU3
dvVXV+/CMs2/HSzUOy9tbuMTkc5FM/bWJlvrLmjs96gyzGdJBj8CwO3bUFYZMpFo
y+8FmujCEp2SKStNDNEcvaiCDDrR7UH+HpmjJuFwQou+j7+15rfrlr6dYAZw3zox
/AH3tXWFG9ULRcgQEEL69fDbS+yliBseBtNLyl/lud8Hy6GR9oUOZp4uOTifchG8
x4iiTKRZy4u3JiING4W/7uuIys2rtLpIYhnio8PWorOh7bZM0fb9MlDmBpFjHQqx
UesP2RXxcVoSxtQ8TawoeZgcA/GqKznOPK1TqpKC28Ks9r8tGXiZpSiD5NY7fo6A
ALtXGiJlVbzh3YjkbTqkxnTuMoY8zexfaKc/AH+ir+uKFL+1PA0bP5c6WK6I+P4w
FOI+0Ez9s/g25A01yC7tXyC49G1DuTiWlAiBcGh3MNJIPcpN12GuN7QJhAg3DnqX
EMlBByE1alQm0rQ+DgoAaI2lQV96nFqf16JIuMTTh06GMizdEvgKyQwN9vfMEcjQ
FyErTTM71acKbHuZWO+3aTYeZJBuaQRYbjZ2OhK9nRjwndX+mSo8EiAJ5Qj1/q3X
ln70Ccn2w7GkMyAkbKXg4vxh3KQIbpoK8UCLNYg56lNe2YBJZgaBSbQMwiJR2Ypn
bGl1k4OBnA2L/aZrKM669T/Dfi+PHiUlkb1mrk79x13trX+fUTN9b49/tyoadTwL
4Mcv5WgZiCBqPwnlckx//fmnzFx5w+giSjhUj3v3+aHjGPO/8+hfB2+o/wzaLnzp
3PKdKRsAJaCnydrV4mbXJ3NEsApnCFd+XbYtCwRonONcUvQ8rdr+yeYGW7QTGLBY
gfFHTz162mfIY/F5K2OWKlp4RZiolmY0V8GgVAcs5u2l63DVraPL6+woWlrfI23f
1vqwzEBefcAOVvFIyBPMMSQmjUhYzkoP9azzR55xy8MzQeK8NpoTzTledypc9ShG
HLD6WnMce1Ad9YQ4yU1QLR8F1KWCK8njydGBjoEt8va6vvLsp8rZzMnDCKAcpFmM
5JgXkWAFc5dF+7OL+s5tq6VPpzqAHMjLnRr9oVjhMiAzhcIlymtkHe2kryXRB1Lo
RZDrWYxrre+gWRNgrl/o7HYwWUl1HPr57dXQsEX7dg4cGNGoLYDl5n+X3srSdHZi
LeQdhllEx8Qz8G32feBbxs444nlQl+/ErkEsbFiTYH/dnAQSx2Iim9bD6suu+AZ3
ZpVv1xwcnwSDXuAGQtLJ/DbR+395Pzu72jilW7FuRWidi8/v930U8cDkcU/t8WNV
6T4ZxGnogUVoqpPGlcpq9a9ZwV7yTo8i2VNdZP0IwTr7ZbULtG2h3Yk16ePW3gv/
xYm9u4M/1PEg2NekAFf6r7F5lmV8ZDq9w/7fJwi6ykRx7OF4T+fV5+N+jh7IaoM7
RIGgNadOKbuhAF3uSw9g5TJjc1NGaulwosjzNIj4k4bvRaTI5AZ7QPS+udEo10mj
zL/hGdFzBZrl7P77O9kz62MR2maXROzmzfHmggak0wAtZHCItE1EBmEumH0iA7Ni
xFlkkVFwON9KacW16FyXszrWTxi2Q8GOMxEZPEAyZjzk3roJYc2sIiNK/TVWh4Ut
cHLhGSfT4ZjA6p1eSg2Nw/OaAxs8tcaz4eTmcauKG6b+6iK7lzXF3iczqj/E+Nok
Dy/PMCWLUK0jLpCOlHmygnt8eB3ws1qORwcB53wUXX6pGbO6VE4eMjTfabD/SNBv
t4Qb+k1o82J/JsOdK4ew6kGhbfjvkj5GywmAbaoYNY+Di+hiC+lK9M87NxZ5ekTU
drcT6TbT6FOPRLp/Txk2MYCO3KPdPzU1L82QDoE8xcZCfImeFHoLR4KGVqiupQSz
DQbVKzVwJsO4KXr6ARkBtMuLTiPDMVduuabaKdFLUd0ML9UxEvCQvi998oyMJG8E
9L4NHqASs3hrgxKdSjnAtpSvlfs5Sq1XK2XDNDuZHmnyNbH0k5qlSclMBDczQQvX
WAwK1PHjbbi2w3cmaBAdKtjJurvEdMe9QIGrQSdlVgODKZkJT9ONfo34nYjXvY5J
RdcvdOoQZT8q3nbjLfwygnIoTLyqXEn3jL0a2Ut0zCfI88QpkNiIVPwwdzXKSY+A
cMDSIlMsyP5KqhUT+ISVFOejH83eirs0ll0enW5ogObp2QOSE5SsOL8IwQIVqRU4
Wq5gGaGLFz37LDcgfSw/PHttKsD10VZqWikpESHtyUNijqaUIxGuoykf3FbgbmmX
i2muFPl8dwSTCQL/HjJ65Rn89QAbPRUGLr2UMyYAUZ0PqtG0sW/GEJj78eUQopPK
F+2imoMBGKq/hxrxINMTtcz1l4apZW3md6QJaYAwWz0a2k02PB8O9Lq8etgh2i0q
h1/NIvEs/m6gzklhsRqVbQCiDowCmNhj27QPww4KhQiFy30DHtKIAmIpoWSOstba
4+3+SZorDqwFZLL4oaZBbHTDDs7vFrAvkeCoF0QwWwMntJZwCWeKJksGH5/kNq0/
0uKVmCUOkmlPZCnZPGiYF17lRjZIgkkv9xopNUG3oUD8Ii//8ENipVX1HULpgB3J
Gfn6zNFe5LDNr64IpdCZGxq3ge4xOTggwvMFU1DHQmfD0UA6Ofc8Kj/oYqO1Ezy+
Yhhf3WjZRqunHR1f3tjJtPay7+CAO5AsUtBJ06Z5uyEmLK+PVJ0gUroA2c0g1wHS
Mifbs/9FWtKQoaTlSlrFQH8Quhlk9uJBLOrNlr6CU7UqTL4zMUBInc9veHkfyAna
ltK/iL7vPNUZ9DrOq/N2PoYmnXbgw9Rp25QqCJBbjl4f7hk441deb5e10tKhGeaT
Kfj/cK4wUAoDXbtSJBgCXKNoM2fEpNoWplc89DNggjKnyl6M/9ngW3U4Z1+/5eDT
SKRD9hXY9pABgZnWalsNmpF588M2re142S6Y7Ufj+n8LJ9gRcqnZLbt+tICaCHJD
3EZPuGArl6iNLCZSAj++2u2JlNlZXKmI5xhxfvHgbrYgwtfImrf7KNhdrVXfYgBE
WBmAk0LzswK+UKy0I0AZBXFAtINGlbcelFjs5vEKNRF8Wl81wH0dcrsGLTrj1WEe
r6jTDsA3eRoW00z1E9wywmFDMIldBUsFxCQ4v2XsXcQAQoMTwdngzBS9YlIkdZnv
884qPw0NYgfyKBOcJ8rlE0cuKx3QlSgLrEQrluzEzm/GCzMZz+adGcAxjkgTl3Hu
3W/hOKgkv3acPF4LNbMXY6Iv+vR0PEzAKe7xu6yBEGLtmAzwGcYPw9cWz2r/zLPt
UfVbSyHpkJ508ws/vJj6H2s5D3UfaAS2dCRbasPmteSPqjzMfApQlVNUorD3eMK8
TugPAbcePXJVb3byPR6S6YUtNiy9NkvLfVlOGgQr27qEVqwXrw9KZ1TM4Mz0QbUa
0U2piu0bz0+G8x+z6yuAWY5YE7SHpHFa4wKt7u9Uvt5cPV/CmCLTsznorIRJcpPl
hiBogqOPajJCaQqcnmRgdlfuttf/ry889uAU0Ft8VoFEO3ZckgmKwp2vPgA2Dmeo
e9dkjk/Rf16MPAc6omE5jHiUirZsxe8kWhWh8ioiIbGAlOTQqNQBJhuk092jih3U
/l9mRTI/ju6o9dT7Nlbx6Y+smU+uCqZFs9/w8z5WyKKmdK3wNtqOO96W5ruBuhZw
VhNZr6NM5xuYYDs6fqw1f5DXbTfsj1NRyU4hjthmMixje3ES+myh0vaqOq7bNWl3
6e80QT9uh+1zqVVDihoHySWQECMOgbmYU3puWEF/SiCIwcCkC1fSBTplF+LcR5VN
YOJG3u3hd8lYHr83svaFBX1rn1nSk39ES9tzM/WB9P5PHGi5RbSjwyyzd6bc/WLd
6EN7WdhcVKW507LghnDgttKHvbJgjkTkBjzImoZuQVx9wqXOTgt/+VoEIh1wSuON
ULGy0fXDJUjqYldhlmx7OagpDQk/noo1aIE5aGd33saZE4fkcNDwpVr5SjyN5hRr
6Rh2IxeyAi8TSduWNku9O7D5A2+DQrkouGrbDnoWLfLyVyNnv4Vs0406RTfjo0td
Q7iNn9VaIv0ZsqmFFWCJs250YwhTDrgzc9cVpFeH0VXzsedzgMfZXMzzaRRJ/Foa
MediEv9yr2ysQYNgG5jEXYU6FeE5/arV4o5uzbRtOeqvsbwvUscdIAbTSqUEZxRW
CRG51m6MJadgEcRLTmFuy/WoS9GoPTJUrR7szGBebDSPc2IuxRTbQZAAyQTIlJMz
JrykqauoL2FcEy/9qeLintXajyrfgKf3p/0PHhwNHdtNt9Y0fxnMqLY3zV3pmn+3
cfDWmk0Myp66zb3B6pNPsQ+/WoW+aBE1aQsVy73vz1fYKtknjb2nLGIGeZGYJ4ka
QLCbM33c0j4aTxzHbKmzdbCqvPGZ3b4uxfAlb0y2r14LU2aRMl61meZbsiPEsSvC
A686J/EIqyWkKTzo4Bgc9KBjdVPttLR7PCWVycuFYnkp5JvAkbe8VqoY+avqq4wl
s+cVJ59s/kMlMqd5R1Q+ABzvq1vpIjPTrY58SBIjQTwWOIMCKSB+HmsvLam7oe1m
a+Cww5fg6K0rGq+KaJcA8GfvI3p9SCqVP6fiY9imUyGsEdUUL7+ePyNQL8Yf9jfF
ufAGnOosN3CNNgfflYnROIPXBMemfIlpzbAJYKo/oNVXqfzv+Vxj+rAAKucvFSnV
+HOKHjcV+MB/oNPJVsCKrCJZdAk0KekhMs5WC3DwLHtftruhWTqNkXiZbz4v21kk
k+3ov+AuFNjAwxTiRb7zqSX11sVeI7+SsXWBWFR4D29qU2D+PyQfYB6WudsrM2nK
utODJSZXpjCuRbOw//GZkQfDF7bKvDEJmNyykpr1AFGAcHlg36QdUrtbJlwsEKSu
Xd/4GV459bce+963bynElLilMCP8mIQGThvYwZMHd00l8VHgkK+MvZvS8N28WIAG
pBZsyU0RraY4jYRCoX+PnzljX3/CPFG8jvNkDnvVhxyNCMvfHUZuCCKfQ4qgTwNy
tX2PwrFAKdEVPcksjOfqE9xdQQ5SFBCHN/GQjglHAxWdTLSQxQrmTdzu8tKvU5Hb
GfxZK93iCjfhDFWXMyBh2CrsjlEAmTvR7IlDorRJw46mCfaYkLnn4vqGd6Zhk3Ki
GlOuS6jCx1RZC+E/diW3UOFGg+z0dK2mT4WJySBO0cs04SnLr/2bprlIkEhkDwEm
VA94wiiccwjZZ+BEGW9URz9j3SGnGVixfX0Ij7ITIhiNc73+3c1eZdxxy4Xq2LcR
qMvOFpFhuDiser3hXoFpb8YHQ+Y0kuVNThYQNVC9vVAzYYs5KI0yHwT0Luy4rdiL
CYgjygmZ2eT/G3I6dyDXSBKqQC1gJJTuSYYmcUG1epbOeIUJNjsioznfGlr3+DGA
qUQ2pmR3qQ/onGkU56Pigg42zjm8TUZHOqn2hhbB5sD00/HkkLGQzfEe4+SuRT8I
4Jp/1t8LlOsXgTEv0TnJqD4HzUuJIY8pLDb2aJXts9gssSj3IlGuavUiZRk8cEzw
UOgG5/twQpONpgE2Ll6KkBuhIh1uoFJ5IJkPMr6iMpfXXWlaqXGf9bAC8xKHRDyx
ZGv6sdpgT+24v1wekxmeervw//UnIB9AsDUGXzCCuLJiOgSAGJ+2qRoIr3wxdm6p
Kmb40AEfaDgo/AXiKjgIIwnUnhNjaw2KNtrBY9gfMU2W2rcVmCtP6N4/TbglzQ3f
SjqiiCRaGAAnEyNrUKInv1DFj5RV/e5YDKO0bUuHspkPrhQPz4Ia6L+PvtoP4tpS
rw2gprULniWM/JNSBF+UZEuDhWG+SNkMKIBaTsHHQ00ff9s2SE1qSLxsM2EKhlBa
U4Uoz/QEf8WsHOGJ/spyGcBhjIYPPoMFEZWQmcc9Q2PKesUly/tHdG30R9uxX4Gy
8xEsCDyHHsrrwHC4W/Smz4BjQPnyDkn+SoJe5J6uu+evgVeoSDzyjjnYOCmJWzet
SrFZKW+zuJmXU5wHyq7h0Zzk5oPW+Nf82zGTyq4nmJ2KL0JR/fMVMK+QKBifkizR
Bftn1cqJqNCA/D6Va4XS+fsbU/WxwwNZLmehc/4oKS6xWWwMSkVX9icnQrJxvmWK
Fl9o65uTYbbYyHu0kny3jlaJj44tsuh6JfLsn4N6ycSToTdLVav74Zo9qW6KXVau
LwoqguqwNwKvsRpCn1R5NMOxBScv8WoTOjL/3QxBTkVJ/BpkK85fZKH+JMs6qRNu
rLVVdrE6nupZwffw0J5ocARLjNexivy9dK4X87w0Olx8YNZMZQNVB/JvCEAN8ZXV
+yfBtOIiM1gwi8IRBCtJ3mbcUc5CV1S3TRJO0LwC2EQo2R4E+iF71r34THwUEDer
/qq9MiE0oXWv31sVzmm6CdaE1Shgh+lrBZayutKUjKXtiz6I3PEnOSXqEEMpgwSd
Nrp2+h7FfU0SDAAt7paxiaWe7iQDQAu9LqCTYhDIuC2uhqgCkXb8FiA4h2T/E1f9
pAub4oEYbD+rAWHODVm9fQ==
`pragma protect end_protected
