// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
P/PCyDHLshw/RmkrRZdmv248PSsKM/D7d+9UGpm8ztbOu8teoz2htMewsUUM7ym+G9lHrrWwFrJp
8/umY7PCRvnsam65v7kpNBHBzikfpSOrVFniQxy/YfAP4Ny6bSsNg6CPhXQsGFe1gl7sHI8m4wGb
KPgTWb7+dExtWWGmRLUyDtMiiNuFMrF2BUwMYnHD6bPNOfe6a3+ZJxsvoyx9/aTAoAPE4SbrDcsb
3mehEIfAFcRyccJGFK+DKrQKrp+y36of+Lae7ZPmvCdw4Nzdfhlh0uxVz1JR7IBd3/QSR0LdU1Iv
G+dWvSHx329bZSwDK+AUT/jhiWGHJwyB/6kXjg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7040)
bNie2PnZpOV3Gib6qqtooTfZBkpU+f7yRx3LppBHV0Tn7eVNNv4YlDMNgS+kehkfPUzNrqnc2khG
kTYTo/DZdLUP/lgVFTUgw3WZat3xouzSRxxdta2Nn4zA0Xo8HNxvzeUrPYWWUpUpJ7UCGlvQzAma
uxyqKA233b5gMYyuKiQhq8T14p7zQGYj7XM32df6Gew7+Fv3JDdVl/1SHhyih9lhav9NF37AkcL1
Q4zly6R4Dwaa5H1HT9h2L7Hd6J7GBLFt8bhgb4ktiZ2edeYGqzQUy91gUKo+lEsRTkj2dtEOqbbW
g9cUu1thSy9maSLJUpwbrix7iDLlF/yB0DJVIJxUCb5vpnDPTLdzOiEcYRcSEdIpUHX711dfrNBs
jRntPVUq3gOgl1vP1fwzrReIQrt0hzjYM/Speyq6KhjGVR2FwXV79D2yR9qH9qEiAnypBDkXiJBX
H5eubMQpKrhnUAislbIGSl0RWd0m3Ke9LhGPLhRoEZYMxyzRx0MVO1UC8pVvPl4pxuD8HJZBt2yC
qpkMdKbcM09rOHUgtpLYOPu/ok7uxPvC+7RUub475F2Yy0fNmAhpgNCymRa1AASWb0ySKT3rFZvN
NIGj7VqC5y9vr7LabK71eguXlIvIpwHU6NNT+8wvEmwPTdaWlXKCUvV20rzXDMdATwMPtBpfLO8C
mD10JpFXdXrBS8tbYIvxFAHVZuKzIVeC39tQqiNIGhMztZnb0/J5dhRtxq69MSFLeXwM2JdAO+Ci
UBz83X084r5hGmv1kHK6zekly70VidcvTqBwzYlmY8AnyMgaxodjpHLX8AP3SdjhxJeX9qIcU1f1
DhGe2kGQQIhEbq4LL/sizZam+B0JG47UBY8hA1V4UOvCm+w/T1a1i1FM2aaj1ZFrj58hGM3z+qGM
5C4GehzuqYaCJFk2TCDJIRor68UYgJFkJN6cq6orXShHsZrgj7Q8t2o6jmM5jTvJgKi2oFf+KeOv
wCdh7zUdzDln+G3FywPrfQtvHbgtwe7ZJ4xTcPDLgP6AE5wkXl+awuZrsAjHJ4SPrmFikY+nlRhM
AqRwHPxpX/tV9f5X4pZg2CcLg7SFq96vIgZ7IAlg7nlQtxqIALsxwFOmhOY3AJmrZIHdN0hNtrrn
8QRbNvhErU+2L+cu220CP8TBqLrYKEoC3hXlYOJI4J0awXmrQJ72351bknOYaDZs8ux8AAbBPNXs
wTFSlFJkSRPQ5oumDbeKIX2gkIfWNHRC9ViKWrumYGvmNkt9HPTlRyxkOdXcT6FMcxHyYnSN8A+J
HoY7JpJ20/u/wbVgo1pLJcBvSgV0p25xQVd7IAhTHuWqOkxmCqHecdEXfDD/USszjNOYmHeouybQ
qHTPMzpQ33yZiY1VUDy6ub18XuptwwY08Z3johggDmIoEqUtuBsxdaMsZyJxkrXxpmflxGM3AuiS
ViOYa6vlMJJPva7fhqFiOGf9y+8AIUkGLVEI4lR6pRie2zZXuQmOTLSiZyiLwH3UEdQCBAo3YXOb
BScs18fePFRVEMpVIDNdFSYCqglsPtCmJMF1GJFhqeGP/XB+G7CNe6qNA1cR1w57Z9x2HMs9h4vo
FU53g9xysPir4iPUjSRtoXzx/W09xjSQ+MKvOyGO163IuwyOitSgVmQAp0sV8OUKUb+uwRWQ1WNu
ncAAMPvNugtv0qgU7vWzNKtxBxIORujfD9iGIrXtIF6hZIHKJi1q29VbPFJ1FRDEDl12kWD2N9b1
RQ5S/cLtKalH8myyJ+e+hkthRxWcxFySM7NDg7lmDGny8x530aFWEb2UC8kvMcuDVluzAC/d6tmy
KIGYorwQpD2+aESk6IRL5AVuwNcI2wj8egwBR7/X5ERE/hq2aAXSpORsLaHOsn6t3/UAFb4KwcLC
d9lgwmEJGwHPR+YEZogWpW6P/Z+JopXPLKzUwXl3ISUlDlfspZmXcLPSACXEfxUboeI7oby01SPH
WFC7LnacioNzrktXSuGxnvExSzLXoEcNKfZ+OyE5uHe+Ire3Vi+enBx4GTUdb7MiKSjqpAN0YeII
qSaQD2XBta7uYp3PhkOAfBZXAiRP5jwS/I2N8Y8kdq7Cu8bJziZKRJ1cXCxpf609lj181KOc7p4p
ZtLw0UrvaxTW7Dhd/hkwW8Xi7EgEhEd9+3aKqT+HtY5T6ixQpy2tIDUAtXRp83fBUNDcCdCo2L6w
KD6NINEDs/D2c8J0ztqxLDB5RiJd7X0M7A8f1GBGRByp1j8BUvLXDvd2z/BjMkHtrWze3EXVO2+R
Nu70IP7tuyOAl5x96I54jFoPg/HgjyuwG1rod11zp10HJuVJ3MJRQmT8dnMPt1evqXuAm5wkSnmo
ha0PYzqPSpW363fNgDVzvt6GRLzG5p2GzOr6qp0xpePhaT6GL6V2idnt21cSRpBaP+N5LvR/Jelo
cnU7+Zj6sCI88Ex6NUlmz//y2KSo7QBZ8kayDQ8DqmHk7iVF/swtNd7C5o/2oNEIRiCm7HYduR5z
oKr16n7TvbgmhotLEAG26sMxh0LC3oQiiI/1GwpxyvkCHqyQ+Auy+t0+b4KsCS/ArhhWwIlAY5Hq
s4mPPBHMpZaRVurCiFa2FqwGeWjWSkvyft4aLWdLYiaWzl4sXkAWrBvV0U8ci10bJlYGaxMu8gI/
nB3XVE9/cuM4mr7or3N4M1WUTWj/w4OltbN3BBx1X20M9av42cvrCT3V9C0yOzz1wx6iZVa0OakG
7Io2q3qoKKASpRUclOwlVHRhcjVnX50oRS6I5lgr+1sCGAGJe2zKPPKmSbt1NVokQh/DElfr3B5N
REnConmng3mbKY7w2b7qtNaxcJzasDqlaI34YEVlzHAzBW4iqwR314FXIJUkSI73DiiLUeshyAJJ
JkTb2TYs1sou8wGCczlPBmfZz6jadanhZ90Qoj4qRwriL6bx096c0kFx3JCnDw2sCBWMzAZk0I4p
CdRb2IXGYcM2ygDsZ5FO46ZqpJ5YRnq8YUjh8675hXe3xl7kmybqM4nzT33IQ81iRKssxyjX8OoK
sfmNY+3KQptSni7t0MDQzYGjavdWYWJ/XliXG2kTHb2ecqNT7J6thydyLOvDmcuan1ugVX4Dan4I
IvkXKy+EPDLoalIya4Yfd+QG0SNRuHnVc5PNxARIagRaeTurGg3sS9mH9Lt6RT+qdZxVrOOaZeOJ
6bDJFS6kWy149Jw7gmvHO752o7Qtrp74uh3q5NCi+rBLscDz+DVY8zQiQ3CTf8Du+TXYVTP0+AcS
55OH0o5E37o28g4spFec3XhGMp+IjFJozxV6YxrDCe1LYLziWItn8oDddhMVe8O/gTgh290RmCIT
kUFX9y14d+lzaU++hNQReYfKNDcGSQH8LtyOhwvywjH7eXPaZhY5sYwZqPISQ/+y7MCWdbuvAERp
xxZk+0D/yGgpdjYUD3RwDa9/0uELmHqTP89z7MgL8HLMfFGt3NQT0/NtWouXyFBwGjJ8XfAkTOb5
hd7teWKn6W3svg4azpYJN7oQg4fTUo93B/YkDHwgb7k5HfCHGwrII4xP9eUbYi5heQeOEHY+z1nx
/uPzNA+/zdzcX2nhdBxIAVLZ4RUtYsMqBArgIVBQRwYiCvUX7zaBBc+B8dPnRrNkXIQkXsrNoDuW
tCr46Fyfx+aVA6LQzwyqm8Tq0vp/99gjzEK6jNOcuE2q/D5AjCoynatCij3uauLBNIy/Ri8X7t6M
EG6C6BKqFD5AOVahwX1NJuU5jF7BxJRGmq+QWDLKNQRgrvsyhfWqx959VD7JbpsDfO1N1bqeUAG1
NGmV5Hnn1y8B6wdxmRXAT4pCsgImOff6oPWGrwMhZgg/jKWzIxOywddw0tegr703YRkfUNAB+hwF
2ZDDes7o2nBd4dTpg5gNUI7LbJXuokE1airVivrXRyBEtrjFMLz637/e0xubKodl3Jopr3Y4rKC5
sl8toBaI+sNMVYTyLK85qw32gwzP18/3vyP7H2Oppc32DhYMoDdZcJquJdilCpd2R01TBuUXnETl
p2GtPGSg8UqT1r7/wSJLUoxEN2WMH28rcjyNvPySaQpxzSqRmNnkSxo47vol1MBqOFbd7TmNhwOQ
gO4/7/4LnKJ1++/ow9oUZbvyfWDDsvRUjJHiPcpGmVxYj88czGsuf/RPG5qSVg2OXb7Xuzc92nBf
/Os7ZOqN1ygFjV+TD30t06R5Y5t4xrMREqmIQI7KG32Hk9QZVOig03h7laD4KV9MwwOYkPG+Fcx2
VLo3rXASuFLoXxbs5wuV9lAvYWgjIMv9Lvf3jX4mxyO7qcYBlwAu+R5eS3vQYY0avY1VlTS1gHoW
+Mr14wanor2G2l+NTDNSqO2L7i32BzsK2X1Z54RXxXB1V5nV8G1Li4g64wnN2ORiaPhDwUhGUCC2
N8m4DutWEDP3yXQCyw9uWb0XOcO+dHnVxi9o0LmWBTyhZaz941XuGivsIUcTJdnnWXjI0td7dMeC
ocwDsUV2IfoGM6OBhbuP9xQf6bGgIc+QeQKhmgEz1P6i69SlnjT9F2ni/Lt6lhTQMR+L/DwQRU8Z
nokcQMSX84lGP5Pg54C/NUxYoc7JE2xuu9q52HD+iyyD+fEOrcII8DdNTvU7XayU1B0GJoH+IxkR
gvFF6Z4xs2KyfQUDY4qZ7japzssXolNWvblfZ3RmekT9IHnXNcLEhaKB6U795sPSAVkCaO05nyxy
9QWrstkYD0B7Nlu4DoEQZTCOqKBy7TqZyX/9YqWJsgZXifniazEfYsmKhCe2KNSljGK1RSWoT+76
7i037HsD4JmQzKcJrhwCq9Jtmm4bIa/HAvzUM0zx0bp7qjTxTjzw5k+rw/EAssc24QURSFT2dzo0
t2fhY3oCwqmVTb6OTEVuIE/WL7XaIyP86ATkNaIvjAUtqNgsDfMTL1ODvtsj9Qvmsnqn+MhQdfCb
NSRI2dlsQ+wYqFbIwFNBWiWDjhqJdkA/1FyP/4Apy4plsOZOO0qvkSOg+QSoTK3nuaIUEWF05Y3F
zVZm0n1r/5adQL3Jxo4CssEdEjqgzyEOCqCEq9I6AqaA3M3+IMIlu1GdocNtCLUlS7oGTb96VLEI
fx56KofOgbyqswl+zz2/tKep1RzGW4fbESxqY8OL7GqIehf49pJOHkLkv0ru/JVOxWlEv+1wHTb8
euo7wKEx6uNF6UUnnYy9EfHSojl2wTjqAfwCMeJ757SBlr1WgDbbY2fWpXhUTapfKmNXQSyghzmV
TKKs+mFtziNYiBGY0rqJT7GMamzEA9kdmaBg4KK/rEc3+9b7JKoWJ3QvuhMKXOMcNWw54R2jPibM
MNn0D53b+7GorIxMae/BEWade3InXJHB065OkwsKp8TotiQr5afXV1yb9FqXQj0RPG3vGnKEtAD8
dviAY7ZIaCHZuqqJ5W3vC5uU1+vyahVC0GrJQIoWRKFMv593oKbjK4G7uRrqM0DH4bDKSLvkcoek
0KB6z+wRVAZkAcscFDS0jrnjkOPWA90W1JM5Fg+60GWK1UlgVdsw54Hg6keVwPrfTaJyvhGTo8I+
hiaLdEj7NVvV01P3pukF1GPlb2V4g6RWmRszNnsIikCudjTQWoUy/xgvoca5imylMUPEyXXMhSqX
JnmvOuLKH4hgaq4KFLSJiBUXvVjWApyJ9POh1ifMvRryXKaKrsNrV75VuUKJJdShp9tL1b65d8JR
iO/P+MeAXrKx71d2i0WFkP9XAz9HuydhQcbcAdewqjOuvpcYfmcr6tlrCDEEeKanuvOlDGEMu0ud
iu/6WJXRv4zL7Nxi8rIpWKTomu/flaCDLecT3B7E46IO3Nzhbdf4GCcXv2ZmxSIJYwSM6pNbYsN7
b2vZd0MCoCe69Tvsl/YyOEgQRBhYf4ei+HFt9J3OF62XHML2J2l6hFkOrtBPQ9huNiJ+jvP55Ibb
WhV0Cb3fJ7wFu1E8Mg+B1AuSzULIYprcRK83j+EtSihz42WLfeB3K/xknl42tOnN/cJ4RiKSU4xg
A8YHHJqB2qRFxzrPkSnCfVG9HvsrBg5uhhFJxk/dyH4y5q3o8yQk5vep9h6zW/qayFLQNaxvIbiR
K9FFAtArMnkcKzL1vx0Q+Mr5B/RljCxtdKoLWPxSXTmwg2o8hpcWxbVrnj7NCD3Ee7/HRlKaIp5D
5djm0NeeMYt4vmRNDDasJY6C5lzZLjRRo3MUVfH1UF6qCgpfLUsQ/s9gpGnorO7qmn2Rn5xx8BZC
ykO2bomSiBF6h7sorbF5RIgC8a11m1S1rGo9YcUnST6InJ4FUdyAYUmogia8XVxCYxS5FX53XrKk
/pHoRdkq2VpaOrOAdy6PAunECDUdx1z9C8uIRK7BiHv34mrIfdUiuJV0cr5CWne+/R+GeVCPcEJd
7TwPixK2VS/Y0q7/R4YAeYoa7uKzCk0tLKROvETDJOfw35XFiZ3XtjR2IKuaAUDq7DWXvR5S3PXl
H5qH62jiUvXQK6Hh/upe+i6fvdtgXmag8muHoxC+N84oqncnD2C/8qPQQn3Of49Esa+oldCjB0g1
zfcmXXPlYRHeTgoNu6RI/bZlDZPYdxLJdKNAxsTqOxWaYWofkpHUQ/A13hV6Ys9qfXwgsV8Jrj5o
YTjQpU1t220XyZjbbmYNKzOKKdZ41vJDoLORbnwvN/gzdz6fmORWf9jfTDa29+/mvj5NVi/euQ3f
HapxxQd+PU8Te1nKdC7OFlPjlJbCZYgc0v+KrCLi0HJbl2lRJDJe4aaB09eLDH56c9FAsjDbNCa1
qw1/fp8tQZivWybNxEty+QAm6MWnKQYESBliD7erB9nLKGDIXm+3nv70I+oHAzN0QmQi0jS9h/X+
eNai3I4G4xvwhaE1hhLBrrE2H6/PCNkhIEejr9l0clgKjL/U1/paV+RYYmflEz6LRQaXynnHn32k
QvfXzZpRf12Ry+154a1AfIpwvQou9Pnxft4dxAGIJ2kN0RyCg/0HVbqhaB9QBFVTD/aCy7SdBOc0
uFkBCrSd1PKatMXycVRDpdvZpKjpARZLPsmNegGw55ZqoPY3dOhpWS2DbU9KcDVOttVmym6EP43u
pF1/qLSduC5spIy726OqbfN2BtjtZk0/QISrMRdxPV+WGBvn/V86jrHk9QEeQbTLHbytgSUQy4oq
0eXx0OHlz+FBIxMT2Qivz8J8+wLzQ0soULEk/giGMzNkKfk9nCTHBfxbtVlO/GwUYtbF8JNKyYqA
LbgZNNnJ6IxFNSB4MMeSAvRjrutT3JIQKiKoyxpO4wG4QziKNqLrQsTOVTYSZjLbuAEIJZzBw6pV
h1tx+TxkNrVc0wpzVcokE/jxoEK43Lw0b6mUBUSAubhZ62B7dKmFVwMMcbWSXvc8ixUChgS8npS5
QSAujonOzEZvTxuZYo4kkhi/0XtPkJcL5VAB6AFPmkMR5Y69bB5uvHo2N9gA3Yes+BcHHTXdZpQZ
w81irYZOP5Uo0ojgVF2G4njltyfsAQsqFBus6ekhaRB1fdlfM82ijeL2ZTpEmzoWbeSjl77DxUKF
RHFVLuyIc0A/oN2hvTkjr4D9Glp0brUNkmdy0001LroO5NFq4sHc+aIHNSpjP4znjdZxwS2EuKRx
W91tNqR9vbf6A4yaU3uJikpJ4Il6WRv2OjGmYZh0cHrCrY4NET7jPfFcd0uoQle4q2op12EPTWQO
1vmMIicvyvu+V1q13baEHIhWEclMER6HEIRnnTdTstL24dq2XErYq5VkjfZOWi7vWIINvPBaN+1g
6CHEgWikxmXABPuCguSHP40M+awE0CxmY4C/eBPh7Hwfxze8fWQoOVA7815I1NZZQsESLqDdRTWm
UZe2m/5uyV4DPW7LNwiL00B5Z2/KGCckRO2DxBpQ8ErpKQX0Y9ekqCFifnITyViniVAfyveJUNFG
4H3t13VmI/QBmdeOhm411qRwyb6kdRaR2ooVEcrnyh+XBgtg5FKHE2FQHsDQyLdCMiOHUdHNoZC2
ctfVcQak4SH+GHUH+5w16rFnImXz8UakXbfHxIVqTG+A2a59hcEWfmohnlSGHqssJ4Ue1ejFohqX
EaNi8samrrsZOhITlDc1ODbQPt46h2NAzCJBNJRpnl+9CU0rg7prEBv9CK71nuKISqrLi6XGmIHr
YmQtEs65+bsZ4W7pgN1CsirsCBFVu+uno1A43v6lD1DEFF7DBbUIQFxnRK2cjcNasYOoSRc4wg1Q
/SCptnwcTO01UpFqLMd4tWxbaHF8//ZxuMpmgZK3wia7AnHdvojDY6+1fSLAfBP/ZFKbRZ7sYVHh
1KuiK9I5Pdec11YXYfavMycnU0UqESxxPyWLAe6jZI97I2Hxa8TcnLiHh5llG1XvZNXBjL064FgH
zGKXrZcpGcLBKZNsGEpfC4Y7528XbDzmjAwOTlJpP4l4D/gOUeuouuGX2niZkLUwIn8byV2UOCCu
BjMvOSZ6J1Se+RMuZshfYwBOzzPl45LyBeeNZ2VKkbVZrUePTJnXZbAlkPB9sOe28Rb/cO4cqQbh
ceoINrePbmBaYGx3mZcRubBUkLnRa/WWr2oYs5emPqlASuhfj1RCRBZfwnL9FSZt+Y4H5KKl8bam
EwFvGZpk6P/zYqJ8zIAM6krS2odWHmtK+A8FoRF5zNU6zZKCou8nfu0NaZv6Md/HuOSQ7O8RHAR0
aMXro241DsNidNHihI+JPcttrRvsXASX0jsBt0jGrJZ66oKr660XvAmzeCti/qrYnl+uagfg4VPZ
Q6uooVaS+LyvuFIzWlIMekLG48qCdK43t0kVfRB3WSbM4p6gph/i4p17UeTKd97aBU4JpAPTMS6+
1vTMX7Rs7jabgpEfVMy/IEOsW1Jc8aHFWC9lGGScs5X+tlHPfVUojv4WCEyIZWbeorZULFKyNgwD
D71IjKTxhKzpWiiRmI9kX18AA8Rx8fxfPVvXZbEmuSbwr18lprx8Q1ScS9sm9OD2eMRxtlNVhX4M
e0baInLdntqUUudmfTVhJUr32xw6fcTWtSjG/V4bmmQyqhqsgwyMxh8NieX3pUrhLDTiM4UuM7oz
xYfRMLxXUqiFKrF512HmBkOG6UzeQ33gYr0bt1mom4GeSCRjjYdhq1qLQm/D9026L2v/vZoN3pNr
C93LyNOCL7zvrQKpX/EJRfffbQseYncM6MEkbZSXsS8qz5RmLNuFDGNxTmE3w/PKXFHE8XYLZjBq
AqSJBdyWmx6Q4Vwkzd7H/FL632LZsGmv3N1oBzVvgTaTeo1VZhCTcoLgound1cLEIknU6GDHpLWW
JRSTvR5V3PuPCpqy6Gk8pVf2lsNlqGsz53CpVUzlYvk8aERy1cCE/WXzhOdjjBmQoRryFYBTKPV1
lV6CFdBm6pDidVF0F826nlZkMUrOoH6wt6gHzVU=
`pragma protect end_protected
