// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:16 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SoEflJ0pH0ayeGRhx8ZH1p1SyyWOhlBr02LQ4oHrEGq5HoLsXe3WILPr9w0pLXy9
/Y0qQ4zAUANEvuk+pDVzZSH4ZJvoI/QUnfIHasADpmyVypgGRTT0uNKeHR3YC+JI
AgpM33HHgfBeds4tHHy2YCs+oAK1keaVWsS9NnKhZDw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12960)
usdrbvdqxkGOLsepHn4TUjby/Tx6JozdP5F3SCVVb2+CsiUY0XdGuD6ia1RDvMbr
ta5W0O5rT5cyqczeHzcyz7y0lLxakHBcmvZE6u/adYPb7h/pBt1xER5VKb2V7IFE
eLTs2U/CnNLCLyel/BaETSPw5AMmOEuZ98DUPJBHpnyZ2GqyzS04yvNc+o8pY1IT
BE47PJiAlvoMBcr8tyb8Jkisty1lQ96ocYntgzauT+XNZd5lDmx0f2ozHHOpnSiL
g0lF/O4wAVsuoh14/5pPsRbYqWU9oEqV84UOw/NntqnYE4PYNzPyvoXcCP4em4fD
n0yhrP253HEJk1RNc6N7hPx2vj3fHzUL16NYMtQvEFGHh78HoPTP/21MYSDJDfnS
AO2jXhY8QaCr4pNAoRtR2LcCzCPvZqTgvoIUVZTtnOlhGC5Mp0KrDcyzqi77Vji0
mNW5gAHGubqmH8H+ejqaogmDssDW+bku0ZUkEGrCIIPl9UOspnBI8FAaappS0oX5
1519uXH8aY8iVZndADhY33/UHp3/AIqRtlwKH42RA+lOvMzwjxrwlWR+LRf96ygt
gUqfVwldTkjmDLwJu0vMz5764FxI/MYOIydjClnfOnskdykrF1vd+A4s0Nzj0eGw
friweiY7sgfliyOAISag9NaWBRaY1FIQGMLH+eHtkax1vrFUvMR2n3b8QAkEnyJh
Sj34ftCN4gRJat3jjrAT7DUYL3Vh+6sMpCj+AUlMqqmlaOpZQDBt1s63cCH8Mqkf
EIWAIEccYb7DfKtESOABjI+K9xFNgxkZHwpcPtYHDkxJRQc9vWjAPnXGO5fr6N+a
86m3LOuj4HiJArm5TNIgVYxV64azrv4l626meZsmnPH/YSQdO3J96zWRomkTwIdn
ntFkathLdCxp21wZQaet40jI2bJAF/cA0RqGgQ+4vlWUOWcB+TWnpU0OHtUDwXfG
78OR/mkRTrqoHrP05aD2hmMMxcLY/e8BE3Mi0ajfvywNn0SQuzlP0eOzUPa1t3z3
jPULny6fU+9cLVFGQ3sBv6hIF9th9MrUuMMY0oKnTE4qNxi5Gvyd7S1huDRl5+pi
bnTyZFixhQl+nSzhIyOeibbvc/70bb8duy8FHIlADMbFVuNK98a1j7/mtxCalkrb
dGkDT93ksCErlph/ZyBgCTD8e/ywpi7iNeDUgj7w9SdZhcObcdb5zjWOjmlZz+GX
wz8pDa81QrWz4AoUbWFOpl+20pP5xIGo+uzRjd3DMfuyG9HpFKQzUv6Bdi22Q5Gy
t4x3DS7EI1sGQgtqTOFBbXefoe48bA7bWiMYrBBzwhiC5WjQ0Xium0uC9IMbNV4E
osjo8hzy3h0sSsPO0nk8F9krA/3uP7QKQPf8FRhJhaJxrgoiFR7Ylm7eUXjXHIz7
LAn84jHQKhV1xDllCNKdYC6aGYVrQc8M5J2/Jwfqmy+cydDPXbIq9t7Tl9yVwrRq
sajP0qDwTwAeMtVHiDBhu1AHYObhSGyLA/0jt0ku0u8wFRQYF4E/MvjiHpXNdY9h
XuBtROrsR6FBLuIOyTssDNnn3X7tu1Pho7rze4475mQs6aUR85o8vihLTlQVnGWG
wrl4tqUlkR2kavR1H2Lb8hGlx2RfxXN86isaG2hQN3hIYf7hqwzYs5nFkAKO7ALT
SWTEVMhF9NuAcV+wdxHxrC7mEOAWaENHyRnT5LWS0C+NmLCmCN4o7ujTmkvklNWq
UAg0zpj7iisRqbCFZ5IbfegVp2g7HBu90BBySNRiJp7UOs8CmhpF7rcP+RbXIf9f
jeAnp9c0DKk76c5JoGmSFy7RV9kTkmG317DvCMRDwx3Xvp3bqaBOk9KQVKd646XK
omMQRuosZi9ZXnSDM6kNLwAfV2rCZkxHvf/KW86yLMtFcGj5mecNRUrvVyEn1gTk
FZOHKKy500vCy7fuHlW3qw6oOU4Dfw4d1D2599fwDZRMDLYy+RGBDWqggIEeRKDT
qcCNJlaKjzNySX0whqJ1lya40Se75ofo1/Wsy0+yCnmAQkUe32lV2J8yFYghYn6z
y/rEAuCuLfhvKEdWYtMnsfXkEglBDuacrXC4MIczV9vyVh4LChITvREwQMOa/sBy
NAu4QtpsuxyR13P3ZzqrC3IU7wJssX0pco0MZHH8Qx+NIKQif+ZgNJrf6S+lSwGb
WCQfdVHUQnzNvU+lvGHUg6m8wBWY21kHUGpSUw2w8w7JiVZXV2VK7bQaa7ASITC0
3Q3oCfLJ0OlCg4lh7BkOqx2kw90erF5x35ZECuTlHoJYyRW0ajmoVWxrdnPIjAuM
VoIJIC2OGDHyl32UZQGeuAJ/AQ1A/yoDFptMSW9nD/yTGfGTHKpJ7f5I9Swm2DMG
7E1v/obmYnx8754wrj8wVlek1VN+LtQ343aF/QyTzDhX6Lsp895LHPsIr9pCX00G
hWiWx7BnKmpXBOopmE7yBLiFhR+aCqvnb1/7HevKj8T9oUx3rPrHgvRbGm0fY13S
gv0GQ0dKvd6s30KGrTuV48ilG1xT0ZxJuy+5ejZ8ZP3QD1C+GR0gCsy5rQAxhHZN
1tsJFuDF/i2eDtGDsL5IzbpDZPlnJ4d5ioPkLZsrLH1Dh8BD5gOjrrtNRPv0OKiz
lbfQnlK10DKqncEMXMUoDbqAGcv1pLdbNF94c26BFqXT5XdSjqV9g0Pz3IekH6ZC
53JH4gh2z1dZGWjuhA5k83oVycUzTHNdikyAfbSQ8It5fAsQUJiJAtehKNZb0oi8
FfXuQA9AeFJN6CF87vSIXK+yhomusWatukXruYliEhIadHl+Jg3fkq7dmNS3yDv8
J1ata8uEarkrH8pnQRwtP+AYH5vhQL6P8bGeGJsJ1FKvNefghPe0UGr5EeVRMoLu
6tFVxk0ZG46X++oN5RqH2hJMP1ejRdCsRoSKmmwXKUF8UPe7/W6/ZLgMkujcX0xU
HV0Jlv4k3jnzClk3Eo7B1S9o8OiCBRgFv8Lc75Nx4zGKXGsniK/m2oT2ZoDEGZlQ
95yrRu6ezbrbbYWcSWCAb8OTSMV0mdn+s4MODkG2qWKZ+FGbA1zZlvVEtj9XbFem
Jip0LaslnC2VQ+JPOLLpCMU/xULfiafwapAR5P+RvIIo1SBLmRKKHc4nTzPrHzIl
aZP0bJ9F9UbmuIyuO+7hAn3DL2WE9fdTYfJpb3VbNFCqwJqrHECPrzGx+jlsM+tr
4qEtRgFQjGCQFl9jsXWDVYf1TsBuUvDIwEZQON/gkO1grXazgqac7dw0CN+yqKcr
xsP65LYD/UQufHv5tI1vNtrOZQLcpG/hiRLbCr7ShHZZNt2q/xa72i4PhOqNjz0x
hF1fMpKu3gGYuRj1p+fAZ6aV7/Zd0meUExCc295J60Y+UzxgR/0AfmXt2UgSDA0N
ZIRO86Qx57ym2MK4nhQLFWXLt3ClMb0t0cLKz6taeWfErMUIu/FPNxgRxv5qcc28
AXgYEYOg1pMoFi08gtghYg+ugyC+vWowVOKeGDVIObo94WdNpWsCjmr7VV7pent7
r8Bo0OVwRiCFJoNEeoK5faSt6JgKGmcRLVLuOEzDDnu5fvy1AjWNE6aU79Clbtp3
ATys/fJ4TaOIGDdrwiWfyuKlIVjIZpml4ngD9n7ZChgAyT27ZdnRmx6L16fnOkey
1N84nGINnbC3I0wyY/beMWayUhdZH7mnUioeueWm7grJOcQIp8RWEYftHnOXizhY
sMxIA7W711/4SyUJqJI+qUEqJ3aHxtpkpCRZUrUP/6yFJRltWFko8BRhEOKO9TNh
BX+m2zKW6L0FzhSl7RhyFM9pySehwiAhtGcTSQJJMnjXnIQ3UrB90RVw+FXdTtXK
5Ij7DjAV3tJdP8YFh7LAT/d3EpWBZA4bgeyyqQTrkRxpCWKjIFf1StHIgGNScxQQ
wu0fEV35v96Hrm12WUkN4YSMULIXhOxwmR31cFqPxlcsUOe40j0M7syz2NRe9Mbw
0rbd0fKJZilt5ofILevcYFgLgZUgkBdwuufZVKFwse+MPg1VfFQn7r9VDw1wyv9m
3NO1c7dYqA/Wu/x/ymCyiT5WMvLHJ4AzkLbGkvKffhbBANYUVQ8/MmlwFNyxgy4d
nOl2+amg7gsPEI+2PcABu4qrNVFaAZ6dxA/0gqD4b26VPTXC/kOot/Rxpam+ds0Z
il+ZsaWvU1KKBnow5ZX9BGIbSiZ4dfwVcOxVnIzevmDOTKUmIh16YwCcBvSMyiSi
0QgJ5j3XEUdBiREiqxHybHFyr82U09e89YLbi8kCR/93j1ufMAt1yFIK7khN1AXJ
0vH9qs2Kup5oVysQdCbAhel5R5DgyvEgZzZjG6vucAZ3r6ALloe/sgpVjeqZB5En
m1UAQkWXR619GAN2zYndpLc6dSadlHueEom73CnQpF8vYink4OXEeAhHV4x/UPkD
UTP5/6jpXVDmBhTS1qPip4bVDIA3ljHPQFcPgWqiBQ4xY5X5wyLj6dc5mtwsJK3Y
swZq41SfVqHoXPksk8QspdrRPdFbHIr87cmCj/fyOT/qhleKHm1obqiRn/9plghm
LpDzR42MOnd1hBJqEkkOAIijZiHDGk2PowDlyBNMvTKPGPjy5sv7+YgvIZ4q3Hb2
6mFpFQChS4Ctzsyc6cWcPmqXwjjGhL8cRRCBZWhcghTYqOqdLJHyaPR9iZQ8SotS
H7PgCoqARfh2WBXdxgfhHU+KAFoy6t2r/fplCfwnrEt45csber0wsjKBI2xAyTyg
PByOJJp9L7EKdtZiHreLjeiAd8WV+URTD3EyJO2KryI38vneige+M86MaS1eYHV+
0jz5JP7sBgInvgCwG1t2cMvgPBgxgZ4WuLWiUfsOwXKn9oPXfNd5o0jL7o8fbXFE
KqhPpclm6Pn/J4A4PPn19jnxaJyvkpCu13bjFRtsKrdf7WP9F4NaHOL7gnsMiR/U
ld5qPPcQ3rfHEha53lxESNgPoFJ/BAyOwVH9kjXvSkXDfycw894ec0YeTpC+cEY0
hhnROLUlHQ0uRjW9dssEkfNVA2rKQOAp7oHpd5XsZbWP4rP172knC6eK6FC6HY9D
wIiZmY/CB8Akp/tEk43qSc+w+upbgtS3cImHEe8w77LtrhdzdoaXRLhiQ471aeh1
IgCGz8Vc+s3C+cGJAmXW8ZZS0XLL2JGa9sDUXDjVsxjlWv2uHeCchgx8Xp+g5Vwh
X/CoiabfEw2p9pSQdokAt+XUBHb3AsmwhFKw6kxt9KHUMxATr+nXz0M6MBunAYGp
eGPgWXDwwcLcdTooVUlCNV46dAe0Jgy9Gdl6epoeKhe9Afw3Vtax51uxMBeAGrDq
BIHTZWs5R3G7nwZjrrm0KqFq3nlWiG2aTlx7klU90Wn/sfV/QHLtzKuOBNQMicpF
tWoM7ftLllJXtPj6llLeVnBGC44pOO152tBX+H5afD4bMeoBTxkG/ezSR/mQcrp+
B2GlpdY9PNZBWx/4kb6eYP8geC5ezknFh0R33/6NnQnvWAOqW3KRQpoNxf9zj2h9
rAxtf602QXLWZinWKjBswR1Cl1BFubPMz2o7nKfWqz6fvhZEdO2Ido3yLU1uwEbA
r4IzkpXnWfRe5RCGGSdhglowQKtaQuzms2LuqaIFgbUnmajYanxB+WgpcQJAxwo9
Gri5H6/DME5KaiuhIYl6Ey4jSh7Udc/uqbIUmWZzD+ayutry/XumGKE75k0YGfYv
NQgIKqqmKM9K1JAKyOef/IdhtrBdZzJ6ZsI10sr8W7C3C8HjDSUw4otl0Q6AF7x2
vRKoH1NojxtnbY2PcHQMTdDeBl3xNaFBYRhL6iWHHu8vuwYGMe1gVbFzTBGM29cX
QKyhRlAztoBGVlqGpIgpR86Lsl9fUt66wHpmAtNB3SqPqiTWh67BqxKzjtEiUZqT
PtnrmGfBT7BLYDH2V8ZG1WMzTQs4NW9cmwb8x6mV67GUYEhr6pBTmAe6AcgGXGwH
q3Thjco4LQxXypc/N0FK4DRKOT2I9Ik83sjaMXpj3pDxSm5PRl1jtbpwqG1/ya/o
R9tl8tC0U8wYpVZwMgdf0lBbb+GVqRo/wN3KGroehgZfbtG0ORaV15cgyUH2dBYG
KTZPBR64Cy450rb8B5BcPkuoNz+HmhqtLmgoJRsOz1PiSjUzq9WdQmoDrf+DpkBT
XGOBQsFV8HrshKv3XPSXgi2Hp8p5ROjI99v5ci6uS9jYij5tUbS9VN+MObEnAESE
6MCBbCOvO97HWj205Cf667No9eqYdaYZSKZAI/Lm593rnmPShWV5ksGOZfVSLNFC
1OrthKAc2qU3pm6RTdveDf8kbGJgYs2qB/091/ZG31Bjhy1RHUbFjewCSXCBoMgj
7NDFTTcxIZIOajX+buQF4qMudDDoNZnhhNWtbrhQBUXeAxxuVsgN5HHWDpuAQW3i
VEP8NaIGZsdYXJrtjk+sEnnL/IjkBWwohk2Ilc3qKjUzRLUMBvly1265dShWHZ1X
aXGuqEnkGgOnvFRnUg3TASl6p+t1kKNZSXt7je5mkxQKDZs0RTdZkXZ4r46vVxHw
5f1lwnxrA5UTIIfbA88bW/nDEQDIqF+wLpnG/wv0fJAWSfWAAqFXk9vo5jtMKHGj
U9LHDuT7zP1JeTVYSyu0cfSASCe0r6quZi2im6JsksHmMkf33XSwYm10vtJgs0y9
dH54gencmexZx5njHEuIvqTYOJk6q7bAjDu0oWqNXNTKSL3y7WhaUyDDTc0pmGOF
QvBpjeh+5GtoL1SzqRVYDhReoiqEirCj91dQUTlLe3NihR9Zi9GFZ17womXDs8Dj
Yp70rew8cp5QkzKdots2NLq/k3Y5/dbHUwZ2Pnjmg0ZOPAzJZrXyZX46pbrIpbMj
Ijbr5lTjGEXm0uQqJs7k0v5+r3SaFJ/J6yukQF504G6EEdpO3HtfsUapd3L+AE4/
fjGde1laP5TZvRZgzGgShWgH2d1fb6fv07ZsI/6q+HOPBXxGL+2kkqFWEPnRLsx8
sWkR8bEEYt7BMfnfBgfqw2qhFZ7qT66bcMU3ZYNoLtXA0HixUW/ZhgzbHt1GAo8d
EEtlJ+OXsG26rAk6pJqQP75JHJ/FLdgKrFUdPwjXW4ANvtPTvuRNbQcp3IJ8XNz/
H5k//dnvvjvf3NySdNOZ8TfRSS1EuRRyfMv816LQl81KckVXWme6r0mAayXGLO3+
eLF5UpEt6kE5otliBsZ1/FRjSJyNFd8EUfT06Jlhhyje4uB4gYW2XngN1hTK9DUX
P9SG5Am5X7ehFIkdx+NVWVdngl3fJcgDJxO+3JUxhswi2xkuPb3b7j0CTTXCZeWw
Kqtq7tB0d+w2ZeVou8wjxcKJRkYUjqoakEFU11V9EJ45kjESA+hM3yuE8AMncBBG
DgKSSUiKhzdxGIkhX5NhU4F7IFBKJ6OKd+FRVOviTFB0JqTsAAlznDCzWSCLZlfT
a2NQ4aw1oJBpNLGFRiN4sThFQ0hTg7woudbg2mLyKy0BjoKi7iIsYol6s8lZvYja
mlaPOYRw4GkjLgUoayL23YGDdWLCoMIOLRt9lbcbHh6lhMlNQW85ypHlep5kXcgh
QQW8zKSM7aDCw2VcVx+khggLCBid5IcVjSqWS6/SfnHRS3liMzDyF+pT8niwv089
EuqPeNZDVdBjeI3LUlBJKTCV6GM4vtqkB1uh/S58dLDeOToxNqkJv9wRpjNzOnOz
b5KzH9B5T/2BfGRumk0jyeleNIM741ySxSGA6Q/UuHmZzWXCCHSTy+zpw9+StGzt
VJZPIn/ZfjqUilxjfkUaRAaBqL8YoQDs56lu/6XoThfmC9lA4XWja+0FroRT1WHI
Owvql039pXezHb2SC3r6uWjvu5ite6VyLpA+bNM02MRgwq+VGkvz6j/4SaQHkWyq
UD2fR+DU+esSZJEjCl9zuWtFW5i3VYywBYTrkpTQM9nyb7NVWQLy2lhUtBEQD75i
8NcgNplCxWOfUcLhTGC44EbFG/6KghwForPUjMC87bnuEPddc2uyfq4TrclCKENu
QBV3I75Jsl4UIfXY2VaASsoRvrh7JpyQPvxiQ09XYLikmxCD/Z/IOLH4+UGYQWt5
rfz0Zrp4vlLPzWNsoa4nrLQfTMFHyer6bhR4O2lgWDJZEa33IOL35iwKDeusNp5Y
kh2G6mXVw+nbxa37taTtskdZ/aFf6LvmoOp3gzjLbWdqBrXsrkHLDhXIf37v3zC8
3NauNYO0ZjhwGVqzdxzK99Hms6I1m7R6SFKYmbjcg3E3F5GH0wYeYMiQJf215Fxr
9Ssj9YSjuPHwbdxOjiFsEDgpm247oaXRvAI2kWv/i67DBWHCo5lC3NUOmNbKc+dn
tH37e9lyw3DOMdGjzAtQWokUjnVdbCwcdjgmKDbpSLHI3kLKgV4dkKc8aQXuLDR3
6WoahMGgp7oCgY6YEatvCEFAzg6rMxz+RlnKfKxzQzUKMFva1Aze1m4FNI8jhM7Y
ctisSpYJL2kUiNMBUFYgX5w7a2uoaCVk1a4sjttgYa9ZYy2lh8oU7kOMN3OUK8ru
YIXI0XMRCuPATvtuaX17TOD/gmIQ3CwLiaYfZeUjPTpviLpmbAk6jz9HL5xpQL4y
0+7WpU/ctYpAnc1u26LjHEzAY7Fd/HZyrjyitYqwyzpZNunri2qAa2H+kb3ksXgg
boqjLsk5wuGzcXl+AY4dVZjziTAUx520KSCvVBgpMQOWlLHreF8z4Mhzso6DrMvz
vejH9fcSzkqVxEjfckyZzXLFUUxQAJlpxtqmU+45U65AUOMxFsyoPSz3OKbRV/qf
nmPHEBI9A1s06qpQKgu3qqocZRh+isn9kZBKAanPghDHEqlPR0KIun0h78foinQ+
so2UdvFcfrLmUQsu2B6Qq25qP0xc35pzmOa/LJp/i85kisalMaIUF82tgpfQdfLH
gUFstuE2NuvKui3QHQ7APxFG6+KmqyOfo5sFbd3vnR+CTxyP85bqZmyeBXd7Fq2n
i8a9xfEJAd8awqyL9gP5ACslugFGdvEwZaJ1lgf2xkVFNh6qIxipXRr/DscJW0Mq
55BkG+UeYhQUGrNMNQ5mPEFlSjX8k6RLVoj/6U4vWLcKTc78NPhHYTl51spZTzpA
Kb1P0VffTZQlcayLqEuS4jPMF1DCeU6sQELPymLG3NsAuoeLeIJSkGlp0n2bHvtu
UokXQy1AOcXmaqdSGLaxZm2GckRH/0njbN16e1DQp+7fXX/Fxu9j7Gq4lySUyGgg
UMY8w3U60RmDAypJIC1ExBuKwzF3gS9pBXVDu6a9pxzjDeEUk1u10f/oMnU7c7Qs
Xj4FcA3Vwy6Rc0wkj9xvQeYaYkW6UXaSXsEaYmW3vTlKmNk0HDl5FstSoKA/ydrq
3rFwMKq42jHJMd0re2d4dIBLauLbNLHhDrZ0/EuEiUVaym8HG14ABHLz2ZRmXFJe
IFp1xxRM9TztywYNhYBMEIhPrAUrlIze959ims3JU/6ANODClctAcY8KOmsiC5jE
FfJN1pbpCGspK/Rga/HBiln4wNI9exyzu4DzD8yu2QxIqbh91owdmnx6bLRCeIsL
fPw79E+3eU3SrkKpogLMyBh2qimNsteBApcBacMEQ8qGOVPRI4M+0eozr1kvVdSj
W9bEbZwrMVeVQaK9u1NNTemwFBpoXG+PVXy7UGHtVa6Sjk/+Lg3A1uGjoYIn6cGq
Cwz6WPSRwUrU63bRJg7Xq4iBAlWzEvbqqUgX01ihrX1NXy4tseqD5ElehFbnI1Ih
NUOFqCXSuWQZxlVNVV3XOlSf60cfosDXWNNkmtbBOOTc0lwbjUxh7BEZ+Ny1UGtQ
sXHaUgWvbwcpegHkteLf9f3nnBxVtzX2D9lJ1MFuHbkU8JOXggy1aMgvOlrkqb5F
UBBxxmNOoeZE1HCFbvDm0zP/YeEGeZci8hm/77JZYW7BwOX8G1OERfnOXj2nc/OT
Fq1YNfHmyRaU5M9+nyqrSDBUJUIgqlF9yV1bKtXyLKqtMxKfFl5G+NDwPHVZ3eTk
DqVl9ig/bhi6/I8WEzFIvwaI3wdw7nrE2/gT4pn1tFebUVUyupwCJM2acnPLg/W8
P50FfjhltgGRfTS5Op9NKIkSgJfEblfAwFnQYUJpO+qjpVgLz3PD1S3qpFQ1Lecf
7CYaKeg8elkA4vL1hlh3AdJ1EaFqWHeChAKsbgYzDRTBGe6O2GX7lJ4Xym+DLrM5
uD2wVCSFAEUsSuobqOSchC8hDETiAI7OB/S8R4sKuvzxTxGX2KZOda8m1ZUOGqTP
RoV/5JflfmsLv5ZEXKxYj6gjHL3HgiqYikAghHbaIxvVwmBir92A+FW36aY/k+JE
8J4xlHGfncxzgJmHrbcQ+lEyKD+4E1XQcWyMjb4kjg2GldWPD8Wy2uEPLIXmHtH+
8NaC5cb5CiUc5/3VTYbfCB8rPQQNz/lPmWBapIL9yrBafoaQs9PZoDovyfuT7CS8
MGHQrx4jg+s8pujPhyH7fIbMHQhQJXaXX15qFzSA0LlUpyXyb/HTiJJlwJTOig5p
T5m4HzqqO6KPwsjyTZhRhX3+20w+qGradQ9GZFZHLHYXCf0S0QJ4G1I47G+ZvvDL
O53UCGofrcbrBAY67SB2Tj8J7TmRN9IWuJ6ixwIk51TFVJpKqxovdz8xflijlBM5
0549Ck4yHHZiFqGRIv2eL3bxvQM7Pjgu1FCAltH5nyGOfUB5zD5AKIoUsIlG+5CM
cZQn1f146TC4YZJMH2GqvQA7NvexNmSR2sqgfK3Lxm9MyKqR95+Pk8WOYv398UA8
vleML/46GqUHE4vm1Z7G/j8uy+iEMM0TpjPNsQp7atkRAWOjgEG1d6YA5beEdKrC
NES9SexL2R7Qy3Am+qQXRGylY9B1M6b9ywrZAom1LRyhc/nADCs8KDSRFK9A+X/f
3wxtlbwpb9LO8/wSO82KDMJteOC10tjSRHa1ersQizFb9fw0AgBmhvY/Gh9AYtAY
cI2u8rq5S0nPpeDmGmenm/6dxALIBtts0aVbMrU9zE2rjDwOJ/9pzYH81+E+xEbD
BTymcaOMAKs/SKpfpa4tAg3ZK64Ud5qczN4wqT8ogihYOITE10NgrBXIOmo7ue/Z
wrXZIa1LiewZLEv+9fHzpOJ54ZNtsn7hqwHDeYhtDZ6ildb27amslCqJ0I205/4z
u6kUs7p6f7X65JsdYLbGIe/fw5HBFhqBqIfKFVw2Wy5vzlHJI9cEVgrUKSkr0pvV
qcBwhHgALbRdTi852jl/eg8de0B10YIlY+mKFF+QugpZKZWCmV0mBhyk/ceixxWS
hto1yuxgE5Nc4gvoTDZyF0EeQE8NMrp4IWhOb/zRPBHX/RuD2VI62wqbfSLLaKoE
KgawFHZFKxjNY1fATTXbljaQ6HmCXiv8h/iAEGvupsOpLIlWBisvbCveq2wIFtBX
PJqStaVywSEG48LqP0ZlNk7g5Hfs6uOqWXS+1y0iFtamM2mrcLWYorivMtXRPmoZ
gAr2AH82zCwsBRvpAm2F9hP6QVXPwabU/4NW3rFO5HepfY2OEyZym8w3Tttprcmf
+5rYCrAWepMYruw4vjbSea/1HuOqZX8R0oEXz0YFZ5wFsfkeWmCNEFxT5/zF40na
0DjUF5cfSm8ElgiZFZz+y6/nVK2PeLd47n2AYWU/PQPyhQ7sKwDXqKLOxg92F8PX
cE/J4mE1ytPvG8tJHbdjmy0b481jbi5M72pHoi8SEQPURu4+EtZbiWgej7vA5O8B
YYxB+G4EXpb3aIyoqn5MkLzXC8kmIJtV90recVvP0fHa4UOj5MshsvBmIjqpHMxK
Lpybp1LO15Du1bKjXvpE7OGR0lMbwb+aOsFHA3shH58PjSi4RxddtuiHViDzOWEX
2754LZMZNvOJFwkiFbTGSwKXPqVoXnFUryPajZS7ehZVPHsMoNPsdRO+gb317SyN
iyMknZnoUxOe49+o0uGPjSO0BXbWFZreaK+PajmMbOe39vvmVGtXS8DDCKM+JJ/6
1x5I8rbpmwjQ07YWpuFem4zVYyKh1VzkOt8Xyax+SPscNbome4gwdnXBbtc/MvIw
0ev2beck1u7F3zcZZLmNlAVrXXuk4xGAPUU7SNh0p7/pwAoawc7IYLW1HH9cIIJG
m3UQwpgudpi1WH7Oom4Pm89EnIfemq/x8Y9VBBlg94Tw9B5KoM9yNW/OlKpyssiX
hb16OAT9GNgfJxrTkkHzbFgxJmSbnZeX3sixugZ/x25xmU6Z2ZpQzexFfnrG4EPF
gozcEEs8pk5xy85IcT51921pi8uOdGJI+F0qVoeMbJUNyORLVs6QpgDcZ5yJzvlc
jvM54bQ6PQV+sPzDPJWipuoZ6uRuo7+nmJQZnpHukhR9H8JymvCu0OS20M/qz8hc
pzHLgfbdlCapGtBmz7iJYJ0q3ufg47ARXP1jnXJRQ6Bgbr/HEA2J/oOYSgm4nIk/
s+mFko21C8wmyaZFN45eFI4AZ9r2Zo/TwYSYLaX2cmRYFwmujdOCgppGV+7JtChe
nnVa1m1zpB4MKFg5yVbtqT7uyHyeBjfujiK+pT2wcM4x8jM+0dMH5TQ2pp6bMkVs
6Aia7nTQNS3lO+8mQF+4/UygY8hI+76K4nbmMh9VybpyCoa04kNkBhg82fl+amMk
NRGjXxdPzIdQOGqfaOhWzPauk0uEvVxivZrGdpJNjzR6uujvqDER8XHh+YTlySFd
RwrQY2jh+O7i5qF4DmrazL5U/Mz6ISbnQ6GnKOzhZcfyHZsFud+WlASVIXxs41nc
C3bHgi6R6LvIxtF8tAgWOaXctEPHHs39BA0buTr2t40OQKiks9rLNabrMrmwjldK
+xxY3xqdr6RLTSloF8mOWSOoxjluZtnFY57zuqRz/d0ksiV3HRRp3ZHz2ww3fFCS
AWQAPonC38fYQFo8m4ezdUlXy1CLFizrn3e/EXv9TxGHSptTRjwd4KQD0GRKXvIP
ic+JvWPxPt9lizyeVVJB71X4DGOmHx3GTn6BJIKVhHLnHNPMEjJx1emAJ3PDckr8
mNCPw/qse28gWmTXQ8gsSwKsjurniKaW2W8czSCuwLsTpfIsfof2ZSO9jKZQzjwm
MssYr4Rp3Tyt6mfliMyaiHBLqfSFXvHAkNWEd/PNgJjIgvUIqsr/De7muacA1u/p
T6y6DwQt96WG+nPq84Qqjm2igJK00z1GsUyyNAIjkY7olblJlajiIiCMFHhH9ZAH
cHvF6SEXqvbglDETvBF91W5rY81Qb9NrtuaoSVIlUip2O2fuGmBQDssWrch55l27
2XG7IUN6L0OkwbsYlQ+TyUQQoEbHN/gz1N3cqGeAQ+WU4VYSPVGnSVBHXDLw9Ogg
phyGZ7/vlaOAe40yo51UVkZjRKgFYEpfPCb4QdvAkdWElLyBY64Wocy1n5qe+Rbl
oQBU5EousXASD2/2pkRJi0SaKHo0useVy/xM2eK0zi3YstEcWpMYm3Ba4hQBdr4O
hbvhKamADmArrj7leis0VetgEwphJE0BX6e8RFMPn3eQMx7bOvmsjydXXA2GL/o+
unLd4MmRlQBdaIZp/LTPkO3+OK1sGy9FlI8MXdJuF75jKRBdZwwf8eeGtO7rbvnL
6Tf2ogNK1/C2cUg4Ch38tNbgeaa3MTRf1U5YS5SJcufHcBO3Gzl6bIoZDyrrRiO4
OFAYHNvHNWHEJwN8i+ZnpevA76ESzaMUIQtv91e5REFOs1qgKdB/8kzpMhJx+8TV
8Ivja4KH+xrgFKQZC4C/4LGwB3pyF1iGa+V5KfJLPxjA/um2LiDtAdCie3IjTOUK
DS70XMmAdBZbve9UJ23JZqVEzUW5jsIPhwuyStIDIHgMlCDiX08LMxg/GYZG8LBI
ek64Ua/M+uhBEzaWcAFmoeW7I9UISNg+o6c2D/ZmpkSgYo32UmTVKRNbg6snVEb7
inurKui5M3eNonhY0I0NDf2TsThtTQ/decsS4YSsxX/rcm5Oyjm3Z4H3O/cSLzfO
DVkmkwuGNt0L0tZUAzBBq3QOjASLMLdAGHZkCFIR9WvsG/Gtz3fGIYMgEmFUORQ2
iokzwZsJUu6QFqATLni583L3vjbgu4Hroy3bL2mX9LKveiyT7gAimtG0ubM69t9o
icE+9Woj0m451bAF28Eb/xjjF+p+FCKaak2HQ1/yZ5nOgDg6SrR8opgbmiOuATVl
cZhVBJCMTGPoJ8RUsoRS8Fxg6K5s5mt0D7EjlkzEN6QNvFiMVX6/U6umnX+gZ5WK
viGySR4XozgoifaSr7KTjs/3WoDGNFqjdtBXhcVkLA4YlM8dJ0xyJm13tyj9vWv2
9nuOifAlhymUcTyGobYcfpl9RTEkS+FcbDrf2Pokwtwgp9w/Q2Gu+AwFPpirjYkZ
1/jPqADfg8gflXWVTFeJom7qJWJ8HChhD293m+Xt864H9HilHCWOam50jiLMkh/k
tTRTnv4gt737NPnzte+GVtgkTEtXQJAzu11gap0M8b4iy5vwqVGRt4qYh+970mbf
cSkc9XdE9KvUQPCrEHUzjmemboaRUK1mQsyFmQxk475LMBEoLiyHxQySUk6agoZ8
l4nntfXEXW7cj/O52DeNPq9X4vHcvM3Z7xA+nZ5T2Uj3WDxq8gJgXZiXpz/77uxg
UHRlB2GPNHNUgpTZ/7vzx2XhXDZH3vz4kyglXah5q+DWWVisVTYvYpg1GB4Xvfvc
ukPahkekfmSbEjR60rTPwyCXD8DoHA94vUCMHyfw8HGW/h/Gyx+48HhEgqx32wx1
sZyGx+egBIjZjKZBre8fyIK1fppKvBYISgz4CuQYoBGDweVuYb5i3Dy1ahVd6utF
Ckqzasqg52Oa+7X4kYyIk0nOSp4DtsrwLLAbDywsERHufX7PMMx6hKXzUOoZh1/Z
mH2CiNRKwRYOomeRXKx9YjgUrCzKAIpiGDmqjTGEpc42UNhGLr6h+4hP2AsJ38uo
h69gPvBdCmYVsrnplQb2YPu/X+GVi/wP0Iy3J9YHSe9GeRk/S1VCJhCjmFwWZgXB
fuHoikofrFiXr2Pwms0t+jPtKlbeCZTJg9cisvLMCYrz57zrHDt7vOahZ2kcG+HL
FjdPfBFVPTnkVRHUi+9We3oRA5r+GAQxZl4LcGZQNkW51S5IxApZwUYgdLMQPggZ
TU1UPlsSi39C5e5MUiFgzjx/o675Z+HxkXxyiiPnyZdjmIBRFEDYXafuOsv9f8Ed
JWMNqHnlBjJdFvdpvck0JE7eUuzevmWq8SgvIOxms3944R/+ko7/Vmqxg59E2+Ki
Kl2u/mBvyaMxXLWIwlvb0fIYXSC8IDvIOFCo/ZcXhT3xzjIwLrvFgBbL7E8LdXJC
ThwGz669GOq16JA5n0cbwtVWl8tYyCE6Wi4dOu1EaNqi6a1mhahlw7H7PNv+vYj9
6+GpHEP/8MYrotzkHkqI4E0x909Bd1PLYN1IW39YvHCW5y0WLLlvtbXIaHDUnMv5
s7/FMm+ShRrDW9asiMZs+TKsBZN/khZoy+RsN7enzSsnPu540xNK94eQI9F6KcuD
V1tk6NNzfIxT7h+3rFSDbgLMpu/+xHXugZOd8uX6ZecPh0vn1R3mw+zfiNk1jZj9
COoOyoEEVi8kAyx3aLSoFSWkyOhaTsFDE1uT7g8+bZ8dn2bPRslIFZdh3nQ0sBcy
cUflc+h7cswzfohDmOJ1mY7xTwXQf1t4RZC4+siiOhzBxR4pwszPph9hJ88+raS7
Yyxe3dTPHu1Svoolp2s9jAo8qIrxcx0PxmnMQW5Zqyb8sqtgcSvSLQqilwsiy1D7
55/ft14wnrirLGM8sm4olorYlRB/mMbwIQ56pCKd+6apo2wxqrGdXQ6jzHom0ell
LWIc3GcfH8ZQ/jqypPYfy37qBqzKNLRNdcLKvvMUYObgxIvZn7FCLzfLf0VGuGjB
o4G4VddW7UrptfAByAGpUYRO8AEeZv5U0GTpOszlKpUIGYbe5V4tNBuR44JpcMqn
F3m6t4VlxvnWTlN85T2rNdKdfeR8567SKFqLVQ2uiceXhYuw32QwKLkPSpqRGj+i
B0bcx2blQQzlxNFVu3Q2QWOjXn3YzCHdwtMOz2YhwNfB8gEWkC5+1NF4mJvi4CYK
rxxR1zjB5L8OP4hNkyuKw4+gGbA+uMgTmrf+wsDVcBKtoKseybHvU5u6iBl8WvC8
0AjXtvC0KJfGW/a4APh6JjZDrMoYOMjAtunkFcNQeJ7qEkkwLKDBUp32EhWUwn0l
HsQysPcoLo8ABFwjZ0l0Kwx8r+DObuBfsPF/NT1oPbj9SfBmhFltQU3cHClyna0q
0ZQ5H7ovsbblSBTqW45IsvzYbOiC6k5toKZWX32xzpWQoqq9uoyLk5QC+Kduo3Mr
rg31NnvL/pUftgLaaeQY0My3ulvej7SMhRUb7oYOR8zXNh2vBEr0Opa4WC9JW838
ZIUe9c8Sj6g64xhTfv5XbjllCPxlET1HDyF63SPwuA9GvClnvCI89VKQQ619QdRC
FV0W+EuopZ48sNuwI3jgy8R5oFnS1OzmG2YQj/4bkEytwxuLf25oHUy1qGcnL9ux
KUpK/D4WRm8+taMjMlGP8IN0ti0cDhMgm0JKELwHuJmPY2N7ir/035y1deXyoSd7
sIvsayAhjetRTikng6HAPLCLaZtRbrcup6Hlmh2gtUAQjNrzM4wbi7sFT51colWc
qoe8Lh2fVjsqfD6HA4STYVGNz/ZhxUblUYM7535HHlOgIQ6XHLNOS/1vb+ZJUXPB
45GxqS7RVvIX8shQqUPrQakfN1CYew529mo6eA5N5RwY/uPh7rzcsqULElQYXIF5
Dbe3ayMiQ0TouyT8KVowbsqFbx84hdSdvCGXLHuf2AoRFcuWDF+a7/I5Ooyta+uZ
MFEsDZ5DfhoQsOunALIkiMaTAb/Z6aDuV5WgVGQy0UB8Fc+riRcrSQ9UURHtoN2C
9THDVhRNTXaW67MQ3s4dxgvME4VNQjuejDwe7NRxMvCc0MdjqXij5l/hBhhpKdPi
3AZFQcxXz5VVytuxJPAc3AJ+yxVd2o4gzrOWJOjrDC8y2j2vpG45e1jAoWmbMbVD
w45YA/fU0or4o1Y0MQW0KSbb1tPnOinC+obF09ZakTw2bdGeq9i99MFoOJnLeo1N
Z/FDPdFRgSTBlWn7i1ZaamHxZG16jlRZqLeD93uAS4r+cUwTZpNIdw8HAUW8Ht34
D96WTWaBx3QSgZhF28GscPViZx6VqlFdE5pukeigm9POR65ia5jOrGU7Bbakcfnf
AzCazLOoRbQ6AsvQRPRwt7BThBbDM/RJkCM2n0u9fLo2cnYAfY2/6UsJaQ1t58Y1
`pragma protect end_protected
