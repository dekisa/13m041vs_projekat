// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:26 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gUR3t7HHsqsgX5OAmZBE+1lXhOlkHD/EoFuuwnZb0QBpGNRnAUQtQBGfFpDZnq6P
1wAtwR6bPpQicaTZKFUFG5qfvPYRfup5FblDUwTZ/OVnJVAKY8EZgm+GVmAvhttA
Ne2Qb3j4WEidWKUcCTWO0/EHF4uKDJcZI0o1aWTZPFI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25904)
TlNupNDjHaPGRSEcJTnSSxK4s3/+xQt+pkegN7msxGyidrB3xZW6odZg6wNcd9MB
Em6Y2pvwCvkt37OVt9qqvHmo4AU6g+wyUPHpP14y65/4Z4vmmSZHXKbi4/ICz9Ae
0ABq1+zykMWSTuUnU8/kZ+oDR17PwmQTX3aS22598n/P/lIpPncfUUt/dAxAk52Y
A9yyoF+DQFNOBVZNLylevldk6vnn+iK7PQYlapHAfZbm1iG44r9H8p5tmXYt2wo5
+4z0xe46TVxhNKjlrLzem/pzysKXg+Gi8rnhZ9vWuZYnr5IObR3Q/VTo4wQUdKA6
SDiPwZp9dwj/e/HOV04N+KhP9ZTL2elYdzIGSSAsS9ul3qm2D/lR7j2DpAqz0/4q
g9zfc4te3/pVYz/VteMFPXQfRTGhUpLeJ3IrUJysOCvAKGanb0+8UOpL7bBo8SPQ
WartO+yjewDYwb7gW8xRFlXDu7r2R10JR4LY+eqVYrrp91G8rswpnh+WVDaf8w9H
0ShTjkg4+LT5MN4oWkmtERSdrhY57UUrssOOpyTZ9fVEGma5WFd6Vwr69oN/+ho5
cAA/uO7hAUgP1W7Sv8tBea0n4bVkAVQK+JatlS0uUJSpka+WBOfnYMfw4KTafsPe
dXg71NW03yKjHPOgi+JuzIhGvL9Sc5Jlso6yLOlQXi1F6jQJxe68y6GqvNALdUhN
gtWOM9CBBS0axiuwMjnJBBAs3iLwKffwopKH6Q8P2aWQlpA3SNiBX+e9dQ0bx5Ml
Jpwg6QOA3TB3UPOQqfv/qv3dAXrrTFVvJAdzQA9oUXBDSjAp7IuX5jxyTptQhl1w
0NwvPAgYzYh2RNsr3dpgDHtdBk2Ml2pN/UpFgsf0fCZLDj3uOyekQTH5NsMCi6jE
FSDtfFz7+hXEWXEhgvg6LvRv5ncBRkT+0UQTOTNGaxv1JwpWAvg2L4tJOV6+ZB7g
Z/mJrCcXSNSSAVDP1F1+oiY1m274VeBI0Bk/tdPv2lWGk7ZlFW9X7WHn9HqGR4DP
3eAIPj4m7tKyFm6EIUGtmkS39XFct5df9eP+ERhm8IyVRjZxt/ImORaRQ3NjYMzS
5JM+QizkGnSZ4Hdv+J3JRte2DySUaMvg317cUFm6fkN4uEJy9bl/kNLlBb8s3pMZ
MlnE3Zx0whURlBm9lvCE2nG4I0n81c2x/tviy90swOR2F2PQBmORYokIIthD8QY6
JorrGJy0GHR4Pv5vJTG6LPoc4hgUJW/oJB9AUcN3GH3ggdzvwWAoEaHlb8y2jkM8
RhfM04M1C7AMnpdzQwqIx1S9HmIHBGhh0HV8W+hA6NFTSVWSORs41Omgwydr6D9u
Mg6Ki+myPMizMy/G6fbJ+1wfNKTNULLIxXhfX2WFRk7TOUzbQKl0tANHomhv3ZWJ
LFEtPtN+usqcsM/zLCvLp1Ma8jS4EtZNdC/Btv/PtKlKJTrraXw+j489OfVokYyg
8OM6/hMe/o9vj45HB3l4xDobWgSL2abt039Fyg1FCSGMuO/NL5jiexh59rS9Tow0
Y5TUc0AsfSZVpFKfEdsfnEeRyxQdUzyD7qo+8NG3aKRIBBKsxLpEKMM+X+VoItMy
WqRBhsQykkHmcRMnhHrBhnM66XU+Ui1QJBSoHqNQuUYzJPt3P6jxudy1LUBub1xU
vXIMsXDUEdSBIZCBOLgMALIUKZoFFgMeFujg6Cikk4zhWwwZqYMVObuSl8jrUwbn
NnVowJdxRxlHacg3p2UNtt7YH+Jx+Iu+xyT5Wl19v71BQFq5hmz6lGkf/o8tt2Sl
DGZIvMeMsi7+Qi8LEGlZgc5U6WdpvVwo59kHIYVG9LuJ/QpCsO3gcK9XzyAdfJSf
gC708KKctxLdcPDTeyVkD6C5B2JDFF8yB2mPQgifXH+kUTd4YJxh/OZqIr4U54r+
VxjDuK49FSv/4fDoB5z3Ov9aWO9FD1z+aVm0JEwLxO/o9ly6v5dka7svAznzkm64
uUeq30V4uVjMrTowL5XpLMqw5P5GIqz1uRAn+Iyoht3T3E1nWgrmSIg7jvLWCNFb
f06zKIdUshs9BKrlDFPCpYPuBfDU3mcprrWSUOC6cDKrMRYjaJPU2t18eWW63i7M
PTy1Ck+wNkcmVZgLNAnIvAzrXEZnQ/EshwM3xYJm/d510vlBBWjz4HZyetPBTCh4
eZ5hZKWADDVC8PG9UqqJJPf8knuipSGASyuqJxpeDxMJQujvVMpW1CbX0ev9O4BS
gJ7++BlcQNu8I9Ug1tcE0M2LZmRcgKEeEElg3+/kKPHQ11VvsM2sfMnnrB64LNDb
Y5vkXGZrRr0IFxepEZCeYgU5IITEBcvnFMCf+NPQlRqAzbKgpk3CGHjibknOeEvd
1QGt9sdwhCtnVqXVvLVuQPBJQGwOvsxmAZfNave6htF7Y2OToiL/sUwOltgpOf85
t9AXhu5lQsKGUV4Au48YH50Jnfk7PsUavzVPS3QEO4WHLtS5HVRp/7VtzKeyEmBi
XX9uN8Dr5I7VHy/JOZmagKOdHz9jiJarc5DgGYN9gR/OuOzi4YAVi64le+Fr11k/
MLgEYfNpn8yKp/SwEICyDUASvTP1zIioWNj2xtERmHiRSLiidUAX87YVs+5y90pc
3oo3SGQ8HvapOoL2OjnGjBPa6vCPi8WGamvZB0JuWj5ad6czpee6T5sB/yp7A5iL
6j1nSqi4X00tnkL4Iv/HqauC/bWUEYeOttec82WOje7sk3N8JfnreL3sk0TLmQVn
Mra9u1NUgAPoI/ls8cqc3eA0NU7I2Hhbeb0Nfw4zzyfsG4EL4tB14AkCTTu1JhWu
Vlk1y+/aVuQoFzoQs+U/gVIeKembKoO2qXdxBGsiw3d00kXCoI7RLtRA1wuxzdMN
MclKSHl0TNPnWtsMCA6mGWrf/rUWpT3j6BGR7wpz8/S136q0YIyWZwTl44ZcjjnR
6M+Gdtqdc79hufObcEysEGuu8jxmdUufXKB8wwUoyAmVhgiw7wDdi2Edxo+dBqSS
88rVkDnA5qllkBatBOR9/ZdicdNGsR/+jn5oW72E6mzK4yKlGCV6Wvq7+KyCEphx
aZhYhM3sGEcoP1q4jLRqQwcDjAtGVE5e5CEjv07GfT1jGsyY00YlnJquqEqIB1+i
Pc+4jQWaSWvsncN/MXJAABLJJsIV1qwIvbe4FJEv4tL2+/vQPDQ3ooChccCVOI6t
/RBVn6oLoixcuCEkepOfa4gIe9iymE4lVMwCZS0Nk2xMnJViixDlXP9ppZS7Ney6
Pru/dV3C4ZRvqRpaQMQvzBtE+5feuvsoGmXKHB2mRfVAbjBjwsMJ32ef0zYBN/iZ
sWXsagHmw4tLjblzWjZfUdZMTAqO2y+0dWXPR+0wv8UFUmIoWUGer+vqiarFH1mb
luat5ZbNhFt1JzVoyyh8HLljlGF/PZPgCfgPpMk7MDSaWnYVuwiikuGm7KijtFCu
NH5Wv/s1G5+Q+pfVogvMJdJWigLCnssmy+NFAGsjDzpVHjjIvvP/Xj+X36Nai/sF
Vtp3Z+wIFkW1NCtrqRenaAkCgqZzJ840ujLoddgOXIC1q4mjmDGHoaC489UGU11g
LJkJdT/sb7ThArQZs1GYj1qDOgr3zYR29UQCmx4jXu5YRd5RBLIKYCqYL9GM6LU7
73sKl3F2OpbWb3O1QhQEf2R3JiDm1ZX46JU+aL89mGLFjvXXhbcUYYOKgIie6hgE
aRH/L0zagQ21VATWuVqoY7KXvMIWBksBssDY6oON8+V7vasYQMwmJ6DXvCO9Fkhn
6Uebe1VXpprLsmvqbnYMg5xfMxiGhAYBI1tUVTSYZmi4Cb0L4tNXtJgd1c1SPjzN
JqmEwfeRs9bukOvKwySggcJCqgd6n7FJ0qtyqEVfbHumOUxZVxQfjmU/lHAXUceI
X+gk5txpnLOYCIvsZ266QfiVtrTQ/C4cg0ULtjp9/b+/BWybt9cbXof5ei7yG0Yx
XAkYnvyV54/S5tcY9rO4dkE8iZCgKyd1cj9fw70caG4KAC2cIgg5QV8mNnC8bOgY
8d5eZjtVHRLzeBBWmoCpbqNtIwYp6fFx4y+Xt10Z52kLwF05oL38WOvVuefSa6sR
V61rMVHiN9prvW8/cPKcEfcRJiMclJtUJW86mmC4PoMHmaMz+OW+zT9VFd6MTNUF
WHR7dagRWOsO8r/SKZNCpbtypfXBWE0mF3UM1j9O2BhU5nR5ZyQyeRYJ6gRskBXQ
Bdm+WtoFnF/JZR7TWBkXau/Z/EN3wHmYG0IQHnin3HdvpuaL1AJjHOyA4QXb2i/V
SogrMSP5RfsRSK2RE//RBAjMYINE8nmmHJzZwosdslllNexeSxsUc1W0u7F02m9k
vp5oS96KT3tb4t7WGUOD3m+UKEiXhGDjhK6EB8nlX9NTreb67vcA2Jo7ZPeLP8+q
vM1EDoQNruohIeVjDl4BJK2u/Ble4hWjr+uhuiWzSAVQMhHe7bV108dggP9f7n+f
27x22Gd7Xv+I6P4eGnJ2abG6b6Wc8GUpdu26Rg+2UNNyNnj8oDgwL0otSFmgNDve
+CtkRGbo7efjElbrgATCgafcYb0adgPv9ei0sIa2AI7vthPLxDU/NprD5sOyIWSc
luuoUx6rjbuxhmyX1wtY+/AARhQzwRuNnZ6ffVBThVv6CGU/Y+R6+zkWK0aXrCQH
KaXCv7FfFguA1nSJ8kATlqmWpj7jC5J7QU1K1T7qjKQ4RLrc8d8v+wxXuo4ZgTDL
qWnodY3u7e0p0ockzD4EtFtVfFRkXONhkR1LEm8MdLHv6NDvM3PQJx0kmvYjpfr1
O7wuPUfeg62Va6RCTcFA7h4sdu9zdSsFCcnA8jbc7Ntt0MlCHPlKfVWVy0yhoKxf
g+KAlZx2ykepDWHwpkQhvE4Bx/gv/hi166bNFwkSzN5nPzJD6yqicrP9HzYEhy9J
SZcYT2HxW45cBc7T10qRxmNUQA3xtALG0mOpmV98hDrUSDAPyJc6AHcCk6UrRxl7
ndKaa5A18PljhRA95P0NXDzzEGoMqddH+GBfQQ3Rd3UpHVzFK6WAC9wEMjJECXE4
lYvn44iwhe9SC1AquglqkMZ3zvweQnkdySct0VMNK15Man6/vmqba5o/rtSpZ2jd
T3Zj8h/DEiQYW95zlg3mir5Y47L0VVfa+5TddGMq+wgxXgR5OjSc3gO2eeVdp2MC
6sc19lrbLZnfurzzgrMDnQJPFwFT6w+aVoNoUzc7vnkIzgWyu2oodRBTih4tt3t9
m0W6s0yoJ+TmRGijEtCpXvSOuNQOHbiKRb3SM5MQ6jmUq1ufnpr5riMbQx8FSR+1
V1GKNQj9ypQnAdD4Bx8os/PzvCPrDSPEpbApcdxDjjkLDYT0SdG+4WWj2rZiJR88
yNmiW5TEN2gRdTkt4xVfU0L83lN91zb/yhIoSxnSzPvzN9ONpwhnrwJLqHuc6zF/
qX4R5St1RkSw5kzv3m4/IkICrAeR727lWVYPb93A1FOA6L8SRQWA/CSW3gfFM6Uj
b8L0pYtwDw4YuobsTC+R+O1xJfnDjv/2o0OWyRNYb38ymZHQMN+pIUBvhx24ELNV
HuhzAdP9ZsQzRozeI1inypIGb85/7zUyw2qfcM7+dCmfcIjXhlf5Z2LUybRtE1zC
nxTEIZyOiDyGxk3qQoedoOaD/Z11Q8FJByBED8H2EB2AUBlPk9dhoyQoWa2fEF93
mBb12I0uEZdhKKl75yeMwo8pLDcfUlav9M2eqnq/zcsXo+2v8swlsU/BxZC0TGLs
8CvTPJXhQowElik3txYHfIbyHJrJANnyVwfQt0Cwj3FX4F8worIJ6FAZq76sk0hb
OFR/wJPT1OnQpiSVQbwBF6+LfufGLaHxOhBoIm7xqMIyPYpf0bPYgsfbReNWqbnS
JYF0g38DZhwwp7AA7xJ5jdJ9Pcc7bUfcCr2WXTbighq9xSQDMrNP+kHAIqwF5MnU
CEwk/8BCFofQWMFktkJnZOSNUc3TnynPJKOYwVb+mDUhNG1ophY+Fb3iOPVQvLfQ
8XoQw8iDKlew6G/Sz2THZFG9kAMD2o5zzkVivdi7rp812OGQk+J9eiVh9Ga746R0
qJ4PYyX+j1oAGnHHYbJHuCbXP8fkE8O2TOfzBFfo3ZC8cG3UrmrvBkspomSQXxhb
AL5jpAg4Madvb3ywTSSxqR8qyEf4omH1nnRclxwinUQkpkx3+BBnNX7OYddoeB/0
uS4MI0dmG12UsR0zfNKbIl8VwdEMEMr8xjTsaydYhClp7WjQqCcHdovmdCHx7Jqn
XGItbZYIk2GbxWj+IU87+1Gq2m5zwzoWveyGlXujoT7sPUcxnHd86dvdq5/tjw9o
coUhh7DBcZxJhK0qlTZ6oWSwrYOC+Hc1FRF0tPX2adS3PBNVFBEKfUpxdnyLd7PZ
0s9jNEPvLas9SorulPUBQbrQqr+uFG5SILoinYzZRmwRaeSAIhI0MXuT6w4X+GD6
ijKz4/d8bIEqJ1wcp0HXcMyHr7ABcLrXK3WtPRVo+p46uqgG/8tfjgsh28G6tCgL
26HIiO58NGxFQfKyHvYSuExNP+HP120mCLygVb0wLZMmWUYaB03k9ME8ZqoO3XUQ
dhItG5UH9R4gp1WNVDoUjcyR8Iimg/tTiUfBTo77n9ibcgKK8qTmpGdxaUjS6I/1
Gf4oKxxv4ALwFBDTOre7mCKNfb7HPfA+obUCfmwSWUBWpxDzYLFf2itkPhA9DpMv
35tahGTRDmtT9eC79UexamUy6X5V9XuAm9o3MXIFwXaMy746GbwDP6HaEmrH7Nhj
yOiapzRK+D4rXrOeDRRvqP3Gu2m//kZX8BNyHdPfeWYlAqlFsMYM5t4HWW8GGxkm
Y6XCWvJDzVmNf1k6KxnQhzVPf5l7h8JiolUg6jDEXSxEwnqiHRmlYSQKHr+sSKgH
0It21vIH/fe0vyTgnaa8mKnxE3NLV3XYL4xEqRZZsHtswug3a8NUen16m2GUM2IY
THYtBxrv2aUItsA50zdVFYYu7ZtWBa2HD+t72OH6M52h70XTdMqSxIPf6cavuOUi
T4a++JxQ3gjni3x2awcyv7RcFucS24czSZLiFzn16OP5kl9FFz5Hhs0CA5qYBurX
sBjok9GXLZXKiApgyaWX7uKay6Tz+w1a9m6ylFY2cVCoq0KYO0iDKL4q4e3hQKea
spvPHZaozchCV+Mk+hhqp7kv0kkSZK6R5+tz61VC2q7uCprN2QiTkT1ukTbVQxcp
s3r/iPOSelIBYkKXxsSroOoBG/Py4VSa44hQRjosVc8ms4u5MojrHTs46YtbdsJK
4kBxQ79B/cr0Eaj/4h1RxuZzZU9KcuvO2wnFWyZuqg3zm7+LEeh31ldgZFFNsskx
FaWtrXI9+hzDL43OmvyCyozoV9nbDNjuFfAqWZvxBMVZ7BU6AcAPE934BZbbFbXY
EVuuK40lqA8s5XgvR0M3lPlT3HciHJF/xU0lqX9gfZ+iXZlGxhACb+L38oz+DJ7i
hVLi7hhWHmRLTd4gmu0dLp3eEqN2bbb+1TirUjPkueptD0Fb/dlkWkr12MU9b55a
GxtlhRTbV/6XBIy9SBh0lKTsFjJZIZn5cL61KIf0g6xoe+dZMKKT1wBnI0yQT3Sv
TgbNC5u7cYAAGRHx2Zphh1ldJhFkuka8vai80sO5IXZ6XaWcIgohjmFxbLBJv/uT
D+kdS+V+alFZkGtWvHnYGOvfABxR2hWcsJ0DoHEeB9F9puHyPQG+k8b2Kp7eS17h
crZJ1kJqQ8PG3OgOQg+7jVJUsUaTztVMozAvoynMSIAQUFbw1uWxzqTBaMoVYSeO
z/S4lvoJkzyPJzZISKXlWfyPMMht+Yaq5DRF927aCZmSrCv3XCntLltxQ2tObvxM
oCJ2HyDNCu0nKAI1hF/QkDk+5EHocK58yOZJI7d5ag5Yw6ccBuCuAqMKNMuK3ZUh
c0VnC3HwHAS3UFaaora4Pf/iX3T0nHtcLna99nBjFPtt9hIXt8y6AKcbHAman/De
9gZNAnrm5FwX9Spq8qmvHctZZ7eN/ekuzFPsJHaq4hq2rG1BFAdgV/LJTLhvtcJ9
+Nj6wVR4G5VPuz7uViljTv/RvgdvaeVds6+TJ0HYBNCwXm0hwy2Bq8I+n5BThL1W
688hurZa5C9ddNEmD5pIJ6treWJddcmmljP7YV6FG3bsUyTkAX4LI8Mh0juoxv9u
cy9fZ6vWdlftTWIE/nd8kIfNqT4QiY+9Y65eycO9CcS6dYPfSRWwsgPk/uodEOIG
4eT4id5ISiLraVdgVEaoBANfHiLK3Pd9A6WcK+g/AZBpdg5f521l91Hrt2G7MAY0
V5TDF730B5F+0OgZIg/pHJ7NV4b7NHOuAq0s+v/M+P+OpU9J/4otcR6Bw60OBjUK
Y3NwUAIK8I+ZbyjiF9BWGXOIBMPQE2xhLQ+af/KsCQf6R+kDs9QVrHegmRHgH39W
+KqRCn6WCHnC2gVnKnLspPo2yM6vijYKz6+FcVqceTQv3wTjrVI/faSNijfEz87u
IJWVcHftbnLjq9cdnTa+9LsyHGNRkMbhdP+M4jdsULJSWrrPDbwQqwKlsiynbYKb
dJImfvvNhjvbYi4WcME+BfyuUWuU1SBwyspQNbe4x6uJKs5rki7jB2/A5KAu3FNJ
an0y5ljQTWeM1W3dlzUAhMQj3pEUou0cJKX8reKwnzpCLtCFPoWxChQnJRAE33au
BdF32LzxhlI2djPrPxwOBnWBYDnTipdpivTeWo1n8xfF9yVWFLoU2pwfiuvDjZx7
dY0xnFOU/egl/z4qRL5r1wkdx1sPgLbT3fnUZFOkj2n96KG3ppBX0ahCgVwfurh5
ayVRw+EcXNEt8UiF3KBIHjGIO+Yn4q/R0LomIl++sRuKP6Il3rNJBASU8J9WEkts
rD1LBphTXD3j3Bk6ZzAQ68X3kpVCYH42uxuqiYz6aIWoE63TrT1WC8smJ71qa4ai
ON8+tEVdOKtocFyOvgtVdcyPJkpiVDWejOYwHMoOOF67VzYhx2LBtDJfxsb9Zo3C
Z7JBjh0ShHe4BBXCica1wAA6XSpwLn62ITrm+wQL09NmsdyjTr+x0efMsiWzmiW5
Ea0WmJs/mX0uLbS09+7LuNvtzB8D/DsUNjWAMFYJYbTQUF29frHautWGAh4/dIoQ
7WI12Xmmw0rKjJNqPNVA1EpWSawWmzj29B8gMXsrNcxsj1edvO50aWhq6JmComvE
MCxfXRZuN8qHkC+KHbyihTNc4dCPHjt0zivwOstTGhQeW3J9ByibR3hHD5UBjDG6
I5R8zUEeQS/jocNxKC69+MwKUTLZkeDz4HiAinqWS8eTiGpyRdan0lF7bil7/WkG
Zxd1//a8Dtxt9P7KadirwhDUhOmUF8SnnFow6kdnN8WhT44MhVGwbbjDVkQNaUiA
vDkiZsH885KCIjolte7BOwJCKIcQTt2Q7Ks5wUFRNTslWFJPy2uSV8xk2me+Y5KZ
Lc6Bgah64T+kra//HUATvcHwDs0PFPtCQrhEU3nW+vv/XI3A29yfVLJZCTXEK0gc
rDxhqDkoXI0qCvO2oMEcQUatNRxpiaJQl9e+O0wVIsDJRamIGGL9Av0rOh/KNCqM
5tKTKlUdz8Ff3jf7o7WFwRBN6Ww5QEhnAQY/g7YiLQnFCCIS1Uy+VNuV2/ARf4aU
Dv7scBmALTYfvMWuCk3sZbqMZ7L1H42DXLGKbABGmNo9vajHl+ygRbWNEbMer2UF
Vliy2wAfjVmxdQYguipsDn8yqnsWyxtsFtbp0mAhyEFguQI4HHB6jTDFcAJ5tAP0
C9WvYm+hcayFCKB3tRxzhQeHnUDrTRDH2uprGrtpHgA2J9VgZt16mhgCSVWwVosf
s5VZDYcgCnw/8td71uEyVYPWE98zccbWV2vy38sZ8eNfjvH1C2BUAXcIQ8iRiury
TZtzBANPga1UTjz157CfMKIDUmVk06VczgosKuD33//eqIwbVvTPRFBaurhcgdZj
DJTlOGnZinW23gFdbO8pm3/3F9AkvVpvii7iYNDeQhqesg8nPSlE3EdzpbXBZqlF
DDqeqN03pv//5n4RBe+NhnWmqs09ofKQeE0cWHau2JPOqhYB7VUFQ0CCp6zEpuwc
Q0/8k0Jbcl0/FwJLIWqDB4vJoBxTzR8ErQZX/U4f/v4DNhhAn7BAyMGUkC6FsZGy
xnr5ixIufYlWlRZE3JhqI6aApv4nBzRKl/cpnS+VKX5HM3QHbH1LjQMer5F+lmSN
DiGYR/55SP0EoMKspj2+2QdqcP5OqYqG6V5cDEywEmrpVCTpGqjcGjEiAuNrYx6Z
DTjtq8LCGgYhe6hHZyGavEer3Z7ErkIPKzfUx0hx9AptgVD0aHDF8Nm+6Bg7+2Fo
MauDkiGfIwZaa9OLBNpta/hL74e0XwfDSOAh2mcG6mQgQDqg+liKKELaKozG2HyQ
5F3o5w5GgGo4rQcc9ZOHQd27v9vImthL6YkJWBrmAUhY6ZXaci9eBc/VrcgBwgGX
+BThqPSM44k0H84nIOkiViwLr0AhGdAT7u14NTARr8Jkd5+wA52poHNdgiSH3sbe
Kl3WHWkIHtEubpd9+JEU95hgaSSlhcH7lhTANefU9LpObtRuoWaIKWP/NG097++I
+tpzUWg3ZQ9hs/RugtYCv/aVdpEJWVcGUe7NazKkM429HkPUiqRcohQSqpwTE1Wl
Xb5KbCDl0KOi4lry3RyRBjPz9SvvS/QlBf5j7Mj5xHJ2/S0yDq8PaIEiVJsoJ8xT
9lZYWcaKJNr5i6+3ipOINYLDA8bwIWMfPZWl8yXyUNFef5l2V5c+7I3oifMISdN8
SFbaZvpxu1/FpX73r5psN+I9hOgfSJ3d7sZbqp9LwkkVV5IN6xgfGCKHCYfMqWqV
47b15+hEloov6Kmcd7/GNxUyTbxYIWfqnN8dJkkgWW+jxMese4DGB0NuUly1vwYo
2OrIdx81uLmSKiwP/WjFnRGA1wZbM4NKYytBKlOXEx7JJeOrBvBrXfUC4E6zR9mn
3MUzcHot0blKI3aJOCmuNtAJcAmeVl7Ze2UjD0iWxJRAxuL5WFxBAJznYHPxDlY7
PKurGH5I+UykSIC3W2wfcxByWquIYzckeDXhf4kbq1FQPvTQthRx0zs/L2ZYH1j+
OX7ZyflANIA7GV1PJQJpg8m8S/6weK9iQG3B2U64y3GUmxvvbykC1WJoffl2KJCV
8xFSGGItTScvoIwJzwofyzakyoGx1qOjfpemtGqrlhYMsniJH4vQF7pqshrtHaMs
aNGc0a0OLAPWBpiqdHWcKeRdUM2L5SZsSfD+xz8KPBZpmCnZThckh+dLpJV6UkB+
xtHnS36YXSOZzd4dnliK/ugje0FF4uYET978A7LOtYF2lk64PkzU/R9mdKkdFb3X
1dwG9DBnrKstTUFvpABL6zOXadTewjnmjxhF2USDxCVfnr1A0VYMqZPXcADUS0uK
nYyR0+bip6GFpZZ6/rNXVbbSju81mnx1NO+ZBJ4fLa8aYmv6BaT20WBWNY8Tz3zN
i5nZlWZQg6A/QER4WaXF1KMt8f3DWIDb6fVSSvx6ARF3N5k3Dl7preS1vhDsfqDu
nbzS6i0jS8y7cn4ME8YGrmKeBnoqdCfr3Fmo+LSdujrw1I/bYNYcT5kLILlJMqIZ
OVVNJ9p4/GzO2PiVwA57ps/WkKq4nsE2EkvdSf+hGefkMjijTe/BiaSkXzIStGgF
8X1KS8ehl290kjDm+OZDhNXray4NyvyvCDyjBKrwOtXMHvkUXfXjYnScfqBBN68E
qUs6Uukhll3fxplMejpRbjtJshY1N2RIRnbY7RxiRW5ym59Md1FMgusPCr4ZdWay
mMLiIl5TuWsO78Qumf0LiK2sQio/k94GUk7SSUcvC6+2n8yquALQ/oUIyLyH1/R4
1MkEmDX6uf78IVCn/Up5yWnXF2PB6B6cxFF5211yMJPNhMXFid5Cl+9vuPvjPWUw
kaX4/yUj3dT4ueOGo4lLGOS0hB99UckdaC12e4CpzHtu9avExnF3v/64POsNrKiG
MtHIXqEQiPHTpxM3B6YP+znsmHOLn1f3uEThEC0cpCWLR6l3az4tHpzk3VXUz/zv
L9ECvpCFKn2VEcuHntoQkLrE51M5NQxeU53zABeTCwYt01JLv7PcpAtsXOUgz5j6
/8P0nJqHJndLD8qF8aFFWEssqmhLeqpf6plZN/LU79QOXRfNPt3HmXoxD0n8/7X2
cyuPm1hnKCfcWlsXwAxRCf45evpPy/YyOo+q2gWLfVzj8BtEgRq72kYodKWPtDcy
31EVLN2CrK3HD7RxAEogLkjSxBx9FkxERBxeMeCBVxMABMFP+2ReRoIihkw+NEpV
k3abzb/lkkx8VZ4358BoA+LUxknkKTPAVwkORWY1U9WWV6DNsIaULxTuGruaVfs4
KtxU/AmHG+M3RD4Q2x/va0c1dckw3JAIfHWD0xm8v8InkcXFOlfGjkJIFTCYjc+M
/iXMWS28cESh9sQWhkS50F/vVqV5nd4rFzG80F265VIvDFOnk1d1yBzCF+ArAEfy
D7OIufBxV7kbm6Jf4yUVIRWJv4lChJyd78Z6SHORZ9QZjfzzKr10p8Xszo80ZRl+
8Hg2hvHirEBHWV2yEbbvHMaT531Xl2OX2sESE4wATr51F4Dujr778wJBGfnpf2/G
56p2FTIg3zR+qw2xNWEcy8GrAZ7oL5m1EF56s7SB8lTn+CQOkjGZ56nX9lguJat0
zA8s3fAq0Ch4Orm27eK7k0RUcGcQj33Yyrm+KDQ4vMTeae0pvQw7xd0dtwK4o+7D
1tSNe0gGolkBEwy2CPsLDc+EEHX4s/kbSJ4WP0MMTK47Bz7h8aOOtkQ/cbVAQbPZ
McvzJjy/jAQYbAEh6rMWpVKgLHQXnxrc6F28fx3RXB4Q0ObISpbDhJfljbyFBgxK
URS+FLkQ+PfBnZRXdlrHYP6sTVVWliH/IsQ+7bOjJBxVI+thcB3jimKM/BS9o8GS
ZxI9imJ/qVDSivH9WVmm247XVhWjUErqk4UaHUE9iD8Zs/JC6gQyDj9VfNMsJWJG
aySxXU1qgU37FQ6taA4zHr5RcqiMCeL2n4Vgu3MqFB6J53ghBBhrb7wz0W5pUAz0
oXohJR+ciKcWdSJUZGjyxIO+ylkSW7Okpm4YMi5xfILqbA8Ry4rQ71eUK3f64amG
SF5tTAYcVj2BrgsUF7DNwz7sIDia3rd7u+CQsNODCWST6SIXr0uRDjwp5XrRiP4I
zFpBqkO73d4bVmOPo5lM8PNBvD0qwW4VziGCEbfv3XakmU4lifvf+R8iBtMTee9f
BuG8yATp5Ni88CWkXRltIjKfkhVd98cOywDrwUK7fRncNDekwgquKxomf3OPe/Wm
fCbfm90oT2mwC+ZVNESfy2X4/+tnVmQ2+UoqtFLv3mDvDo8sK0LKHsLXi9HDGlz5
FNYZ2ebElHuMwdxACecpEm9vK0sAvMnctaQkVLdRtQRj204bPlhOJreaibKMTARe
BLBMHTtO54Lx5AMjTV1APMqyIsTh+72o4/MVsjtSwhldPHEvkcUxNS9LFBXKPJvZ
VkSYJk2IeQFpFIbwnIOIavdXyMB6r9YrqegpBRXP6CclE/UmFJmAIQc4PZ8/761+
rYWwirtCuYhM/dH5ZZxTm+Q+pH7ITbo+54x7PAUuKORPhRHQUw8x2QSaBsSgchE5
tNjEMvSJvOYl8OuEn5jdkSXHiLkkKANvijmsLrAnpQzba55hDMFrsAFDVs/ytsQ3
DrbcuyoOjxBcOvqEs8lxMLVc9wKGGi7wfTKIh7kBfEHR6sfK+4tClsiF0PSfoEO8
JT6nIz+GxXe0i+xVFeeMdKayHmTyBpUL1TlIQ/G2Yp2FITFLClGSkxlDmTbEUFzl
wQLVV1B2yPNS69ZfjAwbbAWbnbNu6Z13UkChpf7xgwUDBiJL9ykgbgx5nNPcmqse
PTvdUhWdC9TaimCS3n8DMiO7xTMbnEmu5O7WoEUT76ResQcMd3QqE3KQdjfjQ80c
9r0+2Czp+dQZCHGBbRRECVO/f5LiKkFagg+0X1aCFGC19TdWjTOfhvFCbmfxGkGF
pK6w0p33siK0ADGaFV9jCyWmJvgyHbP7JS5hdepaCbCjRAUog/avkpMVAfCJcbKp
MT1BglGS1V0GIxqo6rG2ynjo3JajJbLcL4NPxHIC/M0rOYQxei/Tf37v8kmhIHqU
XxzZAPJKjRl/k1y8KWai6CWdE5uPXtqNshN4+oHtwgxh7TsYGXiAZIPjqbs6hshM
+oGbBdtYZXGqQzgQH3Cu3i2K6XQ9unOWgN7LA+w1p2+qDMEQho6Mk2NeiNaSiFXX
AOu8PqfhT1KOliTxzcK6fa29rSfaGl+e3BBBoxg6hgk43u1DNq1/XvWpkhMfZ0NL
x7+s/T6lDl9R3Pfq/uYZD4HCBKvjgN43pqRYLKt/7l2XPhLDmCPylH2RI08akl94
cCFGDDkpMgrnHEqsqFMfVi+B1GPXdDhcbM7dOOyRcjYXZ0nk5Thh0WfT9Ltz7lzA
kmvbPZ6+sp8IEHAxP+/7+wL/f5QQPYzIUFMN1wlyw4d8PHtKpmOE/qUlYEWVyr0n
zwpeceKRdB+9wMjKaywgfr+koD3HH7w6sx9EH+ZBPHsifhrXZFDsYkSPcW92qQln
2tOGVcj1SAq7wKmjnyTv+pBycrg4HW54iRGjhVSALhGgYdNI81ddAQMLi015Dxzm
eF/89/7tVRgh7D2WYo3KaDqS4ebFivFTyo2E1gy1HR5QiJXv8oUEPrBM8tjur6xg
sgqz0qPBq6MYA0L8I9PaPxfYMnbfH2CBwB4yJrJDJtyleUQff/xI2dq/tfof5FtA
OdxUDAchPRiPz2GKFW5UxzWU79nMUdblT6OHuXzCH3ogZfe3hO2juOGuJqcHaiBE
SkknjXmCZrE8WvR6qcDETf/ITlk38KNc5taAafTAAoNtKsT1Bf20VtYlWEX3yXVP
bR6za2kicBuLHhiVIgqhA1hg3rfQXeGznT1b+r3CM42+uKVP3oFQQCHJNObiLmpT
sS2tTYnp+wlUdjKh8Po/pEXOZ3dfA8qNDpjpDYfC/qO+gLnVjcshtKFn/v/dzHgk
lLN0k6ugGnomybffOWOaeYozPaJ2m+stI/oDpDj/YmtgrJbFZo6Rr7lm1Lajh9yn
b3eOsKKiQwn3P2Ky+2Xup+fPLQTFspeAzVi3v+eeWLmA1ARRhM5d+3UO9/mXGgUJ
QRl+E5qr/WMOH1/EQWZuoc6yk39RsJnmw1qZfdjNZFHfkaDQu0sPvOYf3BDqoKW9
+WqUljkD4PgiVIZVNojSaot++Gdr8bYfikh8TbSajZ8wn5qaFCWEERkWWMBAzcP3
rAGGr8umUWqOXaJEDy++5jse8p/ZDP5GaRU5E+Vf1Xv7Ld9A3d7Bp/+Nda5G5s6A
i8yTm1qFDtjU5hUFUgDhiCVzUIvktcPSAt0ztqfzga3DaAsC5z+Q6WK/KW6/x10K
sojNpPBS42rf4ORKStEojhKoIs1u420RcBnKbI+L4FPZQlQJ6TRrp3f78VUhjKuw
MKs/A9ATz+L5bFzgNXSYU7whyVHc3nXpuY1Tebb18wiFvoZYVSVkiS+3cmiIr936
MPkf8htR5tN1Gke9vguMZKdJdWUWidWFnqfVGTQvFRN+SavPhZmzxQLoVZZBGd4E
KEKil6J/+cRHBba0gCMgEMcZVXSbhJRg1jy2ZB+y5OgTHRFalR3XSRit0E4DxPhb
Ka8/hthvfQx1gTXNcOGR3WTFc526EETIf1lpYQRQ8H1RlgvQ/xn/AyE2QmSmJLXc
q/U29KPWO7V8HUamcBYKBLWDlRsRtqw5/k6l8y4tA5cYmkOORyxT2aN6zG8DG1Wg
tKjRmMwQANZ54k/ohloUxHyVKZVtcbswgmBlTVwUMXyEzqwjFJ0+EoXFm/VmSsvR
GyaF2H/SqCtfPUp37ES7kbhBt15W1GoUJTb3DvoWweIxo3AJ6I59n4c5Eq3uSEWK
IVD/4cGuXxPw67438BTcaTpH7pSV5o40aJOL1YrdkqGH9oIWL7N/UIcHhmBPvnNy
NzCzQngRaXOTsqNM9Jitzq6lDRRHLskUwfrUk2x7wAS4PRj1y+5exK1nlM/Rpfc1
w0Em73aEX8WXluvkdvonstCiZOeWWffdcHow3JAFBvg5/1cQZcE6bIhwDLMeURgr
GD36M2xDfBEthIehqI6xRgWVNbzsjk+U8h6poAYUs4kOOMzziSkkHH+ViRsYQ0j0
9l5gYp+6UBYmNWUJ3Zh4rO3N5EdOLScdQxiGbm9LbjJyDOEcA5xookU4jXOWeF+G
tb59MmxTsbWVT0dx4SSQjsXNHOGFlqpbQ5Y1pgR8DJJ5cCXmgHvST9oEUf8v5XQ9
6wmTITi4v7zAHXW1G2EElALXQjlilxE0xdUv3i2LJZuoMroXNrZpSyzwvRd54tJr
Tzoza6TwOrCHxfWgDbwdUtGoHnzVf9nhJKfc4pe2riuEJkHMkklxJ+wxtE8kywS6
M6B/bKKCBTCl64HyE+OoNK3Kqtt6W0S/VmUdiLYDgM7HNh50HGn+9u0XaznsqjVk
7oJTL24Vd80E0XAQczD7n/Vh3O5R7Pielq7pCVvjN7Z3E/Rk1EsaHETNOvu+syY0
xfePySGp34WJ1Dkh+wCjAXvYEDQ9S09J//eQAo64+JRYd+220lXVPJYpPpiM/PCy
NQv98Hfgj/ZjrbIacNeMnSkjCvXell5pab3vjDXGOU7e4074KMFOLxzIgwZg4Rxw
sz88u7Hiq5rDDA+aAfR6pWI7UcDvuxlOlyH+AxC80cCbeyCDvXGLKEBhIc66rwCb
Fo0Ss3xtOzLTp9vgGnn44hwgSAHeMOhIrkRC1Reg6dW7Q33qBeJPA2s30JYA8JoO
hYwMizUh+jbD3JnLtP4eCRtvlyQChI2olNIlz3V/Kyzuj4ciXkG3f9meZLm168cT
ozAF9AzyGDqj4ttwSB7dumCPsrBID+y48G8rUIuC2F1ba9kMYPH0RyL4nhVJV79i
+M4XjTacF+Nd2DN1KLzA3+cB1SiwUix/fJS5JgKYafO2xmhhBVZgU/4ebIGfYvus
ThSKqxtn4nQcpHKI7UXnbgpHAoLh1jWUVlnfHRjiWuHBdI/ecbvRCoOoSRI2Dau+
oXM46sEgD+5qxHCv0swHaV6W8wlEIbUkkxhTz4B7qbq8s2qnzYhDW1YMALUU9Xzp
51wYSvthI+mMBkRyFOnYuAuGx8Oo/MTHeOLQGUcqjMleSaalAQ1/xI8Nd+z03p0M
mpLwycR7m6hTrwE8D/7UUzG47UrDXug4Tb4oi8+etAMiygz/WjiHpJRNOvtZWZKg
Nv6VjKCLgJ+0/80qp+4t/2jAoCs5AaRd61CQInBdCwRO/DRKtpBXUXgJu7P5XeZP
hV3Vf2QnUL4iXnOphsHC4ltFaVl93T4wpqgQeifFv3V47d6ZM7PL23n4OG0MwSlE
Y8RpM2Y7PPTHJ3fRsz+2HsYnCJnRH2N7FR21okl60dFrfjTldjfjjQmf0i52DaDa
N1qxkFZpQRAE3CSqlJ0tv7e2ibwPrMR1WSepPIyjmQ3I62yHj4CeIhNhNgRnKGH4
jQjzeHMZnIVC6TQiRLoDDeSSaC928K9jeychQwugxx2Nc2unH/TEnZT0Mr4hqAdE
9kLqULtnbQkGGW+stx8+iiWR+B5ch6jst76KxZYjTm32botiB+q+oA7P2GcBGj/4
gbLBiwPcdeBsd9+jdAzl7vmhDEuRf1y9i0IYExW4NZgZ9prYDrVq+2yyj+4J3dq8
tZzyqVtDIrDUrKcLvtlOOVOQyBr8+ZqcKH+mnZvRMspJBeQ1aNqYr0KVZxKBQIFj
eD9z+nLViAJ/254/1BP4SZsR3zxvR5/f0DsiovkcqCdwum9anutS8F5cecqoWX6U
Ev/Supax0arWKLvUVWryUE/hGU67s2OTh3w8wgWXJhRf84wOB7VvUyoAk8CnJxyE
dDA5Fyx75Ey4iEcDjzfOpq1Pp+Y7DV/dzYHvEK2mtOJRrParHAMPKz/DG4PXWv0r
BfJEkjE98BLanNgcnPcBxVCXzXMdbP7M9xE/QljvTvjvCJFr6Ovw3GYVmtoWfYwH
FDMTfBd7PH+7GkQjbamSK3eDT2Odsh5Caol7SUJIDN6WYWbGTwTgPh2hjVCJqnFf
HXS3Js4Gklc2EyF6bwWRLQW+3wyK/DIhC23oCu2aelp5fH8VKZH3ckQIC9SKfkzz
r/xjhAw/xqTm615ZOxa/4n9MmbvoMlL+livg4xIJEIHkokLsy67NRB/SUXegSVBb
QMWDnIGOVwKmq8fEVNJenKq3lPeXv7pYJw2VjAAOIdIB+uXWEaPOp7AOo5r+Tg71
9VdR5naMUJF0ooV4zmCREnJcV/Yg2GbCaQa8Xb8T7VjHRV2J7Wngs7tOlYRwui//
e80Bb7Vn49O3tuKUSzKD7foCxZuoK0xmBjHKbP3GE+7qaGsNy9cnS6OpGNUSKYgK
HP7HZwb9JwEFpVTlDvD7EkEdsJZHNAui0iy/aGnHevecgHlQNno4IaybQYow19bM
tOL5wC5yYQPGoL6EoGcdfzThc3ixrjhUO9EBU3KwaJ+vVBFAnr+XlAt8SVG2ec0B
X2G+5ddJG3blC8H8tSWIsh9CEX4G/DMKxZcXid0pQPJXcrwy9AZh/HQ4oJpZj9rE
HYGo1MHSv7Xih2BuZWnlCZi/9HmwOggxKnPDOfGiL8Yg/qpI8+SCs5BAfXGOIm0V
rlECgL4Hz0Zm12+FLB8UodZRWVV/crVP1UqSsqzzpqIG+U0z2MVJTTGsgqB9NVI5
5iUoj+9PRNkb3Rm3HrrXbCPEE2OQB9h4fkWH17GdWQedB+7jtPBStpElWq6/8LtO
Y98ZzNS0xN3wDfJ95JTx7lqe0m4zZqSAVI4NTf54rhUGx6gjLQuvEbxnD2DlB+8/
F4ictWJdNmnTjpCNZCVeO0UuEMKfkJf2pDxDuhim7AVdGhD8uZCCC7FzEuj+G4rH
ykh/tYkuvNb1PcjRg/gXn2Eicw7nkSHyPuuXOObYPogg+gzpCZ5BzYoEHpspaM04
291+KZlLpfWyOjyGSTu1j6ml23odnJhjmADh1RZe/n+nLj7U2O/Z/36k7wb2e2st
lDjJa5mX/FSJHEWVPO0Hl0KiUmFlQYgSSd3wjBsOl+7sOioJ5F/PlBrgV0/rUhs5
wAhC56D4CsQROiYZqidvu+70Sj+i91z5iqJUPyemV9+cM7V9uVBbsETD2Hmhh8ZZ
aOEWZYA6dXRP8E8ARYbnKDPmS4EuSbwBFs4dAjZ3J1MAU8aDf89/be+T+aIpx58A
eBjCZYDkosc8A08VmRqZ4zAYZo+6YQCt3j7B0M5vKOlsXTGqVW99HCQWNJlA3vRJ
vKVng78X7TRwucRB2t4HsQBS4mG7dUlQjb8BjfRv6S/cSi4U6bdBLGqJiaM886fD
p9TmhMfBCRcnmzreGhQjl8mCp9inGEP365S7A67xe0PWOBZZXjwxYmU0IaUJNvK1
nU/kgz+xyvhq4lzgjAvx/2aqhw2xupp2zmR6RMIa2cT61fUm9RqKzwDgqNbi5osQ
zYomEqEpi2ifG1aeTl5ibXyvlu8ha41eu6Hsne9/8fWREzncpAf6okn4FPLyfU2Y
a8G08U+9spYO4P/su+JqJRi9lxe3y5De7g+CqDPveCHHL+VKDqMw6WPfV4+e12Ty
5Z/m7Bs6mB2B0OmTMoDEuB0Lwt2F1mDut4WXzsiL3Ciav1yZnQKAacaA9YGjD0u5
Opfp3yRWF2myCov1h3mFYejadq8n+lrXkcnIzp8LGNDzM6uS0xp9E9/8GQLq6GWC
F7REx6tAsYNnTM9peC21KkCvsGwpICEBgflFE+jH5R052abmiBCK7CXqhLqp8Rdk
v/G92sPeoA/v6A6OFaRAj5ELa/YZEsnq5mu+JZyH20JSRF1kLR/5ZU2bTf2KCup1
dhtak0FXszurzi3kt1kLkkn/WTV2wSHN3aWz2Hf8JcNty2/50/o+XfAFRBS6WFRK
/jdMiezFutNE6+SfXcnoIt/+EnyLB21qlTC4n//NPUU6GXo+nhm88kLtjmCyA/mT
zesgJ7TY8tVVx6xuzKVuf6l5YFuPPx58IlDyBKHCMUL7e7CPuKJhbERH/Fd6+Dt4
ogmQDv9jJIIB9PwsW2eEaqCPskpbsPkiw52Jgh3GyP1hIioBo2zQ8Lmk6pS4LiEg
cciw9rRO5r5pPh7SZYTdtq11dbYgY3fQTgL2g9s9TN5CpchgP3ObLA3B/6P1N7YQ
R170vduEqVJYo3EesSNUv/lghBhFBzrng1SrEkpJAKh5S701IWC3ufHATVb8qpHT
W523HMxBbpM1pbzj9cqcQydEACSDwq35FZrciWmlUeCvKdw4SLPQxCbGqQwHhVMu
0h4MpkHs1qMdSe1JU1qt5upMyLM/KBOUapO4wBWQTQsN07oVU6KaW4QYc0QVPD9+
CmnP3Ngc+2TABenutA+Uk3ps/o9gAB0vZoRWXNo832L6TjI0BJ4qGaiTezMXBmjP
Jq1BR2LzvLuzRLFQlJXw+jXmLP3sYA8QCGZwJej8MUaNYZS4kBZN1rXzq6vDZG16
5KwEC7yVlOfxBnLzUcH7G0XNrfjd1ssHR5GXfbhdHLP3fSmUDuSNsthnAUHpaMeW
zlIip6TwJuilbfUsc35KTZ1jdpsInRvdG+3+FbfncqOx7YPFrPUyv28z6TKCYjWw
jT1G7JlJu0dIP0BgV8Fq4dEKGwUBbq95KCstKS2Xpo61YEhanWRbhqRc3bDdMoHw
QdMZFT6iED1i8vku/bF9MmdEQ86HmZf4Pbx+IbLzzz+45WoVHdQ/fs51kkDvjtcV
UJ6JYjV5P3vMEi7ZVMJavNp2NJk4MQuNWENaiiom8ku7HCwEQvl47Fnzr/ilTxnf
E44LXpMQGKpyXEol2t5rfX8hQB+REP7PZ4Z764u6kcFaCma/qg36RQ+lBuRastDl
o3QNNN8+5s/FiQNHhnKSANTRnw1H0tNB86L12jamaT0nNE8yIMfJ9f92f61U3v1k
RMElN7v/aYWF8J27v8cybI6JiZNhKgz9el+M2ia9+IOsgr4CM8KEnkahfTNvh+Ov
sOsBVMHdNaYIOEGwCFogl6pB5+E+0iZSMi1ZStU06fRba6TheR2Y3TL3ExEE3lwl
zBv7a1eHW67RQzZ8o2ae0Oq1lelMa9DLZ9rYEXDbFJTfK3lpJfszt/o3bJdulEVU
0jfIDbqaFUzq7GWkf1V7YVDVZNo0YZcZwgz9YqWxZa+cZtBOzv6dT9hFsOhQ34K1
9E4eshHuaObF+hVumvbekX/uuIeT6HNCYyhb8lpPWw1BwHqiTc4ftowAYXX3BPMa
m2gmcfHaeZbGhsyifd7jMVX5Zk8BEtxxtUC7UDrPOqbn92Adb1myxgOANXZKFrTg
tfckkdcY9ZPkb1oVUVXL5ky2AT2kt76HRhnezpi60Oj8hrTe3UgukXquE9LOzwOv
w5bcJnISRlnk9ZHjV87wUw3ofJODzvxSV39AaUcFDiuGnva7WWvOtukoy314kvFv
Rgqda2N23mO9vMuEeVEsFXktPolJugORgOCLgzp4wuClUwaYUt52uOTbPEMxtGPh
H27td0M2BvmfG+JajR8DUSiMf5W+22iuW872feQ36YBZbdaG2R1paFp+2iVO7qOS
nCG+JgPzVoCzzqMi40yWqeuFe4tABuLm3eHA57gcgaofnODiIRCo5iGyNC+JGeVj
VetkkHDpiJYlGO6VihxDQuapqPP6vC1ADtsVKUeCUS1ig8aBePoytZRXJu/6g7SQ
7F7M3z6ZpTs4odtw4U8KEZ6nD6LEVnhfd4ns+UG4q9EU2JW3I/cK6eyQ2qaVpZqK
ZiwR1yepjsK2St5zdPTY3h+wd277tbGn3YwdBqcnlu/LXgX8YIokAWvPj4HojeKO
X79S5WxRgnq22lW+nAdxOqc5375nHPkAHlEnMAq00ONU2VUzXaJbPwTsPmvLpCEn
Tg3RjXHIOiD0/8Z4sdVztfzZ2ucs/nBY6ul88Io3WtsvkbmgC1AQ6ahVfs0VQUyW
QZuU7ysMVXEDp62nf3HjaQH4NApku99r/cVC6e3Vzvqs5ODYbi7yuWUhyvAw5xlU
rV8rmW/fsTKxc0gRO+dgre+1fVE0aXWtMVcaGoak3KBP9R+eR7oAI5vWlbUuKQVC
A68HP/ghLxBtKHP7sJeQe4ZmP35dGl2U7OHG7eTTq+aioGqwDso1n/cFOL00O5jN
u92Z8JFBGFWuaMDLPgaQPqUcciXYsJH0OinWGhb3PVV8dkeCBqn43JglkTbHqevp
XW8qPF0q4Ctb7gRGJtTu07dkaPEBYoJPNbEYuKqxcTmUaR1hxXUFnj1CNtZGUDYl
yOazGiogceRQ+u3TOTpNbOj/t2SM8vNzm56+mbir8I6HJZHYU3NC02e8cmsuSvSx
PDnLQOCxLdHNEJ/TU9wY13LbFMF9j6zZWlBA7mZ8FAOdv0AQ6AtIkjjB7KWHjk3r
DpgkToYR0OYO0CxmEX34lVcfadQbltwFNWdCMeKjEpxSDxcHljk44GPVB7OsHbhC
FaH6p3eid26qAmXvoWY/EsBzkkqqODdItT/ScrMT5OJaAQsZayp3UbSKvFysheAn
t8i71lX0Ag4aGaUWsZuhHJDZKR5xLd3HhS26u3j293aANiqPB5e+DVBHq2+zJF4D
56XQFRs2deghRatD7/UtgTtYYhHY/DArghrci0aV+f2AO1zt5Yh6IyjTffwsUahw
P4eIr0cXa8UcIUubDocak2NfH+DV2gTwpPKCueFe+J+KD9gM0ms0enXKRvnz5vil
vqj5hLydpIhOpBtHyRGVePC1+HnXkB5FnvQa8EWBg6QAMDz9xwMMNRSif+6DX+/W
ugs7NcmXDMHMNPYcz2nirD696Xmh5I7cYKAMEBGzXvMikEGU69blAiT7Rwg55xC6
/LsACWZIdNUhvb/CFqxNSqKmsRrlZw7p5IinKK+BcaCa/cKARvITIn0qbmP0sZSh
Jxrcodq8AiGj7HdVCmlgbVm7+1FG09qhlK2PqLqsSAArjMuMfP88K2HIDsFRdDcK
V7Ea2/eDTicQ/6WSbOwWnz1TDUc9PD9c06lhaYnALnMu7YkwobcBvFRYmL0Bbs9g
DnN9uQQX3ivmUslibe0Ox6t9GkFJyWwl16IwB2yRgVyuDUTj04oWBSSZODcbSo02
28PCMbxome4Hvjwp+Tra0H/g0W+NE5FoQL+lC7U8SOuGDxwYpu/FX/rKazNZK7JM
L0/rWXqXgb5l0rBW7aeGTHLwtEKwgNHXAT6XZ7jvQQiN5dQnHX9LKdXnx8bS2/65
uDKSqq812lFyGnElfGsPQ73BRYN3xkkHolHht2fiIJ/gnIBl3XqnnHBk0PI6rmf8
+fvlmGtO37mVnnl2be+iI0ZhGrcgscFARj/GnilwO9szCkOw6RcE9hlf1DqESpAq
6m6xJXRvnSYkX2zs32NWw7mZj6n+A4+AW+uq/GX4hTlLTV8wZ5JsQaojAOv8mO44
ORU0sBatqstVkNUyNzwyuTaJwNL3MUbGkKowgOK47oXzJ/6diJT4F2EonxbDi9V2
D7BY0FlktIdZgSIuCusqkJIGyg4lX39s5hioXQyuK2qTAKKwhqxRCPSHEdIXWYVv
ME3BEa1+kJ3zJDp1X4cIgZEFRGEbuU5GqCxr7ZDmTmOc0q96JmZ9ukDGrvBDB7vV
HHMjtB9YW60ghwxdY0k0TzebjC1M8buCc0xGwSo9BXoRIhtcpZJsRJw/oTesizQd
6ePvHpeZyD//oZojxoUZ7A4cQVQReV9HeIV0NdNdb2rHWShGcG8GSmF7oEJ0pr/K
jE4alP3RxTdxQWC4HMBHPlw5bKILVZxVf9B10w7FK0G5VT1uDYj1zr2l4hX9up/g
obPODwSHG/5h2N0UlcdIrr+VYLDSQunSU7Hoa6hhqSj3AO3kJaczNgRsw1aqKoNl
oRf2U29I7d5NR8KWS1nx1U5OBjtqdAJVbGxmVNDPTIpmcgLX9LnS3d31Ryr3ljZw
O7HxqMK7CNPigBblY+SbwK46doSbw7sZo4Fv41BKzq2pCRImqyt7NreccjaB2z67
geLcfMQcJZpkIAhZCTR7Yxh0D8PoiTQdcS03Nc7qa7pWEqwZJz78HKsCawy6CqtO
GZqPEIiNSulneaXMOs1Qz7Mv2w5tbSQFx+ngre+UDaCn8UA50Y1qtmIizNIg62gX
ODp0ahrj6sQJklrkbbrpaYDe3bEXUhIlO41EI2KPrHwi7XtB6ujuFaAYm7+j1FYI
ZSijviEO0u9rkuaXkzQ2rrNlD1l9CL0satYBRgBJyIh7PKm2IZDEBwlMapMHKyHn
hVw5ASSZaUdV34cYBxgEfm6H6k2aLsyg1LAZrcnjB/jEGW/N1c/q3fG/KQNzIhFE
A4OkB5hR2ZuSRn/5eE0My/fQFMzF0qNm9ni4S5ZTWYz7AcywEz4dkv4Y5+Z03pRx
Qga+H/B4HrF3GtpuUN6Os8UypQzAPwijp7C+psmedh8KAQbtvAKiWh3oSvg8sCPG
8IaP0UnwA9IpnuTZa4W/zn20RHN+0gnQlgdpQDgVYf2aSopjNJjB2kGCCNiP7efr
Ub8W6uqHMxlaOISvl6ZShqBirsikTpq5XYeJiA00MVxZQDibMw/aGrnQV6cKNAEq
NvPHMd9osXJIu058MAC8v+kb3FJsoE8XhtGK5ZCZSoVAQUDS+1OqRDaCaVghWPb0
A9avjKgG9UQi4AwlLe3XSfRBle0LLDG9VLv0KmOfztzY/9LftuDDFVtV8ALx1cMJ
MalfVme8rUdS0t72bATZjpvYmkbCvrfziRXWIMsqpb1FIP9WPfJ0HcbvC6Es0kpN
7Hc8Hisan26c4Gnbh733lkaqlN1Qe9+tUIgnbuTWOdeLg1xMFw96m7O0qzuQV6oC
2nw4kU4Ytrznbp+l/VN0yZmu+CBZXCshCon9/jXgkhOMHn3iCynViqFXupWfQGcq
Y2YA8xBv+CuuVy69zGmTszqz/M95cUU0C/wvXQyOt91mtCc1yfR9p9T+cG+/r6Qe
zQ2OPXYTd4oc6ppS9LxZlnSoCQ8IRABGGsn1JRkDKLmS/JzcxPLy3llwzW6wLQ6I
/pZxX5ugjlrovT5LV3stPmygacLbwiuGlmK2Jg02DqDJ8GKz89ELjkHe3jkfHywy
OCIcmZjZM1sNfIHTbyNH12Y1hKBRmYEemeM0Ei6s8sV4NbQQjlPKejb9TviP6DU5
GxrNXXIdOa+zVSpZqrY/hgfX1PsbLIDG4OK/QAcRVubLsCUboPVwFLi29ZyN3LTM
+cCsZYfcsgH/iyTAZqMysjYYMZwxpgXo2eKudccWFldpOlNs0KYfIqrv6JnMGSs+
ykNkJiyhdrBANojGqxsUbQ/4nMJwEYjtqHlezxH44ga8o0kwLM0EOs97Xy73EGLq
hqYHVDDOOJ26K1uqkGKS0UI2rkhjlNAoFp1nbZvC5k7FzmVwhgdCDa4ZsiJPQqdI
c6tZxNWga/+FpsAA4Zap4PhtiKNdyYS7Bs/PRsrRjIuM1jAyGzxE9uoCy+CxDWfY
cPTh494iiSiKzuBPzvwnHjTfeJ0LV3sPzM7TBsuVh/+MFVK7npPnhAC+x3IW+MB4
Zcmxs+IgfKSB46SKXKgnCOSYL3cbslIWtWOBNOdBbOYNaXh1/+n2wlhx2a70QQbo
rN/caRXOgifZx1ti2mMcyXN4pCKr88jPyhohemqvUjAw0ADAeHXL6IQNkzyGC4gp
Aj45XvHYRtfsOBjBIxYAOZ5TGJyZShykVbJntenhlCwAwPhI5pPTq2U0RhwfRUSS
PlGbF1qo3oiqAGWlWRpSFul+s78+1gqbuy0jEiubDWSDSm7CPvmHym07+/1GBL8i
Nx/nUQQ6us/VV4Ai5HPt1wgMywaKw89IJDfkD3227cTpCUjzKMdOZcwGvsflGNog
e6/SURfzGu6QMiCyfVpzXfKN6bmdRGUPLeobdfdKU3/YmY9Fxl+EvDFZneiFDLIU
5CLveKVzHynO8imOrPg5YiEYJ9J1m29y0kBWHo4y1Ta5Q1if7VE2nmh/knXGmGoQ
6XnEYmKDb8nxIjuhuZFQoOSwJDmXhxvyik5gqwPGLpU/eh9pDBKoJk0n4lEPNbHm
avsn5gJ5nmaiw6CdfvGHEooYBzMF2w+d1Do9aylRG6lwSE4S9ePDdGBXsHu0dNXo
7c2VSDZw1jV7yZblRjLqgpW5bkeaAaAj8N+fk+orKc4ijIu1tpXzlnyH0onDXAUx
mi/K4+yQbkblF0NjrbB5fHEDyK5D9nCmFmtyVo6PwFY2mBuPgJLES+Du4RzySGTf
zw71tH9ePfVGUT+q0gJuepzo2NERH0FUMBs2Mchm8BiT2UvrgiuOcj5pkOwL/RDu
immkUMMGElImoRblvr7x6yQc8+H8gKrbE9GEglOaYULtZvr+0Jvdt3Ax1eb+cipd
zKFQtNFUxJdhqfejlshExvOiQN3bvprTe1tKHKDTAU0rQ5xhMZzynzgN8Xj6hAiZ
g2pSwmVwZDKOhP7zbPFyvBZ64WDO5Ikif1mOrvZjo2onbv35RpExUff9vIgjAffl
ymQXujEO4cjXD4gk3dSiKRmdrpEE6OiNJZNegj2IWA96vw0x+QI+ZvvMRIJtg/iI
NEtarbnotind4lIFqAfX4IEUaL2rykwFs4KW0troHwEcgMY2fmvo7IqX/kQHtXqr
hwcfmdVKwd9uR/qvgEaWwjNnepAsvK3Dh9i2P2xzL3YZcRyY2iuu/Se0SpH1nv0n
5QwatlsdeC0Du0CRdE+4cqhhgSDoC/xm9uGLAaFFf1C1/v69f/g68QZEyAGCt6NS
cHBlgVaC4CxfkV1asyLaFbklB5zfMgLic14PNdDwBAk4/jfzzntDQ7ZkqrTs49AR
E4eSDk74aYLCSTy0546p5R1wqJ828VMP1R95plHCAQsBTrYsVpaN41jn9kweL/Fn
gugmM1vpwM2aIwfosmt/huABi9XPEUSos62Phs5NFzDuSxuLEInHmfmRcq1PhB85
DxPP++wTuCOrgiEB4JfaBYnNrr6TVFzHOF2oUTfJHlk3adM7sOAEtkHO0AMidX/U
cAogR5fHoVXq4v1kiScPY9bXtHEczq7iPwBhqvQ9aVOuCNyDUqAmJl/YETl7OzdE
/vaeSjEs8ADVPYepCSpeih7Vvljv9pRc6bw0+5vrPhDcDfoVCIwO6JEa4hDvWRws
TDJMjc4pI8+b6b04wp0juSZAnRCevc6RXOCWk1P/cH0SRQqIjuysV0knUbW3qz61
wHaad2Ouu95mzOjhGGiKF5sf452HRRBvbOSefIU64mQM9UxezE3XHc4Kswn7y1/B
RRivRR7biB7fkdF4KE5KsX5bb3briDf4yFz7lDsm6ylFvukHQiZyqMERudRezKAm
1yRInmBhM9672v29n840ZQWTZz0DDk4l5FoizNbUzbfgwS4P50c+dvFfu02uQh4Y
3BJWAWh0a2kBI7e8cazQmwJfYDc5flmzf82DS3OyHSTkOfAcIY79FKdwoNIGQrAX
6nVH6QrYgIPRKjtMR3tBymetV9KnWAx6B8VPld45vY27S53Dgwu1wTEFBmg0H1Tk
ahW/+P/8RkZcMJIcjj+sqetNE+F99Yhqa1lEkBaO0oo2ZfnNTdyWX37C7Ljim5p7
Gfj2MRubPEAorFaJ85d6N00qj+WnO1RWPXi4M2pBaOheNgx69TwKNq8KVHBsoRer
/3Cp6xG1NF4scrfUhdT9ISI0n+X6AVa8GmCbqUann8shU9Ssm3TLK/3rKPAK7Div
Ybu9TaGW3yDxkmOsKmKBln0ptVP834Xtbrs22Qg93DINRlyWUU76DpXO4XTJdoAl
Nnd8W+ti1G6GFNQdk484QPfWZ6iPmkX8Qt66QTFRW73QzsaZQpbnoO7RmX2FUIHU
e5k71D+h8Hxhv4Y3oqTr0BlhebyCLQ0M9zW2b6UpS8vZiJ2e95pnRXrMWEEUYIcY
d52PwqxEymU0OJFl55gz0H8rGJPxh04Yg2oAv2kOBVcodqojcEcZSYojr0Sevfqy
GbMtTwi92mxwa/KxpTk2e3OJ1gDKF+tACEaik9/4vbl3KP6yCETcWiaV48VLu4b+
JsJANfeNg5sWxu/fW9QQ//Xs+fr9j0ycLWkM6/eJh2iXrHayzqeAax18DhmQQU/O
wTq/qcv3gN0Z6jwsay4k84AAsTiawZszolo1/3HaXXcTHsu8CqIyOqjaUcdy9b7n
VBDVb6/d0eLQDNbYxcjli2BivyYN72T0XdmaBdxeCjovtl/7k4lMOXDijTx7GY5u
hk4DJtJ2AEjHPP4Y8YFgVx+wEkhl42M5uNBlGCnPmUg/+kgxk4Ivh0GvhwGpHf4h
DBkyUFXSKCnHL5N+e+AS8TGHBT4CHIbdwVBODlYFdKjoiX5G2iMWDF0d/aFFxQKb
SqcK2LgTQuDf3LbwdqEPqd+SOW9+9R0yH0WrVbmbbfHTA5DgWAQyl7NuKNLP2YQL
DK1tnZzkZ3L3zrmc+seOxe/JTtnSP+D0Dtj+kNErwvJVr0M0RaagjiYBAeoSCeTm
RVdYh/VQTcuiURzE05yzlvvDLkSgjRaTY5ESxnS/NxYYVL8UakCyD1vtJfDrnqX5
rEEWyWTZBsoix3HMzHJYgbi1yRhJJgN8x3wQqq7qrCGpRLzdh8BPG0OUF9n/sUOU
DOTfpPxtX5FXwHwktNa8MuH3kAQZNIpITWOEiXBiiZhy2QvCFf6eeHlM88AWK2lM
y7tO8g641avhg2lpXkilDqmp4tc/9+s5uaxBGlHK2B3qLtMzbIqTstfUfvI24obX
QeArQo4rsNSqorZEYIQl3YBnUbV26nkq0yyr2T3p2TEjeP+qIWperARP8oGvSwoz
b5OOok4fQOgt/P/THAiP8q9qL5dBeQ7R5qvPkgFvqYCjPPTCuNLcWmHpStiGnj/h
MDZpbsSi6ATAX3bSiWEt8i26hZ38nr05I94p8Z3ktTy/n/OgLlIFqjYHaTCOPf3A
L+KlGdt/K4PPPLfgzbF8p6TzGYrF+Mk8HeUAXdMORdULhkXZp+ImblL1ANriLH/v
xwYvcVLrEHqgvfT/yEyOaVDXc4PEJ6Yz3zY0bl5eRfJm7rbQdGOkXORY6vand248
qzaSNoT0HU60vPk1m/LzFEr2MT0MoE5MZquTaCbf/EpuyHe1Hc3m1OpqvULIm+KG
Y5qEYirJ6IOAmHiR08J6ni2xiCNrZ+NhUM4f1dmKYUStdkpzR2ZcJHPBFecjptCM
slzXocZnoOvFoaHWfVQ2Atjq1sKq7ZHTSLyZjOad+p2hI4UrUk+nG8Up8gOTpmiL
HuZeMBagPb6UmKtOZ8zdpiKHs+pH9gzG/CDXSu/HqrwBGRmJYbNRypxdKJrhqfDt
RPBF3OTHdNsej0NK9UPKvv7OQ9D/IvXyAg20esJ5fw+c9BpJ7eHpYuOar/r/3G/q
EQp0ee4+IzOxLfeqiuHhI4omnsm0aTjLWYCyvz7d5m+DqOESJi0RUL3tjUQtxLXo
mCvRlHGg8t35D3Kg+wTC9kudEEnIBGmzztVMLf3lc5R9Ax5ujOstJr4yBs2PEk/C
PwhL1eEZUjAAI6DMYfuJijYKeiKVxlL/IpCynWyhTHcDNUGWPyGbipGJ92aCZCm2
ayLSPMgYc4rjpRdL/bXAzJd4kiyC7/j3j6K8q8T6Yz9BPuvsZgS3yEgUeAvsah6u
U++jhvJWvJdNT2DIntuWKSU5uQy7fE40RNkPvaDA0T3o7mTvDY/dZIhyUIWpXbBi
nX06x4wRS246Ab7DMMG7fWVNJKn2G2VCp/Vsqdp/uVHoYGbNWBZklB0wbfCJDFVn
/0SIWG6jrdpO8zrExIjeWCN5lqEvMkr8p6R5NKNvDk5OGd9fa9oi4L2L40J9Nlpg
k7FU3W+iowtXrk0tJIHJu+z4S+Hb5Sk3W1fVVjU9Y0xQVKODgQh3904aoBbylFwT
0OfXm3vctLODD6/vGhA+yaUD1a69/2wEsRvfMM3+CdIXGB570bY6Cm3RuzG9821b
6JYOQLb69lblYOFFZy0ENxkmIgh9MWfiDN9ichP82VyFwnGvHldb+O3s78sfjLvU
kBRZHqfNDHwQc6VH3KAmffVmviTUMfDcS0omtIeGTgM66XgSDWE9eYmPzP1NtULq
TGNHOf4hfjxRj0JaZG1C56iSX5DZuqIaai898Yby3k31ITvVOMhaZGTlC/6WJFi8
BKjbV0gWWsZui5CaT392QX8DkYnoHpcVoEf3WfGBRLcE488KrKv3YBTdoJKbikSl
WRdqhcMTrVrFWChUKl/wshS9S7FET43kRLpGCqyysBt0h8sQ45e2l99t9Yi8oiAo
2o3FiP4xreD7RY6XXN+jq0k+2rMk8OEafRt7xWlFjJhEeanVmyZoiEUinO+Cfoc/
STDpXRJhUqsXv/6JXwlQcA7pMGO9WkVf8mwUR/gQMKMovicTQy+6+KJ11iUlwWeX
hc/mz2pUlhnvPttlhZi8sfxmUz5UsbR4qnt61zq9grXSlXnJcXJS6TlyzmMDfIV0
YBMpXzAc5QWsawaDgpdS4B3MyTOPciBz8zLxcUYEG4k2SphYwmIEPFZ2YPfUqhUX
GvNcreha1ENZQ2dRrXI7EPRv3UFuehiPxszd8zGAIJrPvFEcubKsk0l4pxIzqbBi
Rdk5P1V3q2gVbPdGhjn45TscaQUD3LM/p4IEWuneam/G31uDkgXbPPZ4Rc7VgKVh
1gWYpNI6WV52o08TGHu0Mz2QtA/oQhBDk53m8c6sXgC6InvlA87QL0sb0Oo973wI
uD2sKeMRuNIaGIR/x90HEkDZ4K7M4q2mYDst1V2rHFwiz3t5pQmQZIRVfZ8YjOiM
nJwcWT+GqEMLTorTG1VamJySH0aG1TSzOHAc8OkYEGwlphZmtygx+ZlqL4cNFv4c
KCZfcjYmxboudFHxjOOa8I5gZlYsaG/NVwvBjzf7UaC/FybAqZEPbRRmmsjyzYL5
L67JL0NyLHqX9/wCapbfopcixBBYc+BZeygfz0TvnBWAnqWbjNUqSNn7h6ubXDmY
1HYF3sCOhIdRf0tQGYI/KV01KTJAmiSdqRd4oBaWZgBQWwyOj2pm3PocjbCweSQT
Ob7T2a3rXZ9kbnT4JhT5oUn0L0MEBWtHujb7hCb4TkXCMh78B54ZzuScnqLriRw0
Ojc08UJjDqcTtOdiPfkK6hhs5rtw/BsMYVB659QKLO60g4wVds9U6EzEDb7QDq4U
VVKPxMXZa7Utu+8cmH1gFinFd8SepbpN2n0qr/GURGnoZXh64+d1BzpqOOL1yvJ7
QqKnhjVKHN54SkBqwnfY8O+Y3fh+Ca6HxeoOn99/j2Fx0BiNCzEAfBSklHiBPf7y
VIDp3gWf1cj4VNthOQb3tNEUQe6lLGePeC1pssgGq8BwrnIrhazFIsh5WhIEuhj4
5ia5b966gqyYpc19KCUhrpqPifKI5NMgot96uFkf8TcjIFo/+wbZ9JCuDv1jfe3z
0U7Z6bwlnFB13gW5wydKD7b3qJ3gL+QXjevrf666IHh8rAv76M7kiBWSrc19XEGa
Jia6X3c6GAaZ+L6BnqfbvBDU1s3g6Sx3z8pu/T5BZxpMR5wKXdolnZmfWEECNlAU
3OumdIc74wzxCJdPlPebF/2beXagXtDPENibEhYdWgzI3OaZL57ZGZACtHg0e7iO
ikTxVVAxMEJg1QNFyjX0c7nly2TZ2MuvwP85b2gaRLxqPKralHZ0QP9oi+8tkchP
8OKVe5PqZYpPBiDpNiolCMWBYLoITQWdZWsSGtqcApdisc5BG1u0l/u2QDXFJuAm
6JuZ1aB2nc7SwEiF57TevfSnTqRyL/63ndvtzXXw1mRVvH+ziDtfdye4WWCbYqND
ucdJmZXtx6yUKFzbnfijRtLK0hnTH82xUwa+hyqDxwqt394IH6fgYdsbTqdOCp8U
CuJMZIBeopHht05sznQskzxfxR7hyO4lE+w6kJCLfKYVyvvuoiEQKR/kUlIpb8xi
sYFrroK7DGPHulBaBXPTAAdTICwcKbSpgr3DXGrNBG4NgaiKkCdB5Ik6dqASyY3N
LTJQBWZ7B/2wGYKnHd2ApSTsEtijF2RqArFiQnhPPQvsd4gY+hvH2Nva7wQwiivi
Exq1l408CauyxpGvgqW7/hQM+OtcBJGYaKNRVc4z6PckuPYVUJuSPMxw1bQMqGtj
amQpanXswnbdj7MvTaqtZ5IEnk7V/SnaAHWPZwx4xtrwnYo3xXtc9x45U6rgUeu+
bnouhtko5xM5Y39FO4wPj2F9mdVXtZQoI1LsRIJDrDlJ050GeE3zawEmYCPBtEFm
c9LvdwIWURepKk5nmW9BeMby36dXLI9ftMU+1YWJdw3C7C35S4vo1LyknBmFjSu7
1YpKLWsT9VMsfG5hYGIT8FgBZGckNsjqLABmMBPbuF4LxIbLU60pz3jSOekKJhY7
BE2VU+ORWAhCFPr+OaJVMnyXb+cjTzEoZBzrcQizBK318/pBWfktayv0aBhN4xoh
Zwc042YWAUO25L2+Hw1+56mwnZ/aa07yhP/SC9sfsdd5UskrwxwXb9a8oNRUVpWd
kTQLr8LCzcRwxemwYT5iPmNUvAY1teLtpH0cJHx/9kC6kCy19vUOuA57vcYP2OG+
oXUUQUisqSQyhaLTncPPbBaDD/HMFxdzMsTIlVFviKBlGC1cB3KG6SSSKZWkj6Y1
rgL31a/FKxT5IIQk79v6IBdBPJRMKn9/JBrahsZUNhsnLXrV9+MAWMMMDKLx07N0
56oL25Nd0kbyekHbzd0wVkWfcshXPNvpZ0jkKUAaPAsFbhrqtA8BYu5zc14rSljl
swF8GBUFuc0dyPQImE+jOxE+o+ngxg+oyTMCxFKl6vmZ4ehReJljfV7pd85b7sop
pW3KiwODfoYa4aaPsCSXmPxU3IyuwIKy+EUF3lIN5kEz9zw5L7c5AQGSJd+BAub7
0TNeGFLvy2nZZav+uJyCoaPrVrJqro32YUNE7NWbUbpkNjWeELifo1iGVg8PLMGi
wD2Q5XV11xGQQ0xIhhOOywe0y0LpiKlchQ1c+ZCgaTf10aOMhp53U3xR9XzdEbJp
5YdPHc8fSLFHHtck6IE7R7um1lV2Y9ngfv6gE0qBXsJowaYDpNJ1K3z2BPO1lQTp
nAncG3tAvFVKgjMIiV62RMLaoalMPAqkY3aAHiqEWGijSLop3ewKauA5W8iIZPKN
AS5t3HP3sKB1Y8QJTICF04TvuazdZKPmaU9R6Ecij3UTOCZMybMQZdPYGlZohnXH
5tFEtj9kkSqksO1RvBTF/fgDTFc2CytPl4YcgQTs2ek2gunrAmRIqmd3cr+bp70i
WLRHcJuhKLhjybW84CTKO1N+HJuLqfaIlrruymxh8kHDR7Xz1l+wUMGLhDsos0/R
H6R+2t2BAu5PyaDshVdJiFuMzJ04wqCp31DiAsHADrTKCqaTbfQ4vzqve2/9/HHI
Q7CikqQWjN33i+K1pGlKdisyDQ46F1JNLb2eA2d4CYDAY8AWoD0i/++mVpGcFptB
2hYb9qyX7WjpKXQBD/KbGbNE9QMcaV6Ll0bUanGxCjDzRjIb4dKbmy1S2FnvbSgX
IAzEu96bAwlJbnrJr9PYyKNC+yUgOEJzT2in22CprDoMithPLlAtoiyeLWiIufVs
sILId+bKuqsDtVYy/cFEw4fz8Dv9FMHLHCatb5HwakWwLmgYL3BIiZ8GCUB/32XY
1Nfe28+dJayf6LZ+LjMlOUAL/028HWXtViDiR/LoHnEHZbEsahU/XpNcO9zUftQQ
tE5F6EtjOaTOfHPEnsO908+K8qD1Ug/1Z1XHjNUXN1B+n8wPQE4e3t2N7gVZNs44
oCXGGlpDQBmrNQGZOvI8cq/CZ+SZ29q4kdTaVTv7O33JgVHhTysfGFZwjHoJZhX8
3JLQ0ykywVVq8Vf+or/SW77sQE9Hdp07akIaIWlwoYTWQ0z/QpTqWtFBpSzIxUsJ
KIOC8nN+53MeRQ2DxiGkcA9TVe41elGVURXt+yZ5peVzHyt1nNfCi6avPE2YC90k
iBFseuEsq+zsuc/XZdV5zCM1YLAK98aLv2RtkMJO4132pjwN+mtp7NgA2B+LYiNS
tzbcefgPJYkGAcLV/6g8MZALbYgONpONN1JvTHhI6UTDBxwoImdFLME82X7cAOuM
4j/NHRqFJI/LwmgfODjzbZZhEjmaiPPt9ZzOBOsji53W4W0ACWTuRX87PZzc2Rwx
opZjP4242d8KcaceYLEj/alyzCJ+Uo21ahiVLzq3rjcmgrZyofyECpDgzZQHDvdz
LSh3/rvr4LiWmz+ePlWykvRkht4B8LMfGxCc5Rit7fNz40efBWpeDC4La6bZ0Jnz
u+D2sl75yU8lYjkt0clbTQqEPyzKzsW73dIlSwOlqR97LSw7+JrTxWG1JdJpwe0m
bTdT+Ds6pqICI3tLWVlEAhNzpcMTbOfFVmGZ5kh9m2k=
`pragma protect end_protected
