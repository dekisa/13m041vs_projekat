��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P�d)(o�J���
$�P<:kh�㨁���2�[s�}���K7���[v{� ɛ�Ȕv��y9H^� �H�{#���ȥu�D�o�-ٛ �l���>�Z� �ev�#�NX}���eo�[n���s������i�&�4ca���|>�*���U����r���ۢ���7Ww�xjj�웦Y�V����yx5���bjQ�X�����!�l��w�SV0����Vi��"��g =���W@�E����g��T�E�gy}��Р:Œa�W�1q��|u���T�NCAE^|Q��l�z���L��a~\��8���+�;�ӇUaJ�a�#-������z�Yb\U�Q�1��Y���n����>jEV�0=�<�xCuu����绠T�:��Y�5F��.���$#Dgu�b%�9�����>N$���GJ��O9Ӣ�c�Y��9q��Qkkޥ���${���\sjג�`ȷ�	��bxE��kE�u���ɓ�5 m~Β�5�����
�Igۍ��@l?�Iy��*���Z�����лdAM�Sٿ��������gȉQ���aHu�AL��G �H"��#��0�n�z�2ƪp(Gq��%I�J"I�9��l�OR��>�y��p���$�nJ��Jh���ʂ���뮰������h���5*���8��t*���v���P��xI[��F|�
�<tM��;�m��mI�Y4Xs'x�uޮMd�o�Bm�<���D�viw��?h[��h9���D`&�B�=��`���Φ��x嚑�4󤓼��/�;���豏q��ja[K'O�_҉0MG�z��Һ=Ӗ�+��Ia�E@�z:|b�P�*`�y�(K��:���P�S�'�d���rQ�6��qj�Y��[֯����W|�����ь_'N��R�U���=-.���_������U�4�
8N�c�l|)s_�"F} x���u�$B�����H�'������Y�%���t���c��Ƃ�uַ��s�,q�N�׆2ӍĪ���uh���/A�7�$�J`���%�0��v|���������M�r{g���?VJc�w���`��_��ח���i���Z�)�5��H�!����u�i�b�J���x��z��iNP�����g��������%�B�<`d>@�5�S����Π����߭(ØO)��-�n�q��8�W\��^2�ڱ�QV��eH��v�zRz2I�MYA̤-���+~�Ʉۆ���c^XNk�A�*s��޼�-�`���o'�ox��� �=t�x<�2?x�O�ܥG���^:e�����;�F���ܡKE>B����
��(h�"/O��X�%��$\����s?u��b\��"f��3��F+��K�����5��2é-�ǥ ��%W��uC��<m���;�e�����]AT��)qi�2:r���#p�_+��� ��r�+�kһ�Op���(k,L�&K�̉'B;� �n(��+1&I����Lh�N��CC�J6.�������E�]����� ���I[���Ws��b�z	�d��P0)�C^b$����l������{�'"�S�ry��8��&*��3��YGZ�Q��0E|��:���2������].?�
�� T/xܲ��t0���&|�Qggp�Z៥����������Qڴ,�`�!n��M��0���"�;4�X�d�����Q���6�-���yk�����p�y�T�6��b5a�1d�d����an8�w���
8%��_��)��%V�����/�<�ϴh��NN���fz��3������Ť��5g�Qk ���1;M{�ɜ{3��D'�����i�4��99�D>'$'.��ո2�m��7X�r��`����r�m�B
4�c��v���I��s,��M��D�]F��ݹ!�3�_^�rN�W����[S0k�&��ݧR��&v���{E��2&�0ݤ]�a#N�y R�>� ���	7X��q{��X@9�oӇS�䙯�ZLㅟ'��m��1���K&��A���D	�_�)܅n����R"��dUW�_��m�JQ�IͅZ{��<Jg�X�o���s
ZI���'�� ��.XlS{;��I����!�,b��������Þ�'���y4Ѩ*���j��؞Ek�����D��]ʞ�^���(G���_�{���cmw�<H�J%C��B��,��D7Ν%�DF�}|f}���1�	rY�9���\^���V6+�/�u��!�"�rm�fp�ƞՠ�.r-v��A��n����{WX�����C�-��L.�����u�e �N����Y���|]5�ð� �s��e�������
����Iۘ��;�6�X2ͯ��4I��H��^(�C��=��N��?�Kqx�8(��
����� ���ߢ�{�+4���Y4�*q��V��k�[p�����(���LF&�;�kK���k5��l����ZwE�r�������޻��_ﴰ�T�G�a�%>:�m���Dhx�dD���Uuf�8�v8*�J]�d�t� �lᦥpl��[LN�V�Χc���4�x/�QrLj�B��kt���[c,Q���s	a_��1�H�N3��29��{����@<�b�X��e%v��BOjVeV{,��:��Ê�{B���\w�u���a��G�����;,´�UqX���H�v��|�}�[�Pв��"�z�#����A7c�@	�)��=���/گX+߸cubu�;Ue�i��;�H�I�e4��3��Rf��� jjo?
�1:7�=�w�z^��ߎc89�}���w��r����1H�8oE>i�����S�KB�xB�R��|����+"����	�jk~���w����c[Jh�i�"�>�\��ܓ�P���
|Fp:Qt�:\�Ԏ���B.e�u�� �25٤�M�qfw��Ҧ`���	5�|[�Q���>���Fv?t�JS�GU�����m,?�[�g7��;�¼��]�1��B9��,��TY��%M�J��(\��Wc�r�Z�C�&NG,�8�����{g����8��@fHL�gB�1#���E�E7�/�Pl*"�zq������ ��Q�y��Tb�~ļ��I߰%�HO1�iU>��N�� �lg�w�H {r <���^�>0��^�#k��GF�f�=�&�S+yǘS.���^=䄬�N��b�H��gU.�n��^w��RM5�f��#P�\^�H��~Ԥk|�k��(Z�ؗd������f�����T� ��aR��Lp!�����YU&�r�m�8�ll��sfV�mt�g�q���q��%���[7vl3��ѕi� �CzT�;? ꄞ7L�0���\[w!�T?[%t%��-o�沚(N��9dS*h�0���FkD�/��S���$�����?�eVq岼�ܰ��[C{���x��l�?�r�-��y``�2ݏ�������º^l*�����ِ:�Z��Ʋ�)2axl�sxͰ��� �U�s��W2G�V�X̏����n��!�K<vӮL�����C���O¹�"�9��Y�%T�nҭ���>�j%
k@7��<��aB�ܘ��bB���tp���k�D�h&q�#4r�"z�a
F�u�ӟ���G�,ˣ���.��."OwZ�n�%�/����$��xh׌�o/Ջ1z5�z⍳�n���bڐqN�jc6: ��D�V{��i���w�$W�v��j�7���y�&s����C��T��٨�$w$�o�҃�3Ŵ	��V�Z}�� �F1����K�2+sj��qo�g��e����9bV��Ô5Ft��'�Ab�X�\y�u�a��IM���-�z�*Hcӫ�H�Hㄝ�����wd�}�C:����a�i�r����H.�����tעƕ�_����!�a�����B �c�����>��vl�Bv�a�N��[����}�%*l>#	J����K����u��hN��~�b���%c�l��|�xr@稡3��w�3�664"�����U���`�b����I�ԄLg<�*�ƿ�H@|�� 0�J���d\� 4&bR��o��f����uݲi�b�+�
�e�����kF�BѠ� ���C�5�c����.�:���ԣ-�.˒(�gh�H15�4D}	d����V�Lϯy��0�9^3��JЃhC�a��6�D�]�����7�l����RZq`��p]�\L3�����.�6��T�T�BVǛD<�d&����*R��G����2�r���a�R�Q�R>۝]���A�U��y������Z�Qs�p��b��}�$��B�G3N�֜I]ڄ�D&�sgO���w  D� Z�F�G���[����fh��]�V��d�zEP�˔p�V]��I��������'�-����l �`%`�$�՘o�E3!,���cK�2�~Kg�v�#��<p�����h䕦���jY_�,,�8j$G�X����ڏ#�JW��%��eб��Zg��;�W��7)\�?GT�Dl���>Q-ƕ�Û��:ڂǼXŉ�:dY)����p����ha�z,���	�>��x;��9>� )ؑC�y��X�]��ue��G���b8,�T��!�xs���:h,�S����
yq�>�6���	T�� �'��O,"�u�/��]�����3!}�?Lc�}j_.��q-Et w��'�'Y�=���;��x�<-mX���8��.������������Z@w�&�^)�Q�ag���Z�0�Ӈ�?�H��bZ-f��tR�\�V�6��2 �q�
�g;͵߶�s�e�k`�{3\�*�8AV�ݕ@���S���ш�|�.��u5,ˏw�k�X_�=is�{"i�їDVN�O�sc���cx�o�~�PɍD+~B��EC���|(Yʲ{���]¸b>��Z�xR��-���	�M���߻.���#��mn{I>�u!}̑��"���[0N��y�3v]{S�X�B�@�i���V�9�B�'<%��I�J+e��n~�f��^��
��;��1���3>I;��o��)q\��G�`gO�SR0�w�@>RItwP�8�{�/�o��ٿ+WCш߁zt�4荃�C��j�}j�?%渱�����+a��H�]9������ǲ�<A@O�"�9�\�������xG��h�����ȃE���7��7��m��ԯ�;���ƃ�.EX�*�Zr1 ӥ(zZ�8q���Y�v�x]i��#��
��;���`��_bw<;m�E&�+����0\�[3�9���sH����u�;��78���|��e,�p-kfg��ӑ������޶4ʌ�����L��>uR���P��*ns�U�Q�Q�'6C�6��Պe0t"�*ٵ׃R�v��
 �Ꜯ�z��dSer�>�WS�+�ӱ� �l�f:�M���fU�A&��V�ǔ��I�ڔ%�/)��3M�g�zewO��k��+�.���ﭾc�q`� �¤������� =������V����̈=A�	�[������-RGC���l�������ޅz��r��kTjJ���p$Z�"Ǝ��F��Q(l�p�_�R�I���;DT�$��2:�	1"S_v��Eq�Q��,z�]�����-|�4��� �P�gg���y��3m"N\O�!s2O�!�@0p?�pj!�@ZK'Z��SЪﴴ5�YZ�d�0B�2T�dKJ��{²�זx_�7�Lf��EuV%�rmy|㖲��:����8{?�m@$Gb����N��yWnQ`�u�8���ڇ&d��! ���Єb^M��J�k�K0Sa�k��RU�b�|��oں���l:Di8���R���aV���{������m�}��:g����Z�TtB4ʨ�P���o���6�䉺t�Du�xXSZ�]~���Q(�d]���Z̺�
������'��8����ϱs�ʔ���F��B�!����9��Ȟx�C��;����zOD�]��:���,f�+?X�.��>�:/�{���Yx{�:'�۔�� 
�>J���:���h�u���$���^����H�R~�O��X�A��o�)��w�N�>Y��]ǧM�����\%�iU7	E���}�,b�Wc�V������f~�dP�GF��������9ʟ�P,���mv���������g�����t��s��m�-���)��ՓW�<��r���]�ݏ��˨O��_�*�
�q��޲n,�gH��6���<�0qZ/�����T�Ex�LyN_I�-[��2��)�n�Krx�� ������?����^��Z^��Z����K,�E֓����LSH��5���P�l{$��>�_2Z�L��ǯ��^+X���u^��j>2��9��k�R�D�Tm;��I��J������B@���ޙ~�Ew+k+��:������ڮRu��H�Ͳ<X�D�����9n��XC�o�΅=����x!)T�~x
M�j��k6���@��*�rb�����?�蚈_��� 8��¥��a���I�����{�S�?�_[��}̤CI���Q�0���/�H�
�_.]7������6�d�T���hX�Y�n�=����TӞ¹�s-��L<1dE=c	�#��>�vZQ�mZ���7 f������1�2�l���
�4���<�d�R�����6�sX�}{���,��� ���u�|��K�K�"7s�*��c�EB���g���@�	�ӂ.�B6��<6΁��~'�r|<.�s� �'��Tt�a��5\1�7�A(\�<_�	~�Fg�V'���RY�l��0 _�*Ij�x
N��^�v�I̱0N��Lо{�/GL�3�K�)���}j�I��[FI֛<��Kh�._3�CX�
�h\:��@6&d
�Oz �Op�9;3Zy���v&ct�:��wl���+���bo��~B�������rFIh0X�%m[Z�V��HF<���+1�)�dcX��U?~懱�]虪�s�����Y^��7��3������5��jn�Ԙ� &�����d�q��(�i|��MllJ�$��O]�a��z�Y�;8	@G��;�b�GC�d*ŵfǞ1�z��+O̺��,[؞�E�B�k�(���f������5	���h�n�Y���t�~�A>(�h�6b���_�B����L��U�z�8�]��r��-�}�i.�`�QD9\�q^�J4��~5�c2��K)�u��Dʱ���B�����`�q�t��4~%AD�&���?|zf���+%Ȋ�я�q^�B�Υ�fD���SGŷ�����p�B{��&�c���0Jtŵ�؃��;�����l���	\v|Q5\\$7�����ęVW8���h���+�qz����s�)_lމ�̳kX��z�"���2@e���\��b��$�b�{���¢[f.a��Oy�$<vL������bBy��Qަ�ZoKލ��d,�2�K�y|A�k�펯�M ������o$�m���5Ъ���$ '�i@�Ac7�p��e�n�D�:��w͢����������&��S���T2��b/�Pu ��j(_�2vM��܁[�Xa�����2�kWC��j&$�ד�ˠ���͊�����zI���d����/�ӛlu;�71�b��Ke}��P�
Qv�zv�����ʱ�I}�Os�FW�(�R�*���P�(^�C��>	����ܴ�XT��Y�[@E��if����Mmt7��4���+ϒ��{��EX�y��}��~1���1V`#��2�2V��������[~�؃�28��A=H:֌#ӀR"�	���R��&*����璊r_Z�][O�D,mN�GO��}x���teS�l1Ȥ-G���7x�
�ڈH-���xj� p� �;/a��ko� meg8M ����p�������.�*�3t|ס�C��5�j�7�^�u�T�䗂	 M�)��هUT�����2���=��=Qw���[��1a���+B�΂��v��/�lڏw��[�EI�m_�l����x��'���� "@v\�9�����u�x�T;7�l�X[�;�ۖ���	�zϱS#`�pAj2i��4NB�~�dH�2K��O�zUQW#uT�<���=FETmF|����c�Jk,�t��/Y,d���� �yAa١{���x&�ğ-Q���Wi��N�Y��%�%H����q�����U��&��S�V��ܑ&�ön��*#���.2$��0Н] 3��6���	�0(��e����˨e]&Ae͙cQQ����ï��&��tl�5UJT�7���=�>�����8ָN���%k�*{���u���X�]�k���ᷢ6\�ra����"C��f��z��~.�a�q�&�"�)G���RK.6IbjT@v��^&���YN����-F�`~y~T�	
��.��	d�g��5� A��a^:1�
R��F�E�ڙ@6h���PE����۱U��b����k��1�ȹ�8O_g:`DE����Y5� ��s��ݗ?Ƅ��C8{�)�[V��;$�̏��滝OAR��l���T�s���A����I�������GKO�t����s��uf̈���u԰:mQ�P�g��� �%�er�<ބ&b�޲c~�_L�nDG�P���n�tf/��P�G[�10�:e����e�;[,�.��44?<�x^e���"	�5 ���������4+�+�_��Gh�,"�{ōl��T��:�'uň�-+���sl�WI��m��K�S��g���_�P��/q�k�ˊ�gG��w����T���Ů�-LxZ)����5d��%� ��an$��{�;l0W�4l�D	���I�x�����)��v� �� sX�@^ʹ��]GW��,��������$�<5OM��W�5(.��{�ejv��� ���6�hIj"~,ֵ���\�1z���Mlk&��0�@�zcz.��K%S�l���-;����V�[m+�J�$!S5=�H-az���7u�r����w�ԿX��$����h�G��뷪��b~�_��j�����0�I}r����Ĳ���E)x*S"�����i�̀����ʿz8&�� G�M��&_a;$�m;b��K ���dج$�uk�����q�i��pj*�Ky��nn*f�O�6Fł-������Ath*ԓ[	̶Iv��~���vٕp1��b��}�<p�5�R~Y~���#�b}���V���!��t�HB��#z�Tt1n��e�����ڒe�ӝ�zB ���ĩ0�ǐ��J7vH�� �@M�̻7��cE@�G��U��˪^�9ɓ�g����Xz|v��������u��u�o]bw�����8`��54���#��B�^����k�L������h���D��k/�r{���E��'0��B�;��'6��	�(�f�y#x=���̯�9���WbIe���$fQw�H �.�a��W�t��&���6�M3]��b��y��h��)��m�hP�g���o�t�E� 1JOC��dE�p]
ڧ�#e���5pv/e=Ix�tj֎���ָ�l�e��][c�j���B�%�{�L��'%����Q�,!����#�5%�9x�=H���)_lp�I?�?�x���P�r&���F�o�q�#*CLb�ޕe�	
V�*��Q���� ��ۣPQV�%��z����Yőus���O��;��)?%kg������g�,/���T� �����{t:�/GFXkA��B��n�>��i�2
r6�t���'#6�:��]���b�GD���+��{�Ɋ���+�v��{+�9���j�I3NS�i39��B?�턌0Lٲ�zd�X逥P$.ш����`g�_;l�ř�� �(�A\�@�orSR�f �M�+�uB��̸���2AS\N3�IUݵY�R�$~D%9�# �\�����e��g�����/K�����Pb���g�(<�|Z�K��x-?rw��U6̽��d�'���Fo�/ن�K�Q��L�[9ú�ȗ֙mB���f��3.(�_N�� �������A@	�pD��_��}��GY�(|7S6��?���"�	pn���㳱-4O��h�A>�i6������O�u��"F&�$��`��4\�zmb��3�d�<�(���n�3��h�g�	��ox"y8P~+*��O(�X>)�a�O���;��mՊg)��C��d��Z.IY	w��0��GSLe|3�cU2H�mZ$⦮���0�}�L�£xk��i����SxK���	dd��:�t��>�V�x������vb[�ʯ��e�K�����I�1g�aa&�ޤs��1�{W#W�G?Gr9�wx��_��psd�g�A� T3���v�m�X�z����ƷY��t$$4����N8Z�ʑ���~>����'^��z��bc�9���o��n0j#u8���\�!&U���B|�4�(�a-d+���d�\�o�D~[�}������J�ֻ�T*-�� O�Fk��D�_ق��Q��2�	�{[����`1+�\.��\��K'Z�)+Ne�*?gd�PT�7Jv��^z{8㳰[P�$��b,7���|���A�\S�|5�0�6� ��끎ߵ�ZA���8��H��.g����T�:w�#�D��|S�r��R��9g����ǂ�O8�h�ŮZ?��!�k��, �M���$����D޻o@>^��Q�ks�#S���m�&��]Q�L�N����s"m��H�Bm�����T����O�O�5�?�X�@��7p�����gD1�.?}N�X�����駴vM8���"�$�9·`�o����)����Q('arN�A�O�Y-��z��{�?�=	���R�����b�ҩMS���Q�T]�P��b&a����g5{��A�E6�׳I?�h�Q��a�Q$v
���'��@l��A�z�E��`7zH�S䴽[~\)Y��!b�2�-T��3j��W���'���y/N��>���-��@8\8���s��'R��<B�|J�šJ|f4��Ŀk�<��vq�1gK���T d��%⏨��<i�-x��Ji��&Y{��ع4��C3�H�~o�1?��Qɯ�R�a�{�a�V�<2D�B �_� ��4�\LT)v��?�3��H�Ď����Z�Udp�9WyK͌E�����9�����C��7�1��,�π�qE�� ��6��� ;�|����j��CW@���D�y��x���F�M�G���-smT��wq���U,�Q6V'*w�lǄ6
���ψrg�������`���Gi4����x��Zi.�SK�Fx^�4�� ��z��զ��z���ж��5��|�F(T���6n�@i���8|a�y��B�`LgL���+�v$u�6k���b+��Z�ڴ1L�@Q8[���}�7����C}6mS�������柜�A�bL���d�̾|����W���Z�]��
�*�Z��Q.�m�C��(�6� Ժ`^�:~Siv�Zv�N�s�_~HgX�f��(>��m�8���m�kR���ĎʖS��(<����o�*�8U�N[x����G�c�ap���S ����rA��|�Ȯ���� >꧄�wZB$�H4��ױ��<����?��'�+�@H����+���,O�9ǋ���q�t��3}K~���#�G,����_ā<�mk��<��͑�Eފ9����@kNH�B󚀭���܅y�+sv�}�v�ekI�L�ǃ��5��
x�>�FbG�^|T+��l����b�@W��k�k��(,��;���p~m8�ri�a�����P' v8H	����ge�E��t�09���{���rp�ۄ�1�����\@�O�+<�\�z�%�]"�i{���ӪE��4Y�z9@�nW�C�ҡ�m���h�Y���c�.'�Ӣ�ט�n	�)�?�S\�mܔ��RT��Dk��9o����R�JQT�џ���P3~%��C�����͟U�	�HE.�9�?`˄����"?�0����TY�ФZ�7��.X�"YL���T�-�D�@�>39;�y�n�A[Ͱ���	CV�`W����p:�/v��#�͍Ov,�w�fU��W������LS0�J�I��+Ǥ�~)2�|_������i���q ���w��)�p�լY����1�������+Z���<�����e{��#�V�(*CQ����P��}be~���7߀���fl�dx��1h����)Ѓ���L�L�5x�(�w�vMK�y̡�����ȮI�=;0�)�K����`�/��WرAh)6���EI�M}ޮJ���=1�,�t�B��+�DieӞ�w-��e��>�z����U�o$�Bɹ�[�Lt�^x�U��㙢$Iv1�}����b����'\��T�~��si�>�8#e�$ia�����-��"��$���̀����y�1��_���ږ'���p��-���
��Z�Hk��f�-~j|�6r��i��K��5Eq�Y����Qv84[�"
����E4�Xv)�ˏSHPR�Kv��/C�G�4v��
���]~��kr�B���%��^�/�1��r�L���v��z���n��W���h^#�͊�׋���BqWO���������]*���_�YQS�t��J58>XR$U�Q�kq��F��,��E>1�����\�2�K�*��yD�U���iG+�߶0����fQI���JE�� ���`�2���1�D�����p/=�����T�����x߮�|t)�����Ds���j���נ7:�>�̓0����%����"qٙ�z��#J�jH�ejW�y>]��0}aa���Q�lJ�Ԗ����];��:O�8x�a��{�&\�ja�qe�j�3��:��cՈT���MB�^f��
��Gr��z.�ι�`4�b/ .K�5�-r�����wB���<D\�������7>��+6U���4����2��,`r�`9��K	�Ͳ