// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:27 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iTuyB4VIrVROuQAFlZq51jOm0pHsqtD2taGSjIIQ9v46JDd+WxNUTLAEiHdCxCEM
vnzBdvyY2YO6TKSBAXIqcYfQt/6pFxvGB2sMhQpMTNeccrsDCSifZHV+s1uFORPy
+QcLC+5fKC1LB9kZR4NdvamkyFkgzk7JC1Gp9aLj8cM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10736)
tI2ctV64MeRekwt/bOIbz3Vty9Kj6pVibk9HXLMllsmu9QNq1hxOZ0gVLC2wBudo
quAKdDZA8aOeyPHa1DoBOYJ9ng2+fzA2GpsBHiKcnr/ExSQu4VyKUkdEgGSrNjy+
j8XnV37Gl6ku7r47cMaBQjnAZpzeot2rWxoRZ6gVHidbpRcVqnRjnYI6VLpDP13x
7uXY39ud17CWmzs13LHWZIihTXChenh67uc8qUz/XmwvAHVKGwjlR8ZobdfUwxLn
aGflUz7LHSkaQiMxCOwAxnWXK7tRcH77hCQZv5Ha+jViHKPo21eTh5SVrw7ZGZWQ
2HwL54MaLdYBam3MhpzZ0Ieka91sZp5zAQeo4j28ozDhM24AxDH1p/M9V3sKSP6p
r0B0JA0L4vzR4O7+SVMJ8PKDbr487BEnOyxUJ97jdGaJuyxp2FdE/4XRSOaD+Yhs
omwGRu8iYD6PeVF735ES/oNXqcFdbmwYKH1Cor+25hWjC7+0lmJpfvXlTqLsblhU
WD2/Fn/RkgDb42QugEB1VcoSz2X2o+NrYPO79qd855zW5Fdkbbuip6n252UZu2fO
7HyN7pKHEB9RYczB4X55IM+/P5htDSoYY2brxjiwtB2m8FtZP5A9VHEvH6tiyTTw
z9anWVNGSLkNB42m1CduCGV3otBEy9xWi5VsTFNZH3oXDVEAQeRe+o4nE3Agn4MA
yDvChakFVRYsPA6RJ8W6IM8Cu7Ur7aEu1To/Ao+3MH8qEyuqqSMPctjSAb8KGl38
8TI+0GAqSYWDaYrMpBb2rlqUZSX9wyaLdqyBDBz/mfzvbhr5szgxruvVKRqknONX
oDpsLUMfl0hGtgmtgEVmToc1Gf4hnAWSYkGfHd6faAwDWvdrYmOiqkthsoVhMuoN
4iRb7TR4hp8VVO/cR+Mzjx91F2nIfcekYfdM4s1zUNXjIK5MxXNv3CQDv3u9yryH
9GkS5+6Y1/8r42+/bmTMUDd4ql5vKOsydQ/Uc7h7Vd5orhShttq+Em/THF9vAVNW
nTc+TDcmeHbTB5JTOH8DxjOUIuTxR+JRnLqWDfUTsSIWpUH/YV2yJBZYlOGCElIN
QeZkleNmtz1rXqR0p6XzCywJGh6x4wRjaE+9GJi5YYNW1YNQJPp1teoCaW0dwf9Y
ftyHAZOsCWqRxzM3vK9kontVdmyfmxwOaBdNGQZLMm9PAAfgHISkinMcB+twvfMR
lJOPFuppbE1FokiFi6w0vPRzyco4GvLJF9qg5HsjFW1M/tVS8XZGUEehid85s/qd
M+0vUuhFeQHsTmoFa9bBPkzmZYcZpw0jHBTEDcsoJFRWeQmlCCnqDlo9aEZfhKEQ
LJOZzY52uM5UZ7z1/Q+Q8ACtKfUUmuAETaYWxtYzkbilDbRS5vwfA+uxkXmUNTXU
7kamHQ+5CpnjVBi6flMqpCQzBGNd4Hs8Ru2WpKsbCJuIOw4+3i/KzPEyfbOL9Abm
9zcm7CFXRYmc5NMELEfml1uKmfDHEzVcEvICSc6ZEFM/DApnfr1S/f3yVMggjHCJ
atOmUcOkgz7hzuiJD5VIX49XgeaYh1D9Y2NPdPIDPNQZMhzKOd6ke3A9Rtj+DuNz
7n69aiUDtTU3/H4z2w8STmK8q4ad5mPYPEFJUy8GYL6ti6bNGeD3StRvu/F6Y6Mq
6Kqpe3xDkwvrcSBqUsaDKu9WjpCXfKQkoG/2+Bv8wyBxDolTrWjYm9htH0CC37CZ
TZm/N3EtUx8hPLDWqVT6DMctbOam0CeFdTPTZg9En15NDw3UHAjbonW1sVLx1DB+
FsVEuzWo5HUxK3a0LV+wFQ8csmgeDY9kYldeyHjfMNt8xtpC20rMzsDZXhCwCuxm
t/8AqzR6HmmdJwXnFuXldGSqNjrJdgMCScwdrN8Trk79QxahwzFNRqlKNkm59nJ6
+heXt0B/Gd4zP8PKbSvdzN+Dr3lGd87xonQe08tvVoy8sHKg5IcepM3fUzgzBjy6
CRqGFNYLB3X8gXbGCk/mayKMlJMOLIdzXoSFxOXaE1WsZHIhB9GpTcXxjBgZibln
1yIN8LqZZgtn8klTc4qOI2xYyVAnzxFGH3Vbl5l8AFoG5xFQ4yK73dHOgZDG4fnB
wtHX0646YxplL2jxZVHcH7FfkuguAEJaQNuyFrtJU0OK8R/iq6NP21GSWDUx0ytx
KPcqfQ0A56Y9hkjAd7y4cNAbmFpb2jBRQufaOp0EI8+Ef7ALAWFe93apj/mAvA1D
CoURprOKz5fu8+Os0FXLoBeMUnJHmDwHgDMxby9qT+fmWrRifUwifB56ak53/HWk
hT9tbvSQEpc3+ED4fgyIF944k90b6XDSRtEMMIUHIhdQrirT2/6oxFy7CbNE1Fuf
ObUCEEoJEe96KHNt/14l/hatBf2mnzEqc5qI0VsP7SOHG9RpRTtxi5qmFB9MObX2
5HubWhdSIgf4Mp05cRREy7n9qYOknvU0PLckalGSuO1Uxt2GFnHa6a97LpSiI7/X
ne8uF6FygTjAuMUwa81Sc8YKaKaRVyhfgxHUES4JtyozLUeJXmkQwmhiyAHF+1iL
H4TVLfSIkeUmjH/clD2s9v0UW9tsQcpXtbrs0u3+THgSbD5XAkDnX0vznjrTBoPQ
O3MHQI4dGLxK1tyZxzR7F0FvJfcacuVZW8wv8bbxJ1uLYcMOasfKS2bnuscDBEaS
3IB3oQPmvyh0zkAlqOIdbuaH+hpWdieI4/srI2zI/TJSDi3FNUWzyCKP/DYPWYQc
KaRROQFZjWmit7OLf+Uz/lj02okYSkv6vrVrcuCN//fiO0yyA3zooh3yCriefB5E
6JJIIMKzL7P0priSDU1m6c8WX9Z0UYU0TjZk0SaXX/K22h/dhFnTYUQfzYa8WueF
1oKY8LFDrxJpCOLvFwNEysRK1HCIPOkfTO+syc8sC8ELlM14cxAbvSL0qorWVMq5
43Mx8qbIJhIGa0zki6/BI88m1//ZiksSoK3GWMJdtELZxwRUzTjkElxgRQ6Kf0RL
CGQUp7j8cZk9AVe0eu70CFS/Op5jA0tT9YuE3vCTSWWFWk7x016Lj3Ts26XFM07u
7zs8Ww8/KYW7U6Py4kEymLcsHT/B9nVT0gUa1nTChIctM+zYylMmJfrjam7YPQtk
vL4t3/jFL246aZgpBwq5mR8AgnGhmAsI7008SIgijAZ70vq1FXsnDd/JTz8542j6
fAQmR+FueYzfDZ6pN5edlZOr/EnRjupkngF8umfQ2LsKDkIYG1LEhf2JTsqn77bD
QJb9zQdpd0zXFrCHpLnHrV6u2diytgJmJ1zUsrZwt8fmfxIU07F0nuBrYpGhhXC5
8y2+IdFy8VfrClEI+lOUzYhIWCqWQgxUvB+733ZqD7JwRvn+RDte1Kww1Ch0t56k
q7yJKoKVeNPPg9HMKTYlauY78q67FrIhyJ6/D0KhlrhGtIcTVLs4Z0xM3c8RHAH7
z8vZ8k75DcvOK5oXwT7kBlkCCbV0DsRRb3DRqg8AnIkjPLnpAIFfbeE4tguPfUsp
PRKiy4NPJED3SrRm/shQPrEYhXVH/QWTs+3OxTddpF4abk3e68Q0gUj8jE/IRlS3
3UPqHUQGL6wuzCp1aivf/w6ta0bh6iEcUqUheKNA1JaT8PwHhuWrkVeFYyXmzK7a
bn/vR5OpLiBTwjLXKYznQg2+YQoEAvvmPRKlh/hkbDppWuBCSFxFZjzrWbXiMYpG
CiHxngKqGnmGV1wF+tNvKMx/ntEKT9ss+AJYbOoW8xxqtja2T859M720etKP49jN
EG1Y66JwW3VhgJHRQh7xelMXJwtpIEfsRtQQM1lnjXnFGz53BWbOG9yurqwVkgEb
4QX7YKuqkaoHMpbyjlF/xP2xzhMgVioc+sEdwSKmI5IKjV/pTrLX5I/GF2zpRW3d
u0Tubtk6D/aISY1aonuao/DQE9Sh0uxST2Lf/4hwaitFC7GP2J0VhjhMLhkMRUXi
fcGnLygMkn1IaIbrJR/d3X3aV+UkGetr1aQie5GvSFX5SgqzTJwzE+63Bl8UZxSO
9cHJx6Z2NxidQM5xh4P5yw9/fW3/MrFyTDh8w/bfmkPB8XwbxwPS1rkw7FVOoRqc
z+SxX/kvmrkAgTyHY0v7gqLtQOupHXeVZV0aj+GB2ZbFqhdGBBdF15TyoOjc3Q9q
MnzjYOh3cmKy6W3SEYQzyNfiAtGviHbo699fCh3lz0lTVM9feWmRidYInQ4tEvGq
tcMwT/AtINWe2fgk1RIMqcxcfOCqC5cwe18TlOfRiNyQHhqA5FyxVIQyp33hv/vz
lUUUMeWT1zQZZaZyDMiZwogrMsJV2p5T1Sm/r7D/ur7cq2Vn43JcbghtCDHfJzVn
cyRF6qgBqzuhfa78cKJpaZ4Xx9LdbqKxaAmHpheDDRV9tyvTO2CVLksXKgBXjQWp
4kfKTAQFT/FK81laPEpGCfJrmqgUh0QDqrZL0oxnxAF7wGrOs9jaCJHcSCoSEzRr
y/BclHOyo+j1BPNjoPX0SNur98YdcOMSvCHqJPpA3AEuqlWwFP/BcnvsDYRAD+Mq
gPZy1w0aJgavYtqsbvMPLTv4PcI3r/EaIP5SOh2NdWBDfNtAv+D8Zl/NRjE8El+N
ZXqrEBWEVATvr2qKyBSdG7t1yYwfA1mmP0kr/ZScxdJkit/ig0hZyG1CE8V+vuMR
JA2AUn9Ln1m1nHh/MEqo9Ew0f0hhp54Y6fhVz4Mv0UloDJDJu5Yk7Mx1jhlBDbaJ
2Ee7WUM3vQjs/y+2MG5zlH5hWA1n+ettUDb6DXpVE8HgVzI1cJ4Wku0UZbPcBP26
ws0QAE/VsrXEqHYOb3RSs9K24VkCjJjXfDf8WvVMHg28I8FrcY0Nbpu4inDPjN1X
8UDKLIyG316zS014Zya9Ihs6RNY5zizqpgGP592+KGGW8MUNE1AqLkEK4leDXVHO
/uQWP2+kbPJt/vhpDhQ+ldby/4vAYmAETLPG9q9OJ6r8/LhLn9/drefHOrwpSmO7
l1f6IqkV0RBQ2KmzytVE2IU4VfoLNViRsgepObmcwG10fpfNC6U8JdjfRnCzcuZ1
cq+z/utx5PVu6FxVzDo/kkYHN6+C+0pu72pOp7LNijjLwOQQloVG5qnmvPpSRJP+
JtkJ5j1SDLG/clb/cr1GcUL4wTZdzhfuWJGUpEQCM3821pjOsYmlYrJF6dyJzjkm
MP9hzgG83CnCHIPp8kDt2mLRY1q5XhdqKcXIbpIfQcvC1xMiX9NgTm8Q2v0Aa2T5
+lRzbr9Zmkg/JVgdqIq0roKzsHGlxUuL4ogaHu0oqM9JURhDSav4YSYpgQqmuJUH
h8pDS7Nt6+S7z9vpUKT/oMp8JtG8OCNDZAEQwBbS5Km1C1RLikokLgvIK5gLM3GR
vr5rQMoFkL5ORh5qyonwwlhEXgnP0H9JqCfzDA18GZ6sMDJ/yhpwKzIU2EcRjmZ6
pnvAkSMXIA3aGEHXAKA3VmZQX0eRDu2Q1G6M+HRcUNHkC3TXtPjUDUapVmxNMCBn
1UqRF5bhvcW548u6hZsInluWyDPwFjkLm5yH2Z0qNb3FD6s3xZX0mJFwch25ysTF
C+TcPoMM7HscqBnXwAapB6GHaKisSxGpmbdoTTxOVfGBRcKwsmkDNy1X55KZmOe1
fsDJ472zHRB+npsdC/vUj+1CGuIATYs415QzHqgfQxUfFee6YtrH5kvoBf1uGONY
W97fUcbVH0LAJ+flUc0LvTEoqD7wnplFyf/n8zOIfQ4JxPhJT0bDuJbpjmQl+aRA
Dj2SwKukzGhwVaeNQ94bQ9PMLaVvaIj9aa3XQOxwgs+U0hURoGT904eEPRQNTZYx
Ib6Mbq5Ht3ypgfsSnaWv3RY+DwwamqCNK9FNwU1+OeD06llZRmoV63uzABpEXjOO
cC0l6Lo32ZzV7nJeI1eDgmu5HX3x2ygY64vXszFdNW5T2EVy4yUtNw5qi8BoTjF6
CNQJQAHLbMYmCqNq2/kdUnYA7ADyzE9947BZ7SIM9m9UKFydvZpoLSRO4q9ri+rb
4fKVeMXNufde9P0EhNUmjcWiJSQiicstX5X8ha34xJEuIHNZ5sxHhi9FXSgu/Jrx
UYvkFY2cq8lCWZY9jMHT/i5/IyuzUfSeCmh/85dpJYLG0AgpBu8XQEP93b1SvdVP
H5uSy1qJjDlTLo+Bt+29GQSHYqJ3FtSQqlwDTTn7IqWJoc1eG5/6RPdYYKcJG7A1
DlQ3cfyeqdbfnCb5Kkw2T2Lz+ZWyQdXDiU6vIzINn053lSpPcnillyZI9trsYiCo
/3ar37GtkWQO0xmA79Ui2Vo8rLzGHWlH6H9/oGJrUoeDUuFklAk0vWv6jB3jtfiD
3DMoXU91s3lYn2XWiDlzSg7py0k6LmPVXL0Sxiab7td3ApDc2cwHzOIHu4xajdkH
1aCJ3Ku7IJUb+CFT9CWqldB3g6lVq5wIg7MI7FIKsgKxkXt7mgPpvyNoGCO81obp
LDO3qv7xVkFZ9OkDBdasuhm7cBmFoUu8e0TfmtqzpkRyhdr3jaAxAE2tb2FWUc1G
GQxLscmZj+Z5Y8QrHILH8MXdoJb/aBkmN/2Q9mgnsbxsc6XZ9hKxOUGqAbIZnsbB
HTeUDgdKMIaufLAxqHMXsTWy8iHfNSyC5t+G0Xo5tPEwWsDHukez1R5Li2grHIAN
67bDDXbyD3uUIFvesyse1E/OQyzdZzlPNIVXQPmbpgyzHcWnTyE1tZYetuJh8nCM
9J27clsD6iXWn5chS644vz7Nw6bQmFj+KHwAhkZoR9GRlCEG3gtIi4wxkP+V+IyB
ziXDGcJFTWeBtbRFxECfOcgYKawWgJG+yGBmGbywLkB8pBAzaqBf54TMt4CcxkEk
Ik+5uSpo3AcHWK4Izg7gjj1VuxVxd1XqGdcuSTKFSDfk8awDJF/4LIiwWPTfUi+2
amrxixQ7bNRFxHcIjhDTaBvK+seLuDOm4faCGtVrPCiSrX4Knj977J5VdrnnrVLi
bAGrEWfsFdp83oibX/6F2otKAQ/ZdsURYot066YFZlgj0S4KpCLymAeXv+MiY3jF
FcQkR/aE57gKO7xOQB+gSrlDeUEc0jm/aBGoEVmlbj8H6iHd3NM3XNCtKc7ccfct
2z/g8KKBCamlng9lWVXhrw3WDKuGQ48JkAwFVWVxqSV57ExvWgFzMtDfO4gyFiuA
a+rct9kHIOmHo2tgQPfGfR42hOiPMLcBc5oIumogbNWGru6w6JSYKPHKe+UJ2m3R
s3yCK8KQQTEEcD7KwNjGhyKZZbplAh6IK3+veIxB4AKzCLJgY9gJ6W0lZPDtBX+b
w0a5XSjJvaxd51GQw6WCZb1yzuvuuWnZSJ2P9QvyCne764ouvyEkEcbPYQb7KU9f
1ynIIbANAeRGmJ5DZwZMzpasU3sm4uLdMQs4sUMzHaatHYKHbHPDGXPDylt28aZa
fc3uo9oLK2gIuukWGwhLO89lKrBxHuJSHo8jcKU4D3J5RzUdf+9Iovd9LvqVCGC1
oszniJu3bpei2r2aRLZlUITWIYDXcnUHgTK/3uP7BiIJm/Z/YWxVgaGVcJ6nCbKP
TH6IMcntLEE93iD7ve5vwpI/XcHpoPG7TwnTzc0JC1zbwxVFGcOzYpxApH/BbfX1
EdbRakh2UUdTQSMyavZit4idbXlBM2IE5+3ai50EyaHyiAtXOpHHVzf4YIoEcQdK
KK6uehIeJ37YPv7R7Rskw8ReePv0rQXQ/wjcK2kbAFMkZoqa29Eq4lV//NpaSW3W
RDLpce6c2llzdl9yiuwkom9zoiesIeCAv2hBz8Z7P6A2/1Rjm4C0Um2GQ1qNrub9
r82JYEfLoOJ7ExEl+K63t7Kd2BOOaO0xWfPFa53ebXshJcJk9dGMc5bJsjGqrToa
bgyTEL+93Oy0ZoG3aIZirsXAdOSxqCiZexRVfrMT1gr+Ah9nu0OXBhqXaKIq7qqd
JP4mnhR8cnnV/8pz7T1OPs8qBv+zi/wzR/2bimrWWD8Nsz+EZjL3AG/DWyYgBjOJ
Y+gaK6rr7oQPHb8+wJzDxWVSecW6oQJs0R0YY2ijR//u9Rif98lJpKLFyDqqx9EC
+9WOZGAEC2Q4gYkDoSwVwPby9sjjDsxNE15f44UzalhsThkR/5QbL1NJFv+13dqQ
iEy/XhVMGThKsoCP/QnVUqEdaNcGQ9+oLmdwtFeyi78jiYavLe1mKhhnAN8U6sLY
LyoR3rGNCP4vqcqxmku92TCXtYdvSvC3qnBVAc1r9OHAcwQ9L8ZWrBRrGP6w3EGW
POxHbs9WkUVlMweNSNAxYezEuSrfPKoxnTcp8RNBwx/8TEi1nwVe0htFz7SYa9RU
dcp/Bj4JIc4pejWch41+KV+yIMoXHsQtVuAP3uP7xgIUvqlwadqrOml96I87jarz
oXGobNL0FhfNybmtYl8xfw5jjiSct5D9KHapKs4lSyrAcMoyxfBcGIgSdRaE+WJc
+raAgNIOg8ZL6GA6m9FmG8N8kfmGaeHux9OCuvyB2wXcoIyFBneQ0CBKJ03dtydc
x63oZfl/qOSO0wlFTrKW8z9l4bjdd0e3DByv3a+9MXyTG7T3+QqdUvyTLsOk/xYl
ONIBSRAgQiUWmBPVXj6vdCTWL63Ri9ZKgQoa6pwnfWlIqm71LrNPeiYErRDAlqIB
GNfns66ZkuE/GZNLVfO37r5FgP7+woDHfRgPZ07KUE5zcEj2QomDrEcC6CqQ/MHj
URa/naiV9btlk9XtqffiXzZin5oAIEosy5Z6gcoU44fI7AmDMjFL47p6UxeBYLQL
Edy8O7U54J1iRaq6d1frNa2DXQKqYRYNkt/87yAMWm2fSBa0lSz5SZMDy0HbGXhG
OnxdYJ2w32Yhg136WFOLWPluO4S2AipzfPYl7VFcfA1lHTyZ8rNze5CFUwtwSWMw
GxA8rF3b83/ieO8xzsPRmBgWsMhyJmfBf4emR0v1P+q7RE1P9FZ9FX3ZDpIaYc7T
/NysnE5fFZHs+rU/YM0f41ASaXibo3hjXAce2dZRfU7McPyich9ONIfylygDWYR6
/VsWVy2i6WctvEjpBHXjNNW318GtGiaAE3uZ3LDm6YxU3+BQt8wh7bV9AyP9q0gv
GmJ8vZuhldDt0QjtgB78QyL9kIz9oVqfHPS2bDqdfwSaVjczws0J480RXojgiGhk
SpsAJaOsPcpgcCDD/ejPKtlvO0JizN7Uv7R0scOsu/oFxVACTdRVWw7+ke4iE5zI
5D+I0uJ6ghBFJKF2e5ZVz+roCxSddM8f0otR0oTlg3akOz0rn5XCuD/fvZu9Fh5L
TXNczCGn0rjkVVQJ/cyTYoMEv2/pAyF2fjbXPNZaScheLbMbCvHjDHpjuIIpU0Jp
9kNCaPcxulttYqbjZTSh+fpGMmwZzzaImeVwc+B+StjQj6gLayixJX8ohITwTzGl
YcoZSepyODDyCrY9YTxnIR11KgMGm07ZbX6pC7qhboLjJ4+eNioeiOQcWpJWk204
FgBLdDBMrEAp5RWSowlXyvPyl3Q9O2JeNYYSxB+RVWQt0+WtbgRwTjo4c5E8Prb5
jFq3KIKpTsBGKRgeEuWAYzFJtC3uH6WMSg4VwDOdlKpmNbGNq7se0N5Z+hgphF7K
4CCGw+t445BJDQh1LeODXWys9ubIgJEW5Kp7tLWnIGmN5fzVfx4Bt8Hq4SK7hfUM
EfyuPQsR+CuzhFzlrzVs2sZXlAqy0kWky7mEN2AErDreUNxahG/Aj61CPaok6PxS
uNcXTaoPrKmhIrtPM3+g+aeKzLqKpTDLNeVF6CvbV1smqoQJKeXTw++DaSewW9wq
cACigLFTqiYaC9pyN4eP7Oq5Vr/Mx6N28JSswF3LynG8DXdm4/SzcSGftX0X6C2T
oePaVFytg4G4aOPfgYNgzBK4DSk9LAnsmzVvFjm+V34boj6/XhJq3+n1hlleC9vA
c6xJ7krLaf/nmW4bLFntpHSu1fSURv3yH4AXJ2lluem9qmB2g8DHq+hMF53w8pLM
t4i2l1TohKVzOWPK/jrl9EdKfBhnJtW21h2xm7HjEwrlhijd7VAypvBNDa7xwVz4
uxHCg41LZ80PpWqHxDbpUou3AKH3EZD2572oVN1/UalXUWgpHLyY9UyYomHoMclQ
cSOFg8pBOOjIQxiEaykvLVllW+gflTWxanMRirt5RCIsq8O8s6P3KCQllHaL+7z3
WJ9AMGSMyMj76/fF8VhSaOXNiEDNw8besX8v/VuuuCx7CbkvxGgt/d7lRMcxL5qA
V/MTGF1cr2BdkasMWa5fx5tDf1sXz2McmC1iDGq4Cr0cejiCgmy0qRUvUjZxhN5V
FaHvxWrtcVbsU94W6/V1ii7kqeNZb2bXQRoededyepAx5NYnmIlkEFFlAhBVnVjt
Jg+qynsbCmrhx14zvmzDa7jce3TzigpCuTZmboaRmlgKdE6dbQE5ycBHSnfts8KH
6ac7eoVIyRYMdWwC0qUd99rM3oh8CA3yqDTUtmkvpUWUiGZuM3hG73qouqnB/16u
58H0JJzYrAl/YJh0qSXZO0B6jMoOAK/oIgUGHzspsNfnH5451/dk3yp+Z9hHKP+G
FhwGSX6zbvMbkhqONTJ/iPFcDldDCYYr8QuXLYWRnXF6TlRhXpOV9VZHu0m4Mh+m
FHe7e7zVJ/AHwUjkjdDeSxTnTjf2gVy6EchVN6o7SKux8WvXpiwifGNKNuo0CRww
dPf/IMyYyPkuk1X+8/2UOoGMA5wDD0Bc38r3UZ98LU1S6v5uEVplTaDB9vT+fHIz
8fsXDvH2Hw+iU6oGlSYjBZOmZsBGxueYJIM1dAgpQI+kKDVDzHN0vRDcKCAPBGbs
5OMF8vc0cGyZb1l+lU87GMaqw5ivzI8zaf8bDZEHN4RrMEg6Ew31/FfotB/2Ivav
IhiBz0jPV2rsKV3MWxhGfBNUrm5JIMJwbuhmdn43+ka8X+fIKRbZdXnTwy7LuRNz
Zd7al2IPe0g/pCNMgDEzxXSz2Bfgtue3c+fhK7e9qs/BodHdqogmsHb9oyf2qfGb
JksbT7oOct+4OiWzJeeLwxCg/5BVP+J2tv3ce7O4EhmBPCTgM1Z0qjimTZshgcb4
f44suC7ylIh0WE5EsBgJdJykvILxkk0qrn16252aN0Diys02OaHfUWLzR/R31jMS
yirIpxbIXnJV1TY8YraZgp1r66U2wIpIcspg3U+Sd0lu7+n+Qf+94rnKki/34oBE
BUUkPwoLzPIQgqnp10OM9fqsozlSuQTcB+T1TuB5M9vN8t8L0puYImMmo84MnDC2
6ZG0r3TelfKj1ddM87yL8PjXTT+pzNi8B8BgInBjsZzLZdg1n+KAozrqNGRxTNbI
ueBMwf2/x8CbFVraeFw2tpi21qB8p/scU7f0dtNiatgmTMz59WwRsLebRcrO+K+u
pWrjbka7lkMaJnqRAuaN2iGNfZ8XzUXna95KWtb/1jymg3zzdps1d1GFqpP9QxIc
Loj4vbroSKUUtXn0w8EEatQxuMgYmqyeKh5XC6TyPnkpRJI+cpjewZs8XDzn8ocM
dbeGQUk4qXNoIKfN2Agnrsd6KP9tEpzTDpJux90bEziRq9Wm2h/VALHHz8h/Q5kT
K8XEhubevYxxyEtthQ8ahH5sPLA1cVigO2D0MHL69XnMx52Th07ibxi0HQOh+W2T
3O5Dot25TIYe7FU/mPUBteB9qz4KqHe/OLuPQFtPLI57UMM9t4dYIIOXCTpvTrod
u9WV1KzJ+HzqvbpOWjwkrSM0UF8wRV/DY515VA1LOBD7znUEinRTYOOGAk2lWyH9
jHcgXA/GFbChBwysZtx8AZbnN2EG7YwaCYtV9NtD4HP+HMt96gCVBEbjG4LQWc4X
HdF/bPcynE8ynIX+G27c/T4ZPgUTrwwCNH83026+2Uhk9ouzPRNqG4jUR7Yw68vD
BPkv7V71H9mkAU1nWzR9+wjQHTw7k21F2A1LxMNvM9teykKQ9q+EL9ogdWZyfbEq
ZdDuk3k7cgTKZaiXNPyOUNtBY0dHUoFfwoGucLs9fbQTLsohkOpTUm8MQ2UXlU9U
KuwsX3cn1EDq7TzZ3icVPP7jLQn4jCS/ZzFeXqvgrhNd8WSU5FtbmggBrEN+NxeO
IrRcOTRQ7cD4714TjKjTW4N2OcDJXIY0eURCRuyzVmhscT2uFhecR0Usj2KPvJ3h
7HH7VnI18aNwCO2+xw8aSw0V9MpkgVXrWDCbfg8dquS5lAT2avL0NYljEukERWyp
x5uxXyKATMKytBTMhHNuNRLzJlAulptoUVU+v2EiWSSWibcrVhGnoiV64rKqTBZG
7U3+8aWLqpiA0R/DB7M6RyGYZ4ZRIQjPq5bcX3WI+vRZP4L2jm2qtH7UMf5URIll
kmi7A4oHWVoqmhvd+4EWglU7UgCRqcx3RlPo47REOexok1iFwYJqU7DOs0FkGuuR
nHBpa7I81xNjWOMfw0Fs8r/PUr7rSQ8tJAI+/pffQw0fdoM8YDWgI8DeqyQORfaq
Q2z/+nnpIGVfV6r84E7TPHbPh1dlFB3Ik6scQHNs4z+9Yj2O+rkHSjCxdcMOR+1F
wxFv5q8f1O1XAgPa4BpBbNP8wbUoUBqy8D2fn18eOQio1lK4BchMgsyWyEtXBYYO
0irsbB2dE1LFbp6tDbpNi9z2RhwA5QapFlhfwAyC5J+Nq97W3CVxPZcWUavnLmpD
kyOAJVTlEsE9u/phmg7lR7GYA9+pxJqoXl5enbRjvBMZYWFXrx8iKInCfEEO+KUg
UC8O1TzUzvuPoii7nEOkUH7p5gLHYYC06NjlVaSO6046YVD79J8XjwtBj+7BST30
emcVoqbQLrYPPAFBAx9pLwCPGFfOPjMCUT84qUeLr8FloOb0D5D0ewJU7Z/Ytzy1
YqvOchCc9yA5Vgop4rJN9zS3yfcbYeZzYYuu5pjVPtOBq4ElB5leEgPBwwdlX5bD
/caUImic6UDo8zZ0w4XQvtuaurCIp1t/TguHigOZ9XDe4miNcZhRM8q5CSIJmKt9
7X39KhYGrrvJXskWTK5YJLO4lIu2p4mwr4nvMq4WG9/agYAk2XbTY+GatRX2D05m
LveNIeGadAfQ8ylCiNzzhzNwmxf/vJ5VeCROQIdarNyLyEEDEig2qSypdMnmWXTL
46yCd6fVwukcQvfmbRKDDXpKFx9ZgY3rR7MIIpRB0CglNRHaC1QZ8hLtt4MMYHid
pjnxMfgZ43HhkpjGoIq0xaD1VP44T4Ov3stsZYA6cX7WCfnN6T3OvkCvOixOcJn5
WdGog0HRh6PQL3OKIzPmzB+BI8ZVPRbzOOjK8DcT2H1U4HXZsTjZQCPyMCJmcZ4O
iI07Gczn1N50qmFRjtRA6JaJnjW5eDNRzwBbwAfxrM0gNW+VgRuiuSXs5u48Q38b
lG+myQ8AE86pmx0VBsEbkT9oXmw5Fjna1kSPO9M3H1afwyUiBnUKW/zTncIYrtrj
DnOIoQO59LUUD2K8olCnijHU6KKGE/RwMmvjFQmw3grU4Ig7W1zS5ve5iqfBai63
KAuzfI2U7N9R2IK14Hm9U7OAhmCJbGsEYRB7tN6gsP010SICYTFAIEXuS2hOAgA5
Rh+8nZMQpv9ssFKqmbE1oIU7PG8fgWFt5CvoYvAw4PUYa+LtO2p3hv5l5qSQSI3Q
ckuxY1rTErYlf2qF6DoBIIB7V7TXVZBokBkxLrt2G1wJd5+A4MkbC9h2Zq2JCjw1
tgkUq8R7Z/Ef+yN7I2h1uB0F8Flkdvwi5yVBd9lXfOp+WE1xpt3M7Euo8x+PUjrg
Bps8p9v/4to0NNKTYUfcR+8CvjYt6NTzi/Y6Uu6wBX6J6803ETw6b7rkOm9EXjid
C5vl1Fy4iwAS2ZfZ6BxRS5RaKpob9tb3wYod78FDfGR7/mttrNw2fDbYEMPVR0ch
JAxkj6XNG9mjE/BzRtclZjeatCtzdFCNUgyVwYciW0phEuwF0ZD9BDOWBtUJjOKT
3AfUobefIB3BBZ2OcgAYj8Ao+UG6sastqm5GDevcVlwIZ1M22qrTB9vndl9hu1RT
gTMTW80b6HLPymEaempNntk6ISiTuu0ezgY4+zA/Jw4JMcA0KLwIoHFb3pvrJ36V
chKtudP/sy42jVroVa+/dyJ7YxJpy9Kzidk8BpVQO88N4HSLS52J6a+Lgy8Oy9dn
9naZH6RbX28zTYbBjlxTBMH59YYMYEmLj13Xw+M2609DB+X2KFLqS/Bkrtrtb52g
DrJZdwx11H7wFKc0e3u2bsErS7rG3IugO8uCN4rl2ZGJRnCN5RWsT3Xc09APMZzw
ndtrEjaNy1swcZd0fdpWOkDhQI9bm0/0pKTATEUuu8o=
`pragma protect end_protected
