// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:16 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QdoNAvkMF+Rd9UDFHCP9t6iL+YxSbpJtVqWIvLLgOZq/enlynFkU2J8seBog8Ton
s/tD95esFGC3Y2GrkhasAY2auSzPILXqI9oG0kUlZ2OG8cEQ/VZWfp1RujFmPXIv
0pKtCilAYdUliVS8vhzfow7grYs5RovFpXAK9Nm47uQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31632)
D2oiES4OY0lFJ8z2clAJOIfWcry6nfMBZmWbIvB+YK/BfLawi1WDXeACoNzvMPhR
CB6+djjqAhW8+27FXRdSWxaSZ5X6Q2CVKCCLfMqCh9udoAacyOHOhw9ZtFcfIU/1
paFIiZhH5fAx3kL4HPzk+o+gS6AnxNb+J4n13Vg03jQ8SSzwyrqafe6C3m9Q0hgM
E6vDCCfY2p/nBOXs+fNvGetCayW6o89unXkw72Fj9kYCUaXDIvGWIEYxZz+PKAGX
jNU9POGCcxK+mrhoDUuNGnB6XkUlJWiBo9wB68cMGVowlzxCMysm/02H69KfBADw
Z1S2fzRlY4YT/vebo5rZcEJ7tJbY2F2dNy0cmh4YSY/tBcq1s2iT3AO2SJ5TbpGv
Ew07zlrO304CsgLGbIHrWT4sw4m0sbSlFveZ3/cjDvXd7q6OTQbd2P1+MSTr8B2d
QanGcNUmVXHlaU4xuGFKvxZiIx+uK04TghIfrc+keQfhbFHfg2FMm+DaDx0ELUnr
7+0Vf5KYeZM9nz+nN7rgO14Dtio1gYV/JDH4+B7lD+UIeY6sg8Mcvo08rcRyt8K8
FKFB9N3sy2uNutdzLUVraNFr2/ubv0ZNh5o15+5x+A3kby/nB+eFWTGv5fTlOHpA
DLhnx+UB//AQPvpTUzot6CmZA4BQIVWlaw6S8IAZY9sJLyqCWJQHO5qE9N2e8FFa
M1PKEtvwNfRHx/5Pul59DNHJrni4xdmlluVJ7cjaQ9W/rkdbZi20TbqEVWKMT2ss
UaDWwhLXnaPlWrqzaWrLD+aNciBcoMYXv4T4X6YNu4JV8ze2WQdzdWVS9GLd0owG
eF7iTAIZDQlU9qXknyX/VVB49r11FJbLziKSkQBu1Y0eWcQuk6O6elnny9S15nzG
3sS79Oqle1Cju992EsCNDL5YeJj7cMe3BUx/vnN1mGiLQTjNKzVCGTIDDIc20HAs
eZM9hOYPLoudreoG2j86tOL9xgg2MPVtJpkf7KS0Uyu2me/JSwUO8acvLUa8KAEJ
d7cbSR9QYdYGbUym2qtQfs2pWMy08QEzbT73zY8VcaoDZn6zqELz4zNK7RccrVB2
n2YLXgng9pV0pDSJHAGDdkl/Ig9EGyPBDJXZmkL6MvO7kkGS3sJEIYjBvdmEGxdG
xKY7/f9QwJL4OFiCJbu9XbU+0aqOCkYRhNTFiteImPws1QmDUForsYufx16rMBm2
nUprZWtH3Uwj8q7g42MvPzVYr6CzqsGv9EHBJ60r8zDg/bdvhcZnh/DGKfU66urc
AnCbcfoTC0/f4pu3FI+8sEzv4M28iGxDCNQSJonkE0vWGxoGHqhVN4P0B0PLvSoI
x8xLC0WGYYH11CiResLJD/2vreD44Dn0iUp3m9rqL0f5FfxOvLNYiDSC0fTrUaLF
DikosBrM84ref0AYpcTSme9dJMgJwjWw0AsWeNKQj4Jgty18unx/yyVO/h+l0PK4
l7rqgcY2hbjBU9WFphAn491bcB3TPyLymwa/7/4DEn9+eUV7Yg5TxdU94Muu8KxM
WwO+dbAPlTZoTfirwYEx9Un3G7MJDqrHFOZTrla7d0oDCglZ4xrb3mfXdLWGPV/6
P6jxgM/x42S6rQFO8j8m8YyfH9TD7zW605J6Yx8i7OFVU8+LZuEKlc/wte7FwEic
BBIyXHaR4IZQKkZD9RGLdDcObYSdxDJzDbziG+JUGR+Dyy3qjEz7te2GrUlDHzvb
NsnMGFWO4qAbPqa3gFAFJecscR95fHryhpMwUo5zIQGjeN1p37bHQhWXJiDRep+X
CWy6pttEVnG1A4YihZ2LkJMukerx3jPh8iBQk350psguERynPKi+N56rYgtIna0d
MAZFZkMKJxG6x+1AQurcIpiJRk7WnP+Y7+in4L93cjI1oWr32KkQw/JlQP1SUBju
tJHllEImN5sJcUk7V5CphJ6cluO+Eem4qWslhWjIU6b7YPtcYcnkyg0iv7lBT0hV
+0sXhZP8FHfeGbOoKXEhyd53qGw8A8P3wN8a3P5paj5ChMJBdTjApCFs1XHuLocc
flwEiVaXP6zrkJQTkFk0r9pJp4fH/7D9lk9Vhpelf9KEKkQiQtLBen/hYFNfxyWS
vByXK2STdYYP6ZajudTcRJkuUqk0KcEy2AnG9CNy5Up1TJgoOI/YiHZpDrI6TOJ+
hiP4QLVHoEeuY+BuwedDyHktgykfeanqflrtMnDc6YjO3Sg1ZJY+X2NzaPwUJDjN
fiwU7B/uLcVsJSqFEL1K/xQiqWNioSaMmnoMbmIurXsxzbpCJTPqfHejS4MN5vj/
/csX7V9Jy4E/bakm6OH7z1zK1Qa54ZhSkijf2zuKnMrsnxWB3yny9vYulBQkvsKV
FCq4TW7vcfYtt0OrE+dEdFT+D9hY9T0xqm/n6+df/wfVrwzoN/l0ku1zAMGsgAQg
jLzxq9PtPtM2t36SqfuH9bnQ192c+8UaltbE2MJiTFkzSl3IyP2WJ7YVaJAH6URq
Go7GE6FccXdXiwktNdFoWwqS/FVTnUVVfQ0A5MJaO2b8vdMbf/6ylKHAIr/3lyZm
wou1uIH1YMlujjh9IE6d2oLBC1ZdZ0O78ImJMs+FrFBGS1gwdKoESGqd4w3SAZMG
w82agvirotRT5TP8ya53tkLtNYkidhi7VVs5fcJBF4vAhnkjclLcRnpxD83jSwxk
rWLtc1QkfXXCNG4vcQFXWLjAYyCRlnzeSSgx+UvosgDorKalDdM2TMR78EzX9hMx
ZdmPdthwIlYDyHbGGSdiX37uwX1CO2xxuSjdG1Q8Mz4IxnKar3c6ka14MTPgutQS
hnIGvyIFFJn10H7BbWrFSjijnrlBZntKJsbCv3iGVBCTRsntVmbDk/dvSE0ra9CM
yyDuBsOd0WzEDKXDXzWyfQmix+tt2w3JfELbRDJcYTSOYv1sUoA+GQAjpvAw6diZ
Jiq9SgBcTXN5c4YZWYbh3rjoonCVFCNUUSUZ26/lv9wBiftnysvowbIqFwbBznW5
SVy9IpYSwvf5Bk4UsIBQn5OgfJNPIq4QQzyLt5l0a/uL6H01gj6EHe/gdaMul8I9
0Y7ofvv7RjpuWgpBmOlhrDDYZB1qRDiGCSL3+l9E9ku2va9IE4kvc/U95rlUPnS9
7+/R2wfvyNZHaI3xCOYt9wkxsPHrRoVQC3zd1WV0HUsaxPls6sdMq2qDeEEVjfD/
6y01UNiyW0A6l1jCPhX1+llT99NP4tjnYJUF2kGXFiXYqtgEPd7HwUbQLoz/g5gt
mrBpuU7zEeiOaITFdJZdkn1nUU38Vyo5Y7u/MyF1a1w2YU/nPAX742meXFu6W987
WKeIEN1qAEjhpu+U+N43R4krgkD7UJFB3Wm5+20sDEdHC7rZnijPryO1egZuMwYy
FkExMk3byHvLkni95QZ9YQtbLCHN7vDLGjclDeyM///sdo9vCR7pgh53kGNOKrGz
iCuZlYTZuYvjudwPtNeG/vD4kHk8KpQCittwAEEOTSlKBtvo4R4Th4uvVR9SWMPt
KFhHe8R8SnbOkXDlJYF3bSE/5orMhI2XRfTyVUSzFpoDHZgtF2fSAze1cFdTqEc/
/gjX058Vmy5zIgI1DBR+gs2QUbL/zsqUQ3zouMtSIt0kLC1jaquksAvjtR2lQoMI
DCuY6mAXMP9n8VRzUKCIJffO2Ns46NA6eV1Brek1WEYSnKYTjwfYnAKv/9l/ozHN
EHnIjSHqJCkvQEAgDk14RL/vLUdkzTPoi+UCsiQIU9hu88qmFRUiIJ8oJX2LePgW
bdszjdefprcTgT1uxMrhL4rX/2YhkzpQwFmBCYYHef3Fs3i/EMFGnRPHteKOSeVW
l005JGUC/cK90RCreR2pUR4skqTxesruADVpRfZp8G9Lu5GpqtqtvMxDLKdMWfos
BJwDd6KvGJmjUA4dRlYWkHssPqVrJsfEXt/HJcKDr2OPTQPgqcdF45uAcKAORPyu
fza8cZweqMe4N0zpr+SZ6ZLeE6ko/1A9wTGPPzqtk2BwdcBlcdoDln0zOcXJnjdu
ORYv7KGBiZjeaOb0fupDKt4686FaA9wttNc+FUT1RR0rA0OxJyWK8ZM3rn+L+3MI
MqbQJyu34Rm0uI9aabdz3CSzdTXkwb33EWGNaK71ukFtXn7VXbvT3sylflZ0cZXy
PLD3RVgaP2RzFceeh1l2MXIOm1URO/NT0P2Vqk/J0NlkpAu4GH5Iu1es1EOWJziR
6ANcI0OTiwm6THxE9MkiQ1FOyBa3wfOIJYNezgiOGHPyipR3EHQfGdvPKcFafB3L
iwjOdrOWaiBSopyEEnrgl8bOXxcrqBDTKK/q2QtK0xn5WWhR6r1nP382QjHNNyrD
QUCcRDH/Iak6xw0CrDgSUsn3M+SU3ytEsWolVObm8xhGXFzkepKaf2Z8SS3BsZJO
ln4RjFswzNNUhYePS+pgAye0psSBzgnMpOGZVa3aSkb92EvPmtP/5iP+3UTi20ZQ
yBqgu60wm0xRea2F1dKUi4szYODHKc10IF1AEi1AcDVo5emR1yQZOUEiZGJa3rbp
+3zsmsnABNxaDsgR0Cx+cN29xRKv1uihXlFyN86qq0MyDKH7Xg/OcUknKKizEUgK
mqfKQpq1nQACpLQ4l9VrEmNhp+JFJRRdBJsa2Di8HUHPwPa2rRv1fAMY3d7ZIElZ
nQuvSud73CtgGbdQ2IH0aZgMewSgn7mOSMQmkmz3o7ol7JG7l1iDWonl0DBOjPto
Vzu/xTWvn5r2ZcDsDAkzf50Ofi5bqqbPuSWfXBvWMbqbUR6mBM+uqO7zL7YWz1dL
ayzzq0dVnZ4JPsHUBwy9hWE7Bp3vv9ZQk842X3zSy0R3oTLJXNTtHxu2TtZoS3tt
5QXbhaPpwUm3yWQ8tL5+JwALAYTPbwPqOZGnIhE8Kjmm1zEY23yqKHdgIDRNqIcl
fmKbxk+/KwvUcJZ7CRIf77l0fxi5aIMnwl4Lpd7J3VusHAEKeV2iYxpzjiTz3IJN
lcP2A1hx7hlUYRs46Fd8hXQSZFekqo7l/wOeDEwRSv36W605CKsCOr1cgiFnI9dc
qzEanBP6rn8zStN6jCxyLnExvSP/PomMZsq9CCVlV2Df6VoeR9TRl0i9mEAk0t3B
SlePwq2hv/dfyiDoFi8jPW+aXaTzdBiThTMwrJp/8yw9lVMhIMFKNNm69TW0urSi
YTl7zY0CYZmSjCS9gT6ZJRgIJMP7IubsM6RNb7hHHrvvoZI8ojl8YCe54/GfTN8l
7DMQnVw46V4UTpMFDGcILbnu/qMGcT5Lzg51QqF3sVkrYG97CgHS6ihvBu2RwMxp
SrtdNsILAq5wR5fXXC4KmoPlWXYzvXgl8rBwQxC2mO0TKWmeHgFFw+LrTZsDRIRT
nKtnBYBfZqQee4nTtdK2t4Cal5sITWCOcqkidiDLpTeV0KBFprHrr1VW2bmhQxUN
AQuRUnE1JUZ2d5KH2VCULVOqWM7jns0DA5ASQrK8oud3i1tg84apbv8OkKaAV04z
/YwUUdrUniU3bCUpjmVit09JgVNhLQPziLyHg7JW1L7TrA+bzF8srjgXdROiUftn
nzSsZuM05ro0pg2nfU0nCSizM1rGbCwz+XacN/OJpbNpn9iM+gWAu2NIQpcTugs9
G+S8h9z4jQnCl4lRLWDFE7hItblP4O/zhrzfHJLGLCEBg2uzETuTJQjhmu1nxejf
srRRYFLqcR43Pe5GqV7p8WKmYqok2wdKNk0zlR8jCN8xiiphiWLtB9AjIxSPDxIP
k7Ap+GAfDvGlYZb7hJGwfBRHrZIw44vutvqR8uH5ab8HfXwgej31+6I9tq7FMBYo
pSbtOD8J2kPAOIgRwrL0hPv3miZt/7sEkWOFlcPTqchv4yiZVm67+DguUUsa/nx/
1ZFh8kR2qUm2Xifjsaw3TeoCtFP0nXSkIC4OBLloZv/x0TsnANf1J05ZLdCWRMBi
iLHslqKGw5I/8Ibjc6nJMnHy9rzwtEO1M7VG7VnCD6ZoksGU3fJ0XaWbR9rHqvpr
BMrXixrOatbiUwBfN7g8cYfxF95JAeB5Svh/pub59KUqNq8QZnQlL8rkZ2zXTEb6
sLHWH5nzC3+vRFa67Wtxpc/ljpFhv+v01J1W9U9cY5V4VH8hPhQzczCh5ArU3v04
7kjdMB5ZAq+XK6DNCGKgeACZ3pk9P34w9KNLu+qh7ITFG86dzCdcEjorqTU79DkM
t184Jf86o3eF7PJr0D3krwQuBrLD6BcsMGXiQ59EQlR2gA1hWb9d/ElVzhphAeyC
o2OYvCzxS1h3SpElNKUAdznEv+awGjPLhIpbsSst24n7VdpoyW/Rpo/2EyFRy0pQ
6TqQ9R+FtsvAj1UXu8GgmkL/5SDR5ytUg3MFBqiTjqxm/cSMlRxDozt5CiVIcFpN
/0OwJ61WOk4qmHvkPxjOPgNeH7MHvpYIMsy+ZmEHrMaF+pucFguDL6lPs5v0Vc3H
LzDGCsSHfFSwUgFulL/LWSHm0LDtMaJ7BNZHPv4w913SSWaT6Mo3R9pdnRhfIE0G
jwOoTS7gAcQv1gRsJtIBKtkbdsgT9oGlSUyX8F9aATce7971hH1saiXBdfXyo7sl
OZ7t3699Oc1TGSCWHuIJGllM0T8hEFDMB8QfPeyVmbaj28XXiXCMV9pTbd93OJb3
q4HNTbKocseXWHd3O3o6LzD/lzglwXysjRQO6fLzqalkl/H9KUzupszV7H+tA/Wz
HpS9zdjZmk0mkt3BHmEo8BixEVjPo3VVeYYaF3/iniaGHtCNiJWJIvU/mm8r0gct
9zieoVfZqnmSS/LzgH/KwZGskqYfGeL1VGLmkBfG8tlqAb8zzEwztIFij+CqBhTY
vOwmm+IrlxChZvwSoCLKVJidQgFNkJtpCIYO9TSzGxalHRwmiGHBI2HDUve7hN6K
Gov+E/ldOyszqPlptk9bSX9CrJREQq1sOaoqrgotocBAxKkH1TIv/8JDQApa6iXh
/nwr+Q5OqGSh8WEfzxomSrEm4EbVVSCQvpIWPrcMMpmsb0PfuteWjh264Nv4EcvB
O1tjbnm0Ff/xSl0BlxP1H/zAuxzI6IRd9OxYp+HELLm50MnLqOTGY9rRMEj3A4o4
uXU9aJ+D1Y+LUyQMtSVmm19jDn3lUJlfYsVgp6smIlr7/RbuL8V0T9ybTH7nAAb+
Hnse9/N+fo92jPlpsu69W/XjVoO52p9V6J9eyp209T/sYjVBakR9gaaXHdLDGW3x
BvLu92+YyWnaRaABYe9haF8KoDi1B+ZBPxono16UCRTwnY8n2pCRIkxnIa0D3obo
wPcE0YjybV8kWrA1yf1uRAx8jY/wPx46B+PKDbVtyMbBqr2O5blJTpFX73jcFcee
L/b6uy2iPJ+JXO72NkO2yTRKYYXqpxM/CYIOuHCM5z2QkZmA9WMR7tP8+OHjZ1Qo
WdAzJP9Kkd8h89yhTLwNZLOrQISAOiyyca3XBX2ae8XUNG3007Zb4RzAyn3thfVb
9zosfRbPb5vU1Kj352F+F6SStJVSmvUBeRuVmQJ9/4Geq+nDpg4SsNJydBjxLLj4
Itkn8cJf0iubirEcnhTM8EPG952J2ghi1+ZP+doRUjzwC8m3jMqBPDWAr83RDM8W
g2QeVbmvdstzDXFfpdqlaJSe2B9Ua5Lm1TZBihCPgOy86D7kDqsF+Gj9nX+NP712
FZgY8jZJeNXeqH5OperJA+yot9iPim+d+xWlxExkzwZgkjpdOJekXkWBHxBXFVU/
E++/vNGoUD2pNWjwzZedpgP31G6Uq3QLZRpEbZ0r//tnkuD90RhS7hTngH/bRRu0
/zEg271i5k2Vjbe71SKm5vC3p9o3eTcjxZYK+ErzuHnfC7bUInXJfwsHThGrbz4u
BthQhEqOhQlaMgvjyMUXi/JTg+KZVZiMT6wRqzBZ40T1pcJdwHABguT3XNcHNoU0
b1vrZ3cE/WeMOfk3KBFpshc3BcBWDs2TxI451e+tVAuc+AC2IMRwSWmjGGgkqP7T
OgeNzlIzHzzAlvIIjmXuMBWk23d/twnC/8NqhfkX/rhs8dhIbHK2CY7dxJz8UxHY
SwjO4NIPr2+O8S5/EPfl5Wg3BV6Oj+qtkC17uUJ334VBEHFnt4OzbFpmrZh/8eVh
4q9vyPUfG0PkZzjyYxwU2eGYMJSmZ4ZCq5sJE0Zv5pEu/vqT6yP5muGu5+4CUl4g
IcglUebbAr/Lke8gz78nwh6r1byJGHvbPb1TWegRIOMJVL236IC9IGNpeRbD69A6
epYY6vVMzvK+kIIk1xZu+pLXSKK6oc45ipE/9jvo/NBpYCaZqorMnTyIlXTjQb68
6XGSeWz7WI6iAn/4zIUe1zgs5Ea2eLBdiKeip4YOYD4XF7f27cxI4BVhF1UxoZrL
iZ81Ps99mdu8zJVWa6vskROywb7Pd5zdQI7q5dU0PiuQLawA6P94WTe8C9zoctPE
iSEECSwmiQEXaYdaIyfOOZ4KI2oT9D5caLMq6mfh9yMT83JTZb9hSV9hKvD5zx5d
8Msipr/atGVZCQT2T9/pTwA+zkM6xfZLlZLWlmiYjVaIR7m/9XJ7f8DAlcHGZJV9
XYFuYVlDf0xncRjELUELdDNhHwlxyqkTjH0XJrpyHOzyBAgF0+G1wSYkGZYsRMrC
3zLZUpsvu1aT3g3DLLpqk7pJlNpux19hRUvSQk4mQoP1XcOLYfC1Hmg3e/hjpJXy
zYmI8LpcpfD4wTKQASrIcon+DZLv2ubfrsefmzHgdVQEVV/BpXbihvAOYLKrgFAL
Ctc4pcXuNvCSETN2Bpcqfkg7fGnhz66hoPT5JUp4NA2mUCpQNOqKNGMPYjjp94kC
RbU2Js3OeDQI29nCF1P05vcuLIlt4b+S/xSPAfzk/g+zHGIXZE19P48cx2fvJpFA
8akg1K/gcPSLHfLqIcETk1Y7L7aZo7DMyQ2FRNgwMLT4oTnxfTMMmm62SBfNX6cV
j2NMy41TCgzzjCTO+0L9RsmgmCmcS/Rz5GSxeUaSm0TFHjDbBUXnkIVc0RFleXD3
1QNfNok09n2TtQ8vx5oco0RGCko5zLAV70+o9YIlTngyH+jff2/Eg1yubDWnIcyq
quZ0LNgJMDU50i1W5o82AB/lk0+LxXqHYkh3sRc2CGshCSbtd4ENq6ElLiyziAZe
mKhRhIc8mGkClXpcFHxBaQ4Ch6CIxKgsgep1oPsC0ls11r/vNvRW/zh1nbBxNdTu
pEF28pnJxdQNShsCxJhl8Z2nDN0vY9Rfrx2a5LVB6N2vlLev4kRxh9oLukrM7mM4
im8muwezHln8JNUqIfnKyImZsrrlJd8b/CN3GReEHOjAkySnTZsai+1RB7atEAS2
c5+A9P0Z4Cwz3G77bc08+0rvIeq9pkUVfum6EFjXL1gdv6gfoYhtFtPL5AUMk+Hj
wL6gXoDr+ZUMINAOQ0xwzluuE+CDoNhDxw+H6QLy6oC0uIhPv3eeFJjIZq1ksDck
SdJ7weGpbdUs7WHceNmNeHbz0pzbhoq5ghip+TE8N0tAnot1Qj1tkKofPjgKD9C2
YDCpHMjVVZneFtVG18RdRTtwvKZTjzUYUenu2CbRqnr3tET9nCenjYK468+0J7xw
vkrtWpADItB0HrucBMbSjA/+1zmhLabHPg2B0yMF9xT0tSxA+etIf2WEZOgGsslX
5UjlsoxiGLqm9rTjr1wOCtvvTWznAWh2QSU2IOuFYC1QpKehdiRb7/+/1ykWoQMx
6WuMPbW0df7D2DfqbtN+WNz3aJobm6vWI2yVgubLDvdqpL3Y/4Ss4CQvVcHMOKB/
0tq+CIIzjdwQa1yG6q4yf0EwSuNbJNftY4p5G/fp3QSvJIXuVlI5dYUB20GxCFAa
nzPgDydS3RfVD432LLNAPJfd9i06hxWaSpyJZUo6bRfSf0midMdFRTL1LCAXNPLX
Ukz1uk0cRITy4DQZN1fI9fwaqWU2fcYA6SVFYqJRMDqgcYKlMr3MJIYRRk1bhhTF
NbeAKwfiaSB46iGuGve0OYH6eiH8NBGzN5C4trsc4TTADIbgOp0GawRNGIo4o4bI
SyJKzQ63QV26IKFWi2M6Kxhzo3VbuFGAtQOghsC1Rt5Kpjvlyc2QfID7y+W6gRBQ
YuMsVComTbXigQ6EUvowJZmByYrdQVzmOg9nAqntXSVlYosAB3xQ1e0kHfZ9UqzJ
XurvAr3rMtqu0KGr9VfZhloHwo0Z/fYSzhQBWKK2kX33O30D9y61tTsZFBg9Z1pb
rKcsEYvQm71oZAFvspYSL43kAxHjYJ8/40fqjjccUe+pgoaHCR5ERNIAbd5MsTkW
iBlUz/ty3AOZRPJpkzqXdFVZh4DEi4T2667DEIBcAu/HpHziaJnzz9xf+q8IEsSu
gWwA6QDkSYE1kIOACqVTZAxn4xFjWgZEJCFqH0Ntu5j2Put6elTHfiFNYCD/RnDh
2WdZhbNyqJmHR0Pwm1rETz1DyF0GkmzUfJB54fDy9k7+qmCRl3BPRPzihJyiJRWu
wu0K2Jl53p+YIO8/JAGs0odptpOV4MMGHmwcLz81wfmAIZfT+NXo+wNnMreNLqbi
6OByZcbfJQIvTWcR87LiOSjNR4Fps2rQ1yNF50BCbVPkB2cmsvRterRBnWVu+bQ+
4PYlmys7fY+3b+GSxf+WPTt54ce55LicbtiODC8boGYHfzJOskX/BzpnXc98coly
yXsuFHHTeLWgD4qFkD4vVQAxjSsEE33cbkn6MgPsjt/uNQMjnbYOHmSI3CHaJhgg
j5DIGJ8CPYLxHGI/qJOgODiwpwrd8klvyQgIAd3Cr1UuDaISrx+hWMIxShaHzdOM
Vvk2+asAOqhsXeuoaGNpreePQmVrvHFeZOl+vr8mkr9rck/povX33IcPIZQqoFMr
7NMR3QjZWjaXxD8f7W0jQBT7849tnPoEiE8sVxF1+Zx/VwsWR0A6Cm3C9w7QChRq
bpE9kR3/fHo4/bAqI/QE1yuguIkbaiu24izbR6cQQ/3qeGetWb+0zVwtX2y64Rxb
t58kXcFoKLFMBnkhn7+oe8/rS/JJWRwki3Mvxjsf35m0s6zzu19+UM4Q+qR9IToN
YpuUlNF8+jjI7oVKb/TMsaMc3JU99Ju+F2MaA0UPlRtwDo5WPvsST/heiGKRkVxR
1fgaY4+mUxid/e/AkSTbLhT987epPGnqinAUDLLvBiCE7zlln+WZsKp/mGy1SJ9e
Mjh0966BqXyd6Mlr2y3HNbKjsQ+5CQzoPyJ5GdbUz5VFVBMalI7+dUS6HNYMZmtE
fLib37XJQvG7pg4olaO+VL+uW46NIbCP5+PbBKinVYh2D24i+uCPCL5CRTi0rqcl
P0aapEwk0yYB3zsAAAFi6qaqh/VRpLh3fYz7LQ6EbFJYGs1+CuySqRMStrQDSsi/
R/Oy3+DIXrxWSzc0aMgXFLiN8pszTrWN0d2nji2jOQoT7qMbg81lLhu8lLRHthvt
RAUZ25qnKKKjdFDzht1eCFXi1I9g684homwAxMLX9Ew45aZSymKCSF5xA69Fj+Uw
87rgva48o3uY7xSR9ABnv+ROhrMNbWowWCxR8SZU08WLnCzkm+2heX22S+GqlNpK
A34Zl5KL6+MWo3pCqZ/SNA0ytJSFpL7yEYLxXrJyLeAfK56BLkBGm4IphyCdfvOf
i2aI03/gNhtJi4ikJl4mWQxX5dtw8DTQE4ynizihWInCrHX8XDBFR+5kOCTxtdxS
SadmQCBHrWaYVqErQ4qlXOHPi2Gm7ho5YWahaf4VoN6oyVtdFmDndkE2IahYE7KC
rHuBMjpi4DGvacucUeA4nK3Pu2svMQF42IGVSYx0Ud+JIqnGRnXZUueEE3cxbzZR
7hOWaaBfhUSRnaHrlGm7l8lRi2He+ukFOio3+yMX0HqWSYKTDXzOvnJ6MEILMMD6
cd3RJ83q/vvnWVDhCn2Mr4/PUgNKjVYM5+1c3X529QYN6dYO3LzViRRBQknqWQxU
2BzQyWJ47ge9hpSzAJrgRuLHsiuonBqDnrxD1X4uLCUL/Lgnfv2c1MkPIP8QT4Xz
niPHR5VVgdiDdjne35gCbbXGgIrEjiA9dSm/m3hQZXZTsvnFs8Nrpyjww5Pmne0F
sEz8iXUBotE+yPt+5C3V8zJp+UEooMlQqtKXuH3rB4tPBYfFx6ZkGLwCsVr2MBYr
Hzq2XlvcEyjZNKMhAxO86wR2+UPYCN/ciXk9QI1c8fgtF4bpcVUl1Qu57IJ/wIa4
4c9Duz/E7cz1pp7AaXhyUDP3foNfsoZ02oli7qEIVWm3XYuN3eG8B1rwAjHCh46G
3/umuVCAOpExgooXl4QZPzpWsaGubMfTOwz2RHNLAleK4Wz+vcYY1027vvZHZ8UI
F18aUlX/PTtBYEhu023O8EwFPAFR5MrMMF5nz3bizmqAgWzVULRK6pun+Wj6Dmbt
/v0TwxjBjZSSkbK6bQlmBTCvpbTKx7RYoCiK1TQPlRast7MBaatROCZ/Zm05b4Fq
NTtAYcKKWkw26iyhxs1lajWsdmSV8fjwV2jN6bRN7B5fcY0dz2rg9zUoY8VHlmBy
Ft269T474/PqtNH3LalnQeDBdfnCyhUHs73oLdAy7AWmmgBre11Zb9EQLX+Hy/Di
7BG8cPzM4junDodBmNvmr8gZ8r41ei1IGraF4yunN36PyWDeCAI8MsARcjH/OskO
dQZ/TZS9r6HVbbLKydbLSqXsqMm4BHU02E0pzY/tvO+WGHFrDcTsZD7usE21lrJ/
9xMBRvgGXE6WV9Kq/QKkCZhVGsYKjkjy1Gun48YogePGlKhlnfwEg0c4hT3kZEk/
3jhehjCyJOLIhrqrSGMZxnruzaJjX8URmzN5PJA5L6ZXxoI1Zwl7eeRJRTJ7Uv2o
IPx5KZUV/DGS28xtZ4qP0+hx03iBkxsb2OtS2B9Jo35ymdY/0ipxnBC+F9aFahz0
9xL3ZGvmpM6ZrBK7l6mbT0GvQgVryS8WE0jam84bmi6AAOsmpH0779H9JCChtJCt
jLqB+6VrRoeicdH+BJE4EXMKQiJ0fkpdHU/iVyAFKyK3Ea/GCWzbqLEekbYKcsfM
aiCehYn+U1UA+aMsCmAeGxIELzAk0O9kWp1tCCrOj8yLO310n2sWnsmD2JCqkL7Z
kkbNiR5CjqW2KTCtRPdBzZmku9lZcPl32js1CsTQQKbXXWHZzr0jfK42rks9k5//
K2eTkyz1a79gfSkF5SVIkgJBEJI27UXM7HIgPu4kgHU61Op1UoteMdXgblJFxmcF
Y0w12DjLyvQyeWuQkH3SQAWR9mpjzqWO6T3hgvVR+cwumzno5KmfpOJD5Uq4u/rS
Nv1+P1owN0rS+UHsE1ATO9BuV44aMoRj1EyAIYklbq8X5fksrMOPdL/Tv8zEwPrH
3gDZka4G9Wub9z8CS6iXm7nOi7DqUMEb6AvMaEuWK6TTd/bLgnhGcsaeoBwg9zsz
qQOSctJ6TZX1brTqHLg2lx86VMxwq8IKHT2cym15zCWEQYoe39dYtvmPqvqaQsKX
U8YlNjW5r1Ph7AqfBXZSe8sj+ly+iE7LmmIMt0gbURHVVl1n2bi3MPiK6BdDnj5w
mTzaa4HvkjFB04B9W/vbb7+nda3NaFkf81CP71Fsr3iI0AIOCfaTmtQrnphWOfsi
3gDlemzP83AM2Ac2wrNXVDn0si1YcviuMgzA9/wbPT28V310zYfih58o5cfHgyiD
xDrrMUKN30VQQOIdkL5XiY6/zUe5EMCMZlm+FpwHY/Z+Lw+nkq3xJB91efMHII+1
9Przf643BJ7OIL1NwVIP2UEDESYDa+d5UdqJ+09un1Km9nJxp7DcCtbPGsTO9QvZ
6dzx6j6LjB83OJTGUR3XnfG4/sK/3GPoMZ2pzNRDPcEz8Z95E2GvGIR4k0IOEMVD
igmX8bPi3s/YHkgqI6wm5RMmdStFTaDTtAcg+SiEhoawPV3Rx1LO6mR1Da382/MO
QWECxWOlchLFkHuxADXdm9uKKnAFHSGPHvafAITI9c6WbkzPaFHksmg9inpR1LxH
2mAgWiBNxejSse5tXSTNWIQqpgswX6P+niAF7TxewrcQVotwf9FGJcU4innYa3/e
F5l1eQ1rnyFQYOWPuCbAHrhd7P5xuwKPw4H88exTr0wRg2Y+MDoHJ8YnvyiTaeck
a9jhjRHCe5a7T8CbHKF5Ap2K9UDmHccgURIQnr6O9MrfQKyECCQbK6sTJzYHvkOl
3v21EbXuKR/4sztMY0pLOE7IzYbOFXS/fBkELufFgr+Hj1bi1Ud1YIoHH84QEYGV
IzU7A63alJj9RtjnFM/kOVN6a/VSQmsIfJOJaQ5ZQql9SzPlewn19nRg1wb04JMB
9L3/w02xKNaf1meSJkSeEtwwyTdsnKdbImS4LU+GfZ2c6qC/72oBZ3EW2u8oWpT3
dXR8mRHnGzjhJBzp3Fv1GQH9nyC6an4aIAyk4NpkYzKMiJmPZyXGM8hq7uKSnn1W
fIvPB7cNZu2kUeS47OfYXgGy76Is53NAaHk28hEVtQfwtvtyNVJHrX6MT8HscLsa
U5+FIac4PsZDNLWpllwVuXJSCLPc6B2vshHR+BERSHPaMzY5mRievAcPpoITyrhY
zb1Pik9QFEr7q2YlUP2y642bVFnGa54pX0DcGmt2WbMYSW9MlO9W3ibaJ1s65MTH
URWdl9whjXlnWENrZAA6mMvDpdzHG2i/VcCKEUt8qWsTtNwdPjA1rHFxV09QIlLn
Ny1tLoLDOvptgBQXZpnHpdPDPBL9qMYM97j4WXFImJ0QyHGr5dkz5vj2Gnul2Qmy
+A3WWbTM4szZJlKW29AcI1ajTC2haEMi60QR07QUIY8/UwzeI5Y6VcDnWpAVph8H
DLEUneuzLBY7Fq87Sbfp+z1D+dCOCyOcfM3ZgKF+bV2by5zfOSSIv2616NmJLj2R
Mr/oVJtRdS/Veqw2MIr20XaPv78+WTiWWwZDZ4Gxbc4qWGVBBOl8TtwlDmKrr1KW
+R66+xpvd/MK0tYJrocFDJYI2rdE/MqGQwJTWxOe3MhdPqS8RgGGWoRfhWWz+VSM
+6cOllXp41Dk+q7TfcaxKoruiLmkWd7SgBw9kSzXtDjIeHiqSHlYm9SeRrEpo9Fm
dOgwSRXzcaanv5CHny45CwUBPbSFjM31LDreMBhvHdrrrcodF/PZGw9OVT2k663Y
LbGXwuiyn2QBs7vROlVRV4ZQe68s+MH2Xie1FCuOYW86Wccqbj8eeoP9L1+pigJe
L27lElryk/xGTeSmfPvDhGT/ZVgs/KNjfRi8p4TQRRUBtoRiQLnt72B370EfRMPF
DedqR+pEXYChBuw7G3Hc7H8P2NvKCWwgfMwSNDHxOk6PtO1x/CMCECWwAWPYMEk1
dhDhmqCHnOuLfI4eRbGDL9hdV/ATucEUpRnB1eo8eWZ/k+mYysMX8KT9xwYL8FQc
0x/Dbe/E6a/2LvvFxhHFF59W0ifRPdGxEGFZfOFPozFGSfeW0fsqsKgINUVeeA1z
eVD1DGTQqTiZvH4nJwbXJFTcUtoHB3GD1XJihMHaLHv3jzW4yCp4ln8AEYGYy1ZA
YbN6QyfFsQs0xPkvl2Mm/FcCK2r232FIncnvJxmHTD4V7vHZ2fyGnroJuA5ITozt
z63yosgipnQ9eBNVH/+szKVq1N5j9rW5g7hRRsOn8+JZd/m23Y0CO09DhjR+UxnJ
97fgerlT4OUh5TkMwHDLUD2RBC6/HD45k31z20geo22MPVg13pmWk5pYdi3Z9rP1
uR0k0+ltPjHgOuax+Ub1jUMei4xnvJhCRvimZaCJvn9nc55+Qbjkmxq08MOpHJXu
aZsUKzr80kLHLuRLqgZBIUfxzeJkS9DSFyofoxO9bbDV0J58YZ/9mDtSa9ZMQlyo
68OecYLYPpHhM1brw2JJEpUH5nASmR5+Joi5u7n3UVIoy9FAk5OsuDO+GY6kILAU
4NQWXn2ShDnzxNMEMHAUzRwSttqCzVAEbRmo/K/0ko+GjL+ilTEKKKtRk5U9fae/
9wPNgxWmQBW0TfCZSPA8jo4x1xHDBoZshvdi491628dctWH65gPWg84mOZ9jCuyI
Q9HwbZLvrUJtubevN3Zcg83rrUavPMhdTP7sG3J3nTPKvvtQgbFS25L1HRATL+J/
O7oTYMWQO7nyuoEn9CDCPVJRmPU+F+7jWmZfqa9GimqVYPskgWXS0vJWjWpdwFfO
XCAYfifz9l3SR5YzCjW2pgOgVtb03GP0wvFzC13Gfff2aw51P9ANOwXMwbYZbbun
AYqOJ69qx/BoBY56UM+S0s+aZVer3L3gbACzjlO98NEogAW8QuIbtZM6aT5yyPGD
Dh0sHCP3sxiEEqxORjoQpCgANiuOyhBAutxCgGeqT3UlP8iPqDDzCEG/gemeBpZz
/PTkQgDHEiVxXZpQvWLZFpBBZsui5h7f48HEt/BWlNA8NSEx94WErsHTwmdJORg2
F1SsW+cqG7RimPihnQFyS2O7Q7mdLGE0RnPfTGVMNQnBuNV9rUeHpqo1XHE6tdf7
KbG+BDoRx02A5uh44RfCGES4c9CidWQaIKgRmNL8bXW8kl9CAgpjEjBiT+WNTqm2
3ZKLIrQmHIn8jgIQ5TTGCnWwDh4757RWoOI2XezEmmZ/g+assPTDBE1cRJIzXr3t
L6c9kpqiwbPEeNnVk70DSP8heDouk2yoznjlRsAXKo5+Tl4S6x58U9x1qDl01k89
XTKJLyjZoZz1oFBIOPppc0dOnCyGYC9C6ayKmizY85B52kbPSRFtpHT4Hye4eyzq
dDFdg2o9QLYM5Drc+t22E/9vjZXZCa1bKN27CqQbbaC/D4gxVbaa+kek06lLk9Yn
vZAn+Iqa3z64DSCyJ4c850sMDIQqo4PfiHekOME1QBtBdS0i8W1G1gSC4XVGbetX
NqZNswhtUCbVTdO95hyl4MhYNaXMMqNrw6PLuBf6dJcjkrnhEPD7L+5gvYVSQrw3
NkW7bNFsiVuRsy8hfY0MrJjI/z2KXmQnwdJfyFEyHf7dGvwm/oVa8jmIAK7GsK+j
jMK00xK/H5y4UVosYwpVqBwGnEbP6uzYTyWAKmcfr6kCsw4NkZyHHuyYY8Mze8Fe
Li3VZYIWMCT73ICMMHTBm2dEy2D86tDYjgSurYfjZgxoOQX21zDh+fMVeS2LYZH9
55xP6K6Hl3DQQE1X4n79pFDMxnM4TB6KakUW88fwkVTPPTl2UFgA1DDCIn0SEX0R
gjeKipzbNljYMbD5/fXIu3fIXwtz5tmXqzICQZJAOCwQfHslB+F/DDXSm7TkmXZ0
iIHnnARBAkI3xw4L3y9slavlGX7jI1DKFiwpAGTxzis003PLgNOm6daLTDWlHoTt
g3+biDwXyCv7kTcBlrsRGm26+tCsvfA6U8iX7cfgn1NU6yk5qcH3yH+n6Ka8yJRw
tMZdSMMZ5KNoGCl/QJJki/S/1CqeBIxV0gWiMWTAeRDvWRwt7CND7ki4IbqzCKkn
+HMFrYycgbeydtwZcYA+TZTRiiDMCWA+NjWdduY9pwBSofl95nGpxzlouxe7EI2x
RRs6AyJQ1b08SWE0GjsX6uYWCl2fdLWiSi4SuvMabXmo9LWVE9Po6xbFLkMka6tu
n2yLOK7t1iryyDBWdaTgYje9P8LM9YuEO1426uYMsBsfK5f5wCvQXLvh0qI/C76H
iDP5iVupxLD0xuGhUGvLloP62pK/TtN+pOYjjVeoSTZAorgQBOVlfqGmscqyfxEO
4XevmtmurkiEViuPQTBOWv4PfsRQPVTCSH/cQB7JU0gkJOTDDmmmTbZklAHmZHfx
PGcWt1BeuLoewHaLlJ3yYgeUL7nFZaxdjzfgT3wmK7+nrUh9Bd9ML9i+d4ZemKU9
d4SYHgKQ+84qT3eM1EWGiCQoBa++cNiQl4VAEnkx499hE6ePpruPJg9neu7aq6VL
mWH4/rD+EvrqgKiUgWK1FWIxLGH41eUGPr29ucAYnIPwHCirmVcfJcwLhwE/PNX5
xo4np4cYh3yJcHB9HMJBaCb+MNOXwViG/fBCL+CBUTJaKOGE+r08IsR5EqisEc1z
7ALm8lTwoV7X8FsiOcPK+J3zEthCqDLKBFWfsY3L9B+UeH7CA0Z8CeHZv+K2uxyR
D7fZKBL+JHYRX2XYNQwu2d3lDcw4vFB10QO7tX3WpsYRDnw2uPTXwJXUkk8K5YWe
/N0trYFtS3/1gj4jgXfqr7Qxa6GeGmPVAT2tFAkzo6gzXsBqIQWwu0jrBM3n1LIf
kCstS3WYwV4YMkjqUv8aPnGv42xV7J6Cje7merK3ZVffPYC6jHl0/0rL5lQktBOv
EksDKN9ltQv8wKhgmTVbOAqFLrA/mrBp3y/2lC+yqyoPAonAVDw+42VjGSW6jhpF
1nbvwzUgsdvtwbJYrUcw6nzQ1Q3IgnXR4Oq6YFLaaBYiQJw/xswMDMjtTcTFZpu+
XpOwb/aBg7FoM5uFvy5Xhn/oQ8LVpRPi7FxwNfd9UTW03WMAfl/4kI0juMOVzv8f
93Jqb54vAf2AEb1XolOAbzauY8tBK5E/oF65S0LVxWJ5zzezDCAKIad0xqEac8Mc
3CCyd6SxidocHaj7Rw0G9idSfbrxuxNi0eNUSSrN2b8drqa6NTc4/+diMbPY0q+9
FbCJ83WtQRjwi4c5KvlU66PtG+9OGbQcV+BQ00+iNypotUVUsb9EVTEeb+8kr/TK
7sM/0GuqKvd/7VPIq2WMp/frjJ0uMxIXiqJCwtZlgF1+2GYmxCRFleDAcwPNYYe5
GpAOWmOam8NAUqGDanzAHrQzCF3NW6jyqS8VVGMrR5GRYW+YZEHKm1AdfaSMNK86
P8r3brWGtrZZboE5ZmjrPo0YAntRY/zhq09YQjcp/FGUAte8EWZ84jqOhfcgdg3X
B66IaPMb9L4dzLcWGrzGJh1r9N+Ia9hR8RYOtBdUv2ePopKAGYRAVSBsSGa4whna
uiGExRHzsEQ3JpU3+xMoT5F1Gi7cvO+QaWUFkw1qG1Ld9QIETvz/HdfcwTUnewDO
gDckwFMYfo5Ck86Cy2bstOCOLWQkvzjjo4/xqB6Fbrn2uATiHXHS13oTe19p9khU
jDbDpqniaimu+OvQiSkCimFALhFg7hQWgsiHyy+wdFZfJNnLJACZC6vqTQkAlcNW
e1GMURv/SJTiiFSzj9Ylez1WV0mPAoMwJ6e3bGq3C0++4M6hjSYon6rugD0KsZAB
L/U8H+GsKjzqN5k1qRjHAOVQ08Im9fQNybdrlgIEeLeWyAWsrbXHn6ac/Kyc2/9g
m/Ttro+itfO7HaFPvk6TVSeyHi7vlD85XJyTo0VuHErEI9vIjbL7mC7FTTcnhLM1
pf2gY/lxZB2f0ZDJQWNf7KfeA7N/eEF4a4h//j9gnCF3AY4tsg31JXNAq9dbMAFA
W6UP9jn7n3lK3VLS0d9ZrQCtoyYCmK3TWnLlkLW27vMZozjaDGOtaoOG5qOqyvm6
OSOomZuXHdtfMAonYoc/MRHhwu++LhJKoMZbg9ycm0E8Sg4Sb8fLUsmTtOJIi/3t
YPE4X4zexr6SM9PL31Qe4u3Cd4VxPfvYgt0EzxtKVIof/00JTaCw7JqdSSNVxovz
kcpncsXUFYtwAius6+6tLnLg8r9lqQILhAB2F7djYneZtiTYRbv2daQYnJpRho3p
EItHwJdufeR7a0jFabwVThly2mVrJLLTaV0U2DLPjren7FbtVd1Kk0PIUFIptXRy
1B5exFmG+5k59KuNpEpl4yA8zimEmQK5qgfnkJ5jILI5PasDpX991V5AI0qwEiXY
aYGS5NVxdC89Kmt6aN2PDZbCcjJ9/NkZ7phTrIi82VcLHUn3IpZqg1W7XOc8hlAJ
wo1blBk1xR+OR6/yuUl5pyqJf7jQYZ4Fsn7N8VDq4KzjZ7T+I9GVmTCNWyyblE17
DUd/MtV8LCZI41lEGvcz1rOEQ+VciDhGn26+mfLlgD5l5GcdCUexri/o7p/L4D0K
3aIioCGMS64zIyVDa0fx4sPQjVCEvRYgsb4c2KYFxr/3AK+GQhQEEInJ30ZqoVpv
CJ/SCopUVOZ/YNP3ZfyPajj/u5ItZP4PEme52eH5yoK2K5bDkJ8u+EZce+bTpxVr
8k4vcsf15LnWbXrwDdRGl5ib0ohdhiAdcImRQFiICCp8852mVckAWh1iRFNqTI3p
QabugMArxdsicT/CMN4g9EsDh4dYIEHnlJgMGswiRFwlPQQYXrlu8b155dQTr3cY
H9mGUVGloR3mGKPFPU7CVbxPD4CN5PfJDKEMmwDr2ZtuMZezmQ/SlLHlp/bSdwH4
sl7fGEvvmt4MBvjDRgk5dA3BGG3mmMMGfyG9BQQwWblIXeihb54s4+Vs3ABQFgaS
Cqni/l+hb3hkylvPNKpDlTb5tcbipcxX30O0PVh+xnE7Woyo6W6uedahyou7eCrA
F0NWRUVnMowJKWmnN6K6BMvdZJ+klJ09Emqbr9n+u0iCGM7ce+upXguGkbE9fyGL
fdHTAIjPm7vsNuVJVYPL3qy5IIOg+statfac8UaXvNXIystXnWriHyCUJWS9WkLt
KdnkzuN9Mnp/hHU406WbW1xPpqJWkw8CemE+ra2/ElCGjv6RemCN8GjsIH3T7oLH
3uSBRjYFPqvMovW5spqVAh6C8CneZR9xf/6+c5st4BHNv0cODNEM5Lg89U5ukRPz
vf9/4FfWNLISR/hpfKZXyKLbsP2dvQJXXGflXhtNY1o49MncIRs2/GM9eldlHVFd
SFRdq0ZK8STC0q5Q5iOTiSVgeAFmBTEHckumetVvmk9WiEFlrGrYTyOn2isousXQ
LpnUFCmJdioBKt+2C5hGa7CCjSo4iWupeLSEm6ADYd47+I9sTpq/nndlOgk/v/yR
1GTa4TbPovia7AfhrY6qLZHqjcl2MnhEFndPTkuaAWzWj5iplV92LXoi0hyHO3SR
9Hd0hIDwwnzDfJajebtKISJxz1ltBYhfKGsvxo9Q2Fi0rb5PP7mSJCjlvLIpgpWH
ZExjFJC5hlpprBxufNwwlNcd3/DVK8qCZT8rVATz1WX77Zzr9MKE9Q7j4uTzOVUR
HoO2+GLH0aT6Pl90brOJ198fIMypDKNqLtxujFySwmqtEy5GYw5BlLxT7tUg5c/Q
4Dhniy6Vi3bKOQfhwayhQOaNiG9CcyWMxNYRI6rZOkw+3A6o9HrBwrBFGjaFZ80A
79lt6CD+eA4av+8NC1W8peQQvx1V71A2HKysYsINpt1pvB/gQRfZiOQucQm4uZHr
Rcx7hNPoG9WErj0ANdruub1JKaHL+ejRJnT9tlx272y/B3mJKdQyR6jcFfXATakr
k7PajoWsJebz55M+CKP3QbrfRY6qOprPTLqiOFM76ktZvYVGm0U9KcGLF6gZA7pJ
K6g484R4fGbI37zqWDTu0XJgBw0sSRjnh7F9+2ZMPh8qHKRnqYu5Td1E4zkdPz0Q
t5gPj6BuDp+izbdS9XevyKm1z8IkgN5cqPWXNt8M1SiHSKJoDf8mmjwqj64SS172
6lXJykgeNVhZOtPlqcJd+XOBtDS9Ow6ehx8wOIl5k9qpZduZejcm36kqIw5vp+oF
qXFn8/W8yNNYU9uISgXcJpOkrOMHY7PNoOXXDGwvhLTN6zyXeeKWEoKOBXN+pPAZ
ch+BPhSFZlMaf7cn5jiWvCy7DbClReFYMz+FdzB9ajV+DBVe1IbiuB6KB7aVisTT
CrHV5GAHLGjVHxvPcUO8IAVIhusPFF0yT/1ZjTDpl01/HRuEzmu/GA305/h3GGSf
KEkH1cZ9BqFT8UGrwkJXJOFxMag+kYMF2nO4Shpc+dsevuw4Ol4ei3ajJq7YosHZ
R0svB0jF0Y7qhNVBFD/ydFOmRrWy+A/N+2fPtYVHVVNZcL/h6Q7pjBQO/ZgQ+xoP
QtQriLOarQkbvG7m9Hf6TbzmHahz+DPa4S5XEkh2o5fBNhtyX8fWw6ZkUzOWB2Ax
mj5r+HovsBWYtfNu1bzHXGOSgDw8WHZDILyz3RVFYI5/cElaXaDXSD50IB7FgpPJ
DOJmaklYvjDl/KyFT7AHV4QQPPOIp2qJNCvlEmiudcwHYpDe/ieHCa9BmntCTqbp
K0efn96PB6qH44hRWoeFHGKybvTrphLem2+MhAA4m8GMnPokaV9e+6iPJoCczytc
sxgDIEDIgSggaALi7J4ORDUcsQbqYJJgCxnN8n6X5H3E+j1W3EKmCXu55GkFY8K4
FPVAOFHAJ4oMLKY/oMsaJ1+gO4zQ2ZTlyz1rRO5wiN8Pr5UhTT5N5rpVNWYioWK2
mnW1jvInzOlOzW5IZ58YidvvwJKuVf0YI57xQTRvM2Oz6yBfoH/Xwn6S93NjxEu1
Ocfq53x6eG4PJN6KA4uYRcZNojbw4I47nz0baN7jx13Gbek4yQOz9L0kU8uyqO3m
IAp7Tu+pAxhRwGyvh3QcXN4WqWzYSWsMgD/7BbKLXwqIICMJaEd6S+cPHD0zi3JF
qnp13ZZ+3cf30dfrCDbT6BtdWDWYsSLJC0x34Mqzm3cgAjRrYzlWqqmkJ/9tuC/g
SNz9J7LST8y7KiuUPtUEoYk0RFqh+oK3IxqkUzx4SB1YgFoMQEimJz47ZtIBzaBA
/oJ2a7eywYE8AEGhae7sY7dMx5Btdoj/eQA/ZUsdPXa/AMeCWhbvOIRxKWa9Ytbe
vs9I09FTQdByjTCRBXc/fMWdu8CI/oTqnNF8xnxeyVuk79oiB3/RcjklhulZeL8B
ntAGFt0uVgoT0J/dkErV+oOflJaibA/xqHxxazrDv0UNHOjLMUyZNLnBuVo5vPlR
sGgshJXfYitBm6YTLEs1XFCWoKK4QPtvT8QTfQjP7myykT9PUqfyrxaCkbpy91Wp
xlWvwXmAfwoRiRxxbxG2JwEDHiZLiXq5qiY10j/SwN3fCfeup656Ctg1ISVmHiPd
IHdWZ4+0H+zpipdZ5z/n8ZeJGySAnchlfDc1Z/6Qb8Y9J+ouu+G0QClfC8pIdSwF
BOC1jVwpkcBaaCdZYMGuSgRuNGFPMlwNYUKswIZDw2xjMhyHaBGiaTRRJamDp0dU
nJHvjUM0wHEmDy2cM2C2wHjFP7gO1psH8B4FsaESbY5rfgfb+hhER47Imc5UqMCk
APWhZEh2nmdc87qXeQrrwfVVP0Ju92VLpeFLYSc+bju2WXs03n3/xrM5SX1yxAgA
843gvj2HtwVVjoeys0AK0ZELo9H9rRiBX5C+09/RNaXpCerCq9XvF/nerwUfTlCH
u6kqA9LZdszGr2P4EmHQ6cLzidc9l8KlonS3Zw2Xg0PCAczo7S3xgRRs/d8DMJUv
VnmTHht1zppgSoWxkRkfGp8nOzUkCWWGDNR0JKdnTwkj8I8sWKiS0YmtkbHRun5U
RIFTfRzPyv08Kyb3hwvk8SBkkxxl2+VU4KOe1olleSdFK9SEDK8wbXcxns9I1I7M
DP5i6nkmRzqy9U+/J01kem3FTkIjLg2E2qIamNx0C0Z3CKotXN6xFHxlVysvbJyY
gP13IzilIiWzRqW9aXFqebsbLn5cpivRBqIIz4MAj17vxevVoP+CwF27dT4L7thO
gEZmydGaYOdv6d4v+CTypNOSlpAOc0vHmiu5ut0J+wX7eMdJ6LbgUhz7c+wMB4i8
BgEFbaYoRdC7+fXEg2zLzyu9rBSPMzLEQqXqVW1/RAZvICGOl+WOexv/MOChq4n+
6BS1MOwHJTH9NiucWzmNEtThE+g1ocbpnjMGEZEC7pcR8QqJXZwEIRg3aVZTWNoK
U1pn8dtJ22Eoi3SGkDHmSpkabha4oOgT1hgYdfrefHf0ModhKh75ppxP2A4kAVZ+
Lq4ZsFy58q78IDIyVsePZXd07Dy7SEjRUvpu9FnpNFKytME77cgYTh/3pPsU7Pyt
PMbLnMpK1G+Vb1KHRVj0FaLNDTbu5HGRoGJQd0AbJC+ImcvF3oz1Hb/+ujDSJZut
QDe1um7bcyj8ohFktA6xuk9hCn3amNdPeU3SExXB+zMe4tFT/zOuljkTqsTuDUCx
Hc3shAMaWdRKejCHVPpdtGvzUU8j9ru2zmqShBYmh+AeejZmKr7807938vBvo+b6
S6vW+r1OC8CycdWl3hp7OzkD9SVv19VXkXiMj6fqHURBPT8HtAmSFs93TK5eHAsj
xIAb3nSaHIDk82DzaW2jLFa1C7ecI2iI+ZmQ8kHXEfMdVzex4GADA0f9VyhRxq6/
MN7DyXU10F+RUfGe5in6DTidOR5dAkEZPit7kF6UmhV3hAogGSKW+BMqOD2wV2Of
6e7AiC2D591XPwOkC6iOGX1kXiW/mKTRIZE0z3W92R+LFU6MOtEIptnFKafn+sYL
HP1an6lv0K4aKM+cn3+cqtfSxy44paflYrwsc6g/EINeKsQMLaSzQA+tU9UZEntD
JpmB09F1DWL8ZNgBChtQhdYF+HyTCKduM4D5FMtiv2RvKeoicRtdmEP6dswkCWl/
IgpUNlW4Oh6iP4UXXAQ4AKiM3jHgLx1qqG6D9XlPqd+9t3ycgLFAVvrubFbcIToh
SkOqvObrc629xEZvxuEF64g+/hNFYM7Mr3sDn6rWlsj8HxwO08ljcAR9GWRvT5qb
dCD0soIPGFfX9DkcwOVLTsPRUahuMEJZoH36D2NQIDmApUAGTiYgUmnOsfuFVJNJ
LWfP6edba/JUesipaHLfg6Qp3ks3dQcR1yonYuPCCcJ2MzfCwJim408Ny2z1kDh6
2oOjENkK6sc2PWUHaDa+1Wq8JB4YrDeVWdgMS0Hzac79XfgyRFhlGYZnTfHrHRO0
g4yDmI0X6XdGLn0C1Nq/e+GDUe0bcwyHX7J7T+/sftZ0+wE+XpDBy188aKv0wupO
pzZbbmwkvrb7q5OINzhPPP8XPc5/UIgLYWybYPmR07LamLQIV83v51koqOtnZy9m
zi2daFX1Z/ffQPGWz1FIOSyv0ILcqcI0Q/yR4cj7oHh885CPYSZOKd50q6+w/tWP
/zGLtb0FwHeYZ62IQ95A3xL1po9p6anW6eQInN8PjDQF55bCILFepfDUGwcyqPEJ
n4Qic7FZ1olYoGZ+IpYaeMqAb13T6dtb1Ra/I6paSlNizpIeXUPasE0FB7HA2jsK
0hAKBaVwu/YRVNL0SYqKQVNBAzr+i6l0IKQ2eGF+9iFeIH7SG1DCJojBQT9Spo1d
31ra8vbYrCCVJVsrci1oybY30EQi9NQnCfLSxKGNeeiucoq9bFd9P2Nu3FyG70nG
UGJceKzAkX+I/mJpVepwYz2n8hsiu4idVh1S4dVbOHdEmfTK/nzThFcZAiZxGb/H
oavfOVkQS2MTp2PyVCXgHNaETiKEnsDOnvmlFnmqBz6OMXbVAtG8CYi8RBZOGcxM
0CqEP8Tb+jq9NFL470PI54yU/PYQFzUXZbA4DrLCItLAiHauBOls1QqGY5TLQO7u
1Y/2ln3GaHZVnkYEvZ78znBv076+Zx6ZnbuE9EY4YQ/M6Lu2IFnZ3h4QgvrLByeR
6eJFhN2hPvwMPwBTp1PviC0Tx6c2UMaSx978Hm1g/Vo/94HcxEwsk9iTG7iVYAbN
d/cQrgjJ8gnPI7kVQF21s1aOImeeMXHdmvgDZEoFdwO/P9gQLrObbUAQly6J+eyq
5Z78OrfMbyAEGLw3LW65RybmeTC9w8qC6zavGCNq++/Mw+oTL32S95os5mwtbAp6
4CmAlbxxo4ki9E9BZL569a7etIfuMiJbFK5IdOEBKfG34wwS0yWKxap36DuAEphJ
1radGUIaZgbIb/YZxlSbYL6qRcTESapTL6Y+gEAvvr/Geuj69QAhvVIQZtyUbPeM
/MjzldLwJ3uYFUcpLIIUVdNjE4DBe8hLgXL6rWFuNSo0zqgEfckxVSaiNhtNMf5q
S1qGxi/C1rTakVL4pFjAvOw87JbbcE2mTRRRrjJ+/PMctwp0gi7gIRstFXGsAzbr
7ENM4Yb+hv7jaWpExw6xgoE1dKvLeyqLhGNlmyXSA1lfUw9iiHB4edU58ZXFBsXs
uRLdDA+gacB3WgWa5G76N8+lJbQizGokOWiHIFEXzjhvWsOkpP5IjTBKyw004waB
wjK1gB/OXUPjMZYrVoeRvGbyeh0rGFfwnQpLwxWzdEgM1SaR7dUVOI1J6p6IkhXc
VGnBi0zII7mjCBGmdSI9Fb1musox+DsMzmQMUFK4cmux0z+vyG9tPEm9WNN4gdTN
8gAXMQESI6lw2zB8Tv+StaIOTGlfp/ddvC7z2KPUgpisW8fk4D94Df3aI1BwLZie
4vLZKgEW5zMu6JyfCOpHTyZn8+yJCmX2qqLJuElc0vN9jrUg5D2mKb/P0cHaWoTR
JKrkge1CJohY5I2GZ2J5Q+Mz7L5ZfQTbJgUYmzLPMIucXJLQ3sRkT6hl4kr7Rwjs
ZoOaXYBxqGzcvo1ZqZiAnfJZ5sZUpQNsaHSrCOfW6KW+zq3jMz2p9+qVRu+MeapN
/9Io3lc7f0FVRsp7oUDu4MR8ArOrctxENzdka103W3xmHlIgB/UUl9CnBnlKHYIj
lVwn6xFB9BK2YX9fxT2TJXFIXsXmY1kTOtS0lsDtOs08hdgTniNhlDunFrLs0Bm/
aFCx9aX8aTRtWOFrnciS//XAQXYx/iaR2X30e0gKCH+NuBHarBcdmszn51K0eMrB
TVKui2GyPKD8ZQYc9wasAIE8GrJ8nWtfRsUgwMcx8ucpTl+AElPgODnM7rJLwVLM
nYeZZDokaUMUrEjYYtIQkymURmQ2ZIdXP4LYJ98c6IphYTJ33IwUuN8KBKLckHX/
0+rZPwaN+E41SZIoAQODHbKECHlWOvd+IjeIjJ1F61BxXk6+Y8rYF59R2MdJ6lX7
Mse/KwSZkwMJfs57vE1SowZ2JEJXDmZcoE3DtVKAVCfi9Xh0A9aoHR8M5ViAvRar
GS8raZPIdSGjABRnmr0GI4xVFlzAnKHGwmBvQJ6etp8lxJ7OaIaJQkDb27yJfXSH
+LB1L48kPS+iTdCcXNZ0ALRCfgja+09aQflnQaLQ+3d/pS5eJUye3ydEqt9DEt9z
fyev40mTulm7mxCynyRNeKKh3dQL4T6SA/lzGEi3ZvVMi8PQcXfEnZWVajIzMwZ8
OoVtnW5pSNDoruSosaeoRFUVRFRk1cYSu1Ww9ZxpkzJymvK4mKgdQiFPwPqrcNjr
++BorNwQJJVSJZd3Gppl6zfZ7/O4Aw0x3qNu170Z/Oi1Jb0BuO2GbsLFTy+kRtWn
bNzThVDO9SCTFV5unNxKdIqCXpmnqEJzOm7rZnSy83IiBhbQj3Y32k8Vtcd2e+cR
uiInk02BROXfSDGg9ClXkcTSrJtnkODmW+rjBJY1OXIWVW5FCq3IApkX+Cku5N1E
w+7T1HyjCXNyhytWNI4OdyObxVA2MkYUBhinO2YaqE4k3h9feCSlOgwMObIy7vzh
mRwNn2DbfOkhht956qa371n3jvhM36ZRTAXzv9M6taF7OqE+QMPlCDNsCMRfRGda
SbaYzU0skGWlWdeapO/2ynzy2mT6AqBNMLR1VuhVnmHiDSwUL1r845f2nsWpwP07
19o9s0ysGRSl/uJNA2piQ3GVq2207UQF1k6F4THB8t4gmZ+GM7JVskcXO10AakvR
ubIcuVX0tudmWlWuJfO0Wio8R0wByRXq5r9Yx+NjKZXqP1Iz4cZwcrr5k7g/Xl4m
tmsmyjXPDzeDp6g6SvS8+EI/CFA/u2Ji90aUDJQXzg4VDsn/uvOP/0vyzY9yBz5N
uA7EqoDcdWo19iROAQQ6km/wvL5LcciqcvTQ121azeCB56OPVQnvpJrF2OhlqleY
ni2qMV8U2gn/RH1V8lj310i1rvqPNI4vLnWymOXd/KAEpnQldlAgDss6OXZgyqwC
+fQ3AxJV5svjv2BI3KMkmwnux9FqdD6JEJEZpct406HPRW35ixZ1iVR4LuNn8Ewm
uBDUa3e2BjJ+p0QwmQYp/gUSepq75lx33dAL0ucikZqTIg4IKYsvso7xsFJ483RW
boK6iRemaKhPn+VmC7qvVkidqteqv3y/vFDctLv5Sp1N4sxgViKd3aAT1w8QBao4
5+pke6RVo1M7BWznPnDIcXukiaUtoNCz8oJzofp/rrRWYRV7+4eDRvE/0pG6ZA4A
/8AEe4fsqV3KFa4cpxi5AOs8tGh7UgG+cX8LoaTkMm/Q9abWwY5HtScEEojGP+XS
3AUv3PConvLaFWdt2YmIVrcYGScwPhJouHVgXZeCzE+h/biMNvZoFPtf4ej/Ugki
Py4L/eelhx9W4I+e5p/JiyRjeY9d/70M6RMGDBWXaJYmXx9cDvs7JRZSkuN7nZxX
OpA9W4oQ5XslVqzfpt4dmMA00oPUp6a+yfR4hdy+RMoCGxbwdrO/JdZLQjGXTZzN
P0DnXe5s+nDH0kFJkczBEz2zSMc7X6c7SrZRrSjS2uJNAhVYE1e6W+uaL4H97CzB
SbCQcrrZ7QCetAHx9Ji/MsqwvaSquSpuOq0AC8T3dkyjCxIt8xfD9OaZTp1hEkcx
IUEqkmFqmPASCTfP0YG++0nAdAylFmSZWd+S+Me9DnOuMJ1VimHTO8mxmggDUx1H
3F/JTo9b3Xe/PWBiY2w6EDdKnk4XVpJWrDfTtRXfC9Mpfnn3J/fnnWMZ3J6QjGGk
29X/LPvEVHcXEyR+Os3+PbHaYUDrWKSAP0FpIm5rglNxuzsO7U4wU+5PHXNWlZ08
WHef8Yibk7lGVBmxF8jyXKvIwidXhmXon2jltD4efo3Z3P348AgSOthsIEqGZIez
n8kwyzgstnLNP8InEQ4awiaBG5tZdZ4wmikzwvj94nTFLOhSLcVqJDEvM5bIQMpb
2H7rAYL2sGX/uYJKXal2KlPieAuXPoA6/IR1Oylqr2UKu72UpNYNrXs801hPKoy7
57MR5q/G0IvOx6YmAlYcgqgpaRRoRbnNdV5CAy8BSfGOc4geqRkV3eYzcpVkVuh2
beCD7Uy3k1DXbzy++pX5wNFgKIBE3bC1hy8Cj0cZrTuNniMBxOowZb7kXh0VSadG
lzh7IbhnVdq+ZkNqtzpb0E+CaNUbWEG1SVoKzQHyVoPqdIA6hnQFsjI0QpwV4m+9
ISmBSqxweSnPoXn8Rp7urUwsEhDWZty/Jfw/kbG/CMPlN9EoYMSBwpMBABJhjIVS
RX/9Cubed5nzxX8tFg1M6e73biO9mzClXrx61iLVECybxWIot2NH1j8t2EzQ64VF
w92DDdEHfKr4LykmMITSl3dInGsy7Zhhm74zc/7fUH6ZYU7S56m2fwhFYzAiw2My
51HoMw7pTWlkIzZk/fZltBwI+8qJdnZfpjnuK3392zQSn1pTDyN90oWx5NjlNoId
ZzB522MSwX+OAQlG5EGy1s/BZqs1RvaUV3SQugrSc5c+rvLIr8iJdHGGLiVAhPNb
CSuPz5bTfv9cVi9KGihuLVfksdDGC6lb3evca15s3AIEpAOo2c8xNSQM4G82pO5s
3f22xMVnX40d8+QcPhGGyowuwy+2Z0DJqxY6hPQ9JKyoBEX7ey0SO9GYImgRTkNc
inxaVeen1uouUBlDZe5D4N72IBRGx6EYqxhtUBdrmHZXADBacLa2fv33UpQVGWVE
ldwRk4+uqv3Sn09LrWszJqaBhVaA90MUGqDHBW40nq0TRk2N7CsoKq7UQWhAi1SX
v4eO1+1ZJcKwdO0ekkpjQwwuunj+g9Ep7/imcIyDk6teg4vmmmtlWdX6e98DBCqd
3w9CbpawfUXap1x1KqWcBghEAaQD+5Yxg0F/7gsHNKdc3S0xGLBkAMxJMJHY3hit
Hq+8xqR7yP7n7X3e0CYHACpm/KtVQeD2ln8hUrFQLWcePsViy2UNVF7dtaMVPWo1
CR35c3SMldIgmum7wHmlr3T4PITWY1TmIU5aRqa8BpBkvNpRWNYj79K1DgYcuyhk
+rqiLypF2rfXcDgwLGMOpyO7qYYqWAbo5waJ80IPB6XJto3dcrpFJzEf4Dp5XPkk
Br//cz7mzHmnTSNFz17W1jJVdu21/zo3ZycBu+O/WP5IxvPbC31qLN1VtnF3jtQS
76kVscjUuz/4K0snXVFAw0hDkPL9YIObNM/GP3M6xzxxIAz6uoeTjiKszOShZr+P
qw71YHXWp655jtJ1cfW412Za9+DNPtRBucoT1Km55SmC/DaDKC4bZfWXKx5JILzH
aBiNVHzWRdejSdNK3hVGJSv16O03PY/V6ljJ2jmZLIhEY0+vFHKCfzwVEIzTRdyL
xecMqfXBVy4a6lMsOWtUJwJnDzCBzOnMAWdVvCfA/cwrx1BjtUZvF5pCKso/DBHr
qX2LwTJXzXF1iZpHIZy27auDDgy4rHTT0gkX+Nx2CmcDQN+wIyaQUBkFvcnthPlk
Eu1oh2uFfJwa0NsIzAGE0KAWKP+nj3MYdQ/bdlG3LK5jJOh0JkUH/HsvTCOS/cVM
5OFMCFU0ZwiDWZM8lASgDrUPJHPXGlQQ8PqAckmMb1ndG81W2OeJKARDxkEYA8z+
w2QzKRcTZ5Aq/G0/Bi2w9dcMq0M31gjuoSDsSIhCk7F8R5c7EYcl5AZhycgY9Foq
uqCgFaa2brSX8ab35fX3i/Pn6tSRJbYHLbDH5uc6BqBHKQCYFuG+h5305/E4PUa3
wRDUp5nTg2rO8T0aFPMs7mwxYF7H8jmO0aLCKOqDZz9QwsNNQMy2NMQSZyuo++3P
T3S/5X2mVujQ896ykCF0SH6TtXh/AZ6alxgl5zUinyEelmwdc6SLRuhlBqaTiVXA
JIJ97oNXIpw1a2LTvdRx+y2yjaC9FZCZQvpm1+CduQBSMPWvA2xNppjExkaMhtrm
YN5HzjpyIXKXa1DBXt7z/sO45j+FO3S0uipdxTq4P5yE1kkfRftCi6nzvV/Z4899
Oe/FiesGaGf7o2+XSm2WN/xKFMZcD9mG7kYCl0y8bxiCcJBmSjTCSL3+BQnA0F1q
mvNwTVGfztgEHh21Ovv0WIFFzFSEQOwI/3HCssh3uUmYsevul1K5TvInE6pqiHzk
LZKsSL6Ao7sjTjJN8T4H7nv31sE48gxTqFSZg+5Ls2F67tycDUM3UIR4cas6/NjL
KfhstyvYrAeSrI1AdpnBcX9O4EUJp5g27S4OycvTkAxscAlRegfccOOFrIAQ3S8N
hhtCvMq5mLb/SwDt0/sx2iwfEQ8E0FPgKW8yz3jCYQkpjUDe1Z4rwpf0IGPEO2aH
8vPHQxEiUpZ12EkF7hXXVcHGfxMds+z5YTyIyBeuw3ekcvyrZkxGl09sjG+zYs4q
WLLKG9dYJsOf5M61ju4MVxC+8YgNKACjBC+FikS+RwanGdbpsmVCYYFuMziAd8TU
KDPe6g251LY63FBSaDbXWE5saSu1fBwSHUGIK2TaOqEnHGftjhsAbCnoUkiJylcz
rMFlm8EaEhN+ai527NpF8XwhOmh2iWOcACyZTn71dYdJQUUFgCv6bb32C3B5q8tC
4Dl7YeV5NhNNiLJgeVdlVKRz2k7GkJq0hT5NJJZ4U4E1ppoBBSGk9chUrgJd4eP3
krdRc7v019+wAbJReQI3J+9E680h3FufybjFek0gJe0BCSex6W+zMA2rM2xDqznf
Bb0FVlKNGemzfG9BvzyYnAEl115qsLWLxWBrC5FQYMPRJZs3v7kZwJWuCB7ilmgF
JRAOM8Wx/yyjAScU9a5UgXCO9YVjJWc8JI9b0ie5PuwYgrLBiZg3shOSKmILjsmv
z8/zExq26+hhHtJZf8vNp7j6GU6MaWtgrTiSy/zbZ72WkaDmSvtvyuXWD17x2cC6
xumhlXG+nurc/R/OVrE3U6BlYuxcp28ew9+TA8t6qffEfbIetcNPoq/LFCGHGnrT
wl+Mvt3mOU90pRT8adHLAOu62gptNV7H9YgFJMhXBBeiieGOlD9Mp4yRBxATIn//
1Aa333J+bJabazujz2sunHxWt8BBHZQYw1qYOMF3mJN06fvkF/47pG3sZeMXJNtX
JDCZyZwEHkCR2ehANhSkKQFy2gOVvESbDidTlrXYOU/2kqBobJr49vy4jZq2cCOu
vjPsDULM9Kxzjqb14oeBksQ/TXsPnRXzk+48Ns0duXutnxU+nX9tl+kWuCthM9iv
usC/AK8weZRgOllRW/Comg2jWIZnP5mvR4VLS3IolD1gl1dEIZtnkhT8zX8zH61E
G2htMozY/xTZ8v/WIHSkIWXqTUeWLQGMkKYFBD8inBRpkIFLrcJ99cD7PWYaVx8i
QlsbHwKEc7GGKyWUwgqtE0HKz/ayJiCP4t4FP5d/yMqJaL25u8bt5l7QOXTfjSr2
tzdKQ382WgBBKA8wMupxy8RvU2FiCZApguJwPPPgf2/AnQFRiHmOj686T/Bz/iy0
1gPbkXuxsx6puJYvm4OlsCKZTif4rFkthdTacea21ILZyLYEVDFCt0oGYpkodu7l
ECsuvz3v6g0oN2LGoP8wUVBamoFECZsvVS7RD4jqyctE3MZHB1v61pDT0AIYBDGt
UjLJ0rOez3IUiw981nQuYnHcWCU+O7MAxR+ejP8jQjiyoV2S6yZCm2W1HlPoQrAA
Mxwi0M3xSIVk64LWutrqFLbFFoLcoBaUVlFgGQAqU8wahuL7C2y5OfFUeuF4xFUJ
sLCDDR/BqCsX45OeJHjvoTk4qQBYQ1OOhFQNYtJFGVG0cySw3R9eIQYj1f0Q4CMI
0mTMGhWxCMcfiv64vOrsLOHryoJLX0CtHw/xRJeVS78Xfk05vj3YFR8/Eh/f6lgN
4SRl5XR6GJ0/mH5rtd3SAmox44TppztWIb1cBoHKTwrFl0XvcHo9VlDWJBRx0bcv
z0ajteHqoWCwaG1hbD14kTDP/WPBw82tohA1Fj3oaNK1gAFig2LvS2Lcq/aOm7Mu
n3HEMKaN/gpBQSpmEEIq+qpddsXqYdmgc/7zS6ZxNp6vRctDY11HoXc3kWaHFPLy
NwpM4yBRh9426cGrtM4a/reuXLhwDe+A5EvvN1c+7PxAMhX8R9bJ09F4Rjt0I372
j2L1Pweml3z4mIdQy86JAHielBWeKYc4SkrSrXQRGtqET6HSShs9FgAIvtW7CWBr
BLg19TGLQPQNB8hvEa2zgmXi9zBtMfxbcj0EJPoDOXc+IsMTc2/hwimG84Th9fk6
mSKBaTvDC7kqrcgGloiR2Bu7qAtlTWK1fxm6i491HTb1vGJkeckRFymzsQ/sIYZy
KT2sfYJ90cEPyM1GbZ2JPFEXg2aMsI2hOszHYKCX0bXTANVP4Tzt0c5pfIly5Z2I
m4BS/g1KxT8x0wJMt0s5vGsE5HSWHNa81XJpdvG3UhPfvdXJs4UohSEVatv3XiqN
7pK6u/glFqRakMVYPUX4qgvvYeyA300w3YjHd0nU51hdMgTVTKja1aL08/nBn52+
0iD91n9yhb5LTjh9g2HIkDD84tVEXy82oCVEdHyq8DtUCWAubJKTrgHnt9Pc4D2B
6oD8LJxvoshRkVsbg+HcsrxVUCWi6hDDhnLa2jZyDrG/i9XReftW1YSz4aP6KaHK
PycPFJN6dudCGH28THoTCE3bp/eoIW1qL3Tq+OxItYIo4gySUXpFdfwHWzF1ZN/c
RKP6hKqJ2benVTV8KjT/COLUXV29g6o8FBaSIvOV4C1pEUhy7TJnuoP1d0Qk07QQ
i3JHi83Ps6ufd4dv5rV2dw8Riyl1YsZcD4QXPzbUzse2Q98pxJQ8JFfM2fddBLJS
dMcGOhi0gcBr/5u7pg0E+Cb7ta9CmBGe3sZ9FYS/Q59iTbKKd8LZTrhbqeGP9/w7
++qvagjW3GtQuCAR2QM+3VUeGdhNqlbmCMk3QVuBdVMSj8zkOMNJbAD4ADOJHOiA
R3BGPgn1LM05pNL2yS8gLpgLqO+fShgZmoyG5yE2NttQMfuwS1lniYIjCB9MTtRf
BkzcnyW2wtc9GhsQebofT22YN8Zfxve/Jn80Vaset6FpnF039IBe9ZtSKLzG/VE+
p0Is6j75mboRCfPv0qHW3iCQIEVtjBcFsIR9X0pPlTAanIv9CeJ4QSC/3cc06tsf
UU8fDi4/1wQ1+K0mluIgTwEyW6vr+jCr3NXwdib15LjmVRFTCO/HuF7NMi9oNF4w
dYwMxsKR+VbbNN9obSRgsDYt10E4mqzVttY/W7f3jgq1me3hOarH1Ckqsp7dUS0d
ZGfbMYQ1xgbMo+sQsHbIqn72FxUA0zQRBb/dPR+cG04ZI65z84g8VnWe6ENzSQdv
ohh1M5I/s3pXWwTKxwm5fIpaS7RRTVwf7d594vgxNIxJl3Fx+fZdKpNzn3KgUNGO
Rf5J1D227WZhOhsCZ2WK49wMDiL4Wdno4KyIoap4n+wT7AfZM59VXnmtOeSKk3cb
TA/8/rxdHZE4L8pXpYPoj8BBgULeGkBaD0DMj5rLvoOsZXMWJ6KFh7Jh8vNh68A/
6e3tYirAXKULHkdF7DIQ5U57tfEP+61S+jLW9JKITziaUPYGuXKD3o6EUEsslWj9
Pd+V4nD9M2UtR10wIkGGP/rSbOAGWRdm2yuhLLN/24ToeRMPnyp2gDrBBOyn73sv
wUzuCK6AoEx7AdGKxChZOV+PgLkyAj+MT06Kr9nyAHeEfIEIcMFGoT5NoCB0XPUP
R6Y+dCeg/nPSxcjWYL26A8Bl5VWAPbbTedGPAnuIm0g70hSpWtwEa8es36xEnubQ
RTUfPuRKhtM58XKKTp1qGKl1wdcfSXx4dIP2L7k1FOTk1bLMQGvmiA3DwBkkCKpH
J3SqTAe0M4JMiGIls4NhTaEd/O8OduG2Bl3FLc4gGqVZKLA6/8PDt3SJgcRshJA+
P1QBYwCaOP+mSsSC2EZhx0KLJZRBI/0SzgwwR5Q78aORQJL70tzhILTmkT3TFUfW
U/ZQ9+L99SdeIfPqdJ4S95v2Zaq7ejhC7ln5hxpBkZk2qwsfM8n6DHX4spux4oT3
kunt1/cu++RgqomeURXw0X81znhcmnKyOIom6QvgoIoOLuPACAOf53HjAMIaFQqi
WbUVr3NgYqnGYjSQFFEmS3hXO0f3qdd4wHQ0bjkL835iCW+WdPHQJ72npK/mpso0
/0dTvA+dQHj7NAN13CJsPB4/MbjAKlQWpohOLZO8YDDJijjtuoRx8U60tQCDABA9
Ws4vxPDQODY/N5riEXXD3SsjlajuXrmcIkRkyjWU/omAk1gXE21wXaAtiQjvBKYg
/chXa8vqHcXcasDFHdjjdtXUWAlDs1vKHYkeToMt0jgsoQ0eVT/XUAzQUCNxzdMN
MbUF+sa6yD+whzZdLsSVz2yFBsFAtlkb+UJnnWIvOz5ioIk6yl8KOxKx0LkzzKzJ
UBTzbPaelb+J2KfPbmbinHDx4pqEdPdtXNHqaD03VCpMFONxWD94aso5Zotb3yg0
xfrS9xTFTTWbr+uCepEGt91h0uslfkVTP5v60XzRkb7ALNUyFgdkR4OJdWBo3Tj1
RnB+xQqNOoeWIpui5Gm38FGD+j/gEpMGfDs3tuCNd1lW+AtJWi7al/t6PZ54gIi9
Gj/cKaVBN0rtJutP6WJrOMCEsbP1z9+ARWrdIchv7WFVWaCZ18ejJNJiR1Xm8aGq
Ri/MSlzQNmmhS+3tH3ON74qrt4klD6rRcgiIjl97nX6zbLG0dWW6VUQIxcFhzmqh
rPKhafLHJGOc/y9xUyqxKy8/nfZQdwtF8B/BW/31MHoiPVNHbSYtoNJUET5A0/u5
8yaXjmNeq8SGawbJ1bk5vd2psfgBCIf64YwAhPgfRACFdc/RQbs9OgwRcNTgXsQQ
rEoM9SKrl0z4x0FT1+GeUAWRDQIqo5HdH+XR8MDoUnyRE4ElpiB1D+rGrF8diHzg
YwMsAHJ1mmThn6wXEiLXyRBcyzqQQDlkIf1UKyGaStOl3ske6lf4hXQ4vZd6BYd2
PYu+QCOqHkbYzq5HGJhXvkEyuH8JvHBxzYbaagZlhlxkwfI8OZxkGFtfdGfg+fX/
F9KUrczMRbEOcP5pRccbrdgpmiGtri9fOScLHvZpwren60OpmZH2ZshKIsGv/3nC
YIHBrxD14AzHkUSM0KmQpVwuxHepcgrF580Ib4skAhaTlQkdgIlxg3lscOaOAKK2
JZON8WVXgS1IphwxCv8B/91TZfqx8POlYl5VqY4TSuH9f4/R395lL7viw2mAPLjF
G6ZpewN5251TO4gT279qun3dqsj2n0+hILA4lzenJO3ff07XmrsPKUVSGknIWFRF
3AaqHoPWP8vqcTr1z/hsfYLdsIJl4x1DOXMt8Qb4Gh8GqgvGMTIo+j8MewIjceA3
VkGenLeg2YV03fOxHOsEk1W2wVF2Dq4pi/1STw4daw0Fqg9JURLyREwQrbmwugQu
Z2hyjiPIcHM2KxoN2X5NzZpN7zMmas8NB0b0fOA5HebPYRJ/eHgyui1BvcrepdQ3
+e9W+oJw34nsVdvclREvj3DstGgB9KmsjaDNiSiNrBsb/RXuzEsoo0urqqlToJvp
Xf9kKhS45dcf3uxv4k0kAk0f/5i4CBgtHXkdUjz8zqxJnkUA+ctaEfm4z5xigEjW
x3GBP/wkOUjJA2EIx4ichb7wlklP1k6LsJM+q25HoJjgIIN78zSxUFTNtwCTmDzA
dcxhPa+ioWVyUqe+yVqoeDGq/Z3LKsOMwfBSqWGB2BlZOsaeLRQFcGaUL0d8FqEs
Ty7qE+JG6b+rJrr879R0B+9ufc3ukXeLzciIQK9sm0zQQGIGGM8x0G441TFw/ywA
qa1xGR2lycSdW0cxWQbZYGzXYUHSUrCNhOunW+0N4rdMMAfrbR7oJF3XDwBny6yC
Q/LhGvsoTzTqxpCwYoqhRqunl8Fotm5IzoBQHTYPp1VQaJbPIJ/DrNZp0ds1Pdld
DtP8Hx7Chc66m43h/4G+gn2XuRQ6MVfYgzwdOyQgppOwGv+DJNs80aTzNnsdzPaK
xoIS4uAH5Z2r7wXw+ZugrNvGPgB8L5AgWNPeHNg1GCq6c8vboMdMS70qo7u5QNqu
io7qiW6RZxzMrNDHP4W2MtD4dFIIsUjjev7iASmh7uytgcB56Z2dSC1evZb3G9Wl
62uWpshV57K4F240vnCH0CKnObQavJuNIqX/v56eYzRoFblPqUwhIxBJuN/zfyCc
B5jeFZjG5Yu37zIySzLh7xSX+D71T1lUTwHGTgR2TIvpfUqNbV6FPwUiXJDvNiZp
lHx7ImDAjMTRyocIfuEri95szgu3MAxWeDoZe2pcVg3XbHgB/Z6PmQr2FtsEQfpM
y18grSs2EGBB8QCtYA9sk3ZeEZZD/lil/D4mkOAS6+14TTl5zlDbdAG61Krthf3f
8J7pG/HqOz4fUjevmip1xhQ7KMosgUKUHLuyz7lFA0rTgw4wZ3ZqfRACxZ2iZ0kQ
8GcyDJoJIRmCbX+khGLoWVaOvkCiW76z0az+MP9e6uANcIwaDqKLU9IZKHaNzBbt
PvH12JI8m4awSAc+T3MBguHw4J7BcePUc8ec22/3C6Vo+8oN01D3e6ccPUZDBHfo
P9DKlOM6y2nNr4OMKArY0yGEz+KgdrznIj8573rowQu3XiKVkrbhF8xPqkbsG2kk
UEFzUTKampNbrY8p5d+wCKx2wF0WrvjYbF0RROxwg1dnvNEjNKRSX+tk8xEOLA1G
3oZDdtPYfAuZLHdmQu3PNvdPHh8f4U1gATH9Vmt3gFrFp0Yp+N0Y8ssPM9uDcMeG
PwaoJPZZciS4y1yoehTWDQChYw1gzINhL0Uv0zKgXaZ3AnuYeH4ORunUELq0MfEh
lpMVXn7TkpopygB0XtO3Yzh0fIYSK1h9KpbdnnBQXJV0Ap5RyQQB8XIwOHRm1Via
dnzPaj/9R2EbeyRKZgCTCGJIdUFmMtitArp90lynedAH00kSQONJ49TkVzAc0W2g
PRPTFgYJhAhyr6tNfUvTiwokIDIyorNZPoP0z2vlZrwXMTxPjmby76Mh8iKj+grF
JhmONBJ26VvglL4E332nZ2EPgrGkJnFAtG3W/ri0DsMKE/76qmQ5A+j+ssZ+jv8t
tjBx93jT66Avi+zmxfQqAgTILSq5xfY/DndNkYejifX5LSkhOlxkS62PO9Gi9133
G7heggbUDEZ66i2kHn/4CmZ4QLvh6cevIFB8ITuoRV9OWWynVzeIPZwMN6WFPsgx
z5DFOpt8DfcSNI7bNHgn3F7B07Bob5t7EQUvqrCkz7N5sPtjgxYr8MpQTNpy18VJ
6V4reaQdTVcNAVbrT0Z79OYtsXmWqnUzkZgZEK5UIlMkyL53sYKN6TtzJPxduXsI
gUo4MkmHesyyQKp/4rnUMOzWdOpMkEOiAkMOZOG9X2fgPgufVx/jP/xCcj5wOA/f
W6YdHXSz5CoQP6ODUEaNtxZAIQq+FPuBEEatHNZsyUbufNAaxRuMa3H06qQVb2Xh
NPN2wA3ZyEPPorDFd1jf/sgk+D2USgiE7ZktDl8tCXRjNsQORrlSGYERYemSSRdE
NopmLeCJgXp61RWWTjepCogvusCnc8H3iN9IDKz5PKVdLb8etd6X3j3ZQWCXgBB6
JJtYNHblCnrKfqz0vL74q7l61u7scvh2ZLSOw1929YiWkDkd/H5VgjDd+qz9oqoY
RtLUhMzt+PfCkxI+/5hU7eoycu5JHyw03rTxNNJQU47yLT8Co1yJ3xoMOMIpSOyE
Hioooy04vl+H322uVBV8A7dxZ38cQ4kCT77EWvXBobBzLFnMD1dwkuC+fdrG7euM
nkgRa7WK3vv0DGuS7ms4D23iKRh+sdix1qRrfJEYGYimiN85tdR01h50qInHe5J8
y3y3YY7lM/G1fp8/Vfjt5BpRA2I1ylJ3UrQ77D8oXIqboYJrioht1c2i/ELGFvOi
Au148wCcLNhJqlHNojg2essIcXnW0vvgLONGDhqWI8xP2inU56L3tHgU5ucrS2FF
XIpMFz4SiWgmzJkunBGhUevQx5JACuMKrJDd3H7J3MROgM+r/H4YgTYB9ZWGtAZN
480SNM266XB9Up4mTN7NTXtmChURymShOReVSRp1YXafq/ynYObabb62Z2aRvm9g
X9qUcVEPOFIsGMAiXh+PbvtCGikhlqTGVONgWxku/9SjTM4Pvdv3oZsnv21LmH8W
toJosVaW0StiguvFRsKtiQtwaGiMbkhjgPcVEPvcLulW6/Dbz2SoKpw2L3Plof86
By7k7w+FN3VoP6d/GraOcZiLv5aTzKmBl2ZH76q9gPd2v16aELwMhMvvXhNsrSFO
aO9GTcqLvTE1wv/Q6wn1VtdiHbNgGc3D2DQW2J60HUINLR6pUmqZs8EFipdZuow5
wEzxz5PNelxlPIw+z15wVT68bano6Abqx/AJYOP2afIZKXUk2vRyp6IYJr3TLNma
ieVJTXjy/IzoMuk1L7yuQow+3j4vct2FiqzcOZDAEZA3PuNloWitixnqxuCcQmZJ
O3YN0pUYwIMeoWSRd0mq5xiyHXldWG+MsqEaigi0Rqr+DZvLyvbcHxgMVhRHQ1Cl
73Cad91xxF7nMuduUvTtFhYSGBTz3ZxuQgyf8324WRKcrGoMJOy/AWat7iWo+Jru
Tue8Pez5ru7+m28GBrlrdSEkzqbBe0eKSIXJFbJf973HgdX8yM2D2/TNJI3QukX9
U9jt/CIsDEfwixt9xKKXiakxrJOvr3LEVdvZ4kEpvQDyXOTCwzVfnpQ2lUsv2AHJ
b1Egbnn7cLcJF4EMn9qT3u4vY9dWoAZck+vbIRD76hm4kNTagGatt3m6qraUnP/a
eFwwTc6dm3JxQP6lKH4Y9slBT5vZv0bVxIp3gRLFxRc32iq81imjcvVXkMJQ1fPr
shapgn19Lkclap7zbjGlrRTk3tzmYEXleFeDNCD0Yqk00/oKoBrvsw+aXwt+6G4Y
dp0M8OWaJb6AeGfDXzavBpJnsOHNFxsNTMp7Svi7FoNXkZhYgQ3vKXj5apx4KutF
8a3GJvUIRRpaCyfSB2/FZEo7/8lzzw6tJp8sRYWl4LdZlCWLJAVFoKVIlxLlwixk
oHl+rF806jQ4mRXeCWQlmFqZ/A0+F2A8Lj20XF695LmYqa0krth+qLVwDzIG0MnE
q9kFC2KXVu6uLDedBtKeLHiAZ2UUlkKFWdBFC7UFMm90WHexp6lujJLZetgDM4aB
kqoof/tuaF7ns3gr3WBgJHADSTupb5/1X3zHK+7k2tYnQIJ221Tt/yR36+2xocRL
OTLZbMUwhomhIyW1lnLvK61+yNQqF+R8L1Ali9lShUeexyT/rKZUQwKzyUNsrpDG
Sv1N7PCgyQBbz1qyQNd5iaS59kQ/6hS94475EDOOgeNf2TIusEOmWOoqI248k4nh
jQeyXRArLs00c265kfsIVjCSYi09HIzIuT/OVlA4DrCzIGTuMdA8e6qAo9Zg7jBZ
N/3+8rMAEY2Js5srLRUFZvnrAcOwo0e/QxF9btW/nkHtFkHRUji9NssPusycak2G
1VNk207syjqm9KzeWiLQ4r2ykPPvJQg/k4/kA7kvYfWPLgcV4ywxlLU8sLp73Ltu
tauPv6auLZlGD9Knhes9IPolc1YUwgBjhhv9AdVMm0brJ710bHKmIssU6uj7uM2x
KBgwGjnOM1xko+vXObBvGitOqz+EiPniIS+LYY5TQzIlTxEPjAYrb/A2w1Ej8iPa
5B/8IJOHrDs5R+Z86NlAHO9HQspiEcCrk+pKbp8KMvhXvHDHD2hJFb7VVXs74jao
P7u3mllBMDlyayuDgq/Sa4FdyGdiZ1cOfC8VvpFdhaEia7G90MnAwAMZOUMjvtrb
rscRgvhYDvVO+ab13LNiE/cgmoZgbaXrhTYQReZwCNmFXuhMb6MbPvz/0Ifmwjcl
zdd+BJ83M04srWuPLjt5T68Q5He3C9zsTH/w1IHJOtQjAnKbeAKuYKAhw0YTj76m
emuTmqH3bnjkb2XbeI0ucuBmGX1Nv8mHSPvCkappYNcw87DKOvViARcwzxBM+GQY
NcO8WIpUJ/oNaBizo+4c3VCMPyilA662Ljpafy7CSpWrvYqkYRyQ6moGyqiMje1m
U4jKwICIGqwbn6AN7WvcVHr+n9w8hYdC6lbNv6X5LKneC05po6Ff5pJnADrQEQGg
zYNGFA5sVAT20AoccUZaAVKzJzr4aWr8jON+vAE7IPU7mc0DQgT74kK1RWgGR5Q6
8q5Hbr6wqiM3hnNd7Ux7xg+nGNqJQp+yswz+NsWg+9SUQ5T8FzjokKA8ROmb1PYK
PX5J5enx7o6Fz5ptYu/FVwzEoK5IzRkCqR0EC75WIWXbsTKLM8B9zaQ1OPVhujr2
7bZupPLZn9KMl4MdYC/zlVI770gppTSQj/taIFonU0Ficn3c/A+cKZgu1iWNP28r
8ytz2TQg4M7vMd5mGEp+p1tebp7Z5etVMW0uO6lOPuflRqhrQM4y0ZolqlONxTz7
mO+I89s22TlxM/sljLdm4b7mrLguWDM2NnI+8aCji8lBZovszNu46ZD9R8HiuWCv
AFxdHmzrTYL6WNbFIY5Kfo5mox/f1XndN9Nn8p5FqHqBD9v7NXivo1ZbrZIZucNd
/TYBRSI93bhdEYljT/TATJdkd7KjjFnRE1qlLzaYgrbwwk33yjJbapBLB5mqIoMO
Rcidm0uCP/0G0ZVslcLBYVk1IJrLOdMWYpO/hVUG1xfF9uv3y4dgnCtbdCHUWd9Q
3KCFLQAtV0LRWAUreaQDaOG59XB1w8dqSM5HSP5zcwjUyf4y05dFTWsknIG+LDtw
THSkGs2je+rwb/70glW1hWTHrgm97rHKeYLkCpHaczLLVGDo6+vFdLgHBuvBzMpI
/uLnNomRegD1s3mv2yLhqymBD5YMoLLdXo7/Ja2whwF9KCf26fk0pK+1lNrkKsEz
WihJRMJNrB7iQBzrSpSlPoZdy69KLWylwn93SM2JXXPAJTvHej0W02clkqE2uESR
D1XKR8gZx4JQB50t7XKoB/vJTn20xJ/+z1wCoxLLFunF6gcZ/LTGvA6owZDD7Auj
Qm6gYkWwZRdE6E1D1jwE1mLYkC2iX9XHRG8L3GWdlyh/JGPt6Kmm/vCVYkOrycx9
lbIGHssjVIOkZkzs70Vt7n8NmW7llbDKKAdoMDAgoitgnGh0eKW15dOS0FBKDM3B
RNi32uKyT0cIrip2kA0Ijbk0XE/Em8Q/L+H+CwP1YpNufp7kf3vBpDUTeHJ30WJ+
cyBriw4PBpN9NRbGxztEdoAZcjYf33pwGPgNNqrhW96O1uMzpziVIXu44UG/lP4B
`pragma protect end_protected
