// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
m9X4o+aufZcFgU0ZlqhIOeQBhS5fabSxhIKviA8+QwTKbDL5g32zkuPC3X88SlVWAVW+oldAvm9K
mS6TpgRWbkLj/VEka6UH255wJazn7BbRhZU5PXOGdIHVuSDvGiFiLNJt31pBvOykO0/9/bxdHIwF
jr9oKyTSmsZ1UmWd8YC+KHOiz3M49r6krQ0l5vCYnIzYC0tBjYkYX3iewc3f8vvvHYawZvLE4VoA
2SLHF0A1IkfOjScT9dqMeNnpLSl+CF9pOaxo+57ppliuImxzmxcKl7mIbDlx0OxMLaPZncwHhc67
Bx/tRzt39ZKr+M/6G55mm/RTZuNuoFKtLLViNw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 43984)
rk6HI8PhBfrbGJoqK9jFhP7528n+ZY3tm5WM3XaWLTP2nPRCVYrH/ylAbUM/ETnz+7M97DIUw+Te
06w2xHOs1JrVVFXUVYeEibmsisFr8iuHERoYm03pDKLJ7Fkxv80v2fqHTg9pl5D0tytVaNuiHvBg
+4jXXubTHssHjPZ3SlZ/YuWrAGlP99+S1q1/dwUXJB8WbyeYAUz/H6VGkeMRcoyAGcclg/leXc48
GnFrMT6H0wUgIcDdoJInmEwSZbME1IToBEZ0O1sXFAl36bB97ZDJOrFaq78MB85JprO3/Fp1hypa
zA13Ar5o8ANsviEOejy3umSJU27cf7FWmA3LeEAhCh52C5Wco2WhmrTQKH6NmwIreRJpgloWO714
T3y+Ght/FMSlpVRyj1SEJo7WRvTIR+687hLyLhrFwp4smLcTVa1UOsi6/ZhRAjVUUcymxRt2Npvc
cifb/lLq8cWcJ8wHfRr+LWldzQZsGj1j3tTQHiRJg9whSQ1F4X6mx4P98j/BzbZwC+GbMczcAfBC
l1E5YmjuPEox634nGyR0Le5ICFissaVxvcXxVz6BcF4coXtyc4OgsAeOMmyQ8fIPTNHrlm5FJxj3
fSBz3Ntd7M0ISWROv9Z68D537ePhphyJ9MPsvyQET//fcQo1tj+vISW2GpHFwDVKDY4dZa3nTSWe
C2uOJ0Ng/NVEMvnGlpWm9AM9BpvrSn8Lt9sarCBKUZRLDkv1Q68fhgtm4p/G69ikWBDYRUc5Ufr3
Yzy3hPaIHTrlE8Ur0govf2WZDyZ2P9kOlOQQauDM2jt+IjU5lXRilY0EntqdHE56ye6JuUW2wFUL
XdD6NOxBjnnZyVpEP8pSSdWbtk9E8GKbf1n67M7Chta0o6vBTqbSXoorz1HuHCjhiSpKVdQ7qOV5
ZCNEHk8lkrQdiDRShiCIbaFBeOWrbNoOVVdi7uOQ8ABwV/81LeeRltZ6VmPGSqIKaIlgCGDU29uY
i1Om7UmbOU63df3n9FTbdhj2ZRoC//98jjbJddQM58va8br0C+DIKVwZv01xMjnhMs0cbS+7RJep
BdZTJ5blaazU9i/VRWEBWSZAtLUX7eCGE3B+/0J3PLmQJQ4t6I4fA+UYT7BqRwKbaUhTY7+jR3Rb
DJHaKgjdwJHrFA3Ayoq0dPZY5vUQKmGbBrXOs0TxgWjrBAjeMMOk8jTdMCXCaMCDLmgTVbDMF3z2
eQWq5h1yZA1AGoq0OSc8WuINqminvs5qpzDjyb7j3qhQaM4C8FVgJRI47EmYgiTLZ4z2RK0CZLLT
rTkXkP4blMAloBQ/NnuWuBkduxUhy7FCA/8V3sOMpB2vQa0r8ip/uqFEmBA+r6jRfnGe5RRdVROt
dGO/bPHevu19LWCLLq+E6dvkuQ/e9PqOQ8a94upR8dbwNSeZTQYi3f3/YVBrlBouWL95JZXXKgI2
WG1IIjiHkOpvYs/YPpNRRuABk6uh4ze5+6tmD3IyYs6MyJ6q/CS9/G70xBMJPJpYX2jShGtsSt4l
9mAqPJIWLTDFuJU1L/Uht18e2SBY+nlkcQASMGpheHn6GFIcR/gdnHShoTYp4C/IGJwVQzaGJQnT
WoBM4vikYgneBBs5l4ox0ezAydct+MfGQLDxxmyD12S1EtpRwhxrrIs/v/cRUrTLd+tplKuAkW5Z
hB5PYhssFRr/l+gRwDYr6S7r6pWpY/nUMhSblspA09DH0if/n7kOkeYY2yRIsJXLruUSih2tsvia
whjdpjfVUgh0ERzymSbZs34LtnW8ZSSmXKn7xGpyYuIN0o6+3xPQ8FLjsZMZgFWQ6NTZcn0uqMgt
GC3yklKYy9N6i0GCeyjmrxWNcWcykgID1QTYLM48RQJ1ze2+UGp9fDPQsUM2qQxnjLguAkzDh4fj
c1EQtD/DZu30HVO6g5+3VwSMeldRv6USEUqfKAu2Ohrpd7g9SWBH4VbUdMUOGeLf9b+WVBmroxJf
7k3at6LyAyghZ8oi5aUIWgBS01475yhV6VIrpv9vkoA8Q9JyFzO/LNDMBfDZRckc0sP3IEww8ckD
WbtGu4L5aBP5MYgs2Sx4t659TiO/DPFa+AZOAb8Hz8mW6V9NqmBtf776IJk82+Ibu8XkqvSZ5nr1
WhaW9rJwp2u/xy9m+Pe7H0cjWnBXVJWPHKJR0lBqvqPYjHxK2M9S7xdwVRKm0gJ0JP6BKLxb/FK6
ofZBFZQTyxTK+TwDih9HCQq/FXSlIX3TU5eawjvs2vJm7x37ePU0RdeKMB1bh9024vkHoZpQS49h
VPLMmSP3jraQprmrxGcgZSQt7/fY77Dm6BCjsMGhWz+K+vht2mU0UiLFfdhoyoD+dfPGp2raz0Wa
ywto7V1ABNTKf2XD6jR/KlVtUJnLqpCVFZd/s3ao7+DdIC8d9YjRrpGavBzYF/Ad1qZW7oZrnWp2
g8k2ZKMMsd62SpVOGwwqxRwxkbPsHsVdz1O16SoOYjZG5Ur0c/SHT9gJgV3bnXKvCEkVEC3ngUUi
I9w0tElK0A1Bpr57CBU+snos8jd6Iphwb1fnTZoZTykBu/TVZkiIQYDxFsMONAvHfRALUYhTXo3o
dvQHXwCB5gLEc/8IG7kFiZQAd2lFXzb4+kiKiwTDS/oD/hxHXOdoJ2+pFo6ZMpTzPZj8Rb0QEfZ5
OvGd9rC8XOm8ZBt9I71aGrzYh0KcIf0ONzRmtk0m0MDcNz7DQ/i0q6CMCaZJyGbqsSCZHvDMRjTx
qaPaermxYqc2SfT2csJkJh1ft7kxeqNQTlABBmuXa+gU9LHJcVOEMB3OfYh/bgYxLKtBkFfY8Ri3
RRW7UmbkXzy6Qiv/w/GrqcS+8M6+XmLF+8GgnQB1LVVWmPdIfLG6t3lLMUAI73XeaRWLaaJ9y2Aw
NL2TKBbX8uzRtmRr8N9GwOEwqY44VgG1Tn/PsDrIY2Nwo6tVkl/E1yRwTSzpnZ4YhCcBF+lyoneV
TE27RJx74K9LIc86jEDVaGKyoSeU4qjVhKHIhcZV08DdBPzfrMUkdFKYAqZ3zCgIFVjZOKdUigLR
FzGNcKiBGCXDA2noLEfsMt0HE1LCi0HrQYKlZm1NTVw2rzKQohxXyK4NZGb8x/fEgUKECmSq0zwC
dQgRLVtp7S+mt2D5nrJlnLXDUKeU025WssR2tP0fiakZaDm+XKF51qZZZCkj7a4MvZV5LM/afsC8
O7UDClh8JuUUfPFFB+B75mJvQfbypXliDL1HbsbMxiAr2fVcf69WzLo3LJ6LWmZWiqD9uBMVMwpa
AI9kMrFI55jOosY72mOW6uXD+/CfSNns02+0QRuYbcnX7wnF/mQO8tJ2s6kscInHPmNZH+OZH9qj
J+lGD7DuoSLwp+bJpmu24LyzCvuAQ4oZyt3eD13f29G7ldIs7mcl82UBVDuQXqnQoJipXfhLxQGV
Wp9TP64OPrP2LXpkzKR+XrPbpXM+18eB34PHqWV4bQWYlDSDPduPcuNRF8QLEHuWveK3k3PzTAhs
bKiEAlNxeYGXUFJ+wf1Hi2T2fYbJhy6f6WlI8cf4V1KMTnpaao4sgPLvJF828gDAAyYWXuyd+Ltr
QuEBOxPlMQkHo4CV36xhRE7tsPLrVUfi54Jho3LDo3N2I3f3TSUhc4D9ufXASU1ycdrxC3huD39J
luxS2LarQqXSk+hW+yjgHjPliTrMhDCx7lUh7fa2qiU/q0suPu6t+FryIFo1vJ1HK1+NiVEIW+pN
3esFpxPKz9eU6s8I9K2TyO+aDHGvZGmx+JElOvNaOPT8aoKkYDpfl4zRNWE1U7EcxOktMNOwW1TV
5tOUCTjoyr+xaVp3C8O7U7nmRgCXi8kbTPConKQivx4TJ63AXozQmCfqoorG0m+swGqL2rejAtgM
COpRM9vBln1ljaL3H41CcLVACBMl67dRwMn3zupxaClC51YjrbY9a0zFVZKdLNLrQHEuaUCZHZAv
/TH9nAIf2pQ8eLcs41s/lMIk8NXuVApXwf+GVv/mY+5kgSxqtkhnRrgrPKUZm7nxP7QICbtPdg/a
Dy1YsJycfzUYKYyttIYERF8YLYnmieFYwDzyX6keDdY2LlfsFWF+Z2aYGh5vHGehr9qS9Ol9PluN
lxTDQlaVipIQD3RmwBcMwaepz2+VcE/fNvcbSLjRCwZazKX67+5011bE2nBXhRFvKNVGmZtqbSNf
B6AvQ3EnXvvM5APB8bdqaql32X9J4WsZxvGXOZ0/HJ0zgqJkfQzznTm6kuML/mR0hYuh28alHE/e
kypgPyHqIzfP8QtMsNGDUAlhs7FCfmDZbU97W1GNIYI2ggO3sMsGWeVVEkLWVVRGzWCftXLibAeB
/J7vjZXNuZ79i7JXfBSANNsL78cp8pX7j7F4+eJxc9PwapNkHo/VUITgj+nMx07DrajO5udPJt16
/QE0AoH6Fo3cHZwj+gi4gEkmNLZJJ8NP//o6hl6BdX5ImQdlIpKsW8p8TWrbA74kqoIVlyCou9u9
BbxrgWzgXvr/u1r/xxjHX0bvEZ6B7p/TBsk0HrVE2WmvBadJCjGMmOSn++i+E6kDMNV4x81MutaA
XYrrCDeOY2MNrrzmY6pJPm/kTz+vyrNSdaY+jBzmGvm5JNBWBWCOxF64dJcSh9AQ6BUwPcQcAS6i
fF3pSMhGs7IhQegfQvr679qFZavO2TTa9fo7PQ+b/GZDRnIA9ECMdpdFt4JbXOhNRnrqyRA++OMH
+4iVM0sqY1lPprHzJSwRWp1e6O5BDgNy51qZZdCIDeE6J79qxzv+Hw2KCA21zDOs/rc7L2jYaAqq
4eYUGi4eJlDpS+TVVKfcZytQ+DpckdUd2J4YE2VGaR4lRbgrKYKmU0UdaCbRzTfQYFMp0v7krzs2
7Z0Y7fGKw8J+vNO4FZPKQSSQXrAMLBJb4v1H6hWPl6M9E3wwDH1bnyayPsIlJf8hLTmq/+pNIiA4
l97G4SUtzUbkxph8eDi0/xqYkOUdbkg0UoteH2tT3k4dKD4ESfuXGimyGqb9Xp72hkbYY/3FwcTY
8wnZbGPPU5mY74sl1BTBlHCauy7dqNWFtMQf7a050PKU3AK2uwUfjCn6+fvhk/QPGAWSpn0LZrFE
ENh4RRVfeVD21wRAEdysVZZvdnabzXfEjyZenSHsZvNLbQVnUatU1EMv+HEAXstexi+XfFMBPERr
dTtRCg7HnJYJFTzgsgSYlvnWwj/PQ8mAVndrxIXUkMdk2cZYZA+RhQW7pWouyUSAkAO9KPFI3O0O
0W3fFOdQFtmQYy5af/FTilQqwyj0j8iZ+AEz3D347Ckw8kD04LsSkxq9zLBEbfOnyQeYjtyHrllg
DLisfltMQvDD5TC48ufy5/nyFw2vK2OWzikrxih8ZxGeZj0Njrg0axxSz3HXyacihd0KLxfxepcH
b8j2VHpYB6T1Sl/gbRtSEmdVZmI+AKefOqGBEyqxsphbzg5514oh7sqW2hm4Uect9r4uKjhEWREh
js9PBq9skFZwLdcimxuRATjP5aaroEnEwaPny585+3VMdX9pEypcifzdtun43u5HmXNlSl0+8KKT
Y5FlR2EbnmuPaf1li3by08smNh0a2OgAL/fKbR7AgFtKDX1/VEsPNtcB7tKXSl56pMxuLaZDldnk
UTy68qGfW8ezMH9SgqR3izg5dA6jzl5cUj+fzMn7oDs5F09mY9ptWJvxXWCBn48twYi0Aw48rB3v
dKGSQrnUUqMrUT7leYZa88XovZubmtQ22mP3i/COGS61GI1yIBQgaWmqoTHFHUYz7JcJa7xeJk/u
KKo7Fiyiwr2hoaDwek+ISbK2WpwV3gmO2K3b1crmPa47cMVVMbRZkTJu0H3ItzQauRgiJM21SYU5
LOoCPNOEXmgJRGO/tWLL9af2J4C8ZQlQB8HcYM9PPkPpMxafA1Eu4VACKGuK+IJv51WnoX7JkrGc
u/SUvCyyyCfkS5V4AhZvVcAUQkBdQx5Udwi4SZkD+ZtGOOlh9wjEDYyKLyp5y3BadL4WlE/1/SIY
w88jqYE8IXLFJQl5Td4O2pcA+dqvVyp5o7eciiLznZPltllQOSyfA6DXkMSjYpTnVmSqLorkGSBP
fQHh8rhr53qHG3k+vm1ZDQzCkx7ZfiUxGfEgMFf3PIVv4DUaLNEbz08S+b/ixvW8oQuAVFvPK30k
SDv1V+8LIonDCxfiMjBrwKUE+7UWsuagensMubKKiyJyp6UZSATf+hIfLr2IlAqx9radOyuqa9i0
MLGANe/a60/H09cgbecRU+tb/1vMNxLvNPbjel+Abp6lBK6/vKdKtUPtEqniy/I/+q448tLBRCdl
gLG5Q+3Nz34zLDsgMZUjt0wOZIPDTy47CCGx/ht1vWmp/IaBYiKqgDoyMX64QwvovaFxaA4yZ/Va
uy63Swt/ls0KEORC6ODzKKiTx+L02A6v12R3Ong3EWOZrAPHbL+QBZWCQVklG2PFxEDOr0RveyIR
lUXGogElEkGfWJW5NhHujCDqXuyaB9RHLKWUEwmWiTtWVhf0OlOW1D/geOhXP0Kmbo8mZiOg+HHg
JQco6SDVDLL+iYuPQbjbHbVHejMadCo5+694wW8oZmoVWZbmYToD6ZYBHLwH2txnNGRWBF5g+kKx
pk5fJoOmLD3JPgRqjunnDYhQwwAGavaFinB8BzkkocyjBg//WKvydtDpgXa/kikv5xi66dRFDwVY
O859t0BMpV7K2X8hv1e9RYscMMriXBRQ01N3lLb3PIS05HjIAbXkz/yMP4vZGPjTm1hP5sulRlWt
H4yhvpaHxIrNnM26DdKQIteQ1dyoMN+3i1s4CP8gFh3yj6sOE4dhEaQHNjzQWIDWo10xX6E/dLjs
O4py+zOUKpg618Rqk6jXY1kNDzh4JEff1ovsSKYs4K8DL1Hl2jnU8QpWyRQ6cBPMmil9O7pDvAiG
7849pGASzGhaAMhXROfnjxfEHArnNIP4xMdq5Sdc/JeZcvuUyDSVHoIAR/A1wUtXxJGAavB/po6D
MAWcz9ZplPoRFFX8DhdLI2jywr8FjERUKQPP/DRQD0WX6IXCpHeL1Hbiwg5EXP15EuyizNl99bPX
THUKJ4b0hRhOMgwYPXKoJbc2BdIrwVlpF5nMS97UepsS4RMz83y1C/kJCGNGz0GFxd4xPZ6GO7mY
D4BGT90ljEYPPBNbj3NcdJj5J9Za8eNcKhfdVWC923MjfG0yul3DU0ayFudOcBRuLcInY6yj29rq
bGTQ93MV8oofnzd18liDDUg+OQInl8O9VQ9rUGmhDsNceZsUxql7tteHbJPslUNdf0Z8IlO+xCn7
0Cw/1Y/eNYFK0HZAlilXfFaT+F/tALcq2p1L0BExF7DU/RvMMDwKLms5DPuoBN+/dADHho1RIsSx
KCzbLREtFfDISrqpZrMpMpDeGg4DfgNjdXHtIrR6OTj9XH9IElUUSS0RsAlaed6IoFij1dKTG53t
c/DgZ6SGClIHYvvUT18u9xGCH6cFPGoLUQdZ0ZoSLPLiAR+lN14EM8DsG8AoFP+lUhA/QHBuSB3+
mgEnrzA6+AFBl25nvEIHmK2HIQw7dbaMcVbqxk8p6FTz/lP7Xa8gQym+7dc0P4DoAhytQ3iDPAXb
/6fFVzI0XWAgsTdM+NwHhLfZOpy2bBn3GrypLkQb2egqi5LuZp5atpDFj/fvgdfZrDr88eYNTdOc
8ZsvlStSplqrEPISD4j8XiQfButCqizDI7pYYkevuUxEyyMbgBwh7WCuZlE4hHLN/OxG9eveJ157
m6mV4kCrD9V2NUpFDqtI1F+XFWBJbc+ZA2BpxEzW0WJROyD3MJc4BDiNfQ0pqsCq+HJKMi+lBrtN
vLq5+e7uUJrmScKZfoqiYJegNgorcFTvYly0MwOrOtAASLL60j7NEj+8Ccez4HKu2MSzZt01ooDW
otmmjU8RGgces2aVNfvXGlKVQvG8AhjJYcMH4fadLrmgTfcOrzsO/zyG6JRMFRVRY8s/+tDnwia5
quQT/cvu1PEOYLtfegclyF1tH8YpGJJRxarfdY3plUMbFWaOuXhkyu9hX8GjSpuEhAj7d23DSFcH
fnBY8B3MEezv9HO2c7uvJC6dMLPuBpU4DYaL7U3vqSVNqENde+Ka0+nt7mhV+eq9Ko4OEV/V9p8i
Axkh7V57qwxq9i2g2fCRiRpgBOHGxURNL1/kABpYOuZpRVN+kmNH0/TN+xzjjonYeyoflt4BkhEr
pBpd2pgJR4nES33vyKR+amkpSd5d2ygCD6SpE8PnWKk9OnTuo7fd2dW2oy78VYMMCb4bqQc74w7c
Yz/n6Xe4q8YYT5oYjMe9fx5eiW5S6oHn34jZBe2jEzQgx4HBaRIAhfnIM4ELuGaHWGS9RRKlOgbg
j9jOVgPTH3KiZxtsXmA5JvgukQMVoxvqUZgqfEyV3MKKqDum2n5UhYJn6BF3tjJ9eMTa4kRgdIVf
1DmM5xuSFZkWHNuB54vk8anqNYccZGhtBPRJSt4l9riKQ+hsa+YXErlKx9R0+USGkb8FayJbyVE/
wFMTgIYMsGMfqA0Y8EKj7+GQQ5KOc0jbgEwYdliyamFQwQ7iscfL1S4++bZRDZPZ800So6bBXPWt
3+k6wTd+NrX1AWwhywR/Y5alpwzTlkfsPbxB6stchn/euY7+LXuTQeJkAydK4svHz/y3dkNeOBgt
aZclzfLqq6go+xy4MrHnVPZUadHHzHEjcDUFJXgiUqL63Rcb34Nl9370jzqMU8R2jowbTrtDRv6B
WomFkjgkVKIRQvUy9zVqBJIPg8aVXSaVmGY2RN8BeKGnud5WIW264dw0zoYp/hg7j6P0Q9w5Hno1
K2aRs+dehzyUiTabpKXHWbT5AK9eo+dWta68KKlQjgAhBP66IhOdqN2pv+dCcNbso4SG55FXwKFT
oY+ASh/ynQbtNDT33ELPMPViS2T4SW/3KZk2oJTImwDEqkge1JP+7tTu2M/jKEPJY2pghHxXZZAn
/YJsTVDit0kLaRb4IrERWRlYWu/Sip1ONLEvmxKtPrbBSddqfw0XItSqieK8ci9bRPRUcETZDmLv
Muk8TlELhyzhypDFVgGKKAwAiq1nBFykVBmBV7sdyPAulMlWsI5DdYvzLgQxpf75sCXq2qv0w5qK
3gLr7vfiU36H5ABYfHYfwN8uwrN3qe32efNLIDlaa7gCJb3Lr2kvuzWKsqfkeQFrVVv4euI4aDvZ
Y6eot4k0WPb9EjFZyGp0nZjBRfoeMXQfQIPpQ2lrgps19IfSTJN7a3kgWJ9gMyaGgPU7uskDj9X7
zzgcktj/bn/EW9tfb+kMH4Eo/CMzJ+kp62uryT+wL+nvTGOp7EJ3FfiUPaB63qHWsOT0moSUdBho
QI35fY1hYSH1NH3kJwdk4tnOYI82cAH2Ww25zkJ2AlrT31O2qToaOkqwPA+Rbi6hwwumMT9J/wr/
1vqx9r1QLG4UyMN/QVdyWCXX3NlRVzojLy8zBaPbo42lTwCWF56la+RgtcaBTti3MTQvAIonHzFZ
fxWRYATvHJ0yyWmUD+j2nD892K/gguLKE6h05eH6ovj5Uph06RcueX31znv2dldwiCkQfw/jQlVb
YCag5EHOnh2HQQWrMgTpNcrBEDVcU7o5gcJD58XATJIQHvpJyYzhJ+VN5R0ObpMDVCGLpLyY4CxO
t+56JQbP3GXpcJsRjKIaNISQ6Ny0JJ0DOltkZrTCs/vBP/I4i+MtqNAOYBMDlc8NEf11MLCz1DnP
+Tmcz9MWDtULq8qlUAFgxtbXcIEVJaNH/9l2ag72RU8oUiv+TI003FlJFw//AWva/QTdpEvNJ2vU
84XAA3TpDx+frArFJ8bBWP41FEAOAf3uPLKFMxiYdovFtVezy9dGja0yIwsT1YsgF0rZsQ3+iBtj
C0JRL6f1/GCT6Z7ASc2wRJTqFinfRYxAkzlyK8pvTRJHcSt5f+oCjTxQlujOr0ONto+C1c/fxUSO
8QJxPQVYbI4S99lI/ewf7cbrXCKgOT5HRbs1T8opJ/tWgA7VVA35CaPymHEiH7S3H3Qh/5Wq5ehT
U+Wu9+77GBwMxe9kM18JgQU3gExlrVoFQQE3nIFmaYJvTr5GiD4pCUl4L9ewF/oXK6UGaiqAdmcY
dCir5h/mwOglarAWMQetTSdGdVl9LYn/+fooPKzgh6TE8bg6Dke6YMRibZgPAw9esgMh3PPCpnEA
Z23kv3UrUYv2SJJkp4N1OZG45Ne//7uKNjGMdzhOcF+iCC1CAuAGkw/91ZtLi4snr1BMyEYuKmTu
eHCvKWmcjD+owl11aa5cKy2IJeBAA4qcMxaRqGuGbWChOm3f7Q9XEVViMnfPe9Iah8o+UPMHqNmZ
o9UMRWPErCX2aFpIA3W7GQ67vvEH5DlTC+ukYWf2jLQf/o3to5TNTG+Mu0cF4sXcbRG4/I/y2UTh
+l0/DfwDAPtlLlQ/F4AhJO1jm6bHNRzr7CV8VIIdiPPWrtYHCaW6qn3i/FXcQqhjpny53J2xFnUY
Pp3NGqfJuB6OeosWbBL9EBV6r3rXnWRWYAC03dPVJyYqnkktSpAReycC4CDWZb2UzzqxAxohQpdP
x5sQ8U/GGNzczPhNBsVBhTilM+sOySiC9S/VJXEagAnnTy4PVPy6Qu2rotIZ0BN+OZnnXjjUJ4oG
dXUVkNuD2IR1PQIQxF9rz50Zjdm9OB9j2dBzTcdSlV5126fxCD63Z/SJsMk97MfHUROzdHfcH7u5
1KeMyJpL7lkZeF4v1DFcJ05Pj3+1Z3xHQ0k7htp5e28pRC13LY9N8p8sTLYtUfI8xGn9SEmPbpYa
pKNeKuWgfoEPb/8JBohrVYA+S6omEsEHdOIo5Sx9pbYLfujSWAwIT6dMZLqEKjOsA/jI5pErmvI8
cWAEly7X6N3e65XoU5fKzcTbLdcLLCRm8gz7C+J8EgT2Ex9T7qquAm4DSHR41dO3KgQV31vYJX/a
ZQsxq9zd3oMh9r6PTgYQ2o9yVLbVes5Cpkq5e9bjInLlBCXgMlMgbm2g1km3zaP2I2wVW+PcUOIF
QT2eI7iRPI2oyk1WN5CGPeJhlvHJXByjDaI1mdRQ/ZfTFVAKkeSkdsN4DRvnkEjitq9zqVgcHeWU
O+e1qUzDzOKFlsmk8WHCpOQwptKkTPBOrPr0k+1O5gTxRZZbIYQxCouLQq5mFnYQu75Qmin0B4pR
sgHR+6VJGqemLIIP7P5h208+s/fKmGSqKBZXdcdkgvsidR4DYVCgQdezD8/LUuGnU8dXhl0r++yu
2YFcQr2RylmfuuvK/1NU3EVxp5sK1riwEMhuhM76M6VdpFqvA6Ord4ntMxlS/zAOfutjTr+yKKMj
aqNunNmXcNmz4nIuAl3VeK3Ih8t+J/xoaACHMWMzoY0yD8HFgqUBxhxhMh4kNTlS5tSy7ICqkLE8
wjzxMWBf9hOEVJhsMwRaf44ayytffOh6rlKN+KlKY2WnBC6QzP+kMHc3zQ63PJObTv/T3I/Pu1EM
G3GHzbBtCObQ8TJMGN6nFzYsA9PWpPrY2ir30/v0+znNBoOwYj1JKBjds+iHdlJgwPd+v8urhKN5
AxTJxElF6I5Eb2TTala8B+grLCG9PV4QQGxS91WpFN8TTkvhT8Duh6MMKfAUM10NTF6XH0fb7Lso
rk4NM9KCVyNFcNlHqgc7ZGHywz0OzGSyEsF8xmNtcrNvB+CXCFah3d1KtttGhU7utxv0/1V2BUXM
dMWRL7tYf+Ry66LZ8X64ZudWGu7HO/8tmE8hvdkA9Einxjtn6nuKtxMuN2gBSM+/iOxtn/gm9c4t
MVSZFP6meMnDBEL/VdYMQYw0kXugJIcCIqAhPpFLiqDBglSD2w+PHXAIZP1MPZCuDqJvXI0OvQSD
UU2syUHJ691+BFKmUJiL4pBmsa/k95hG+oo9h+wpicn/cfC0gqiXE8EMWyaJRNpgAWIxqBUedGqt
d/MA44e2g4RWETa4+6tYL+1Bv8p3hbuNhWj1NI2wSb5hd/lOAtN2oR7lQadwG7ZZBJwgF0NS9Tx3
RMNgm/jnQCjX10eYcNmKDndpDTr84LIsAj8L7l1FqqL46BAXvKehAJWndFXsqB6sS2msamQXMFgT
ZYjOuh/I+6yrFVQ+UKVQdlB9IHqyNHxANDa9c6P3UJEIpHBpE7ImY3TimQZtfO90tTpONtg9zQH5
ECsL/HOl/4ujpuwdeQVxJ5J4yquUgO+C9Q0QPNTE9U93hLhev5mOqkSTocGJpjRz9Rscdfu3RsSJ
G8qDz4bXRujnVNxBY/qI/dZKFx+e+ge/mcIHDA9uy7XkScq7EuoWGykD0I8tB+k4bnl0PumZAG3E
jCodARD70Lxo7AkaAiKdxbL04nfUUZtmdfHnVeqw0et0jakjT8pnbUwbY9sstWs8GyGVop4h3siC
XqUO9hRvelJIdQqAdfi/abUj7mYGRMd3jRPKlnIGWCF2Gtw6vdqSRKWRnckHyz4pa5Zv9drcmJue
DdDoeb3yZhGg9yHPdD3yHdbeYUAUb0fKr6y/W9mPJ+5lVmAgfXLHre6IOZQtQhUTfbG/u7kdDn4S
UBFcSu3OcVAqHloR8JbHQfKUnFXSOER1rFx3Re3eDDZwhuiejbSIK5cQhpZtcy+BVNIr+pVZpGqX
mLw6V/slmYpkofFv756kRtb4BALAtV0XC10WOIMqCw3zfOfi0/KT1lftFU4yeLDzpYkP7Vb4osHV
TOLFb8LF5ccw79ZKyihdlz1PM6CG1mJzH+nOFeaX81Ll5J9uZhTCJhrDrJkC83IOiW7IgsR4l6NW
Tcb/5ywrohUX3YvfAGnQ87m4IUj/A1CwjLCr6zrC2b/5v+vA/S0JT92Ln4NNcEm04p/FvoPhohZY
hrH60n7YP1ucVLfvHeNbf5oiV2DZjNIb75r5PuCgyMlNa6CX32ap17WSBtX4RABH9ZlMnZhew+FE
IPmWx+duxfOttdk5ONUqa8Udlzt7Hd3je61eg6uNAeLsElUv3VqBDO9CL3a82ObPjcPZbht8V8jY
xGGULuplZx93xv9/DMKNDUjpaNZejQqFkksISydLMibKSZdg2Az800jzbZLq56erwqofK31jMN8t
+N8zrLSqeK+pNvcF72zKj6nA9z6BawkfQLFptBhVhW+ubSEtNPYaZsmzc2P+3hkHhOa7KEjnaLX4
/Apdro5QeUKBMcS5xzhG26J73ztfw1+J3NxSOSGZ8IQPJ2Zy70U6YuTad2GwZ75dzMdsDzJowCcZ
uRwtvULUjGRQHn0cUMn3y3Gm7punTrMM/bAgfhOUjQqGck+uecH8QWZpjYl6Nv43aZ7H0xaW/uo9
kfbROmaWPcypaGlfbBCv02HxL2hLrpkFPvYP+wwTjFw+1u4mU/rse5QJYwcdl3jjuCGPGZ/zeB9e
gW+xgTuCZMVJQZFN4sIn3TCXpzY/yTULYM4a5MhWM9+qSbLJN4p8Les3Q+bmsxsnYzmif4gLaQCL
Z6TqkqBcJCQjzMpUcRsONbDj7J55P0r3dwKp7emoQ52bvkSk/Dvhd9pfa9vS8rMhKnFTuAj00PZw
Ag7ENEPVDmVOlQH1vUbRwkNimo8pxjVPfly53f96lYAxu7uRhd9lX7NJvRlXAIb/hqkut+y1C8HL
gL0Juqax2vUfckBlRRjoBSKAuOH0f24izgP4Ijef+8ktQzJlYCYv/qJGwWkZpMQm7DPDsfFkCWK+
/PUNkNGodsOsugPWfcEkDrtYc9YE9Be4OsM1JyGhcZPtMaDcrzkllF4S393jEQFfbZfRdu7Nq22X
BNSvAOVP2DyB9ovj0ZMJfESE8PgWaQWx822ku4tJDuo7aTZR4ytJ748rF3ju6Qt0YBt98BwUP6SR
BXoCRa+3cUBXp/CEFdcBd5Rx/Be4pHUPjzJ8Ne1MleNdZEBxF0fGTGq+8DTVOaYx+FHam39P9aYe
qmcS1HDk4mqcX6iK1LenhKU+sobIrZWpT7WDQFiFLcYf9fBAmJHwCaY75DeINWKEHWcX8WNZqYsK
p72/hSXTGLWj2/CzLQ7KOW1VDrOBS5EqlM8SXzJXjoNflqAOY+HsMIqsL0HmaUEMavv9QnSJLgye
syeJswcmPB4n9DmVA7a+EJ73QcU4Jyg5Psymg+cjRlIMqgFeEv50w2CrCNmJXx+F8LJAoURXHU1R
GrR/1JSXCP21hQSR1wBZOaup0IeWOyrw7H1RTbGxPxhi0WFPpi/Fy52jBFntAqVGF7hAadRLOQ4M
C0hF5FRiNjswfSRO7IskdmG1/DbCr2xz/Lfz6HhmL//Yuu/Vv0UujKYa44XoTeKznBUtfgw4fVHl
oi32GeYF1tHyXk7AvUkHlzs0+c0V72u8c0saGjMNfEGKJklKJeb05aOjjnmLE7tR7Am2c09czLen
ctw/ODggK91rP5bG6/0c6IF9GqGar1F8PB5y9EKKNCrpXSC6LMSOYqyzwg21w9CRjHrypnrQYr3T
mDQMfe3V+hbNPJyLT2chqyCml8cUVhCXrmfcIuT7Y+o2kRA83HpxZIXcJBDEVEzhehmi2x9OqcDR
LzWTyus6Cbptff3zhXz4eqlPrso9M40W/rJEwNIJdIuDoBHuau+UKolHSVx8HyJq2ic7fMRZDH3I
WMOBp3w5kPW+nLzpRVkioJnD5wEXP1SfgOzgd5SDBdhep+w6a/Btr97rBsiAIZ0RNqAlIlHmV/4q
6qHF64+01B8+OENUxFiYmM1LiCERRc6PxZJXtRvreJnyZUm4Lpxw+w8W6hTtXIe+ItjHmS+vgFoY
nrkcy0eLzgq0gsoBRTf4y4cSPn28/ca9pdN2HBmC8IGLjHrSPy3eqCWaaP8Uk73gMh/fIp/+6FNu
NssjjefpLqzr2adz2Q6tn6lmsZ+tcO/tM9Zq2Kw06xbZZur90ZyTYn1z8MPo3+2MCAP04Vu+S501
F32kDVF0i34KLq7BG6r4qPBUUQPO3HwkOZ3yB2/v7zk0iU50uImJ2mLoTPryCBW2XVlpr/zvhdSe
NQI5vo0IH2up07+m/i5xHNZHbO/d1IhNYrNf8dJdBvQ4JJYR9golPDLCyRBp6wQRCxACSDG6NGPS
e8bFrQk4XOkXp1WcZsNWlfQl/wY9kVRnhu7NhdIOflbegLAMJa0wsVRaMMwEWe++eMfAsRPmhKvd
twvxC6Xol2LQEbXAO+bwMyxBd9nbA7pE7Sq9h0GhhB20Y7m9IXvTRVN4MY7vvCXzX+BNxyytJZju
smh4DixWVBwR7nYTFRC+m18cLtf2lVvQbLpeYaOff2DnqnZHWjQlnya0zkEwg2OD6k7ibIpE1CMm
IQgNREpFOduYYuxjLzvwc+Y/3oBdwXLJWvxC0K49UQevswd+Ye+Mnk/jB69qeGI2yG9u1Dh3998M
t454+4Sw6dSwLbCZD/DrCry8W/84zoSaqf5gwuzc+VvM7N4Rkay2dTCwVPuFDCu2eBLBXOe/NMKc
xMNDKjfZiwdl3iipz8yj5jp0Kv5VMtZPnOgFfYMf6KBs07LiNLwCvENaKA9uD3mzJ6seLts5dcpl
ZKdCXpFsCzwkSVdIidBfKQ5FaU+lwpefDbruGyWVDyStZAoAuLL+Wf+KMOcR/6PzmmjpS0+NKXxe
TiXoeq4XyC3WRJ7xcNxuB3YA7mJs6qIHsPVgvAAKIM0a6MfXlr1qhIpIHkajT2c49ULhkKiT/wj+
zCTVwTpzm3pDUs3WBrxktnmauXgIoS+oXfuIdjWFuHz6ZmDbPPxd9R6YMHO0rJUGZlYN8M+DqDQa
Wd3a44/PNfC29J+e3GMg7ZqQXxzn9nXgZ3xKIczUZ06LFa7E026EuvEc61GOyuGe6afEcr8T1dKB
/IOpQyhD+yMztt9G/7tthOswK0bpzg+5bvNXOPdjIM+V3Ngc10IP7acUBZiQqCzOBAi0y044N7n/
fOj9HrhTI4EbAcmNl+gVTv62JFsjprPXAF7ghlUmD/6FiJo83VdpXk3gNG3NKEU+R+0rbHH5XWLL
v60BABK8pJcdPiIQeGnxU8WdA3uioAYf9Phpm+GtxQ4ZjRztEo252H5jWFZSal0SU10YVAOWI84Y
mbdFlGaPi6l96z/lDxj/iE6WNUg+u9OyqIr/44drmF7F86JvTPDnYlgyVFhZF0LjnH15KFkqN+kD
DGreOqaOClm9rW8XE6yXRstBiPYRfqQZoHUQKOU0lmu1q8An2Z2RJa7Xi94LiQTyvxWuxQs+ufYd
7YcUwD/RWxaBlygbxujkzCCxqbtGP/znO4yo1NgQn5PF1mav+2TElzPcBlqP3CxKC2Aa5UE2QQOl
QpuHP6bPCASA/qivnizDKyz9G/Sd0e+jwUCbR4CC+EUBY7EqydQ36x1x7kcDOAo7cVC0aH3iPKc2
x0+zTC3X6JWPh8z5hqlEuYMZpjIOdjXVIKGWQk3gS3AfOTlzfYzGBkhHDjLKNt3lizEAdQF1Eghy
5LdLBGxlglZ6M63tb12A4/MBYFH10t6Cls4KAtpmWd52GrW+n+AGgh/BLarclbsWqY7tk7UyUKkF
ANy4hPmvSf0UKaZH1NN3tH6AHRJlILnwDr4yh6O956pam6FscM9iFWh46IdVLlfHjnODBGst7nrR
S/At1668r4zEnOR0FcnXu2x3HoSmTSGEAWvPfpVbFI2UURxTTEuf7nyoivEpzLvWav5m709aEZI1
DIkoYlkd15SBxdiemnat9wUecMCtgZItvUf4iPfV2WIQsKbyks+U4jAMlL2sO51ZSEo/lymqOy4F
6J1jYSEz6wzSDEGF4Di6CpDigdxJN0iGX+BpYCcyGodLmzG67BboXZjRM1QZiupe18svEjnOJ3I3
450mOqyRTV2S4yc80t4fF0v/mP4u5lbDYnKJycdTxlvRq7hvo5VuYXItmw7OoiPZFZDZ9+wLGg11
GZnJZXHXDzGEO0AD5ukRj3AkyVW8YjzaBLF3pVBxrv5PQ9km8lKngAA1VG63XpufY/JG817HtKnG
LcA4WNmJJ6BLxrKzpt9pajAKLe5jUQU2jveAAJJ6lCXhmljg3CEC2/6ONm21Tikb7jo97KOPwodL
InX4HBGtf6R0Biul9TNqkh5VKA+Rm7LzYw3ZpE3hB//NTIHbAG1IK0UQivBql1z3Hw3jHNZeUoFR
8JmDXImRiAYTAc2c/J3+3BQdJ6DfYr1e6VupVU5HnSrYIuh45T8Hs+w3FyxGCEJpd5QZCxv2fuUA
s6wRX9PXcXZQyVJtNdNkwfXm1kOk0+JkKBUdkWlLKiepFgEKUCim8XI98H+KxC4h0/Tpt483ug6D
eaRN6yZtu11aVZsUDyMj558YsTQ+EwJdMmxV0gn6VE8LqVOAonxoXv19WLs4pgRNFpVtvrN56xBO
Si/V1/4A/vAsGGv3lo8hBXFIlSBYeaZubpKKZUhHyphrDuHU/U7Jlzjr55vT0Ss/oS2Mf/mziktU
dETMNrH5BKVy166FuW7gK39vCO0Zw0ic0iDvhBjpDqpQBVRRA2dKRj/IXyTudqgfCpveRprINGfM
c818AZJqJbLxd+UvtZg88cdqcJO2Mc6mfWohwBPmXwJToA/wePTFZ2pdGlKdLQm1STPhErcQJ48w
BwX6D2lUL3w4S50ycJLVN5t45Xh3um5AkdzqYHLgqMLDYJ8yfvcU2/ybs5binHpCphS18uMx6S4y
NwAMXSFBC9mWM8E/xvBG9fQaeTAwW4tLD2bM0MQ5hrxfMRtfORzyYw0bAb62PHTLBYBCSDv0Oug2
HRz7YmtxyCC2DDwCdt1SQG9X+Z805L77lcKlWdaetCltzdpcQb4kQrKSxFZ9sWDnq3xuy6lj5XwT
0J0KdXh32tWPGNDbigob3Xsbgf7lYBktjYFNC1agAM54HziE/AkAjUJtUVoLrv5jYzQDEY/XGK8F
pNS14obb4jF6Al831mw5XNvsyJCBW4XlYXqEpiEmGsvdXVYTTFuyGHI8jfAwbpw2vMgW1InyHaTq
R/SNtjW00EQfCMZm2svhTJgXmYgDKdi6ETi06PdKwqVQv5OXyqzl3yHzsSogYpm8aNJf5VgRA77F
aVASmZwH+sQMkIrxudpUSVI/cegBPAaC/Mj7267PZbeoNwaKO5Lh/VJ1sMEpHw6HKc4LAkewuavk
uxzZSyzYb6ugimw+F1j5vGjJ9DmkZvBc9+3s2ipFKDWGQ1Rs7zpaA2WkreY+JhYzrOYEMNdtgBWr
tdvq4XziFDFuVZg10/1czgcmexsv9nEYmXcz9tQBMm2mb4ZOX8maIfnCS6nwRBH0QE6UQxxLIBxt
Hjkf2uJWLTacfLf4AVnK7Ff7yqJtSaoXov9mVnhQQ3R/RmH+2Cj37sUspMcmcP8Cig/qrNnwQl/q
SK3S14G51/3tv0FVmXpuNxK4a5NIo/SI7fbVLgZrsTP6q7Ew40cFkJdY62K5cEdg3u+SRSoBHkQO
1R4ofhabkYmspADCID8yaBC/6neiBpI2ZIIwZ1Rt9ISNN+WiQcuTP8bxzlsogsYPaFUN4HkpZQPK
gEhipWCc5+N93kWHGpKjrw0q+HsEFyzvMzv8IjI+jYYCDpiOn1Dh8MU6YvfwEKe1HPBm/EGtifWK
2zuE0+bAbHdbOJUGFLxu/o6LOcON1pfVnQH9UFJobkER5JQudAhwMYa/d+UbdnYQOcJo5pdVDv/y
kyPoiZvZHTJc2UlqvIsMOuWQ8Wt3g1jLLRFTs41k1zhjsLh5OkPpKO3b31qgyS6rrKsdxQIM4h0W
/68stGYVxzH91EbcTZKBc/0xi8PoJnQBmLDyvOQ/ErvY028GLutjOzvQJBYSue6syVHV1MWvKojx
kbRY0qSVFI5DLSemBHODCWHAZ0nX4MNF0uT9chzC6PQa4HxmxXleB1GmHrVIBg7hBg3/1jkKkxPO
6dMiseMwwosCFln2dKbxskoV21fFSJcKxVpLpgAaiwzZ48Qu/yOeNpDtDczeLYmwyL8Th1Wsb6DG
raZ3rWVKIaZCgjbViV08VWCoqFo3/uYHpzpReTxh+6xwadWt0RbNG8S9qq16P3XylMwmmi8xDeDV
+pyGuPUGg6lF1KjGYXBAsJSv4AJVulCIhu3Z7RaKRpwTBx+cYU41OLLW0x51kKprEQdCZJTbaTIH
IhGG8Dhg08TrCQCwp5P/ktT6iPlsEZS784sq8zgjUEwQ54m5Z7taP5mlmt0QDmrCOWF6pUKYXuFp
01b9AgpryU9/vAY2JBBXtP1AArHJvk42tKJeUBjKOKDTAGl4q0By06za4OkzjxdwQcuoSdd9SGeo
0IFErPY2IYmSLkPWoAjx3H9OsfPi6JM1qS3rwd2/z37d/2xz/zdwGIG6mf0bJ8eLlArYPx9iaY6f
vk0S98PFS3A+wWF2C+hdc/NSWBoIrW44iJTvU9RbgFKSxJEX8gBwOXgIF0C2O8C3BEOw5ik729+K
b25xR1D5zzMfxBSqKsIEL4f6g1clLetImWVao170uylI8+fzjGEg1DsbAiEBZdbzt4nKCDJf65NE
va8WDm7eYycHcG6uTqzQi8/4z/qP7ikAOvsr8STgrvBr2+y2TQ+TAHOQSQPu/c+iLjIC5jNssUeh
KogxK5LnaC830DY1qLLBms3QTXXWeENdXujKVBD9LMNt7DhxXGe5fswFE2yc5p0cK9UK34jL6lsj
g0Yt145H+ANHD2ovLdq9Rv07KtIXxJLzTztuDkjjtv3rA/SAIawh7zj9nvPaMIzwWQ9Hl9uh9552
KVhxMJ5ib1l5h+i3xJ7pnXSnIBCJBogjBIE8B4hLo6KlKGJJmxcRJSOaTt/FpzywoRow2Dm8f+QW
C82hnLC+PctIv0/OzupiTTH4dyNT8QTlEEGJl8ckFoooBcyP7zWnCoMyeyBt6yOp+CH1KcbtXeRN
Ap4BYu2c5A4fFF+GcJjhDMnvkyLdBVb7KQS4vmWp1F4HTDCsP12K9LgKSxpP1fPQp1Rw8sECtqRp
5SbSFiLXXfP1Q6cIVpKhinq5rPirw/+YHOQLljj9IU/Rkvf/LDIC616xTg+3qIl65/Ms0u6A5sod
BIuhM1Sn7qXSo7qZskC05G+TN1mpBMKblTb7sNis1GVBRjoQEuZXPt7Loh02eowwmr03gwEVVMMV
uIHgYbAalZJeQJrjjEaD2BY/A16CB5xxOAGQHcMcrQPQc3jEi+WmOJx2VHRt++v2Za4SICd1FRxG
tY1kp8eNJ0xBKry5uS6ikVE3ZqSiqQTExF1PhvgQGtQFvf4SbOnwvIk8L6GHFApqfC/6JWw43Cg8
R3HDsJyNYx2/SN5hNyPOplSnnP6GNKLdnY/mLPMJwsos+eKD4edLpQSZoL8+tsr5UYso4iSxt6uK
HO18c85iGmCR5pVVIypjoX0uduObdEbaJ5q+fM5hSWQjduGpYeXn5mJPQbSyKpkHO4AbhuXzWA6N
hGkyNKTOwjXN9pblM/pjOkMFQevbBxYvS9Qr3XptzNboCUWTFKjz5f2+ryzQIjh/N/qICAv3osXE
QmLW2+ImoBsDxjisKXIvETY14NAedvRjGoDtXUvNTDUnlAeadcbwGod4XprPB6n7TFxhxIb84IV6
mkFTcY4cLTy48H8XDKQJe2YGNcoFxlqfK9QyrCvWEpfNpcc7cMisFNLn4VScAqX0DUPaGPXVKbxW
gv15kcOOWL5o+R8XA8RA5E0qmRiisucs6ri+XqO/kT5Yxhesw18Q7PHNMhANLQ4vC33DgbR+LvmG
zANblMfx1GykTO1r1a9Tihtf9BSmDp+ImLzV6Ic7+HWbn6bTUwylg5/okTt3+N+Y8aK0jr51TJyn
Ak+F76UN7CAFqfAadegRsICB8lcnSjR0dwd3laUWdZf7g294c5Tqy8gE+3arTVVsuWPwo/zcrdy/
IdSqA27Ppzobqr1X65pn6dYhGQehEvt8w4LSv9qc9lqLUNsKoTE+4k404jRkj+OrbYfwgCgidApP
3KIoda383jumiYxpvd1XBkRwBUzsEUGTwcP1m/crLO2nXsznywtJXnT/hgAuN4LvVDUr3fq0EYKf
rq9qNhb5rq5JGr6/dVeGBDSH1MPHfvKuHnL3Zmop58F3R3g7fE9p6kC9RA5LauTW696TzTsYOL8m
BFGJwaf7qAdQiAcpw+qYqxihHuRAYMyKeDsE0tSvyi9mte/Xi5BgKpirtgM+wBXrn+37niquWZkh
SbWO+Ruq7BA5Vbqlda67YG2L8sGbkD6I/7HwXGY4mnsiEBQlYC2qGDW+1IoHlqHOpSymHKYnG7J4
Sor8Oyoe2y8CNg3HBUIQnu8qTksP4LEe2aMs3uzDgaqewFsO6/M6/tDYFouwZGTxhg8xQu6lEsDX
G5f+Vx7pmrEqcSaULpzT/3+Hts7JpOR5fGDc0S3CvC9qO9GitFY/a659V+YC//hPnsq/tlSfbiUW
M6TbsfhzQBZzH1H8GotX9zmaZnccm7YqHTVkaF4R76DoElKC7w2E4JJl/oHuKCO/28RWmWZnUuGy
bNfERoG6QjJim2vEp1xady06SBYBGoJriJNFE9Gii26oJfzUPyICOqQyoIBsWQsYy8l7RQioyMpI
bFBbSoh0lzHgBHTnzO59H5iNkyxcipirMJsH8BU3WOCAgefjiqghJjqk4cRJkTqt/TX8aqG6a17i
i4vsKOsMTaKSIGB5EC3NR6Qqu1HZUj5hNz3QLWXLjhTD3uHdQvhluzD/LL+AE8qvBVc/9kOhSnar
2Iz46s7ajgK3IdR4BbtpC1LlxrTMnpuBbpIgyZMqrdTdCz+XGzI7STpLzf94cv1LG0mLz4div6vD
5KEIXXR53tkDVUjTi2HsNizyvdPu70m9d2XuMjdFwwU25RedXiaRve0Aiun9DoA/Nv2/WCZrpWhR
Y3Ed36G0vzN4h3cbuQ5ZJIYM3fZyFcnN/QzzteGGkOcBxpx4unuZqtnKedc+fIEz2vgu64KwaroD
KzNCT6R+EyL44q6mvEEFbNXICGey+nEoB1nwHrozg81MHhSdlbeT3WDHSBu9uSP9phKGfoKx6tv7
78i7IMNfR/t4fPpfwUYNtjdGf09iOn8u9WR3NQq5BAkidNvddXhqy4MnuemXwOeBglDceaJpt0sR
uN0yjzS1hxkJZcemSXm5PY0QcnWoF0uW0kqbM6teTasipipb3KG2EIcADyqtFU92gtKcvm74yt1l
y+JyKHl9TcxRWWnTKHcIxj687mSLxS7CB9lXSE1vNktkXv/LeRjpzd6W1QCovMaFNPVzSsHXJ0T1
sIHDUs+GVB75OA9X113BHKu9pVDQf+no4rgnpAqdqNHkcFVLJVB8r+CZOnQFSQhycx7SaC9h7l5w
OCaIRerGq+pubphi5gMHOh9Zudd551efmhnSUcn4bfBltGlR+fjLfXRwA+7MMPybOXAflHivXbs0
qdtUnE7VbBIw11UEY9vF4d/plArSfdtAsqrNR8ze76Yc0e+Ole8693Ird5Zpw/5/GbtwFOueBJJs
HoxasWivPS4GtTmhPqqt1574NgwGZvwOQez1OGmSXEOG9Lm1yTED5ogyrLeqabKXNMKw/nd8b4Uf
QMsu3CpiWA8zKLC8xTKPjOOLgHQETPkxWi0EJi/afZ/xb6d/2O1L5hqcGa6XA1w+15YCqxL9nlVd
WJ7VWIQq4/rWwzhB7/r5H9ovDuTItBLAho/4b0ldEGKOblu9LmQWHD3DOQePnteGzR0jOELg85Z5
9mRiqLW4lzjx57QlgguksN9/mc4klkzIgD4dtMr6M0O5dZuOkQmildOjuEQLJ0oSVlyqCBtnvUIa
l4yVHGOOdbMOihRc00qmWqdwuJ/6BUIyOSzR2tXtRD62we5Ryi5RWPXQjbO4/qR7CLryqRxuC/pt
4QNPgkrqQYrni1k9LJ6YZtBBur4Bqd4U6x4JJJimhs2AtSS5m4BHcP6MNkWN5VlUewt82ix8SsQV
9Pve2J0JQjUsjtCfatCny8oEBi2DIdwGC5edV10IwKJY7zzgRIgOZskFyO68xeBmhWcZCaB+NU8a
TzhTYxHusW1/YGqvWU6AdHGam4DODcvBsemVIMDFq8v8lscrnnrnAINKeSKQtmcrASmOMOn20bFO
BO+7MA4lT6xtlO7DkfW4YM2AX9LlQTnYcCwBcU/50x9NyhFOYc3gJztMPXBGR3qYGRsMMPIHoQnV
E1zWi8Zq6xyBoWqGLFA0CDv3EWiabzStNWtyFGUPBRJ/pTzQXEI46+9ZTAJ+TJJJkuaWJWVN5Byn
9F9k5sK7X67FW3L28TFwlDckMlxPoh02+XV/9F5wljg+idSxUIPojVfg7YM75DIU28k2SDRyiRcO
NAF1nkQi8dpvmvQVAe+gXxbx/b2BIqesHgQXzM/Zlve0u2iF9KQspgduX5cWqE7JVrPGU1C6JPJ/
yVsr6+UbQQ/bPZuBB6FuYK4BV/U1zMmJyxfwZem94DeHgN7upnNLDxyBsEOxRAQhBFNVXWTDEh2h
pxXJR27XNDLqtXn9oDlSCJ5Wwufr0h8q1Mmw/Dd8bSNmIOdNgFcMStbk4nTzRFAlp1YgspV4JjkY
+3DnOnfsJY78NIGNwhi4qvGXIhZU6MwT2vsM3tc8sCYoM+U7rfTdb7TDpoYsy4nWRedWcVLqPUuD
WISuKNjtciebWME1LztgAx0kN3cpiyRYL8ps1PT9zn/HYZrotttKzR1evR24/G7Jst+DqgudtcQ+
QgeFxQYE/OihnqJZRYKlyw2FJfpA1vewPc/pVcIScu6U8eUUUjNDsy0Lu/fm2oicNnMi6zMl3DFT
1COTn1XiksPIHIz3RvJ3PBrVj/WRjKleBtpm+z5keuR8/QgjRmUMaObrRibNWzYX8E48IEYEWvG0
e6rU6GNbtwP7WEWqNXmPsNOhKH5b1bo9SDTo65irNO1VSh9pJyEhkcFquOOP8l4Fr67TkIW6F8X9
iFXaXpRjyGg4NIGQ0CYtPTa5B5FE2sPPgLIn4CGbY9EqjCijHfx+9Qk+0rzJnzPYxGqOrjfPbhqQ
a6abc7rHNHRKwrqRrmemSkLg60laqX4fVjUgNDyrGw9j6upwN+cWfFVG01PRSGvoMzqynoi7lnTC
FLCB9aGG+6cDwX1ajQ/kdSz6S/QNHqRzAmqybyBkq9MfkJwVGtK3+sbQFoCOcGfyRF7CPTxV/yo2
8pZBl6GpoePRr17ciNllbp6JEY/zdhOMeTdyeM8wS03eox9eQ2PWc3EnXRJ74AJGrL7GTDM56Fvt
N0vAJZ+gvLQMQSW9aZzgJQhobvMDIaaPGGqlqEdsWHmImK1lJYrHqY271OtxHDaJ9Ex5R5vMiziQ
17NaQKpP6zF0+Yv2zMgVMZ6fsDMJj0Ew5uc/AkpTXHq0Z24GqA4QpK7PcenTfWTCPQ4sC/fJb3PN
FtvJaS8kIrgBdv9H5KH3pIDJHZ+/qnrb7ywgR3GKdVLn8c98rPMa8HM5edqecbRzwNiWFW7yJ9Ee
ZLrCSi9sCR9Y/k6dEVLOdlt5sh3IKaWyDJIgTV3cIwvhpoEpqkqn+BxIyXmz8+QU5Dwj+UpE/n56
HfHr5ARZPvJMn/0v5ymWqzsPf3HZXP45hgeN0vGS3Lncw6YrjpDem1kbkpwgzQsphU2mAApqPlKB
1G9mT9jZB3t/Pn7RkJeNf2WMi1COe4caGRa14UVP8FoFvEi+3JVitcBFEtPOTqK36w3Q1HyTTzq9
zvvpx38uK46d/xV62vyLClnEf+U1uG4tb8TuqLycPTV3qjuwhFbdXM1FEjHOj4I4C670CsI1Inf0
SGjsu4/+EhAHPJCVGi6UZSfffkUXGJJ4xhgAoezxDdZY9LRGud8eYskDbUvh6CUPHwb+oQom5Tvf
k1RuelMALrhTVx1XZob6ziOvdep2qM3ieqZcqPWkbVo8cslqRnwbd5eW7mf0Uc4DHyUaVDGtWceT
6YqDYnS++uTll+Jb23hx3BSU3bI8d2kwSPXgc1iy2lhDxX+7R7WUGefdRECTpNbQb8qrGzGKgXCt
qBZgGAQxy98u74D2NfSGM3gQAT7xeddw2fS7gz05hjyHhoGYDGrULFnjUzBZChE2PcOo/H+N6Kpt
NfhleON4E05jWEt8df1Cvm4ESwVkPk0zzb0U0NC/7+DSq/ywXT0FmB+vnAMEKDU4P1eP46FzGG1M
Q7sGFACfoOuFjGCZabZlSKOSf5TL9mLtGxAQizWkpQDZ9iEyGEARhhRYl3mTPI0t2nLAx6Dwsq5v
s2xcrXJwO1TnEaxmrXuXJjMsOboG3b4nduNMpKX3IwdnlV3ovjuchEuiuWN9FZNTtTto9T1RL4ne
kVvWTdbCAMsrCjdYf4EV4z/4jBFp4FC4ZQBcQdn3SKuMr+Iy3+7UEZN7hrqFmub2cWW8bNuOYQrr
PxBZb5RtRgANamKbBYkkIEv90i/GrJ4sCNil538y+aH8vsLu9spSvUmGQP4t9747+hDuEgBGgRGN
7tuhFBPPtzvRZCIB9iHexUikDxrw+WYpVcpdb6Ozmthgypp3fSYSOOpCmdL93PbwXIajyJcQ6CRp
sXyRTmJIotS4qREjzrFlqua37WPt4gZHJ5j/MQmNaKaK9OA6/E32xKg2YiN+6lwJKb6jjx1mybAG
0PCvji8mSOZpyg+a2AQryoEgEgdwwppovWmgq+6GUeHENu/5vwD7P0wJhL+L+XsQ4o63XroCh5NG
tuAzRZnNJvxGfK999PBOYk+eoF5tQO+WULoiqy3WlfHvcI5DLDWt53hKeNx3w+84b5/gU9FBkkNV
pWHX2gqjIu3RQezS/lCYbjbRGIHpxBAYtf2PZXirRYLLO8zHOpgDKq90Z9yHHWw0ZcfcVMNm+8LE
QUk4JJkBHbHeFfZfDY6IIgQtgfUKNTjPr4h2PmVqA/HA8b8xgQOI6uKoAUMVwpX5omZRwm+oi5mh
VVt8H3UpmlaEwBlnXwIfrWUT0IVCBv23zCgDX/BhRVLPDRFZ+dIUjMzjA9IobXZwEGq+TTlWcbVu
jVFu7KX9U3kZM21Q0696XZixB31r05cjH+AQvDPfXgIEmYYHBP9rPlvu4i5w2YGoVovdcXeItEzx
bSaZ/OWDdkitj48n0dwJuu4Il0M6gfU3adBe+6pLe5EdeA5VDhMgfBp+0Z61kZ46KqtWly5bfHPI
i/wSpuO3piagEseDC5EziBWbjKIVEi8hmBbML/sE1L2iy7HrlCE7iodNKcM/IBebku6Xu3wh//y2
iQlYE9iRBjqakTw5sqmS012Tsk/hjPwQ3cTk5xhhPNNLk9fm8S4ZKCKJFZMfe23uh5cOix7mVKWN
Vw2iiZ2JG7C7/bU+wKDKFi2Nkbp+/6fJqHsRguyHP3iWEIJZiHyHGIstXq6rRi2ojThtLfdSiVRo
3wKrrwsgKJ0noktwYwolufu0aUakf5dsIjfalEf3xGQ9VXlkG9YCyX1TW7sg4zxV51syo7cP4oiB
LH4d/oith/mowCthOrKSPvJ3JpqWbSSDjfLq3uJHck3oIHbkd3DBdYQjNvIfRFBYONTdPl9GjqBw
Tl/kmU5qLkuJWM7atWD+21f31Bd6Cm+cXUIk/MRDUu9nEJqbddU7199/zAKrbmNBHGdba0ydAxJC
VWuAlihGfHqW8iroQJvUGvAo3geNnmhwYxIa/t9KrEIzWYuFhPrNMGvqA8Br96GJV6UnDFR3Nha5
sVFnnNXc00HOvFjbKKLKGuIcdV1uF3zX7bFtqpTnJS98fZwgCh1NAm9PuE8i/HBgY/e3uPjES0Np
/btvkwEu1yRGYvnY7bjDTHivTgL7j6jYE1dHgi+virP1iuoSkUYy7THmgT5D0Nw3tmb3LA0Mo7MI
N7lJHueSt1jFpzFkKz43T3YRSQKO1R6oR6QeKZvT7bu5ezltmrmUkl6RpZHAnaX2P87+KnoJcMra
llUbm9wnaYlDW0Kl0qyYG5SVw9D5mye1HS+HFyzyBJC2f/2v9iQpGkWOTySy0F+4jID1gdhz+RvQ
8R9j8IAp/xfsHrXxJW7RF8duMRIsDB916zOEsdDwJuSd9X8rFk0jek5uzLctBgrrA+xbG4xCgvfV
c8WZfAXeowrp1Zsg101eqZF4RlQ1I6GHzaYNQ2DUkQvLsoy3AWehnoRazii5yUhJizFt7u1aUQ27
iI58f3qhnxo1IDMdc4lPVlICmDFTjBqT8aX4R8lWL5efdsxcAxd6WQhc/yykrPNH00jBJXnDK4aD
OCDlZ9M/mDZYCddmN4sSqNYDV/cY/+MAD25UGALnQ0pHxqR+X+3Up671SVGGf3SLxduQlNdWvcmo
7iEfBjOeYAJL/7P3oCKU8ACSLQmQPOWAXQCv/ZD9RHokiEujwrT5Bpuu2I73hs0eUf2dXtsdW3Fr
/tBpmWFiU/0uwAkOfrVIlB++MI//Ankz3D/lBMSVR66HQamG6yGzAgycjlzcQ8lUwPQFVm7iFPNk
iGnxjB1wJ8SUUcfO+KWjSYQ3IWEjFsiopKrOQ+gIB4A59V8RZJS+ylMOOlu9uqCZDwvyqASi2mFv
/hmA7JPMuSdI9aWgOTjFWgtREJwzRVR089O0yGtqLh8o74oE58AYiYA44mJD2Wcu4tK4jBVnhdFc
HkpNeu+5WJNRrU0CEhqEJLKeUOWTsCio8uOHNlYfxngg7GSzXuktw9dHxDR+xY0Vr9cWCMbKjacJ
8y6IMyNM7iyxz4BfZ7qjT+S6m+Zj2poO3sICwJEznBm7XtEE2KcmZ8/JCmrK24ImWHrA6jUW38BE
qE0VKQ/Oza2cFWEywOArQFK7jxiKBLW9YKXppXX0DuKlsk4f+3jSC+dEZNM3B1V0sbJhi8HmQ1Pf
RpXK0eklTJ8ctlKwpj0JFL+hedjI5ZPbixw0VY7MruF1CShB2wiTraIEkAmzogSTrGwtTgQieYe1
5/evcYOdoZ95Go0Vki8KeZbjQ9Fg2wV3EqxQh4GG3PT6KIL9riTFQUJgTRLOZnZZFGwfVmwLK+7k
HP0oX+evARShkwb2fIXU5kDNLnW7B2O4lJ57+ESzo1GNZIVcn8DwnUil8VIfNgehx8D2IAlPT1LC
S6civFjrNZQ6rVNWX0XtpjF6GyfuccwwsUojY2Qt0X2Y4f2zGS+U/FtTkg1xDEF3+HZbQ3bWj5fK
8Qm1N1IXW2sU8O6T82aV18UVACalW7TdpoyQK9os0FbZ77G68oCK4edYi3ykLAdUyUHTVdOK3HIz
DM7RqjAkXi3MoLIBXz4fhBGV2qRqO63a1TqH9TeGRk4l0XN5lIvCFaHIm+YuQd4tAKvKhiKuQoAY
S7GkbKY+UCh1pd1IH6Dvpw4xGUJEjc3eNnPRQdatuCrG08kgJ4BLYnSCQtYQdvD1kS2eZ3mgKViI
k+K2rBeRd8a1MniVWLyt8YruJ6EJbM6nVflL3GLIy0ZHvpZ1f2Rt6UUS0uSkuw4vsYgxcEu1lloq
qA5l75XXy5rTRuz6ZMLMbY0R7SocB/SPNJkBRk/m5S5875xMOWMx9wxSHLIz7Kr6DrcvqyIQCMTa
PtXRvOmRKFCq6ZbDAb+XSo1vtVIqrrgZBNTyf998IJ4DL+Dm5WvIjwwjNJPAj0nF6kVxTci4zlNs
2pYpYYzc/NmrwwFU6ChTRyD4dXOVGZyS39nLjmjpP+gUqkj3EccpXmdnF99/SVaukdl7sxBfo4CV
qhLyhf6yLYJZLFweppxk3ehNiOARdRTp3CwEu4yd6Ea15WFJ/mGU0gqYXYHeoKVAk/uuo4S4D+GX
UsH9CQ7x3DNVsgg/Tw04od4kheWKqo650rVKRW8/TmfoI53LWl1DARtrt0gszJ/reVHCpRl45B8f
xRpfRPeloPnHTWoVmqnu97K5P4ue1KZfvfOvw+gauw450HjYnP6Twmwpk/0FlEWmpQV4r/I32/Xk
BBxR/JTGneXHKloZ6e1Cw70119MTtaLkEgM6Szcf75K5ElAy6KMp3Ns82Bj8hIa67nP0BnOqXRnR
+I2IeME3rwMPVQJBdWt/lhD9qAIquphDLcaECXc4ZnyeTmLN+WEibKfQ+7Ue8jOtBm+gz0rCMU5G
LkWIiZ1dC6dBBN2IsWutuMLG6AvQo96tkKEgp/HRRuTwf9B+lB5VAqrE3z+atd/kn7TIRkRwVY8S
ANd64qVxL6gGPiT8P3Nv3rUrv2HUw3BOjNYuXerqCgJcI1rxFcq+SryzHVTf7xqkbCPMYJUZMOGj
5br3+vtdlXEirIbU5aP7IqqlA4ZFmZk1jYTRPVEvc5cd+j+3E1paQEqyp9Y2cN0JO+eEguA7cfzL
byINf24qc3+d0ZX3/dhZi+vwZ35hybBjaZmECPkDgDZsiv6idu9g0SVp4/t5w7lkOBxVrkLRDyf2
xuaq0mf/Okd+y/4ZPSk0bcnrjwpoRXmrOl1Y8MSRKwFwc2HrmdtZXoQolywmP8iv9pwRw1OO3DuC
kW4eVfO92W4T9yeK2XwpBE1hkZz+kPZx3r8RLmVTa82jIrQKkZusn9gjpw+poDq1uOLp/CU6vfHl
Bo2YKzmsOR3L1z467HHwP3ukP42ty7g/Gv+uoGJkQXTzdyICtIrpvfZEsrOvHRKSntkt/K2JqP4p
Wkrigkc7w+n0+zYtMBwOxGahFAvbiP8FYA8pGC2Kn4dfM9MBm7icXYJyTxBAqpPNjjfFjHb/fh+a
z+ZFu764ef6a7HOudvLGV051f0YzEKyjW5FTg225/mM5Yqo6NMAzo5ttF47G6CnZJheWVRUwgpvj
KRCIVKiCoTNM+qlq7ugM8GX+8qpjKUgfkX1VZnJJYzQmItwLB58uhKwRyR01Yk+PHoTJScGkd3kC
2OBvJFXmgaxkDDMJxjzDcVgz1WsTofU8LSX3jkQtIJH26jsNbcIYVMTPdnKK7D2uGqnnGFII+CKu
GN7AlvykyGEqMMgprVn/B/46Z/E2YvFlRO6+PZoGPWmr76II2l1HoT1lt7p7UOorG8A+7Sb/1cyn
wv94LEDyZ0U0S86YrmaFOh4AjVPWUCTVnTH3T9GuhDA33NnV5jnj9d5uwmAk8hePlDMKVeOmRO45
hIob2A1bfeWOfUF9oy/6JIGzEJ+b2RdykLQ94ARJqcOtshs2eAk9ZywUgVZ19OVdqno3eZJrktG2
JhWDEBCwIUTE/KevVlJBZY7fuOLkr28nc21T5q+PHkTJSNeVgTsU/PCSEptAYp+SfQpq3T6zZYRp
IOZKZS+cwmp6zeu3HUyrqlZAXmCA1Srax8/NUAh/ufxbGYTF3/fl0k/7eCtYHhz10ejWnXQGgaOu
ngfzYOAVQ36Ua9iVM4ie2K9VnT5fVJmjwjO9qJHJPJv4Ie/AIuMYHbXpdDne/B8kdw0yBuXgH2ej
NlTmWcCQeO7GbcXQoKVWRUsKLAFYT2zUIbXMpwUhfY3R/xwRlrAFEcf9lWo1AyJLjS5j8o7vvLQG
fuMq5hBhW2Ad7xcCHaIDoWPFlPRJ+/OaanX0UOPs7NNEgfxAkbso8OHv4jOTRpoQOuiN0riIYG+4
hZ7A0Z6ufnayekTXLM5h7p8g4zN/kXMYYuqz/HFzNKGVUmJORI4mgTfWNl1TP73wmSUYCmcpfXBv
c6jHKA45Td2tHYFb9lyNzVWV/IV4ex75pSaOTtXzyrZVExydOOmfZasFRnM4B/WRLyR75hm8zblX
NDZcCAmoRTU+eWZhX2Ot0dKyiqr2wAkImrpM8Xdk9ouUcOvvTYixvZ2o/7rlenTcNIR1hAt3J6j4
9BMRbVZHXHMHpKEavpBEA1j5H2QAQtZ2II8s6RaNJVcXFFg6Jdigy8J/wNiATQUblVl7ZMawde+3
BPQLrAwENvvr1kKT538ySCeGoLNQtz9xFjgJ4Kr1GQh/jXZi3YEgmqtzBLyPrjgq5gFmvWy/AeCI
2Q8uh54wD4d+pMnzYs3Q/YYRiUFXwicvQenO3m5mPEyC0IxAkIhWF1s+p1L5YfNZPuFuZ/fdCj9h
bf750H9J3EQyAM5jbjN2InF59nscSv9qtXdNfDdG6+nbgQa0kMPeiaI3eVTW5Zy1BldIpC6MluPB
tbBVm5Q/D695JyOgJS9hguMH5OajVqS6BbAUZh8xwFOoK6wcKoYU0mG6Yy6U76061hggXZ4IqpnC
HSbA5peGfRbHn3K8xY7Sj2Z5PexMHEBOxYIQWGn+m8v+xCkBbtz2JS/LOAwSxFct3Tiq8u3lbXof
aiSMaTlNiYGbAvNHYknIcujaAB0P48/5mcI0Ni1t43Qs2E6h6f0xD1GXh8lmZApRqRCPEiETyLCG
ZSK0wMygiRIACcdwZJLBp+qjcD2CILaPRJ2voCyBI8FhhvvORsq8QYvuQdn+2RuOvX+zAR/tNqf+
aBpMhVbMp6BIWM8PEZigrIyD9ifhs1dq3AljlCdsvgI2l+8sBS6vvxy26/Tj8kd2iznckZEXN66c
95+4rQlSbmzLoiy/3gGRW0nSgIee5aHSzE8CM4RsVOoZpeZdKpRZyo6ogfljLO/v9hLvVLfS2sIw
yc0VVK2BTFqL7K0q3Uzbvsdc0as9NJJ2Kq96XTujfXLY/Edzbak6kG/A15ev9NnoY2B+ynJpzwEJ
oubQLtCKGaU+A7IqhM23WsfazbuO/dqAVXbIM+FD9xqSG/cgwBWvvA0mD6WEot0OdEyoX66Akxjp
TTiX9d9qiBju7qmdUsmN7eflmOZnBJylbgNnvle159LgJlFVZBqaQwSA7VfEFpBgCkOnf7XLUYtP
m6Xyg96Q3OFh9bP7xt8PZtTskNL9WSH6oIBaJFsDnH1c2gQgYkBXinkiHKp17NCxnt8AS7qDpnZc
JvD7MCgC9m4zZV92u4D4OIHN2Au5nlpuG1lpKIiBFzvYdFeCN97sTlx+yriBoZ7o/C53nrpKlCKi
Rx9IPBZspIPkxu3ThMerYQAfS1gIShohKjIm+Of28kQL046He17AiQKSJSW4ZfRFr6fVii28HmAf
1ggOkyj33y5wa0O5n1RZbqGPs7pnbdS96gXpGrL4qs4QnvnOZ3shrn19oMgKjMe757fHpgfMTaD+
kBZsICOTEfN7FLqs+ffi9pQC1pIQgywToPBkkftbarfOIWzRfHTHWygJ7eqMSIOBDRfUAG+Frkc0
2yu2bErjFicWIXBDG3iTcqMy92+sMNHNEu72HO+aWX254/RrBv1ewf9pyQYXizbhHC4phshj3sO2
bsH0+4ec1ArUMCW4DGgxPuX4boguU7USHXH/tZrq9M8Cu+sXHsUK3tRgfzLPeBxhDoIEOziKmlSZ
ddPE6npOk8P4Et92tZ3FI4GQW6qyYl0r/FcKf3oQL5qHUPHhhCTE6mB6n5HAgU9febGPJLcpm06J
qHiAbnx5aF2l9nfKmyxh9Nj+8GV5tNhidZZfEHwFK1f6/9hWaysGmNXqhA5mdnfwhSoXM08vsdRf
AyBp6WGmU/eVCda3F8YUC1WKDO6fSdDRLOWPWNFQwrcuipRdX8/goqmcRltTtTkGS4C2yc985ms0
+x/MkdyGd1hR3ZQjRHUDj6Dv5PEnH7TQLR3ZBZDIzvRu+I6/EXcMfBdp7UMTrZLY4H4uLnrtEjtS
WpNdk3K10x+jBV2VNgq/+UVfoNWLNQZLDddM4p4g493fjWE/KjAD2TL8I/PIte46MkAaAiNJyaTZ
OHzDKrITTkIG5Y/F2JhtEUxzwAJsx2sauNbaRPOQoK/6/TSxFsbt90NwHIFnPpSmAx3Awo2e/kOu
5Q0VtJuOHJflxAWqqadRIE/0c2wWkkE2tbuZAuIywGKzvEmcSd/dIGTfKzwosag2/m/6NDLVwgkb
iCDXpin5J1TXAkLYk3fnAc64GGtEoUTRFrCfNJMi8+eYWovRX4fXFpOCC6WW5RNGBebuYdE9Nxfs
20ydSjCziDC01WEn3fYwB2uXkv8E9JcwmV2x4CKfDwW09Cana9vE1g5ZkhyFIqGXyqdmZauKKZMp
D4Ne9z6PTe3OE5/802jsTYl1p/S/DsnDTVAD32NxdSpYE5YHlH/+JJe/2/za+ITKlxCrO0JUY2s+
dXRDvgjJ2Kz6YTDpjXS14sK5okTmOL6loUpGRiZDaDZewGJykCOHQycI9JbQJCHNIrwX/epmX6pO
wMRXmOyx8TuFcwgzhCZDfNSfzoxtRBlbdgQwkuAru6+v8i/wCSDWTz+qAZYhGU74XxPCEZd5/XQz
Z0brrxyRe0h99HZ9GCh+tUV/xp1PtQrqY3cmXBoK245/PQRYFN/Hqrap2SEcL5r3UGqaCnaZCwY7
mEVAeWyIP2f7DhtY/UZCnxrTIs4jc2QuPKfqV0Bt8uw8LUenampih+7bDIa6KryQ15595MyS+pxE
MAHG/SZWiyshILoqrFysWMzJqGXl+Or9zJPZ3lmMmJoJQOTbNyz94POz+S+g1/LyF3c2UqC1aN6d
YQl0mA5eGT6ktCAIF1//3crCCYdtAmZS+SjzxhmBJ7it9EO+hiPOHJhhm+H0l3/uOABLHAcF8wq6
/lDM6Jbe/DOKdEgO9bP1P3DP0mky50klzp63Vd1/lSH+QTTQiG9BFxgJUq1eMay8VTGQU4hm2akF
kTmzfkNFGkqAGjZt8fgVpXApny7WOjMCPZvegrHVkpaEXr6QwBRjSaqBuDj2orZ3UEEMfjzrNVCp
84Qcq9xFe3eG0JuhQZ6KaTNJ1MA6NZZ4oFAedyACE3myO3DVd9xOtZ+7eX9GdSvwhq97l9iNYdvM
/oWF+2tmFL7ESMRAWypDFY6gf0JwyYROnrAXqEg5fEUPPE+XZzNJ6fU/fFRIuHiP/jxPfOBUrc3U
d3Qx1xotKeHEzJg0OJ9iREnm/P7OnueOoom0uxfBTwVagQ4TySjRWF+l9QvqkOHq1jegJ2VVOfYx
Uwc7ydsmXZ5PLOZ8CoOjXLy18Il7HurSG+OBqU8LNW4FenqcGGG3we0N6d8h2PrNwiM526Qv8pcx
zNWWwLxe8a6gIiu14nJN7DayA8TW0bQ4Wrvq70xO7pYzPisUj6T8nSbt9ak8Cjq3BogV8XPSsh2+
nSm+6A4VlvT0s3zUL+bfhNGpywju183Lnksx78j6Ekcaj9LCdwmxmbl4wNquZcekF+x7Tybf5z9+
Ss3oPCaExA33W1Zkgx8IGagCAZWtK//hrttymLl19OiqZtQMSObF2EAE+uJIZ55nBK7wjiRyL1sU
4Bkt2BWMQt+MrJbhe+kgT4Vf7nqNl7OhB/IK7301zCFF0GXrgJcDgII/kA11RhsHKsS68D4IUTFy
RDJNXbfJW3lSztI9AFnH8BxlBfKY4Xu7jikm9NqRuR8xpuNOOWnCCxxSejO94YHF5inh12+PmQkT
2AnPsGETAkHc8p8nJUb/FMaYDrzF6ccVzrurvTZCPiPVryb6jFyU7h16eq3km+NwpiC/FnV2HzKC
iXqSu7gnZxpyWyhOMyriudaV0uC7HeOXOdWwoyXVnRbf+rXwqOYqeSKMEv9QsiFVkk/VEsY4D+bl
IA8Hf9UeiHz6D55AEj/c/Z9crmLvPhuz6c/y1RlQYsezivvxcH2Vu78AY5W/PVKgU2NWsNfzdUVh
23b3I7ZF23ScsrMsK6ykwsBYpujGZvHq+LQdvbBUmzfcEAX83J3uDX1gSVdYFDGUhneWgQwpa40p
yPyF0W4nQ4wk5KlLvT1kU4gjWuW0dM13dOteqXTE+fvXWX2V2M08Zachy/R0W8yKvWowuZjVA3YS
3l04Swz6qCWZtmjN71aoeqZXc0DnCktloew0h1M19db+7krRQCFyTpcKSwEjVOKC8VoOt5BM+ebW
mvxL9tGuWoXDVyb4v3LG+cVo3ChzuWMvyXRoBQZ9y5hc5LDrIc3nprtjVHbUsaH7zp9LzW1JCcbu
YePlhOSqengHqNy1wUbCZvNMQQJBXo/Yd0gpJPwLMqkeYRlw8zn8cfXP62ENOZMHRyuaW5bWRaiz
RUIqsoHC8OlaeBdgtJuK77ivLRW0NlDZz0gekBWsPXNDyZ+sUYWGs2KPP8GdCg+J+hOghxTfv0Gw
l7CwRTSKK6nFV6sPv3QWkthhQ/PtFQbA5DkDdRIZXHrFJJfAfCsEthFGAV1SHz8DyW0A8lfgT/bm
Eioa71mU0+NutubqkFNT0BM4G2CslJdh8pNZ3mzUg3Bp/kQF2wFsLo2tlB+IGTyHjQy364L9jR/c
BA3RtplUAQicXMppam8rrwGRB3CH7BhZnSaLKNooKfxtiDPMTP+oWFmqCTc0bPftw63SUnQjIJ56
WqED4ut1OqiWRb/TV2zZ1U3+LM1JBsyOnFlJQ6c0TC+RyJsOFKU5KPSzrdaPRfuS3h3F461mnDmk
V3AzWr9bb2BMnzDDllsj7I7KCKWcl15DL12eV4hVoWm6P6UoBpqsA5vUIYJqoQVwOGrnhcjA+euP
MAKG+ddNr0+GtZ+BmgB2S6ehMEU+jkP1tXb2ZJj9Q509WNjtfof2jMrPFDcw8R6SP29dMMZHpFmq
YqAkxu1dFkuJXwH77M+WBTz27Sl96g+wgSv23UxDZBrT3PW33phPovcP8qZ0c896Zpni7aSqwScr
4PleFWEpDDFYhPumKzbZg0SU70/vql3Yne4IE2CkvRpZ8lGhbrvcd3lz7A0Vwdzw5ipwfVSoNRv4
0T+uZ6qJ7VkchyEtM1K2KR+K2GSa4jUbg2MuBY2PSR5SAM6CL+P5GI1mGJUf4KC3K8QGLlQHsVOO
J+yfl3eWs7wqCMQf0jzq/qpGhbs7k0wqEMtQqlRMJUrIZD5PjQGRnG087OG6/srZMq7QJrRXHM6z
9+gKNsDmGEQ6I2fOEMGojJtCo3z04I4LpzM+ZmGP3ZrkAyHWOH1ptLMF+2FfKWrfVcfUQAdtb1+X
GxUaAjtW3+jUvI03EHWISZn2qO183E4CBbDDPUEhzZn4RG0hpTaQkm4ueXqUUImrty40JuT/Gsha
VW2+hAx2fAbQ2jJPN5hF4/dAvC2b7Z/DK15JomlPiKGuf9MSHLUukYRatWx4E1MSN0maV4Ifa1V6
lBtMgznj0lPDwCB+IvsSrchKvhX9BN8WYALfWq4uk+PxoskfBNJU2/Ggfew0Ik7vjibGh7SWO2B9
vCArolHpqRNM+6kGfmyQ6pN0gqkEZS4R/O61w+ZKVgoDlaHQCd69kBnlePhdrRiA1wi39mB47sMe
e9PPXbJK8T/zMO52bWDdwdL2Ro95sq84Q/qu3pj14DwsE2yrNiqH65IBxB2q1iAwiR9jgTiOl2gr
ieLoFEnkItqi+21H2NznLIhpOSJYurJxvFrk5av2kZKFz2zPgVJ6UDYTExa8pDSU5Aicy/zIEwcc
m6WMJpTwOXFRKrc60jZ70dcZjCefS29SnBrIiPKjwJNPrNqafRuNqhB9b97S3QJYRZBPfEYIayvo
2osT+vyIiOanTVtGt9/iyGRezjp15mqZrkKYWv+gaCMzpUp+5Uy04I5VJXxY0CqHZt7Rv+WKg8bt
irF4rp6DEdJJrXNLZ6U/djK68erpBXKJptc5FlmY87N6Hxo09R9v0/YPBW7e/Sa9TurT0bFlazqL
Fn3P/ZT57ERGhHrd99t12dzLM2TmCF8zpClL2FmbFX9jZ1kRNhSe9lcTFhWRwukdPKUlQZ7Mme3e
oR3BSy666PRTK27FgOVolh3fgmHlT9JcAslDzpFVfvbHkcyHbbw7c7KiTG0238T7i2TDQuVGf7e0
7TBw8NIyLgDyg85Vr0sX5xSj0OmxrlyvwAcJN07lm/HSAU7U/cDWR5ggpJ9y3mIr/LqIGVYuyHWH
ZZMcfXDTl7NBLX0dnIk1rfIC3eu59KBkdGbk3nePZNdGFIDot6zAA2G41M+BPlm9uP8wqbaYDSBm
HCIHZyy2BYaYk5imxCtp1ecItgrKQlgqrZtTrlHbG1XXC+A56rne9PwLTEF3FRqdohZRaFP6GTyk
FhRbOBgN01/IJbYJ4iLgUssLgBbu6D1d+UP8yd5Z9HjPp4zkpHqu+wv5BX3RObM7qF324uVmf0d0
su1psenSUln67h7+6zjZ8S41xtqJBuNdn8dEz9tFzLE9YR09sEVuYGe25uQbh4/LImmcEJfNz6B0
jqTZKqOuKk7TImTDhebxS/IFx73a9oTtuiXZ+5FzimttF1rN1+b453SGG12CD3Wi5Ur9DluiMdQS
ZUH7o66Ky14XD93kR/E4cMAA/G4YJ0tIePkQSJmaxr23IAotMLEnq4hZz5UCA6X1O2LMUByFPUAP
DjIl3nIUhu9PrcwwWAvpFekLO6BRsosaTyQgzedO+ou+bSDMp0D+RHn+XuOL/MW/BTvHsO5wiscp
6GzGVqbkeYWYfSkxBAmdLBzqxD4KnA81XV1q++d9aV9Ia6GynIfvl66WsNJNqro05ECx9n50FJ7g
xSj4rt9s+QPQdSS2AQ09G1by6Y3csvnG+xucscw9UZCA6oboFdEOu+BSedlLoe0m7zcqbbHmHesw
q1w40JqJvs9QRU/kgnAqODNtHIhsVjzGw02hLb+pa8kuzgdDk+6J5uyXxtmGkLl7VdNhFGpOrKAg
qmG0BqxB8r6T4aG8aN8VCME36TpEmfGS9vr5Y2e7cvSS5uHyOwKaB4kIE8pIpRj87PaZu8muPBRW
TUyOb1Ej5vgqMZVyEOWkQb34XrKptDj8YveHamVFSAX0FMC0xk/3pDSUF7o9/COjvJq377sH1mrA
ZCPTemWusOGmBmkS6l3hmkd0HoQLdfLiSEER3T+51YIEIVvP6PXZhEsQhlT3oGSds15aDsbbmh0n
8JDRd3/ra7//agWA1Rr6KfybfYt7WP4UWo/uEI2+q1wRli97UT8YdJciAw1+vuz7kSa6sDF9Za6f
HBH0lhmHRm8u/m1PcLBdna9vK9QwOCRqVhri6pkGri2+XWdLgeSfL9Mmn94VSw4ypqFftzRzHbaP
SDGItwX0FTYvLborzc0MCWFPwth3sZywkW0q44tr2zxfu/zHfF+0O9ypuY9UiPeYr/jtGvwxTQ9s
1KG3DDEDEdgo+CAFEckurizQU+ZJulgiyRN/pN7yKESeKB0ic/9C1C0jZnOxj1MMc6vs1ZEx0pEg
KDKT/1josgHn8GWWOC3En8qaetxkG/VWb4xgSg/JCpjxhEF73T3QJZ+cPF1pubuQ+GCAJzebnLpT
hwIqNKoiLaOClcj329xjdNiR010ZoI9/BeA/p9i6G4AVx8banb1/+KyCb1CgvDGTnzb5CRM/bvYW
PQEZty+29Skcu+ETMRekY3R4Y0LQDNhyTHjqlwQPkVC1Glw0Hr8YgOBc15EJxTwL2jKRpEDpl/3a
F+ErlyptdFSZh9T+6DCaL7SPWiloF305X5wWAVKQ0o1UDhjZV9nbX/ZLbxYUEJ4z91fDjJ5yevSG
fsdxrGX2d6/UYr4jxgo69Tx0Ua8bdOcD3FaK/TjEgm1mjX+7RV0MwVvVXM+ps4RqwY3cU55AEwyS
f5AF0eCbKfHnPsbLK97WvJwWnTzoHLAW13nKziLt8VcYGEnzLwLIXwJm/p+t+49X9qbpqvH12jb1
iEtolx2xNDjtdtXGtaF5cSm9VLkq+OL6eOtaUHc0WBcjryCxYenZ9Etohuk/gErqKc+nVgr3zXE2
YmkISu3NIKz54Mv8Bb0RmqQWghKZNNrcAV4E/72ZNJZVmE//w6uQGKEIdj8hDc5hByckwvi205/H
l3IBPdn/fXHjhEelJsR8iFOGbM+WXqEg8pJkRWVc2UnUtay48OScjJmwo1ozsMYlzhrKbuH/S8u8
MVjnLvikXwNsT2xEohEEWPr0JkTdeqxHEweedmxhhUOlejsi7819ZqLdrXjKy2iHTZYl65n464Np
iWu0a+elKQgRRvsyrEhE0AubmYPUk+skx6kXi/pFrSL4JC/1bi0MOJCdI6lhjZRTYgQfT+tAeqag
xCkdB8QXTSDvoASiU3AC+RXHDvmKHE+bZwS7sJBW0BXePGwo3blJu54YK1LBFYnRsNCmbABfx3cB
NHNQmgCJWRhb+Qe6pUPk5bEuxzL+PPRg0l9eEWqhr3wL33y3xuAj2PQOaXdT6OBRMVN8TNpdgfnd
9HIWA0e4t+zqawisa4uLyiJuzWCTaZyVVNkoAg5ClrXelJDltZZ3BC4oB6jZ3yCqSLGZxW3BJ/G3
iMdTAT/lnhse0hdrouWF4HJynDLKNRTtUVv7Tyc5vAbPZgcPvW4/iLOn6bfkusJg6Ha8dYpFmJnW
otxnkwV3vyNmPjmOuBi5ti7tyPe4J6lc/FvGwhZuuCeZx8Y8nO4YLgu4hwJ9VS0aVZpOmya/PZFg
cpEbcY/H5grIZal5nvCPFGUzuWkEXWzG2YxgsKd2sspdpA00vM2k4gmn2p1N1Vb3fdBjfIya8RIT
uUt+nULWuaMa/2Fuu1BGwbqtHhR2eUUWJsHSWEgGVpU6wSRqjwxIFcUTHs2OBgSm4VWw6lF5Z1eW
OCA/IiUxHBohWwMQbUXEGFLtVbKSsbBiw9wXSJKfonssbSN+8Onl7UlwzNVMCglhw7eOBitzMyAW
mbPMfq70p9OiOaLeuPDBdXoTEvHDLxsYKh/sxYKfI1qrFSnbtiH/cR0VbebcvKMI4Ah2V/sQllo+
O+7dFGoeHhxwJOprfnxAIDaGEbXvm76Ak5kYGMWbFgtILVAV67/Rrb8cr30y7XOIKxWNvGbPJevh
w9jAl9EDYwXw2Wys5Hjo03sVq3BM52Mx44z2ydSlncwy7u8Op0k1UVaVb1SExWO0/PnCYQw750pe
0vMGyzz+vcDWrY5uO+5+EhvLaLxcf51D1tFhFp5JVJ2h+qk6vy8DkrWI1oAPaDFBABI+3D4rIFtM
YJ8n7OX7cJikv976O/wbFqzzqlHPP7QHXsJ06jiWZ+SLLBIKTrFu1NaG4QktNeZcm5xxXFDjKVDA
2eKDOhx7vUQt8PoDpuKIHTQzhFhTHsU4KzQBMO+pygltj7Cf2GjQmqFrl4rp8QyNok9vL+DPRZ6Z
whuf3xXABswzRhJivNxy13jTUF05XqhbqDBJYeUMBkPyElasqd1iCOUYk4H/hvupoA7BhFwXu/gF
FzSlifWNmKKcOqjQDMICiC8ISFz7F1jG8+CpW5dJ5eo7sj5yw00T+A+LCfXk/jrxWKOXYwF1wzo5
uV3wJm7LVUITTM+BtigxOOChcLebk4HyLjWMFbZPqKhqw/0rA3e4mJa3ZGgsz1kw+dECbYxNKCfX
4e02+C7fVI4egDH253tin6XGgjVDhIFaYltjlkpQ4H7ISObwra/qo8fEqAzrCMaqKjQbHWzAeNe9
fPhbqGCcHvpxNyxo71M3bmPKnebkXyLIaq4vVcm7yC70Qx70TNMcqn25DyIALwyPKQuSz8N9StOU
ky1S54546en0tU/7R5EXsYTgz6Z/qQV90g3MdozJfQQLJh1aBX4Z9T7OCJdv6MOT3g0q9AfhG0oJ
Fyb0O6nzk/m607qF2T/N8xUqpTbZuveT9ibnIICN8+2Cu+Q+G/QdrzcLBmDpaqnwViGSpf08q4os
QzDIycIKrvgNr4nO+I4VrR/kWX2PBZbaKA0JLrwNaTXA4PQw4ovL4TaKSEGsXHpXenstCE3YYpZd
/4hIEoZUs3lzqBwMeV5+OmudMsd1FI5XVUERfaB/kn1Eku41S9JtEV8aOxBDXoGZPlO2D3JsDwQU
CxgBe2QJg61MNlUO2nByxq5FzXmwe+5kuZ7SrGmozUsXxMaVFYtSA+r5UjPO0TnLU+8RlsWnW2um
x5pPcMlQIQlTEk1w4eufkShHjRG+lXFRznTstov9qmA2mox6H1IUS/3tmtENpLvqII1thCweNtB5
u2Cu3KpzvTsVCsNMJkg2wzrT/gMbde/d90UCrQ4kegDUPXIYodqUouvL8H2hXraLFOUKutmUS7Fi
tIpWq7w1ReRVtDwl7zj57N6xUSvn5HoAdIvdlv6y5tQgw/yM65NtDJ3UWe+yjPdZhDtBRPq7weSv
E9/pitSOzvmgJ869p16KN1vJEooKpOQ0c5X5YtrR/Wf095qu0C8xBskIXer+TVOH7CeHlluluuFK
1StKUxVRCaSCBjJxt+EJxd8hfVtPyisbf/plKJAGSz9x9m2g/drsIOY4QZkYIT6FskUR50tf5MSX
9bnsySr38j1muO7TC/dSIG7NftlL7GJEPpOs7eErsDQsGgPts0zppezs40wbUo6f8uUkq2wM+4+O
m75hCvUz2P+QyUTQLbSTsFKWIU+WahSTJ+eNAr1dgDLIItHSXnsKfgN1phAZSRithc/jnA4mw3Wu
+58RdSMA62NomokmV7Zm41A4w4UwMDGwFp0P3uAcNOxs9lEBS5mM1C7yJopI5G/vOwZ6nhAEjKmp
OzyBYQxuE21LM+d7TCRulGUzPeQSvDmDkRbHqm7SSpL45iDChhCdlSb5FQv1ST3/2qRWGdcNjEq5
oYiI/4Sf/8z4oRcwaQvWJWxvIr5UUn2SO7CNmmGRrC7iw0Ield6x+4STpnPeYz4yTL4SReue102Z
S4wcmq3IZJCGwiWHy5hyTlqOm2LBJbqtKl63ukYhzbKS93qRkrncTQWHabYGLPyGdFsGl5rIXBsh
nbbq6MI0u32BGd1Lyc7J2VjeQRf+BSp4AuMBzdNUp548MwJ9mLHiVDQddwmiRqU1nJtjeCjD1gNV
WlpwZPWqepKPoflsRWWwWUW2/oLXplQ2htcdJ4jRHyNlvK0cLcothdMwUrMne2dpx0k5HPhxbhDc
WbEW8o/NzgDPsEMUCoY8DkOfAaYV2kQ+DdQds5CQz3s9+hnNo8z89uTLmm+8zCb3IFtyKm8KFgeE
9XhSOaoI6RxfMK3BC2jfnFcooZ4wwUjyKt1UgMF3eoCkST6mHN6vvq/2zUiUPEXu95LqoxffrWFM
XewMLcndn237aPqv9pid7N2TKxy+4z0NBbgAESJvh7r6W/sAMIli60zjQoq7wNHfVp0h2qeMaG1A
KqojGOb38vl8KJyNEUqL0a+PW+S18oj3AazWHvQV5gA/v7jwsQRavR9eH0sn/Powv0XuXiCS0w+g
hfjmnQKJUX8obobvvl4wk7laoRKlJkOOJvNZRtl2FmwsPGPHB6CUYq9PSkIBZ3HTthUu0+fxOn7H
1DAwABsuDc87X5DF5W4+b2xPNp8L/xbzUYjILa60o7LtAH9MMbLoL5yNtgnD3m5NMBzXw4LNEbjj
FnHgnCW8YuUL3hNnuAFUtaTG7OK/1GwxTeh0ScCSy9VXjVfC41Yvy91CHxaU2t7Dw7X3K/ZBfqQb
XFwcrE2yDBi9emcZHi2apuoZqZ8xHz7gOILkjSbsaeeYt80lVSC8tW/l1aBwO6J5sBKGnCEaSZMB
PP+zagCiAwOX3aYts6zkWBqwJ7bRTwR/eOi0Q9alJYNMQ2Re313R99NN063cvvx3h7pKjqscnWxA
Xi83bbcrJL++2tgm3pkn99MZBJsqOTcJkJyfQa389A9WGU5ccqQ12Ph+rj0TSTbBSN0A6ZFkfsGp
Rs7lUG0BC/rxHmPXOqyHPGCgaXfykQEpfgYA3f4LoljBXsbGQ4ecrLhn7smyVpxBzl+XAbyv+KW+
rKozRzKJJl73uukuLo/nmB7kMrWOLayO1j7K9pWlvJatiZwFyVQSorYpDho0miZrU5gs4AGZe528
+/vHSiWOw/0peIswvUWcCXszgjMcp7wjupyqMMqW+rlTOaECDkaPshdv1IxEKNhnK/nZic003L4U
rcjT3OGJJmYHpJ2VnTO3paZvZWTEhWh4cxmgeNCSDhJAwF4U26VQZe8/I4zP/B5oR9qMFK4Ag0mG
idfODjhzthYzWCLWg6JoE/ItdcP+xkuSm5Q/WpAf5oSAASmpaRq8QQ+rMEKDvQYRKH+7fMOaD9eI
N6Wtp+tb9nWiSJhm6upqyM0EQQc/ieFbfPIq3tewupx5S1yRYJQH9Emgipew1l0lO/M9nfp5PPPk
cp/8lltYvpCZsr/0Mq4xbfIurzi4Rri4Vs3iJyK32lIdfqZA6MfQ6kbg7+D7xyUb5mOkycUYDRKD
BtBWAQfAPJxgjXQBgXM6rvyGVZuFD2hcQiP4bOS+Hh2pL1eucPl0qBK01rgUtn45NAyQygzkesVc
4LS7FJ2AR+FyH7XGCrXIA3FqigAQdmNXZrAIUerPETtEfZTLncnx7oSgIl4T2iYk6RL+WNf4Sawu
KIO+wI42oEpP+V2E5RsRiDG6NT0jGr1Jil8K1k8UoOH+AWgY7rf64poEtpDo65fKzycmSwWRHfD4
f3mYddfBuW2jo9p7t5L1MRh1Xtg5kW4XLWesYrjSIqi8/0jQPLOzZUHHXV0UnTXenYTnwpT/C5WP
JLU7P8mrJcu9NKPS/+RWMkq8FsRN8h1QrCMtshDDnQJARuqEwkbwY89cMOxN9Jj1nB8Idurmwg+h
2KfaAaMvs3lLYF5Y0LxI0b1Cdm6cO7vsns3H6rHjokXYZCuxgKcgjE5GmHhG/++lKuwUudoYKf2R
cftRLpQscbEFOh4jPWfZ34pxuRVpjtE8wfKNXVVn+1NVZApVb4A6WU6rXjRvPY0aSIJeacwoNjj2
sS4zm3nf2lrWHiSo+tJ6evK5nRFbsesD8Eyi+mV7LO/YdOyGbPVisrw4Lf9585Ul4uC+RegMlKJc
hWyetZcxCewcekZrVtacwCTrTzBBNVztFMSeGK3RGohLW8G8TEeE3ml2kMRaaoB3uJIyXYWDBnbK
aNsxUEUxboNPf/PgP4Gje5dH4cs/KpKRtEx5P3eZQaMeie/KFuau/Qcu+x+ySqqHR9A3nzuSCwk8
Ud8gPE+Sk/WQ+hMSWsr0qVqTHdFW1B+uQ0SeVxfyGy9Axt38Gdubo5wuyek8ocKc3aid/7UD/AJQ
oi9DqBEG7RxpBLW3CD1u2jo+n+YyGGkZZZdZOvCulwBX5jfbyhBt6QXA1yFSUT0CmNE1XSA1eWrp
U3VnOwGPdiM0VYOZ1UncZihGBNRpSpDCuSIgxUoimnSYJvNrmVe98R3Bgj4c+Ruygg6HbOpQ05zd
9rdTs5k6+NdiMswrFQsB3PRVFBHZDzc6VTzl4+9ywUUunaEdowHfAhEkQ2oUj5Lj3BW+938OuxB6
6N1PXBf2ZbpWZvwn1TEOhavf3R6/RBEkkcLPMA+Ik5Imc55/gesPzqNJoWlHJSDub3YRyMCg10Ma
vt55WuoXwN4yGNRUVPvymWbJTjdH0BJoQMx8pKOR+l0jShBY24/Wub/TMrM7gziqsOjizBr/1axV
zSZqmtRIuy+Ttx1pUhl3acuz5Wc5f7Sux3CX1thxNcWf+V6I8H9Cy+zlYdiUp6HD1FewjXVzRAzP
lHodBzCeAny7Q5kFgztTGEFH7DPRV2hajOQMO9y/k/n0xMo94SJubdVvvGIQ+ijr4Y7MX0UCtWIl
FgibjYSyAVW0Zg5fm/JT4kQkK7JOweHGJCSyJpGqKjYHA9RA0Dj5JSXbaXJ9mDO1gMjMIQNskuNo
l2fzFkGaDKZOjqHzX1hBMBH6Nn1Bx5nYP7OYalgF1XzBjDmjFYAoGBeJfWbjzdEXs1mtMB4h20R2
OhIYBt9tjPsFhsXZedEx434I0SUT+Xy0+u8ZOsCaMu6tYTIPJI6LLSz58y08dwY0gN5xvXKXUD/+
+e2IMjv1AApo6DfOcbNgj3EqtyRNsrUOpOcn4slnGQduvi/8HmgRDGA8FXjT3xHnuPNcrOxMDEEs
ll24DajxAJuO47ThJvEmUbf1oJ8bglU/Tcm+jGZfVXtuolVHHPtptkz94HTVCZbHB4/mNcXONgUx
lWAUv7f5YJL549cEBdw1x+GKNitDshsX2wxslcwMHRx8S6mw0I9UXAuodRi7dgsG6zo9S8v94X3s
PWNombd6J3BDmO3GGQGVP40JWn8mDFND1vutvJ/KlfOLrem1VcJWItMY7FfdD4w8yiXt1Uo4DpJg
nIE3DmnZpEEIFZmrDyyEsqnrceA1GiNutuugmAonWN/9741At9SacCnHInqFe0JRyC7FgIxe2awf
BRPLeaiObIcURybfJrHxI5w6Yh+BoXP5xvFi5VwX/QGPsL3e0yTRFPLVc2fmH/122TibmqqvGojw
b4XOy61DGf9Sh7IrzasBUKXiyVSTlXeQfqAwATdHbhaX/pbuxBTf8RnRKXekFI/HTSElmscWHUVV
Uq0lam3CfZaq2iQlgZ2cbmZA4m2rM0X2uRyiFRynB4cVUo/I80HvARZsfdyzFw76VrMTTr2WW+zc
yztEGXpYpvXF8iGSfHH7cpF317hHkEmMk6c4GSi5U6uAxwOoUy+aTLidCOGtDaYTQBI76L0Di7/s
xe9FeuLxvyrP/tcFt0cQSok2taPZPR8WvjFzF5uV4+R91/lbjK7qoN1z+Jz4cV5lx5sgSL3k8FEO
EqCGVz9uXa6zitChhDk5VZKIrjxDo1uLTijqlrWNI9/AzWmkN9zopDgXrSywwO7H6zA9+QUiHJer
GWhPbPrv2k5vbTgpwFSCQtSMUOv9RZjSCfaPUMmkrzLmsZ/EjGzwtaABSCxbfhVC6OFWgyVVbtx0
hfzI/XN1abA7svgn0UMlfxzVg1Tmt5GePeHLfNZopEOhXvyaPmGWyBiUM0ugvXgMY0xXR2QHAltn
bCCjQKvAscpTXobQSdoGD1NI5lIjxfOJmwYCgvnYyGB5iGohaNUzVcLaTOSeikewBf2ZUwmKe+6i
tv6DZcYCJFEqbFFQsKDwjnpRlTgCzvx6771RiXut97ejdlnvmPwUt93Bm2aTFXoUHWblNBKJpF71
5pmdcG5JeGZFLeUFgmwcpA5Z6IY/f7UxhBym5TC+oOpVbVld3lyZh2CWY9HfCi+F/ZqxqALauok2
6nitSXpVFfZMzXKYo3YwxH9yDV5pSB9UqGttIti9s9Fm6ypt+1+dODbxp82u6IF0B+EqkCztJ3Xw
zDJIfd3HxP9x4WxD1H4GeSPe35Xxo11ND+Zwd4jNkkQTuQQFMQhZZa1SydH+l8cyV9KLYKYuu3w6
8L0UU1DLb2Iz9FBE07jn/EN+zb0D5ev+8lEgC0/RvU3K8Frik3CWCmSMP+WVRcepV5laBBqiN+vx
7bm4joqDci5YwfPjag09DPtoLKUn470RCpJumqbfhrcDMo992pZpm8DRGnMufVw8E/48cKWIaHtv
PvmwuSEPtIZ2oj44Hu89eMS6Av7z4hHrijOtqe9/Dq4M5gKbRZfFPjxXFWfZ1Uonw48YYbjL+ZJw
a0u5hChZoo2V4fnAR1Fhgqzk7qTM3mlvWk1BDoSwY4Xt2D/y2gI2+3N9PPr4Bnqof8Mv4h6A0owD
O3pmR29+HKTdAd67Zae4qkHZGyCdwHmhR0d1AdyKunf1QydojJflyL74N82tly7LGLruFR1XujCs
whR+v5qhYA1+ItmxDFX59gwd+Lv08487nSAZCCM+hb/9ruC6cMVZ0B1le+ogbid+u1a5sagZpQqr
GPOIZfC4HfkVVmFnWhqHrqGbwFch8VlYsoKe4YM5J3QSiwctSh1j3wL6S2OGL4Qk/VOpFQkv5J35
FR8XDv+WIvcQaJBmLrcou7tdSSZ8g9k7Jq5HNpEUqhmfmbpneZ38BLhQmqnCToMQPCRoZ/rZTzdk
v4kU1iSmhMdyZaWi/HB4M6cv4es1p3mA0kfapBgUb2ecjw71PPntfRTivtxMCThE5uOhtd774lnh
LgRoOYxIsNYhBJ1e+fWCH/GZum7T3f63coXpNMFyAfg6Q/jPW1L1fM9xjYX2zVZ90orj2wLrC8sF
9QzXpNjnxKXTI8tD1/TrPrFBQq4tNgX9JN/l86u4m8USoNTvpJLb1Krg7d3Dig/pXYFPzZPvjTMd
vA80zIsb/M8TJTJiHskRXGrq9+4rupUhz+/tqp8JxaWP6Y16mZdkg2Tuqp2y2a/jR3BmQZEelZcy
fadSLb4vsrBditD8RNOMUCtgFO0EF2Vi+Vf+Gjmm+t9u9kwjx8PZs3GZvJnSbWSRYuGNpZ+XeFPU
r22k4kh2/GHH1wyIQZMOHR1i0xxN3g7bexmCT3nfv6vlwN5RKprMARuruXXCmIiEKEEg7OgY7zlc
qc3K0CfBs8IlL6u+aSkxT8tNYL0OrilT2J7mBy1VaU6s1Cx0OOArKwCgrFc288dP2K+dOtxRsplg
k1cNBX/M4H60+BYS3jdvMmcMkM0W3M72/PzKy9x23wwDF+sTzzH6mGEuzJrtJmpc7Y3FDzSLwdI1
wt2GyzgP3INzZYAKuIEV9xN+32RF9rP7uqDIiuK99f9RDzNZGKWuYWcGrYsGPOsWjox3RPgU6dc6
VHFRKU8MJLl38/NFFJ6izYnIRhVqLzqBpbXHOL/nfBtNM68uLLvzsJb8BU7jaZfzsRX26oIDeY/X
0m3DclHKsbPxEnAE22dK7Cft2zQj+oQvJjvBvqZ+AT96HDULCOHwoAYymlBcKvnBuFZOGEPvIjLy
ZZ7Gv57spmZ2X4DGqiSZU7aGKsGbf8S1EHvzzOaqCRizSL2aG56YbrToU89VsYLzNOXwtcqdSdaT
bJg/xtx/Ii5ARrYGNBxHAN1KFejhALS0a28/DRiMS5LjHiv9MUG0rk4m+3n7+FXWQAR4bEaesspp
C0GGL22PmKp2qXABbcIGl8RYzG/vSGpBncpHW5k3JEUML1UMQ/9klcUVFWy+L1ZhNu50QAPEZxcT
e5BFdmtgFdOiM8KI/UNU0VrFSTkjSMrqrBTSecHOTyLPGmkue2HSdl2d/ERWqepLVQnad8kfhh87
PY4kZzuTFve9u9BWrBO4EhcyGivEdJ1ereZsZ6sjrNcCZF60lD4VsJaY6/cfacLSmKlYsjo+y3M0
U19wkTvQjITHA+C30Vn7xWjC2gEwgKk1+3TLx/7R2SVdfpv8OYMMxQynoRHTYzEak7QOL8Lunhyz
t+hExT2NRKO/FVh6DVN0dbgP3MIbdtdZqerWoqeo/JfXLA+hVEAjZfw4xds2er7Gpk80ppFhlCFx
sXyj4FmaeL1FA3veKINme6UWAGqUKjiE0gf8xwtoxSmy5CynNacY5eIUzm0Y8PQ9Pet8pXDs2cyt
47MbkhNlN5uhm+iXn/cvxj7hKOC4HdII2k50QhqGJ/PUXDOWDnw0eU1wTGLltcpSQyPJSw6/MM1v
EmBsCK7ge8IfmAJ2h1hTFWgnIqJvvttpox/rgsUscrViWoboAyZVVJ54NTZtI9lda2Z2qYJd1ZtA
FoOcg3G3m1dLjTs8HSIOcJZpC1yhPFvohR1tYKafPRpJlt9hpPzOdT7THeur9o8UjflxY159Q+kO
ukkcKJCpn+hNe4wUkK5eTX87jT0tawwl14UT6S45R4PKsi5xttfBRxtqlmFLT/Kt4051hM3DnlBL
wxuYicLvH+r91wiTYAi1Hi/Ygzokw7H8JFKulkZBVr90VoGBgFxSg7og4+g0gFif+7QtdadKfovO
bo3BtHN7Smgwrsj4rqBm3SzWAsz7S1jjFf5BM9AgB+X6Ejs/CozP2b4v09MZegzgcXIYOXnjunmN
jPirw35g/3cj7RR4bv8gjrMWkyX7W2OuRI3NuS/kUGxuaISTrZtuJP91kLmYDSjQqz6ezr5uAQgR
HSQHBnhF/dIhliwmJBqnVbKAE5O3wk1oDy9ZFQp6sI/Jpzaf8uaW7L/Ia17BFa6LJZzZnKdWQQD9
VKpbDBqpaz0BBfNgZTXRjkwr38n3FVnV/kVIq1OHH3JLI0uw5OSRLhVY3kFFZBTZeRxA67rd7Mkv
DBJeEUF018pUZNyOlTSSNpK3EAI43nH5zb/fekXl3JAi6pa5iDYg/8ddWatdXLQSAw2KQOCSRuXQ
89LF79KG2/wXtZT/EK++VQEMw6wHc8Q8GTbfkHY9Pv5R7q/f+EvBw8R8zgmjOntvQxf8xsMJ/i3J
p9HgF8pGLsmH+UM21qUlOoiKTCatwOKggMZbgipfgXvO/sO17OaUIDQmNXyf4/mODubLTvi8uV36
P+sPuxBf//w8EsimhBJqGjOzkpo7M/tTY2O+Kwu69kGS39lSJ63EEmomFKd6Y1Gv6JuA4uMgZC+O
MyaY7t/01yRcaCQyn8yEnOgOG65gmMtNhdk+aEOSAXwM2fjqtycbeTq9B2LBjNvRHeLYAZlktgQx
xSxQXvFaQXqr72iq+2VtLWAl6BagxlMuPDOBYbkNOb8SiIOdV3B7POIO33YIl8i4HtgH76iukzY+
TqL51MqNd27Lcxle13LXGqQ0DfzPH1VWZD7eKRKtC3gRZQOqembYceE2BlZ0zeFQH7hqC8+KsEi7
mS5RSSmRJg102aZE68DppNVoME5Ouw1xKejeudTJYy6rUmbw3uij5RopBD7hVo6jOSl6gk4Q1hl1
NBAjQPy45ykt6JI643ASYtqJ7pnU3jTbd53PVxjILbvpytHmp23NuVZYnSL7NFVJ8xX4R/9tbGlI
XQNQCWyjxIx6wFjsItCsZofXRga2gAe3xwjkihdf37PGID/WgC4qyyWbpBVnCe0TpJWTk/ymJblg
FMCmFtSTf1hP5i0wO3tvHC3cynPS8GoaqHZ3PlKggDYbR0D1gtqyItFpZNuujicKDaMwRhQJf2zS
JAXRoJiHSXykpD6x5z2gVSX+y6qYPU3WCubPLoAOAZ+6JwDRxwbVba84mE2ZWyMxxBC2NK6MTTmS
BTrO50/3viZczAc0hm7gD9Phc0yXeajR1/u40nq6pEiigyxGdfUwWwJ4kUg6IWPOJbPx0RtA2p6L
f4W0uV3gJULcYEh5bfRu3ZBLa1m3g11cQ/070Psk+Q42bMPX9T86HA7RinKkxEohjakTpyqRh5Jk
BJEcMP3BQFZ8jCrZaeUEWRmJXG2FGDIuFGU0HorYuQBRCKUHIu1T6bS1DspKyOPMryi5LqD2W+7k
yZjPyAMIPZk1/VYH09xCPFALz2gm4bJwpW3sPwjWOhfwcHhRtkBcfsdzN0HO5RH2/lGIKRsA+yUA
FV8SsO3Lsb+zhHxX6W9eSZ391XsHIoM58vqUi3smU1PgQY3Lz8c7z3/inCrr9Jz+d2t1+AOjKoCV
lOWW4Mm3mU9kGp3/tIt422exj2+h5MGZuOAEEc5p5wQovHipQo/nQ31znXC6mWJcbSk3ITEo2SoJ
PnYjBGQyJAFx0G5FgOaLqrZfmPmWCvns0CNoxWVnj1Za7yhnYe34LRPzuWZAwWpSzi0oaY+cMti1
RelpyoOpiMmTud9RSlPju+EvIut4nSoeLKFR9t7ikIo9bTrUTw0phxF03JpyQ6+6CUeGRLWZrB/5
I5oKhlTdh1RuQlEhXtpH0De5A1pidRxnI4E5OhWrFF3iBMff7BMuDB8zVbk3SyCDOxAjQyr9USkQ
xCu7G3dImgWnYmOTQYcE/I1IiPovLrXArsODEgyofTgb0l4+6M958Q9c3CzQtwXaBtR0zZ4SW+2y
lz6cQDhZhqJScU7Lb4Zx6/3yYiDrNUt+j2wc0HdfgkYfNnJTPu5zNP1kZnY3Aom/y4acoQylgH3o
wevXTP4dedK7Au3x7dsn0tyP7AeANtVWO8s+b/OBmZXuF1K88sWEm08qmR/gxMULxgyssTQR9E+b
ENCAQLFTIKxa3JceCq8DykwTt87IteLSRESVrZSLJ2t3c1jV/rBOZbpkB3f0EH99ZIDK02gw/Tu7
6EDJiJIROYC/snRj4h2r7u257J4PvIm9Jgwnn7Ls/wEwG7Fc2wn3VqLocGcCfppjvKrTXFeBYfAG
pZS3KslPC41sQIxevpuDVNjFaMB5F6+XmL2rTzWsvtfpewiH9jPMW4SYNnj03YPEnx5l8OUgAtuw
hR1kIn6zTl+u/Iy9AIV+aRg/mpWz+PJ8HQws679ZilWxPDlbvbFT6OBvC2QkRcFyVtDshYYl5sZJ
DgZdLDQmjx79+zfCWu9zLwHRYIkBkmlHL67y3fKVFVrq940jArsSh3dz1Tj7kosj8rMZpRJ7fLNV
PbkreMVplG7M1AFOOwPmXutLY45Q0MfewW4aNiVTF9izKE2MaIvB6P/iu18R399ffPul/jHjpipA
zDcKbu+CvNTQ+lP0208Altt9CkP9GWtRBdsBSp1ssvhcIMEE0slCITDWvm5Qn5hnHboVsfo8RoAr
Ro2Hy6HdCiZp3lC6RejNifBgMiX3LUHAQXXIXwOgRhjE4sfVs0aq0z59GaTuidg+Hi3guSn/U53Y
LeFmHGNaxWEj0l5kBjymREfz1ojWMNEPEnES++/paA5VhKIPPNFzt5MMlFgN9DRkdpC4Yqddb9Kk
ggsYQmnaIMDdhDQ/SOOektyZBG4gVZWKfmV8MbGr/NKX0wmrKLR54jWllu9LT5PPpBUtOFe1fpna
gdqq/Av8qZfWRepf5U8EIvBEErg8znOy9pOKzc2hyqwXWiXlJWVAa9AQQGyyEq11I05Y0c5b1pLS
jg8G9JeDqkGFpoaH4WVA7eZuMvWvpNLT21MZsf5voHMZd04zhvs5EZWRZmozCEnZqTE5I/BDKRLW
OIhb/QLxymGV/pyiJnFt4o+BxbMBtR9xwA8xmtun0ZUo7pllANF4xC1YMDYfUWiWegNo1+sW7oFk
aaazc9P6WuvBwbRkW+siYShodiX+djGXFaxA/tlaYG2rEa47zVwMabVUSpj9cRcOsGxEpjuXydCo
Vc6jOf+abg8G5HaVmtS7hYmQE6DAdnwQzuI2u+lozQ0clbfAEXWcx/gC+/NtDCAQyxXh3Kb2VIz1
kAb/5n/9yoJPGpZg6CYXzcaBo6gk31G3w3qyqp+wEPzp2WsvXyH52J89Kl7/qcpMJQ3i4g/8tf5p
H3Ecwk7CHPmj8uMu65U0aokj6CwEcv0YgosrCdmsKFei3F5gP3U2HIL+kn+fxp9627WfW8sUGD3M
shM8XwnlvQdDVJn5GxWv2lcn0G+jQtb2tQ2khCVR1+sQ7KVCDlfpn4ifDy9kVkoNyi0UElPjDACD
TaK7lb148+NPKRUdL0XSNN7LKuYttD3p+MCKWzTkqxhfeMgGhQyNqGG3min+7DGOf3csn1E/A4Mu
CNN3/7N4YKjpr1Gdrxg54WzPDrXlizc0Yv3i9t5zagTAXXd7ftaTr14MP5lMxALMQsj3KU3zDDx8
sj0Ao3f6Nb8wHp07yrLSXCxw8MTsZH9GiwcZ7HB3oJT0D/9JrdKQSJLMVlcOqG483F8KH5AkPBrg
geYbEJmkmZtV8cxMPTMZXX6T9lRMxDvwQNkYwrDIYugWs2rnQLWlvMuImDPr4yK9Kvs+IlF1VPxr
sahKllo3WZytKcrZy5UFMbODXRtb020KTIHAs6VYB3qmohZbKFXD86rPxQ6g63Wx552BimfYdTrt
wUtdGVXpCLy1/+I+Vo3gXd0OzrYcctCZD2gDYrxfOftePdJAwgibtoBi9T423ZYr3t3tGBgsUGZl
3C8MdIHDbMGTlmArwRUy1nGDTof8Njb6iIkyV85/oXM7vV9MnCkKmYgNkhZd8925kCaBBFunUd/5
E+Imsp47GoFyba9VkuiWNFa3ovd/owxVmf6zgQz+pA5IJaapCH+pEx1TvUXeK2p40eOQYBZjuNHg
gTbSG5BwM03IjmNp2GGOulRtc1IdUDVKNv/04fiai6tzgc0Hc6QXq4s5Fm5q3EozQgr3kaPlDY7l
OXS0mkXT9fyIfsrOou1cqmFpzGwDzUiAHL6jU/YmObww3I12eCIqO5E380PmILfkILlHMf3d2+bA
uedYC8DIgUlqZVtX4+jAarW3vRde3s/3oVWG/XWS5A93sN2O8m/a56rtsm37p7GHX+Hw9Qdq+GRQ
t5IbIMjZKrBk1RmbuvGEdT8Ap1dlO9m3D1Ktm4lau/gIM297Ihx7RWPFlQSikIheo3SQ6WVrSAPS
PGUOViLUNnGchpkIptRQaSzVh3FgNxapood8iUDA3HoKvaIg/++MshvyXCUj58px4+4YdRpqjClZ
0CjvrF1b/EriiIuN26B3/xsdDw2/yJOHKBshuxDGRKYt2PhitHW3QdMgw8ePckFW2n+SOfWBLQkZ
qKocvvR4CkRyvPsOzAKyG3TRKkwd73ucRYc2tvaOigyhJyYPsFMYv8kkqQeBigakjsv1weYibv1D
MyoSdUb5pX7g2gf9OJmKipcL8kY1uxuHOpiW22v3LQCyNnUugF/8s5vjW7QUioTeojAb0BAIRcfy
VClTnHD4z1DtU/OeqWYWTMFRV+9CNxGd84ZO+bxrb9w/5tZI2eVa85ZfKSjEiyzbvXFrJNrd3l/t
udI7517oBQ5FPB6ZESdXcVl4gZ2BTfi9CKBWPhPzkAfo439YDFn6VWrDyvdpNuDqJ1GeoYRXB7ow
vF2b3l6qqzEU1wb03TT6dDuGi+1EV7OuYLPl6dz++qJHRGdmyei/t5t5aegfsBbaMQgaf6KN0Zyg
9LdN1k5CnQhWAhGXunCtF7db39987h/yO7xXiAegaID5mXNe1npbMofgQPPIZ/uZ4N21B4KhRDQF
2n/G/PE+HhJYWIE6h7W87lIyq/FCwYiaiIaR32KzNPrmDxPtncaXpcv+7F3o0XL6Gnxbk84wxx9Q
Lcf1XKj1m4CcB0xtNH/q9mVUNF+l5TdM8+xdHDtD9eL3NBcaTdw7OmD/cjQO3OAHEsxGZ3sRzrMn
dK2gdA5XxdJqvgAXowb9ezu2HEtITJIGJ1VSLmnAf6QTKF3uTJaO1fH9SkxZGncu9BD7Kgqfr73B
O3RBwfC2X+MMwvCXHOvcKHSdG65GbWnCJdIfQoRgksgyUerBZ4kYJeQih5TDFdfSqtK5mHV8bFTu
J6aqBpKVLcrF59DV6UnZXwtEoRoqBFyOGEwt5BvwZqF/gBgM0Wu4eR4sbo8EQcFiRIwtVBMzeSiR
tTweDaW1T0PNRKMi+z+ORos+2pmVLhMkZ78jBtSa6bJMdRQI7ybogqqbJm4I4VQWspXbnlkKuO/+
vncryyrGADKwpdJ4w+aghp5dEhtrAZY7hTWTcczQsr8qAqft/9CedMVGhj1yJr6ksFP2zDW/vpAm
xtP/cANbzr6fbvDp2kHY4qiM9mlRE1IK5W8w0UkTfKiWjvbZoRt7TEpS+nNtI2dq/bMNn6H/W0U4
QJt2QyJ2gClyb1/cKXV48kzcMg50B972hFK8FKDBXtPUD7jWPaALCCEqMVFyBHv/iCkkHXint/a1
dxby7SeUkIxhk8nr+FMDJkyqLJnBGTf29LZ+Vb4PTLG2QDHLLbxze3kbOsosuCt9dkSflhp4WpJw
aQ0uy9XVEOIQi6SvNEukweFJXOQY2lYw9yeem5FyV2H/feWbG1vSOWwWyMNz0fhsUOVchuk+olly
Y8lkKcEnK5AFZAf3FeQR7nhqL6qMM7qDOrxNJ6ekKESIJnKgGZQmeNz1mBMn1oFszbeQR5nOkvQI
2+B5sAKtdXX6OrEoIldYFEV+oXjD0zksfaJejRmeOB87KIa+Bsay9k4917L1dSCD7/7SiEIMO6ft
9aAVDOk7DvypO59j5NTFauVV9LbrZ73FiTtpjc6SXeizpOdCzV0HQgAI0umBW2+vmRnFbKkcCI6X
mwBC4jdEvrrFGbpDYexA2WF7PgIVKlikCiJBsgxfAydNJzZXscgRz+y6FxhD5dxm7zWppqTmhkO0
1wasSD28B9dypRUP9viQgCI/LZ1ls1kO2Q47y/o6Rd/VUQksYSPdBF23lOfeWGUK75QWmsm/b+en
zxF8zCgE6zcY55HdtyheqC8v8oZgJHkbmgshUx0ZGdpn6ra9Nv5zu0c3qfcRlU9wevY4LzgmUkTF
tf0nHb/SbKRLNcCbDmd48JMvp7O3mLni0GIUD2QF15CvNsPsdMtxzGr1+WceWAIqhR+vh/b8EP1g
7OR7uH6kiYBOtUowe1ISnW69mWgVWOlfygU7KVhYIRb3jMJt9Db3b/Eor4EmaX5lfqiQJqTHQHax
q2CaJUkzI5+d7Wezd3WTO6cKZoy+KoWhlIB/oA2Og4XXLc/BPQTpwQNKLn8sj23PM+UeK3D1eByd
fVV7dyxCMQQ7WDH+k6lK7kiL5jGsExhoG1KsmJrEBZO6BG5nBR95AspcFE/VryECYX90BloXlcco
iTA2GvriiZZuwhWOcyb5ZV1toWDd+3nFvfG+x2RRGub+S4PMH27MbGCIayF3e73MV5P6SKVtTL0Z
IBH3Hs6nzBei9vfxCoXjUuaYbl1omTVsiJXi3LwhVSBbjA7GeByOnMdOFKYTa7JeDtBdA2RRvUAx
Y74vXj+TsWJQOIGiupMVOruEqDRLGghJ1SKCO4YDcJmprDqaTVIznf1msKJxrWARU5Ouo1lRpgCU
07J9UPSWINQj2Iavj9J80MUe7rz11CHecVV3D/N0gPmZiLOdOnwaMZb1L1zApLKyQy4YTAnnJY7h
uRWEESoTM2zwp8+YNu5f7iomtmAyKT7IHWgshR44+RWXy5wlr35fsKvS6VV3yzY5oFa3q0k9IboO
R0GXDveRMiazHnwWIlhJ7ZaMsRCa6Q33oNM4mynxZJr64I/xgKxovSBK0jMNx1UX5g2SFn5Kqo1m
c6T1cse06/woAMPaP+0mZf0H8r2nAVGttSdrxXhyBj20NJ6vctZXtAZdiwPlHO9OcILScwtgraUs
HKfSVC3EcOwPPUYkZYPMfH77AoW68WPwpxqvn29liQobhnoCj7a4Tj8cqbANC384vxySRmZIScog
853+jkVe3+5B6IIDPuCzue17osQy5mR1uYd1XElJUw3wj0JT+rTpbUHLIlEAYwjpkpHLrm+i1qM5
UJH6h0thhBthdpbpXMNohszQ6tudzOF0utLc2vrpxZzdDNwuC+Ad5u3zzeX9Sx38GyOSY0+DLYMW
5XDzoOwEQiMS35If0SD9ZBXMTQo+aVZpir92h5x/AJtimB+/2iHgxuRGz5tlPCvlVFtTlLTeQTm1
3WSzLlx8hYCROUCqdH3OdlVvxe9pU/9181bKeB3ezgMpw8P7R6XXyzZz3SY0qrPhW0VTVTSE8p69
ERS1vw4gUoEpscPxQG1QrFtE+Jn8rAZjFX+ZbVpBRefWB685X7O6XB9RI88WArq+BxfTW+F8v6aX
u5xip5ww3OWGyHfef04uDbtaOptpkUKmey62005woat2CIUomE+LynFvLM5SXzANJiNWPxt+laxH
i5jedvUca8ApdjJ64oEMiMO4iygyRtZKzBEXU0B/SPViqqEUG48EAlHVNtIa3tHFbRtYrtSF2OtX
jC29kSq42ug5AuwWQvgLhYg0ii7zWD2USot4XnV8/8tZ5CJlb1ca7CkBS7Wk95NS7FG1ondk7kYS
fpka+ABMq6Xwzp97xRKz+7KTR6b/hT/UqQt8tGhF6+GyIoiP6R/X53MEDEEmia8+wPes10oj6+bk
fSPQ5fW0P7xBnN6rr4zRs7pGWUDXI6kC8GC9ORDNbWb0ca2iuyCdCh7a9rinfKc9xXZJI6L4Zd3p
xjW2/r9mW4fP8WLX7qw8mVhqWf8Iv1A4PGODi8XTjqxw3DxZ6qSgTlmDh3q/e7h02HtrPpuRBiPf
CF9Ij3QdSBJpz98/9Mim88UMv9vb1vcnRE+GWQOmuJepsZ94lCzeZ4Z+2vsRj7ph+TtDZZDXoGNi
Bdf0V7KgCtLa1XJaQauDfn1eYV1/ITlu0jOehnU03dN90IfbBaR4TlIah42oiUFGURUAdiH51vuU
iCyzZUHkJSRRRwMRc0YhYCk4pqSpsGR6uegw8zvpJl0CcUX0qVSVx2rYSMeon2CudjdCY/Rd7SYr
Vfs1bijyWMCJv2w5NonkRSjmlnaUMrMW+RbbX/A64QLj5RBurRB8xaiuds2SuxOFgz1iTeytGpj5
h6Cjj6IXbQqCWqhxmqrovmcZZQOUXs0Hea7hJRcMB6BvBBQxi1vCTyJGEFnXlf5rEKan7ILsWcEe
679vbGYu7M1OmEvccX7Z6KhekGYNrDMj/ndmZeNB33saqudE4gKpYzwPsy6NasCUsPqC418K0tYY
RxYtYhCd8r8u8pyF9AV6m40dGSqSj5mbBf53CXEhTEoWzgI2aa8i1iQJsN4NX3hs6GsPs7RroYbQ
Mil1DwNk4v1mssgAd5ZTaM8v7mrHtIhtGx1IyrwdVNMjlx3IxbShzHWz6Un/xAf1sHx2g+2yDPM0
ctKABw7T/NlNOxtmAY4SJNRWthPKvdBb2CPCc1Jy/PyY9D2yQnllPCURHZ7t7Ft65MiPhHVB8Bv7
M+qQN/gPfiJc9wk/RVKP3U4Cu4mXdxbDf+0dF1HvF5MjTIOYfHysR2aaGQK4BU2aT/Ck4LCVcXZS
O16uw5/+rMG/Hk3pws8y3tJ6IyG60Yp/bRLCxrFZfOxtg7bifZm64W6p79Zrs5GVJh8IzKRG1zql
uw7adqlC7gKRx379Ekc/rwV9UEL+v7plZZzR8U1oennz1f1ebzTMprbTWDeX90gfe9hC6cRq8tUB
2ZwuwT+meEk1MesViER1ctb+0OPp1HFeAOhUiMcmlmD8tF3qFUtQr8jhjll2L1AtF2y7HNsp5TaC
EkAGatPKn5x+R0+Nu8KZZhRCPWoedV++99BEepWFKbmMBL3Wd2+aG+M8bYVPWjgxChHKYS3VSMbN
Vb5JbIQOsOBA8xVVoLdujim/zkZrVYbTLNhaEjJUHiLxMdajvp6u793Srpw6zsB4V0GPLA0B+7qD
zj/rWQ8RpUi5F0wFoLSnpGA9SoeGvoWuPXSXQuJ5GMFHoBlvYDibOaHF+rfvbSvXdENrwntUwvua
LvZChcCqs9h2u1lTnPypUE2Tg9L9IXenHbSuaikeEGPJQsM3TR+/xJsVddA22/wQBD9AULg96Ohd
yhC/bpHzqngM+dOMDScVXuE+37upUx7PSpIv7gOqw00uJQEyiCURBLPTFXcr4Lfj/WhJp7+k6cTW
6n/URj2KDl16GZAVpX4drnWy7Rgp2OvWlLqHtx1r804M60brXd7LCPupP3hCQODgM1OiIkzvEE/E
2cV7cX4ykrg2wtJrw8hsma4A1lA05F4K9xArZGx1XjuADc3HOc1bf7kHL/GtnHiPKa91CoNpf711
9HjurbOOsKEjaI5X6hb8Ha4GIE4XRT9DxgoWms4tjlGgM19B/f9k2syMMcv8gRlC96DnksJAWxbL
S3ZrmZ6Zh0ZzZtYlnAEYhTRXWCniclYCGILFFesR1zKR7G4BwtbJmwLl1Xhf0tCC66Aqua3uGNtV
L6LP6tGvH8L3oAmezioNYd8r903jZ0rtrtOAHqKjuYZORwUl5olndFpK2C4lCk6v0/i9xmMabOPD
TDLcMftNQbfwHwDQ9W+NXnSSoc+nHy78ixc3mnvMOnEZn83BCfqTTj78oXmgfItFJWTShagM4dO8
cYcgnn20IEoAdRG7kg4hr6p1JGX6w3X44OXKqSqtmP36iut5LxA36vxCO8SdcY5A/xhw9vC7dd0O
+OgVBinJc6EsgqMESNtSb4xXC/oRUxkg8k7QQLvG8sPRyu/ADY+XGku+ns6hmS0WPEwCRNOX33Oi
dNv83AHsEhH7aUpX1eouzxTkyPX+JYF0Hm7tu82v46UX48cW8kJ7uNAdMvcmk9hPkssC1NSs6eTi
dCr0p/E1r+qFdXu8cUAj01TI5CRyuNwQ9gajL00FceVj8GKKeBHOKV4gL+8LCvzMvXU3VKKn0FnG
RyaGlUpV4ctBt+I8L5w5m3RJsGgeEDdJW3JmCOEW0yd2FTOZXrgIojk7BbcANyDNQVWuM7f6c+i0
sdLOTS31cOuZflpgYWBwVtG61js0oY3Uk361A9eNAtx+EnDOu9jtzpNRqbCYGQvvRGHXjU2oaFkb
tIU8Q9mNAGobZ5pAPGKBfTvu0Qo+XZ1wwMcRF5qxD94lJXYEgQ==
`pragma protect end_protected
