// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
WTIrlrlMeY/suesBfn+URJQRxBsASPZVC7pIaCfLip/51Vn34/p6Kf/VPn4GIGB1s0jFyLa3jasU
iK4Zcj1+sa7WzOjhZ9iBeJ3eNHgh1+8fwKhSC7Qh9AyjyBNgIe9VnzWkD1iMfTtfxy3wM/0iNSfG
6bQBf2+xdNjMtTxpcVYX3YpFPJtZdaRl52GR7TDsfRq/HFP3cUyDHK4+yjlS6lY/7psKBbA75PYL
6kNPnsPInPrriwy1/f5G166XwqZ26el7M7ktOjyC2yyAMDvsYdh04SMXUYP6FEiyPb0kwcV4Y2E/
YTSwl7L6DVjZUOpveSg7D24z+s+OKKw1W0gnMg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 35216)
jFuPy44xs7Lst4awtScIkqbB9sI7els4DAnOPaL1lDHQf8WGjZG1agCT1BxTN9bx3Og27mtU9GAB
Kr1NA3b8WHDkeLPfoPvD6RbFzKS3hZKSvHVGoU35Ydpo5QJ9IHW1pZ9uJq09N51YGi5s1pNQ9lb/
IfT+6jrLMjYyRch59ovXCO12LxbQ11PBRWL4G8K7dkAAq8Wp83aaTZtKtlg5pcad4/XO4C0uCrYj
ETPKT88E5NugFWx0dY2KaPKTRnZk56jPqOK+6UUO0bRRRD7cUXpLLpYj7/dp3oAlsI7z2KrQThES
3+07afwVcM0fkJKq+nUW9W12olQAQ0LbCvmOMOBPXRV0ta93LTO/KTCteiweSyerK7D4+w5Pl+/A
S+eUO4xmfFuYyyU3bcdqAClHhMZwvAXYzdzjhQZFqgnUk5up3Ti7YjlSz34cpFIkJiFe0OLHFQ4h
oeAydRqN4ncRO5LDPwQZpQNWmxMGE/zhjWIqUwUFjKOymKMrBUN5Zuqcdv/m12mJt1sQAp+MnEG6
2ESXqnreLmeZaOih7rabaXOP0SNUAUji2xCyfoxrn/kNuLbBuW0T1aXIH7XQQMqsazCP8wTDiwsV
hOB2AoYI57iu2zk7a6uzkvAAnLO3I8bTpb3seudps5ra18S3xNLS6uxBWBE8rYAhbo2YVI+AaC8F
ePJmZ0z+eZhM/AD9Yt1UIVPKz+xB/fHJcGNf3aJl8m7VAgO/hnMB1mwOCAbLGCPZJScVyMKjZH+f
frTH4SNBAGYxcaXCtgqyuJx/PGJAV/BEdfeHWbuBMzu0TGFEPy1Q4t0F08Zmi0h1+VCoYExDGo36
FoZJH8qjb3j918NFUkEUtfDzXyTXKW0eElUrEnv01LcJGJsW62Phs5+Oep51Kj7v0rOdHOCLjPDd
DKkk/sEbjyh5XbhBYiBqrHzepK8j0H3wRzPJWK8aYA2WJ+elZF3a2jobUTBMRJmJwVefQj7oGeAr
BNyQmGZBpJ7say8mo+6jWj/fzIa9cPsKp0ObEHcoU1YQyFlVpMDo1c6NekxbePqz6CBRAQyV7Tx0
aPp0+hw6s7+Auc0CbFZVjyeQB/8RuDkLb3XJb3YVCqytXxwW3zUUMDic91NG64fzq58yiznW00es
Wq5OGnnPtrGtWS/jw8n19RmAUI0+QNUAtPrWnSGmIXSIXVCG+Ow2YAX4NZs4GmVNjEF6fF0hqVh5
k7qZJf1RW9oOGgTeyy0kixW1dTioUqXWdz8gRzodfLleGJr7eWx0olReBE5+3zZVSon8hek8GTQ0
SSRP4WCPA6TWj4p7PnU+wrZBRVORQyHoWnlcTTWg4Y9NtQ1OifnG98OWg1itVZbNHmLd4DQYcqJh
/tSNhFW219iXzKg7XrQzaGsyGkpfWqk5kmI/zDr2odvQrj/iTTphrOho00TRZD9A/oH2glVwk15c
NiEeVrjpVLM2CYcaiHGxrAOPVH5s2nSwKhw+kKSk/Xrm+hBOsM0g1xxoR1oNFWqK4HFg/evOn+rb
v0uhKLgD7lhJiyzBcqvxiU1Vu7eXSLuDf+IlR4EW9pQOpADVO7ZJZC0JE+yfDtCaoKsMt4lqMAz7
whOmfaZagRbd6TOl717ED4bdlXU5VK+K3zet66upaqOpOBpU1YhaTDJiOOZw4z4D1bnVlhAk65mI
okc6iQMN2/8BBn6F45YYuui5a2iAiOa6FsDIUm2t0gZxY3/CwTVYWA4KIZW5+Ir8b3pPsj04xgH6
whIrrb9y/3qwXdWFCtn2rLRFxbTcJ1NRBGkEPFZANcejelBOjup/lPBkKrJm+9LjmMksHk6Pxo9Q
HGdp/ezAQKdC9k+qZgk3GybEG3SGHjizjUwVxnjMYxEPDEajrw0VcpIFASuhgsO1s/A61Candm/n
j/NMlAZN56ndGyiyhHald9RsxLl9rMgLITYaZ0FkJ0O+hQ52BmKG28J//gcjHCBYLEjDU1ArS+ak
eG91Ffb2kSIlPi1+Q9psWkz7Ei5X/zvYDTqWNFUDweKVuodtWV1sdjxTSdsMQ4kCacjIeIe9OhwO
WURD9YIM3Et5WKHDNIG/OBqeFw5JtzaWlmzigQUZb8Kgt5fB9QH7zg7dQl+bE2eB6GvEEGmOlrSO
SjEj33D68wY4GtDhRz3nhHjkLBS6PXSoxjFnwKZ6T84+yUYfr0EDQY1DSNUFG5QqBXa1r7ZLES+f
a/JiNTBOBvGnSeBtSCOKl43c22+09ghjSP6g997pl4iH/tY4aLEh85uI3uKHS7U6XIYw9Vr0ChtS
0gGCS/DKjePpDsZKLkQEfPouiX+vJIYEMk8iWR05JafIBwKW3/PaYQ6Qlrckz7HNi8eMHTKXMyzD
YMa5zaD/9EVQkOGTlrHIlw9zRNCpR4JkbVsVbysqEeIylrkoTCB7oxiZKGHrgVYiT3B0S0H0SheK
cKBmNszx/mN+zseWgTYIi94nT2OGW8gjVSd49AdcuFinecwvBE/lbvEh06DyLiw9WMOfJxwjT3yL
c0Zl/VZAfucS+83uCtLbtsKbqzsCSzqW2sgV0E6zvoabrDsFBwYKmDChLq2AX5I6ijdcHd5TkBB3
jsoXnxkJyhGXrPq55M761KPzEWQZqq7W1PJmpMjqcgsgCs7bVR1Z2Lg7BTrpPQq7YXPw3oidjE6C
57go5prRB2gFUhQpyKukOw/FkJxAZu8KWap0sf5ymZqaXwa8tiVBWEBEuF4mqVwZ1gDcNqcNjttI
+IlpU4eiUSl+ezNuMyyIl27npYHCtyPNm1jZUhjenqLE+mVTMUc8R4NHhP5RRvogSDUjr2kXKXOs
4fgnTRcIn9yplVjoTLlbu4ypFzxvNgHtg6+ung30/yCDil/TKpfupflzOmqpNidcNfpztxpXp8NW
LtVUPhnN0C+4HQjflDHfqTw6LHmkH9k6QNNTqV9dACWdEyrh/SpXC+7CKzaTh5YhMCpcvgGQW72H
izTX2xJV2sgoRaKstc3GuY/b0PxGd/73X4uBIe7VVk0cMGjFwr340VfMfOA50KsVJ9oBEw8uxAjA
N0TFGBWKhIhBaX89aMSL+8lqDRjx8+AsxU2eiJLFT19lNQSXs8nabkQT5ELt2iGcXWAShP/ju0LS
TuzEZA92OPm361Rnhf3grnMbZUxbZDwWhJSy3zV4RM/Is4eOYw/6QV3FBTyU580OGBm3y8nUJBTw
17yo5/DMzjqo9GlvvDOOX0p8pp9AfBs/1xSxFsQhZKWsEG/PZFlNXMATbRPxbkjlBBVTjIOyxtUJ
LkQ0tASJ1jpReYqgoSVDe5iug5Hi6mkcMryA352uS/HgSF9e2U6d3VpuvRjtaFCd8eUw3pJLCVFj
lmuGYQoLIbEPXP2W7wMjkfXcUSgVdQGgw8MENVDSm6KNUwUs4h655teRwPDSLgq0OKKht7xoaQ4M
CX9u09S7FIoZ5JH2y0PzmpVn8NskMe0cBbAUNkmj0Ncz1MCP+pcmWjuNoBAKNzD8WwEwPd7jB1fE
6TJ2ONzHniqCsE3+Y46NBwWevmjvj8Zsf5WeshzSQcBlsfGjADhrxdnpZbgRKeJEkn3WsF89aOWD
qDhk5XHKnr8I/ACq+2Et43uCj+2EfHdplM7TSfV4sv0AVrfLAANXSTheglnZ1mW14rePQUrn3Y9o
4p77pUiajpj5C1SV/KxhvEVAVdRfGkqkbuO/Edxsebqh+jOxFYNlk9SvypZL+2n70a0PYGc4YPDd
er4zZ1ujaEKo+iVxgro8puWLJhp2BU5LRIASCXzYNynbcIlTcDvJsWkhNJj1WBEtta3JxxFzh6+H
f4Wpw5lc2gZsi15ULa92CBFYtltoZaUxPazZ3Ks3jP7DDiD2o6nsx8Ydv1UNgRIGPxbCcyCmvrIb
hgdsYYivsVIn9HIGVhp/TqGo1JrHnRN1cOktRwz5v2Zxu/djh/S7WUiBHCYkJ6FbgUw9mJhGNiU7
PyCvDlgO6gbtSK/+Z1C7DpErRsk7fsba7XBQsCU0c0NTAes2R1Oi1fC4yHBvfBdlycUCU6RaWUrT
jGDy03jW96BjbL27du+xoKVVYYDBCaHaTp0V8YFuwCvKpTpVZv2KA3xYJEESOHQOuuh7CYLVXXAi
lUgP4qAIhjSuUC8n7vIn8cDi3N6b8N+4uFW6bVAasuo4x1GK7uUDVEO3nhljKg8dopNmXFEpv1mb
em3rzrMZuy5JPYyTgqEwgZvbXnWsInrw28mA+S9z5xW2CiM+aM+n9d8DFUGmaZkdp7Ng7cBY/yII
dCS0Erm6XFDPTV2iXsULvegP7CKjguaAfw+6hDNmBBOXXQ2Z5r8EYXbL/9NvFarKmXe8OmiT73S0
C/qkDI6vbEPgcZe7LvkGj28Rt3AONQOb0dtnjENFIt+R/8K5SYXl/ifV12oH7X6d28mjc6r3aDuF
7w9KKCrUqaaSOto8GhhmPd4U8fsYSR4hRa7MnyAbRIVqGtHa94NDtzhpXQxKhGvdU46wgevNo23Q
3ynVLecN30KiuB1T7pJ8mh4gNj0QYqtCxKqSkt7LKA4uCaN6lSRjNljKtMRBGNldZIJR02LTXiKF
sAwYmJtWFwzH4Se7x+Qa1nqLdi8WttniMKr/7UouE4GrFBziLRtEqqIExui1Qb2eLrymvxB0Wqsp
1C6l9z7b2LU76jhDrltkWNaGJV67SgVojJZ1R2XSKV8B/vb0waugeMSXCiMzFb9BjALhS/9lRir1
4RcqhHSRIqQmIKcD1U6Of7O2OajT+kxkJvD81EcgFaBohEzpR7nyK3ZMhnKTziaX8PbbQ4OSqSqB
ryqzJR0xUYmBLUyJIWvjpdDAmaYKc/ntvVChsc+Io5TCw5gfhZryYeyC9JU6NRMItv1YMlSHrAXN
QaqbntmfCGkRPb3GWAEMnXOciRAsEKHcgglyLcXc7QoDyccdktcsAPvcQuxllihArfEaGm58Nijf
FrX0kfP4yKOmJC7MQOcX9akTU7x75MqwKgxEw9+7qBTviLpG7RYQSgyeK9BJXLW0JcBCXmDn2987
X+5JhIhYXHYrXXVnnf/lWXEeO9zzzttRG+A5VylwQyuf/qnL0rZBxYs/IKLD5TpJ23wCYUqzkzEH
f88ilx9ODQndJitNGCkluCY49gRdZbmGwYHjvn8J5Ett+txM66DodT5UB6rruSrVPRyhjHcGrMLc
v4w9ak0QjIs79gNDjgn1IVU5Dzj7LEEvdXxRpjGy2lLnoehn2MlqfNUI9EscxKRpcPGyVKoXL9bw
8k1zEktAGJ9w5EwZrJoXOzxA0N72Vug9JWURDo3EamGMjQZ66HAG5fky38Ki4jdJosLoVVcjp6GU
TbYfO9YAueWsAQntTA0HjwvlasPhgD9HKpqa29fYRyvfvl7riWqzttAO0cu6ig9VMFnmfW2reL+u
p3pmvzoeAFMeST0EDkvvFoYWBaw7nQ8E9OTd6V9bn496TqK9zO27JeUwB3APLoOyGG4dFjTtIeOU
dkMDLWOG/q8jYNgj6ztKunZj3QbT4HK4dNFFJDs0HEzKR0REmif505MwgeMr27yJpUCqV9S8hNab
6DR27vDY7BXiDjqmZl6ElddyV7gj0Uw/26MrDF8GRcDBekWyQsRQDkodzPmhqq9FvLnjjcsm4CYM
QZZb5TqpPlIMEmSZkJdV/knN5Lk25wc09YoBc5DyCyWabN+0sAODQeBkqLqjsFr1zHRy2ndIFpQN
JSKwjk3XNvQrvq9B1W47eWp9bZ4uUSMeeYguqp3LbloFTFEpMh5gAATqqY1jp7pMrPYOWJmIFeNl
sd6DceqKP+zFqbQDqRGcD+yGOaZtgJyt48YZp1wl3/66JVeqAfKgFx5Ss8Yh0ZNZONOInLsuLbSu
UQft9rEO6Q9cRLSTCLl5fqnHh8IWGl6jn7T8urvhVVlhHkkp9FIr7mc7ROa7kBy0OVMgsatGzJKD
3P+sUG0KcaDUzbR37N7ZfiTS7CHD4DwabY16uy98t8EmDf4OAs08raxsc4/baTtHb4xCLSZoJOzs
PJzH3PB4WuvMDVk7k7tCgyuNhaXszmmFgqvc+u1VErJMJwmhegcmG+GaFbnB+veK2WEckfhQ9qjJ
4Hz7Q55T4LZ93Fdako2XiwgBbbxe/lshw3fnYnU1ZT7qfmEsX5A/oMFGy1mo2orV7v2N2kci42Ku
eTvXIkwW5GIjXAVgftCmnGZo7dByHCs6ecM4tlypSkS2kmRlekqLPY0MN6oS5pZXMnJNziKHMUWH
U7zke4nolTR1r5RmC0eyaHepKhvxnymPeLIOvCVVjBDI7fSW39VvW0jcC0/02FEHUJYIYE0d4RBh
iw7ToNZ81aFq2RzzyInnbajWEdTrgUdEp2hDUc0P413s6fpEpo+Nzs/VG2BCo+tzs1PVaVrMxffH
1uyqn61RR+7kRoHByVT1NOE9z3i/+frUI6YwHiiUoU4+UDzmcrqGl+kAvgi2skO6XZfjRDGoVoxW
0u0q4/opkHYFvhw91CrzcXXLlWR8kGspJyUDomu6AXMBNaRDTaM8DjydJVLBsNsq3pBNJ1q93Hw3
oisahl467zpTm9/5WAnMWiIftrIW0EAqj/XkleL3FNA17ztb/gTNJFd3CvQ2Z4qXtLoFS/jXzIRE
nXmpOw5iGHlqWuiZXYI8V8NZ0VW1wo9a6BRjBzX7qACDSIRqhW2HZGYADS8xb+uY3m5MvRP+v8zX
gSa7ZVs0WxUpxbQDb/YamxyDtNno9wYg3Gy6Tp9A8ZE9huglUzcZfe/3jLnFeSoUGATK3ERaIzy/
pkIso3PWn/YMmr/ClJ7MzH3CLOgLY2S22gg7wYQvb5OoZAFbM6B84dgmbtLG8fDCx6Imi0scv5Ra
cQFd/ThLxcbgb6SzcaFY4Gb8WJ9IhREw6xRh0ojpyPc5UDbZwKQ/mycp5E0LCXFnxmdHgz6NARvj
r80+GVo3GtFFXk0KH46wOI0epWmOinCFcWJByWr9BVEd4Q/7z0h6uXkQUgcCcZZ6MLDAF2wvSLni
56tGUddvA+eHQpkA9BXhuWQZkiHyfd6BQm1dR7AoIDp63C6IvYhcrx1Mb5CrYtGEJeDuB0yJ8zi9
kxC84Oa3KUOiQWBjJ7qh5RK4p7O5Fq/6uWrTmhzgrC0QbzfDHqKZ2e0UTNPQt7brDw4+9L9Yhqud
Vk/77KXxcHQ+lAM/NyAB3+blKJS3SvbC9X/VKpBPt88HQNsVAYleox5Vo6NP81Q6M8Ig03Myu8RY
BZU27Ur6Wmrpqrkm4g/9KzuzKd/L6DpJxVWFiKuiZtsJj5ruZs6L4zVQ+XyhTByUGZvL+oDIwAsH
N3gVQ7GB3zAVmw4m2Ux2MRX66y9UQvuhGf41bZBu1MKBVhYWmKRkcg6/ROSKPayGhiEbSZVPv5Ze
+X8qjKOO+Ud3BHhuh4VtwlbUPq0lo3+UuWJf0NSttF8/1frWDziFgmFWpIvIKzwO7XvMwfCK2QbM
XkQt7JEyWWh77l6CdfjvL0ua2/sAOIYyL19wPe8lV9SeMKZZT+HIs1mAHoCUcLU2ezw26Zm+JBci
9vOpudHMu3Avutju0fUa7jh7P/guAgs7so8HJp256jsGiMZNwkqFDZqnfMAVfuZSgYm8BTSjhaUz
GvPoERoA77mqZQIGIqjYugtztUD+qYtox1duVb+CQ6jlcXpMAiVie1fyaW+AjhuNfcBlmZdWnp8I
n5vAw6VKxhyjgW4moupSFqMnniad90Qo5GBctbysa5wR34LFjpXpKOvSHh6zoeBuHJygwQGQwJy0
Nq60/bg7hf+6SGHM33QMC1YjauuD8zObq1VOHWQ56wMxwNN17qvjACaxmCsBgzRPv+3hktgbFicb
i9G4DVudvJPsK/pfBIp++Y2eNq659XqK+Ck06RNy6NAYf/A0UgZMJqXp1AIuLDsyhleg0wRpK4tL
H/XNfUSRzR2NwYVuOfgw3C0Te9bnB4DPHFEAWGH/AUSgPS/B8KH+J3DMC+ITNhKWKycRrsqsIQNo
vIcqyYzWYOHeHpj/fEFWPaa9vxVjWNAzGOX3BIn/yHvu/qkRATQtXpt3HKBoZYWu9s168j1atOUA
05md1S8lZIEI9snCbm/NmOk/0y+uIIM3yMFdRc2/021QPQ8lSvRMQ+3GwAbkBZbToQ017p8t76Qq
R6rjefUahOd0DyxEzxJzi7CBiUYI2kCumIuyhJr4WYMW8PZO4XDxZFQwWtqI9ZDSXvps45KtKCIF
2yWZbzXnZVA16i+etSGvAPy1rWHL4+T2B4JYgSnAKcZpR8Q9ZEU6/MYX+j5iyPcYfYhgFb2MUwS7
5Ldg6e4IgTxPRNTiSuyuuVcP7WlZGTi/UxsHrb4UygCD0JWcvyXLelAe8LrOv+WWHOp5sVsiZN77
Uub+7oeBYaEcZYK72J8TW8Vif2Q4UcN7UUhPiHKvllxMndMRV7R5C7rJTM/58VBckEjmAw3JwIfN
p+l0D6np48woSAvkrB9+1n7htfxeBhORWovuLn/UqEQvUb8auQfJA1Du9twx9R2vlbrWmVBy1Pz8
67oQ7UZSIWNvIabjGzW2s0hJLH+BGM9EhlFUvfRW8wlRpZZ5QRDAVpDRawkzAURMlsnEWwh/Of3z
3naLSFZnwyKF5SDYHJjI7TG+fiVyKfoZxaViObV4T/M8veBJMpXb6UzCOlR4IjOqIIR7oi5/DEtT
//2wzUiUd5KySZp4ngHd1ngp+oFDWMm31iIIm/R/aQS54LxqNUp19iXB/P/LFCohtZVYNacJEUn5
/XYsIyfUcPwwTrp/v6quVWQ6Ca5eMm9FDVbt04lzu8PDJYKprvJ04ZeXVgiPfy/SAK79BLX3mJYq
n8srzuzCPmFn+UZe6WGPCeX+DIKjzqKQapWwmIWmeYj115EnP/ucTQq+KjxlHj4GkAUJNuhG+ynG
2PPNn7l0If5+IRLm8idKAVKIAiRS3YRSKMcGDQO8XS9RWwf5jCfAHb9ZWI7BkoNYdhdcMdFOAyBP
Rx9Qz3VTdtJ7NBEyrFaz8Pu80hMxssd8VJqV+xa/tgk7ZTSWF0GkBmGXldXpuQHaQv5BKql2+Yk4
36+eX1+BoUNTNpPmSS7KAyP0gR0oUg+RnLjoAfxOLe0v7Pvqfz2rkx+HI8QZM8s9stYwzAtPZC7+
AOfFaEFMnr5fr+JyqzeLgzu6fVG6gsJDrvqcGgZKKKlaCpjJ37nu3yw3h4dyhL+NvdlIh6qYPjyn
ScKeIT6ovjazOphJxmrmTSVrLnt6UgqoPw3iJBmXf5ZCjKzTJqbZjCV+5EXs+DMQ6tIl420y0Sfx
1znflWKMIZkP0+02dRoThF8p4sCLdRbDkMtl7DvmetdQzgIWEZQl2GO9HoH6OdmwpdRHiTLwB4an
HXLtwxcVxOnsQXo+kBbCEFvyFD81rQE8XlmJjWDQiZ8eV4AkubedaiHhDcDPh+s9JY+xW59qSD+i
8iM1CYf/vL8NubAdhdC8nxRpaYGirdBD+GBYwqY7rKKM+DvJ82rDlFiAPfijiftjxLtOjrT4utFW
0zBuBKDbMdQho7wu43GjyrY9zSy6sliLcopbylFj+50HOZ4CcgECLTLPpVj9sERkBLXXdMpvZQgq
ozF3xJKPAKrVdjW0pDaGg0a6rBXOzKKQGt4YZQVToX8hx/gCqAF6A6BX+eZq6+U+AP5BZyEa4a44
tchL6EziWo8jnyGE5ETFoIgzPwYoohQBuU7kMwIK+LqqGItt3wwdC0388boAWZEfiVPXhPV08IWs
sEue0aIQQmbExrD13b0FU4OLugRQyHYGAjZYwH532/tKpuyegpby4eyvmSV8ERFUBWjuWb3JdxpU
GkgWjXtqPFAAi5l3Ag9/WbWxivhyq/WpPRfYYxH4TxvJahUImtKSyZ2spTJ/oI7vk8/Xge34arnE
SbQNsOcfDpyITrf3/1GbkyR9VCFcPAb2nrFNY8K9qpC+xv15i+hB++ng7WrsSv43kHopKHoLyN2M
ZpYB5KjiTih/jCn2mfomyk+omsBDCFx9t++O2r3NEkJqrgp7qbSwm/gOU9stJv7Ff9tdCqRBiJnu
c7zApRBXRsWi1/ilfM1Xy9uHki8sodsfEVYitsdWJNGA1ZqfUNiiFpgimpsINA6hI8ECUS4+rkHo
xMnKqJAK5gIrf935GP6kg4xdYwukqGCy/NnaxJbgmTkcMrbCZtOEwZE2aj2+VTpqAJ7zSteqKhnf
vIAeI3LzRFpY8SjXHZdnq26O/XrKVbsq8skv8pKUOG6o4dsFH/glaGFMXdbzawevpvrFJiM+Euto
nenCShtKARcruLC7enT8WI1W6I8pH/s6cMWeDXUs59C0tTWriiWg7uF0t6KQo5eauZcb91TBVUxi
LwenTHVsqORpblkSKSNnq5Xk5PsG/pMU9iofPYpkEObfUn3FxCbbTSwc29t53G/NXDVCywUqVhAP
n9KGXPv2u6MRzna1KY6/eE5Ij8p8CjPfIaIyBrdsKf+pdqF4wn1GJ/t3s3pDQON6fLeiR7zwMCSX
7Yjjcve96mBm8gE/V7+oF+5LDSKGUDLS53z8wkOghwM5LT/IRGDZ73KzH79BI9JwnMrGJ/juyHvC
O/jLw22cIDUBvTVdwQIC6Ekx+K6/nI/l+wRHED9CflWKCFGlAs8l6BqjOpX1ACm08yrsu8bWY1Mg
Dzz0qgHcIseUJ+2/Y9SGXD81VPmRA8ulfth44wrzUNIFZv+VtMQotDVCXIZF62sdxAtzR8Pn57bR
aoRAEtRLxSs7OgxOBKt2+WF3m8ER3eeIPGCBORJqdSoM7BYIWUXs5aJzhn3i1TE73IcvTWY5u67d
Ds2Nm+a3PZIFd0OGiEQgpuANEtLLMQoTsbVOlzY9q2f2LUOolEm9CtAvu6HHNZlbbHTyKeF09WPW
Lrn0H3rsOMaC26CXdQyM32ABegOgQzqbUTJCkJuhI6Wmi/0oUDQNvBUubgxbxu+/c0VGeYoqFjll
yTVqz2VwKOvZl4zfApsa0hs5nY4fUuUpsf4wVNJZoZCTV+NOY6LHzfVWveaGsNXA4Q78WD5+Kboe
ne+JdFaGrROO8JWV033iRK39AKKvO54/CIXMR1MQS6KQBFJoVsUrDRug2mGqTLV5FOXR/zhnOODz
GgxrFKF8lL+d3g4Os2cRLzwgAzG8DcTslpA+PA6yqeOm1NJy0BZPLC4uR5HOBg+Rp3fmBwijusax
NDlNBJo3yy2czBidbE8cZGPxS4CGTQoCeVwhxQY329Pfcf1Sxe57sut72Q2qXwcq42VLr8DE3k5V
mEWFL9g0n96FFV+3A0PaIaUxX4yfgQBB5muk4zycjg82GoNld0Q08n/QzzVs68fhFti/plaYJWyO
NpzNQZtgDrhmXm5J+aonm1r0NukqX5uobHUXQNX0+j8QXx/TMh7iFGLKU20Rtmpr/YD/ehAefr0c
Agn6uWob3RO8EvhEgBU9dYnTDz7atMdM7Io05r7tBiZnanPn4z2ebVYdKDqIeClYqZlvnBhK+sL6
syxqXfuZckwwv4t0cQzpTlhU/9zrE83n7r6zg0WtbDFnMuYr8wDOBYdoi/JZz1PT8nmj1kkKM8CO
xbt2RVv4kZzVBmhm/Cl6hq/suaWTFLDtfGFegZ10tyqZqN/YyAV+UODUTLDFQWfkAPmsCLPTk79p
ZNdtkuWIhaKMiOOGf2c4roGAdAKboKCp5+hyoZphc+KlvAotWI37l9Nf5yVjqH+PpMQdkqm9SyOw
tIsJi+/r84A3BKreRlqIbO88cXEp0QqK6reJeproynn3eH+Pubx+C0tjSa5e9iG6uuGNuH8NMvEN
VMBtKPwtodYIhGFeFjOydLPA/xY9kJ3j5QQdpCS441lRTBDp/7/L+pUi6wwEJwMRsIY4SF1bGWMX
w9+0gDACZDpshP9jcnC+fdwVk2lzlL+GLUJr5t8oZNmb1vNd+I2T61q2nx+/3yHhgMGH7/fryEgx
91SzImbEQq66q4dODa3Khrl4AYE2zDJewGFDS4cpOtwNkdfiHI+UDm5nXMj9cR4oWKu5B/LKv8/+
Ck3OIWTxnF7Ghy4Ug9bzmPtGkmvGI8Yddbk9/H7Gl+wPW+Hk9t4GVCR8/r0rh6GPh/iDnQVr5bUn
7iQASFwvWQmKAZYf9oAViisnnsN/YTvCu7x7bYTilovXy/dgmdajzix7xlkIw1L1uncVkypKa8PS
1k7Os5eFuNbXLpsv1y4LVWHd4OM97wUmVyHOsIwx9w0Kf1Ntm5Ii3jRmdxjTckMMupZZLG34IhAy
2Y6vKc4qZy50eNlUFwItITkxa6Z3R1+EdJfoR9j8fGDFgCpi4XBsAPeDWI3/F+cMhdXjLXj6JDh/
6EzFUyLVWiZFJTp9ltwro6ne3wuqVSvBRpMDPccHjSLDDHSRDBK89rEFKHaYa6KuYZV8lj/RhhBU
xyaQL00IdTxkr+MAETYGAZLh4MaHSzNzsKcES1s5P/dSMI+CF766nKx08udQeo1YPuw9FJQv7cor
1BRKUXWjZbAh65i9yKU1KqfC9ews6LP5cdJuaUxOVL9xXTnjZwFRRN9pzK3wdlvC+cjLhaJ2T8DJ
Z8Lsri+YgqTupoCxrYHArlKe0Ycb+RN7U4O4sPjjV6tk2xDe/qIadcHuuCNZCnFP/4k6cnK9vXce
t8N2x/dMpjDhIpgIfni6fomnp/R6I3sXxcYqPRXiLg90x8uyidWSHCJau/z3v017SqJBdLnP95j9
7SPS1ZptzEqkolJvAkte5G034g48thzayJLIDOC1zbNCdx1QCsdHII4uFQksNIud0/AmjrpJeTlB
1LpBLtd224YjlyVAUdlWZPph6CFmYvKDDRcwZmISrztEKPBjF62GoY3x9EZECUMIByQc7X/iHynj
npJwFhvdtYOaBPgB3JvFKRKCFv2Of7kL54UWKNIck3XDN74DVD8hUT2YXn8Bz3gTbesgSZmJ3KZW
oJtukWwwi3Gn0mLg6e3DkAXk4kMsIX1ySabl+a53RhE9c6Jj7t6mrXcGUfNJ6n8kkD1EAJxWQUM1
OkenqI/B9fbijPnzgKOFQ1v8GvJsjx6q7HAeGXx9w2RVl3TuSdCL/WvFPaPy/G33EoS8S3Z1uUqj
HESxz+mslfTyVtl1/Mr+ZKAhC1RHXAw+WHNUOqDqoZ5P8+s19EwL4JmSkHnVomBC5lMwmw9/4ybr
D4i+2kqN40mW7t5O8IlUmfbCRjWE2eb1sV8+D/KzHMyDqdhyX4kcm5hZ8vZM0om3wjqXAGaIXQ28
wrDZpMQvjHXpZVPUz9qLyE4fx1F3Ev992qM25sLbKXxDds5vpQyjTcYZELvfS6Y0zru+cNAv1aWb
Efe4v2sCgYy8Jxe2yVmUdHx7pUCIP5+dNqWS/Alb01+ZrCASoivAk4sZAYno07uvSA0Rz6gAH8ab
3G2fA6zkiuhmdAVku5Cz2UfAXkeTAi+oEnuXMS6OqPgv7fRc2yOeuEz4+1ZQUZNvhoKU+LmbvC4M
3V7zxbkGWNql2xEHCx0QZZ7u91sa2UZA2cnjJg0vmTG4DjLBIvCQ5YC4qvfOFR5PS/CX1UpnErG5
a/DLLol2zozzLuEn3RNmhCTvOv5KDJLCsaozxlmI7sTDmoMA46l/bnV2HeRSAqIa1MgSsh4V7EGI
PLSsfNRY76IXFqQoAPRmpuEOXf2Joc9djPLbvd3z3JlryHCj61nolVCk34g9cGbHS2sNYyzm55Vk
WrKe5IZmxIeoyh5EG9GoCVTDBSIuURBMYP4O2L+UHnoTg8bJZO1kTzjw8Z1r2tKQlD4L5yiOGqaN
X/orojPMk4mLUwKJxZz2acMeENyuqQaZGwv2o06Etd5ZE6WskEXYjAd8WsJ8lAQ5X3DqmjLn/sz/
EK5L1BL82CkJZLJruFhdW15BRZ/Ub3sAeCtp9AzjrRTelzslC8fRSA72qLkSjG88VRJj/NhbptPM
6+GX4hTdS16UvQnaAjbRp7VR2FrxMjy+YXHrr3DttOyhGzrzNlbnaBGuFLYbP5i2J4QsgM6/V2Z+
U96Zr9BqfjJH321gO+sQrtdHDTZWVOG4q0uXY8u+BtnKNnJoJ7JIBI9eKgIg+MgKu4Bq2fXkhF4d
TK9ek6dfQnXNhnpcAwLBO7pX6IF6T2GHNMy3Aj9Of/+WgBV4vJjnyUzorx32mdn0pObm2bxNazRW
c4o1A3QfglvLVEdCFPdANHKhKTsVJBJhbebYVOMa59Bg2XXBFxVXhXFCkKhZ2UExMk7hlDcptojH
ailjdiB3GkUm/ynIEa8uY087g8MyMGD6Jww3hsLcUHBb5cRK+qvJs61jp2r5TW6MQ1vH0GfYB7ML
2VtakM9aHk9qZ2i5MzMK92R2wLKGSX71QWzlKEgnDhjfinxriypyvsxjToA/g6Z3b+bYOaE8juPq
6JrJ5O0u+wi/BfChSXSlghz3UPZ1hmcyoibmGhx8WsrESeUXbSffaULBRlsRcr3XxJmTm3xCWcPX
5SuilxGjVkun//dFn/c5Fx2co92Upc+wFA6iK/8xBl+EbpdSeHi+W4R6xaxDB+fUFNaMqMa+fA3j
zPkf0D0AF6iCK1HOyvFr2QRHVvee4LUNPfZ1J4IrHuTZ71oRov0fq2dmqCHUGjEKFoI3TqZyb3ME
yO12NLUi1rpGmS+qEezbeXui3xeJrvEyTwaRsVw9vxuqIkV3G89yViDiZQDFBBlJVSFAFoJGgVEa
1oRf5LyMHttKrY53YitZ/deDsAKsDs0Y3Gjja+m+Jc06SJReoXnERDy4xzfYuiBaRxf2aLzFUHX8
AeXC7q7uJxNBsnES5NPmQ6qm/Js76FqHQVLChpH4vgmEJHwCxUSSdaWjTRNMI+T7yfuy70kglft+
C6Kphc1jDGPVtCOMuvQJZpLIs1prPgSHPKN7T+Pgf9zrfqrlzaYneEgwoGw2zAAkiEE2ELEsOo4v
N3GcGYf7V1Ko5nxXLuBoE4eUOVPcEgbran2rRNYzpsKpL52YZZ5pk32fXNde8RucioOF6HXqF4+A
kQcQefmNXdXt+TOpF+fYB9jSzWjYqz4HU5s1XwZOSIG7ATn1/7qZEsYV0x3LBUEhIFfB/5IhePe6
IUrCnolcXb1/Jyg6C3xhDFr4PRlNZVO1OV7lKIaRYmz3jYjmYAJtItVKjtanG96IbOlPo/NmMAR6
eA1Gvn4p9owmUEDFL7mE1wooHuNWLGJ624D+m/BxfX14OuowF+YzdiECKNF9sWLUMsi99Uv25l2n
/fp1pSx305eqY8AqXjeyxIKAjE15LdgUTtztS1WTV2EbhBA3T51pYIVKkSl20b4zapfvAA/oHnqw
FZZF4VD1zgdEc0yI0a4izDtJnNsZNVk0T6zZcWjimX+NW8Ivi74NXILz8QucFZ+VhMjCsr/XmcbU
8/ZzOiPYcfwDw6fNh7NK9nHn/h+E/RszNwmWz3OoacgPkqMxCJksqOW5InzYirzY3JrWnwMUSpCD
ew1ehNjR8XuLvZ//COAI4b7wEuHsY6f0YZ6Mhr5SZcUS+2UefC/uyTwkg2d6wCQvrhdYYQXeWeam
fRp48dzJdF1kJMTNyF5wCFCBCan2oB161ifWUF5HUSmQPa43r47kMrmlYwD+MRCT6ALmT+2sPWR2
3k2cVLJ7iZPiWnQ9A6cTCJ2X10B6YnrguhFGqefEr9hE9H7VIBma2Cg4jwA+1ET7ldqLtQRl3k/N
VLlivKNSwf8lAT5fJvAZz1NXEVnLfD0SLK8wxPSX7mgvwbOcxWqajog3rYe7/2erGrtdQ5noB8qZ
V7TNf7B21JQ18NhM2boODcKuuLhRKceXJUDf78ZLJJnDpNYrevSA5WnUVssjipmqP3Nd6knIrNGk
/u5/PFAAUX1EIOnXUerXvorxSuxr92m0dBa7GUtU44zjs52Mj9wnFILqiVZSJlgj4cUFlMfzsalV
uc09X7iIFZCPXB++ifFfIX9mWhawREDd7RzA8BxJTi4hlOOofmFndzB/DxbzJDq5GUH1PySgLKsS
0TjNqazf1RlhiPw6zfVHTz0Sv8DdC/drb1pVTKyBAvcInNv+BXPY1BHOogzLQzsR+P5PjHBSwQq0
F0dWoGSaWCIlFpWY/3UuANZTtPC69eXJ2kCptK47sMNWU69jw9PEyHSvMdgoI1+93aIF7SArTI1X
KW4rKiSS8Wpv01pjD0/EVQYb2azzu+blex6cm7JwkBEXThGEkAtfgHhpWY4vqj96XsV5bfZ0Rwkr
LeY0+ezFXDbLxKsTtmgOpJVJ6dy5jrC+EfkMCLUK6l6n+5X65jt8ZEVsroOw22aSwfvPw6mLrF5f
UTQ5im193cfyPTTH+96vmFOz81IPbzvxQIkAxM/pEk6lXkJVfcm2278plDz0e7g9Z+Pt+bdhTNu2
ycMuyjTQuowiOpYNpnS+rXhDCGTTbhmjeV4SeS0/eUZ7HILhHJ5/K/l4GZ5+WkyZ6kfyxiz8F0II
qM2fvcbB3zibE8ZbxHOIwJttO+A6xeHneuTpYbrRff490PHueysIp9JM3gp3G4m1iythW35L/1qr
P9smeFyW7i6DgYWd8Gf/oMO2k7iIW9o7nytwQRZu6hypy+gJCeoFAATRrctFVyNOQ8tHzDSoS09e
0KEk13RKIcsBY8u+SJKI+DrkNP0FwIZMB4Qyr1Sn5dTt3bdtoHPyqRIq2n1DQ9FfXMSlaTNL3euH
xTK5ZnzvNfvjzuM7pyqeys3pfYve15nGlWFF5maZNaCZm8e0qU37mL0qYqBniXEx2ntHvj++YuY/
L75xdY2W+4umymgruGBp8RuIEPHrPhui0ASEUNte5hmu9yFDfR4GeKxCtXY89pL5X+TDF0rHH7Fm
EW1zDrzEPI5rH8Kte2QoNPPqX5e5aCz7M5FF9s6A0py3FhXD/EpAtd0b6slsRlsCnwvtBwjEEGwx
Bg3zhotWr9nwLnfGG1Sftx6612tHTrAIWa0Eo5Uz3OmQGu2rle+h6FfQ+Hm5bB/oLwsCwx/LtwW5
QZ7p7vWeplDG4s7JxKQ8tLaalWnnOo9tJI8E5PcslpWllDq8Kj8V1EQRckxNrWbL7tjUmHZtecLn
Tg5GBVysZiI/X2xEDSRP+AKJwP1IyHkC1p79ROivDqeB0n0uN9Fg6WLo3T4XKcp/kZXMhuOFRIT4
nlirWWEeObt8y1Gpo5Edeuh55VC6fQJ/UZw2MBf7nMnBPXivGO/ZEnm2hnzlyD6ZmixypidrpVdA
qW3FiehKmuOGYQr5aLyodnIevl4pgW8Za6MP5RzbChZMID1p1ezKQnHAFjKOyQf6O7NH01Ga3nTD
ZXLGfMTn1BD3cb1CavYQUzEcVA5BfdPkXm/gNj5csM3FiGHpRLXwY8mpN6HMUqTSfJx75C0GeW9r
iNv4aGk/YCz8nIOYMTmtYcpNEQ6EJTq9J6QUh1C9ew0JaFjZkl68FBpIhD45oroTyaPEvjbBBhcR
s22acwqIAEQUhhVf8hAPhzSP5EoRCUEUJP1ucHVedN/DjlTUIVTuit81WhAW9W9Hkp1XfobKhmBI
UAnybNqt9gH9gP7ZbIVj7UGV0jsELyr3R7THB77TPjT/JNi2RstAzxtY/4ZRw/7m23Oh9DzE90BL
tvjJVCsoK+4tA826xKfkbQsy/zAZrdbkD0bxKW75kxqBRUlbyUnHBAh+43quBv258Ox+Tg+WyYdX
IFENsGZ9rdsv/P8+ePiUl3ekagUDuVMIE+rmvHVaC9teWkt0JVizJeChb1qcfKJhEhYVHuBsr/yx
6V/ldFu2ZscAvWYCIDOa9SmbYhOjbSBDSsr2k0XQNtLwNJKtTKRD1+/0dMCW9WIp86zENwT84XXs
ful018pOEhuz1T34+BYn+MvG31S7m+5TQJDGTo1V6RHeo7pxwXa7B56SNofwFFK2klroK/1vkvNC
fNXmGOy2L6x87gxXvV47MCu4GfZbkaP3WyiHbLoRPYkY5HCNg1mucAA9T3FqEjZC5bmx1Jrx4B39
AHJnvwoN+ldUDe1JiR4vvMzZzEOvXbRdcbjuwu9gPOw3Ex+c28VK7lTikD84PY6lLCzSbmqHpAuU
URhF12B6mTiO+gE3pTGc3Yy7DCr0avFjHYNvmgLuyEpS+bd6lUy4uwlcoj2GF0Au5NEwNeQYNgHK
ed05Wy9lQH3exJRDtov0aTUSxJEuRNaw4djle3JzPIrrTy9ljuKG7jejlgmq8IU8h4IvE7n5yS8z
OnMNRXES876Yl0tL1CWg81C8gYEaoKELmC2IKHzGZ3hJuEl33MImIPfWu3SaqfpQbvJZLOfOxm3L
Hq9tiHeUjW0rp7qSR4dsIiTmnQhXlm7ZwrVZrZWvlVi+GiQMakQqo8L5ySxC55Ks0S0NVvifI080
2nFxsuZ73bgw/0yb/x2VrMxJ/s1DKIyFMsXOxblTyC0BTgdyd2M7hAmTVzjkQzqKH0K9vA2L+g6+
e9LSYkMWu+VfqgTEgvBzN+ihDTQb40+pCipYds2kJylJudvhlOKLdUMZN7OZpfJIQbIAFuVBd6JF
HuaUDsgPxx9z9cW0C2TcrFlIFWMNa+7U8+gxFh3QKLj0AY04hw2w0rese9y1njO4zMx9/iFyI4D4
kblxPCoGIeuhu4M10U6XXIT/4RcNT2aU7D9VggIzjwKJebVyegErbpqkwnUu31QvAFa9svtJWoyu
d0NE7dcoYKwAbN3czZLyXPNlR50MB8jUj3be3Fq2xTCPM969PeVgkU1N/++UdDIVpZ45d3VTDWaV
TcqDgmQl1w2wSw23XuweaT8Ja0wvSQs5AlDQswgMCvp+vnEJ4Bqt7bV5b2dRs2EQIBh8QvgaMsRx
8eSZF2QU+lKY4AqD2vbmZAOx+ssZp2+vOSpHOgC/cu+/CqHIp1DVyI3DdXFhVuT+vY56NduhrJwh
HUxCTqxIHebFEuwmRNWTrYE2xf2xc/u2av/iYyC3qD8AywFICqh6Wv5bClAxwVZnNhN2ZYrs8k2Z
1QQTbXKWZSacWMD0vFM6dnev9m6+/LDsAdHQYvJXHwDS1RYHED7rVI3EcrhojfyzvxUEfnj794he
GrnkiS8QYd3dSvwmq1BUrLGt28Ww2mPBYlmlOK1FjHed4q1z67RjAhd1lNGfzgBz5GJDXYmdOl+N
ahQ6wyne2fh7bVNGhz10xKf8e6NW2KwHkVJ0K2yNBssAEDookymzYwGoRfkw6qH5CgbytSta14nL
VHcn7e0WcZCE2QNSHmauQdX9aIDo3So6J68xgxEIdT656WcArMN/Xf4MYNcS4WkLJXYaamcOdFht
46AlMbb7NodGvscuVs1T3QM0jBFHFDmPYRP+LkQHN25bj3eJyHeRgBXI2UxJnDyFiQnrzlMIg6lE
vwBw7XKeV/3mdMnkEjj2UfYp7PJCfhSahnPzRWzsNGd0kZ1g1GX5VSH0WxuHjyPZksRiUW8RRN9y
IOcrUTVkaDlZBMsQLLXpZD/TlGEC2FWdn7lqMY4SKksGlVBy1++bzOteH5Rv6OfXdY0V6Jp1GdZ+
eRnIDwjhjHc81zTLvWuRTxQ8PWAR+39i8w3qPPxaxplOjSU9npwOQIVWWLElymJKEQgzpktS9n72
8NMMhNTI23i9CbxDN6tOv6+OUVrP/QDUuJrG+V0rtHj1cCVKpM59ZQbIOGTa2kz1swCEv/1EvNNV
JTuDSPLs72f+ZCByQGmC0Qr4PtIuzEmdni/xylb51HQEKd9xAhh7sqCI2eYt9BBQaYRA7/Kgny7V
hzmsrgqX+jsWiPLRsiinBAFpaQKAVXRXTpR1CjBFhu4juop4TXKqNjNfNVBs7VNxKkAbUityIYGw
vELq5dG17WPg/sS9ZRXauH6L46imUbVwnMUEfCQOs+iz/QWUNsMa9NBoh8ychDrZKbciGqLVkcdI
5Ohs0ql80hQFg6A525dFAyyv0W3KQOSt6L0csMjfi0vnIB3FX/aryB4MekaZkVf2gUtvKKvM4WIb
nVM5jYeF5lLWvxlx3K5DaKwuQj9SOrZo9mxRsHgC67/zxv20ciSBcErZrmH5wF1JX6kUB4B7vdF4
mySWRfLs20U9W4brWD/ac72yRRkpTp7VStO4bOp83GACEGntBSQloboFgKYfm5BkIOo4YmdLbQUC
ygP/4mA6kTNWgDgb+0PK1ybnG3aYjgSgvwBie5FQe+ZHagnpzhliqvOvctFb1g5CrABqhqXzitqZ
o9hq6xUVS24Qa+CWaghFsgtj0Svobu73kEIKAZaBoftUmNuH2pry5dr/ejf3h+A6qQsxLtzFvM7/
mKMSdy86PE3XXWYP124MVVmQwPpze62ZHvatnZatkE4esvb5YTHYM08mYotAi1+DaQgj4zbUp+k5
quXlj/iLbYNmg2Lr9oxvRHxwvPjH/UNnJdtAOnTbiP5cd+9qoikeXlOOYuRA5dsDmJSRODxJx1RM
jlKeEbZLMVzguYvDYOf7cowx0nOlhxuG/vY1a+U7aNqdPjgOBQ7Ler9ueZz1XhbB2R9tB0T60mJ6
yXbXGoHISMhXNu9BYPkDvB5GZYN6xV5h3jyQ8tLMLho9pM+BOn8b6XDMSf/zw+WGpEL3Gy7hVzCj
Yrxx+UQc3W0sxM7Eae7MFalgP/xiSJYgR2ynEWTZjeoi9lXm7krf0D8A/LtFrCg0/ZYlUOYe+kjQ
/UIhl/zqA3XYiVL/tTh2GGwrWLP1VKIDeiQdzAJIZwmWzvmNi5EOicNx2aSKuJAPu5+QqQhPB60Y
A9sRkguy0yh1X6t/VaQ25CKhKH28+9fCcYLlNI8PZWbsMIxloUefwxs0X0MfsAH6wSb5RZ1ypFmE
LNq3OciPSl304Lcwme7czSmarlt1dvia9fcWx3T8Am5qirbsnip77WDPSyiRGBstjGURsupR85nB
BkHn01QeV/21NaeeCF+23Um7AkfuJqMhgwEZWLb0cVdmuYNZMDFRgqB3fnKehIxtT/AKv4nr7N0Z
ajD63lPy9X9JtcfLO4k5ECpYfHjq98dVQEOquGBtZyyVq4+JVSUNAIUPX358e5glIxfswYPqyZkt
6SqfYHDBjrz8TCU3vTGXIXueG6jsePobWbBTDw8XCOJ/8a+GL34gJI9Advzi58Wz7TI3bqi+D7eH
v+yHvMByH7wh24/0FFnQrjluPEyifPbl7Du8N60VjozQLGCG2BwowTD3JBUYZS9voFuGMaKdFmRE
yEOFoJHLmCMPIxKGa4qTPhTdWCNnY+Sgv8Hdbf1Q98e2SMV4UHkf4xpB+1+v3jzpGPT3IEY4l1sk
0v4AW8WLxOmNZpjLKy7wlz5jIp7TXWDQ/DGSlL6yyOYXJFhWG8v4vbjwpb4Ay4Ka8W6Fxq/2aUKD
0pfG9Y763+mA+SmfbRQkxS2cvCYkKv64xF+lQ4HFgbfjXozHrpvLD8IkSmnMYMn61w+iL8sMDiqH
8/ganbf9vtIxQoiS+kux695NMf0L1XmdGEl7+a6khH7j1Si3BOwBmQSsFKW043XgnXr362f8VhVD
uT0CU38MPvP0BN9rrmXoZXruT5w5F0gtaCUv3/2mxzD8ANk50u+zBcQOX9/7rG8qgiWeCS3PWGMN
2+l3w7bL8+o+mhnK268kasu8zmVkwPAHezcX7umNYwFiIDaiVJkJ/gyBTgqjL/jkrPDSufyVNjki
XuoRmkVfLte2eOmwmkAaHgjdJwhNQ03ViE9JMAwlVVjRjipH11qIiM+bmvhrsPeI1jR+MB0ERmM5
/+i46R/naZCw8sliHv18Um9HZXkiAj8YsAov5uVxCKdvAGFtFQM88LVeljPwFYUEXontx/eHoTM1
2zrlokuYHjMEwkGcIxPjIkkRLa07wskry9Qq6qTOi0ryc/R6daTbKh8bZ1F6bkVIxq6rvGDh/T+9
xgI7plOTn7AggC8UqM9NDmyGlBLh2MjTGIXFYydGWNijbDElG87cPgU/sCdVaIAldPnUe6XFYRsR
DAKo2Fh7pWXiUwUSLhuGdRDaJTBiD5PRaML6IehDdsqkarGVNjelD34ISA3S/xTUr/DElNlt1+nO
MUr0vpgBsV88exGX3vrwpFm7VGIspa3Anz+Wzm0UZCYItDtcB6VVCmN4/4lXYt2i/D6ZpHg8C8JX
01CkF7FRTXs12WhjDkp/cudu6rOJMNLuJssc4mNutS38ngFQyTl0Jucbwq68KcPKNn8gWRMyUiqA
V6echajARbIaR/Zn0N9GQ5fW7nWZ8Y0izghtbuVyxqyvp0N/aws1YGrUaVIOSULWLKIO1alpqlzF
rJgzvqa4Rl/mHYC3C1/VeMLDXkdvV6AaNKi4aWZrIp5A0CBPSQs/RFCXkrVoezSZL4tP2M5vh+4d
fTcYj1Q3ajVT47pgu/d14bFdIkBwlVnVSJmUs2hvg8E70lBPFzDN39wfSkHQkEB+JTEEhdZ6P2FZ
JRUUroOoj5DxVHDQ1ca3XiNZN25lyQMbdVBEh/uxjoQAwCV4UloYjyN0mt5HzGHthb3mPagLvtUV
70+btDF7mB+8Mu2MglwEPrnJpB3Z0+FgesSXJRVe/1yFAAclgV2wOY85vCGyQ8gj8bDxaqc5AWGe
U5pIgk4JVh9v8GJTszw2xwGY4UUIlZi+rCNYRSeurX6jRe/6XQFUHXjWWhTOs9LZPQsEEuxN4cWQ
K1+N4DQuE4w6vlDkOQS+06WRuekLNRMymecER5/F1pbKKRTnlQmF/HEJ9H0eychOh2rI3ObPec3Z
/Q/CD0heyGqX8hqU7N8hST19aA3tWi1fmLytNl4rkB5QvBXqQJ3d9ZXsY8dJiTkYzEkc6mUO6LUF
pP8G8w7yCWudf5QozhAkg5vUddbbORqfDf+I26JahSYwAGIxtHX9v/q9f25MfVPOK5rSXITvoB8w
DR+w2+0cGDC5q0ToUUPoaOek0cd0iSNTGlPpFzP+2nCvbOnffU9yoQ+34vuNgrSJW0Nt9+eBUNZ5
dxaunBOF/U5AZa1a6Rt2FqB3cGDebRSv5olb4MExKxJf/fF7WMvp9OsiZArao/TMNqYucZpsZZHF
7y7lQFCfrOVMiM8Fzske9V0g8qgc9h1+PBHmMNKYUy+C3wvKecy3LO7FeEuWEf63a83nxDCzI9ZR
JUlk7zqP5XOD0X9i4WaX8OLtpECXGoaahqnv3seXhuSMiXjPX0omT3+bMOvAoNgtRq4NQaoJCIKQ
R3OTuAfcxrJ7Cz3Cv78dsZfoh1hX4rNRB7jQcVNsoPdBIsSbRp5bUGSlInyOR4330vl7RdET9wj4
30s4LomXTIO2BDzH7XAwuJiGRxNot522dV2/OzRXZawFrErfQSIwgmBouji+eXjS9ZwcdMkrHgPQ
Hd5uYkaOuAPMcr8ec/bFCMRQMk90heoj1h2XTCbyzEYA9m4fPJJ6CjRZ5woQh0syBBInrpVgEyoX
TCDoYfeQ8BkLI6gmZnCRcbr2QCbT/xIJ/VPr0BZ5t77VM+So9CbSk2J94ts2gMqNIIEG95D0nszb
xKgafeUsQUTOJ/+13baArgWNBaMjPSqxXzzWtN8ped6mWDzIMY+drLmDqmrCpNupI1Wca+c/ilWx
FEOs96LWCd23wfiNFvLvabCweeKXNatb8ooDY/R98eJdh/yeMOhi01NwiYFHG69agDaHttgd4blp
Fx8vXGbHO9J1ZZ/UsLlhCNubqazEP0Ve4HFRLYkeBiMuAxZ6ZLe13PhXd/fjjmvPJjlityBZUDRd
0zCm0ZUAPwTlXyc3adv0JuTlW6yLIw+yn+RxULBD0dWKSFx0t3LQS+qlP6Zm6dHfSnUxoexXr1U6
vjNOrJ6ljMeuT1uLQC+7o5S7r135hRUgtpFfPKeh6iWAJmKWvVVjN/a1SIZJpnAnzwNQ54w3odQ1
Xmpj/mMUVj5klrU/ryConRC8v/YImO7YO1ymEuP2jpXSwoCGexvaDlDhwPQTKk6qU0u9KmvHD1x/
BiO/l3yHrW/PagF9NUl6l4e3/dL6LgytQEviVCfFpkV2vSvmW82trQCZnxiPwgg99BFyaWYhzrwH
hv7VGUhCIgRRiyGru2iAwvW7UCG/hWZDPPpoRHdoVRm3aWTREhjYt0uC/ModWf46BRK+swLSV+u5
fkdnfKoHWfNxMU7ossHkQ/7H4X1lb0UpMrhIpMWPOxEnzHcQ97wN8/GCStSs39e2pz4ZKm+lipaI
UCMGljxrfMeoxKwpBLIyMeBG39QW1DxWsGFhzOS4GwRmN3aD7EcSSM+UyXyMnE7poKF92gdDsUuq
LOVBzIi9ZobGCF3zFnk93oQIu3tbk5lnjZi3hD5Zohx54lKmRimix6Q/xlbHQDCmzV+6QFFJkWzp
O9o0IKpz4VUGR0fROPVm+xBtoVE68ITlHd4ra/R9j4brVugAKoF3quayk3RqWSGqypTcdxh/fjCL
h9ZeWu/4kIKj8Dm0waFWSrxfHupHh7H4cThUyrWB0JYouigwVNhCU0am7iH0TplJbT1WWErgV+oj
o6QbhFl4fsPvoghlLU8iKDayrnKCdU59Wl2SR0O4o5VhRzfq56sj7eCVkk1Ls3DY6ykjralbs3sL
pwhqz9g6TxBLZ88EgmTqnU5cwhsMrXP2YhMHbCFnfxvRdiUFWFaaldh865RVGg4rPR7Tj1b6AaRT
Z0DoYZJQPJivDPukRofTxYC1ABFhzgPTJ3tz4uuug1ZcVxWEeiWO+Yt3dDuWtvZ+RPUDtnhJxQhy
d3KH4BmFJZkobG895iknOGQLGCGT424LxOgsodgTzrOdFYZj2+wasJDexk8H8HKCLu2cTb055VXb
IjvfM7hVMUU5bj9/wXeN/uu7jbXQ7sVkmCjLFLicikvrq2CP29owAOgRk8fLPMICtnPxGz1Qd4Z3
is+HUvJw6au5WFAqycgqGorShbFAhtwuyBwrkMK4dfFPOWk+7f72uHg4kUs1Zo91J5CcPKOlO8iy
ujklwChKVoAQGfAPnck49gNNr9RtLKmTrWGGXOahAT83pp1vwrnBakMrOUNC1FpCcLcmpBytIRMP
TyVFckAHMSEvA4VmRrmB6/lQAoMMrm6tJEQfvbxIdhvKjWJFLzCCEtrMd7EE7Sbxl5F0y/Dvh2lU
aQaEg1/tUj+J8wRCiOyvWsgIocHK3paqz0fZostJEMdMR/eK4zegY0+jJJ8cZoiSVAvbZf4uNJSO
fC9iuZraJ708GC/5djdSpvaMNkK0xmOqNajVwfanpgvokPwAR61T0+r5C7egC89WXFZ7Wkr/pghE
Dr5tl5KfETjinJMzVnww+qaQXuVC8maC8njj4WFMyTS7xDgxzw0rZoEkCjK+SxmF3eKvo/r8ByY3
GJnnx3kEIZUYp7UH5//zEIMTygX7jBduseYHrMcsbYiDn5k0kjf1QA7GTRaDNh+OXkNrBt9c/46h
kgxHqwQWBBPqOU/BN4U0Y0T30xrbQ+ib5ljdgVSP+N1uVpwqUIFk2GD8t2gwkRf3mNDmDzUlmBCo
McNTTgEfxE7fOKMFlsMbPQldVmotLh9xfL/yipXkW48kTGHVXN/KBN/Kb5oGhyZAY21j21mh4sbo
Mf1iOApioV4BBkTRDz7ewPj/7Em2kaik34/mjt0M4byY+1zJyYg9sjC2/B65Em8+8thK/hHXjEzi
cwcMookI3ZwGZVeYaHFLTq4UNflwpAC5tJ1XVPZ102809M+XOifcpH/mwtvK//dwvliH3shngLGl
ZEbo27Le0ssqPze2mml0BJ4g6XMpAXV0Muqq2BVz9Hpml+/NNG4q1ZHcWfKbEFjBPkCxHzSUP3WV
4u7DEBTZex09Bqd9pZfRx/URRftKEF5P88x0S/Ux7UxOrJ+4AyiMKjI8o9GEdOtfGjr1yzCkJmaW
z8peqosIzs2ObvZzbCblT1gI4VsoKP+pn/sKmS20N860aacfd10Vm5YZrVdQG/1R+bJsH6flUcua
StdgoSRkvAfR9WzYJiQdu31Z5xcHlQu1w8yXRjXgNOPmYKM7Cy82zXmXO9dwWweGYN+y8yQtCFHo
VzRuSHGvQOV8EpTDQKBaHjBMBHFNLj10ay+3tykzFxds8naV3oLun5KRFABPTswT1+EMmsHYHLAI
vehPt6658SNM+qx5R+DdjxEohFAs1vXgsbQbZaI+34XOHvBFE6hijTO9KllIZt2KSAgHG37Zlaj8
KWpzFyi817U15UD2NeA4y5GYBfP6anbE7NMWREXv6fYmdefP3Zab+b6EWc7nQ3WSJJC5tEwkbfQy
G5rKNj+AQ4+i3+0PB2HcJJXOcD7PdfSKFXwB+qrZGHpw+jZjoFFW+BUAW3GzQQBVMsGmBqq2TOd7
bQ9FrJ6dwCHGWRuyPUYL+Ug1/gVmI0IT1Vusqekod8HODzLmyAjnsDLWCDgPbjeFVheUSlBQPpkm
x9MrrIVwGVM5FhkxxsL2r8iGV/huUSedw+8MD+Ges658aN9GCMSNbF0lAlV3iB7wK7f2W4zDPkYW
znPufkvYRIrWJZC41mqRixcYJnabWNnotOlQT7h7b76d45miqsNNu0pnrZkgMucueoMyBI5Mu2mO
8IfknjKVbRvyYEI7aaLqBJoXxexB/3ciH6/O/2qzA0+hKHLDGZfYD/To8Oj7HJkyBZQ4c+ZZYOFW
F9W8SELpRLJvDJ9fcX6a3sSFV8CCdfVf+hGAnuggLAxx6NIFHFSNp5hUvk3dRFJ+PvFxxHZDh3YD
fAeiY0o0bWXJe4IFaR+OHIZ4Etp8pF5W0OvByUDZ6ag6BZ1c6/Hat/iVPSn0OEgDKFN5tW4Q7gWX
4FwkbMrhvkOu6ZMfQMNul9AoanM1fz+hbVfPNbuxE529YCDW0k/OM2zhevC0KLlM+Tl24ybFalcw
X3t0GeqRlwZdXrMiTjtSEJRWtlB1W23OUECTcErYuqd5k7Z0V7hJs0uhzdWCcMO99OpZhQMj+cKP
DJvJMdx9Y63i1CJ8tMBkH1MY+UaIvQeC1hDD6LEfrNEPjMDGFtsiD2TtzR3zAt3zWhOyt7iH81Bl
J/t3fr1Zq195y9xIxHpKnKzb4ZZsbWMocaH2RHtLkz7uMfMueNdDVv35HVj84p0OY6Qi1jifafL6
6YytTU1qfdFBV6SCAQiXd66BAXjUrXYm3rl9wxvv+7NNop7yDJrhQAMl3e1j6XRIKDhc2S7I9uLA
0HjnJf7H0/AxTStrrS82fwnJhOgUVvUZKZhR6S2ozz/zWAFgKlUbZ5VuQdzelJH8ny0y0XvOh0hN
DbS1WeutKyFuYuuN6RqF+d4fFByhfghxBoG2tPYGv5ghaSngb8qZmOHqm4cH61XlQu57uqsp4Rj7
w56WsiDIhDwHoV20zaLgjIy2n9B5mFpHRzBiMB8gXxM2CGDtdtXOtvfcTd6gw8OuVcCSqX94mSJZ
ccGWJNHbAtG1iZg+GnUfv1QGCf0xFRZEZGA0VhCPB6fHpGxFnKQN1R4YpnWhfk0M3AX+zFOq5yed
v6mlrvdTcBVD/VgDMC6CidT2IB/Wy7K1fYtZruddZZh0ZN3fLFqaMLnL4DaUfSUT9AMH/loKI8TG
OCaQJVEYXV5v6c1w6PX9QVun3lL8XavojDc2LoYPn/Qc2+Ah5gvR4dmrKb7tPoxLFvfSGQPkszV+
qwNjBLmTx+QTxbaOEq0G8nBDvbhiorvNcekOv7NJrIaaBKqNtDOg8ArkCwhC8GAKp9efszg6Rgh+
fE7q5HjvzQa/OfTlP62M2+kTYluPYm+aJvLLoqTxcP4PHvinZLOn+l3jIKwZpbXasKU9d218syS1
OfW0f8WkNREaUGMB/ZoMCP7kBd8bgy1thChE4Bj25i1aB5oTGeAS/0dZIvxZXVeLIQwmimWQyCtI
AIR7XCwdC09cQt7LlEe5TZ4Frh6y3a4ACYFTz1mjP8JgizQWw4Fn4BlsVwBJNvELmUuS6q5udBXV
hGxRS3tZ6Zybh/wLpJntgUFrGZAy3TQmyLPY5lcWSZWpljsYx1CgqNLBsoo8+mNfU+AR8scRRLl0
oktSgDmkQS058OzcAF6oB6dOjcaIIdTvF1MdOmtuVmW+zy5jTaUZZ+SKneG3AWDKAxKbAlPXsb9C
3TfqsJ5/q6mETj/sgNhRugZpWCx3D0K0CvSA+CENZIA2En7bf3d38UtkzYtFqFnq5SaN391fYh7i
SHs2yIdudV53+Bq07otQyvWoPa81B6MkbWNev9axC96lNBWUj9l0z83TRxpADg/DbS0EEIxemnka
t9PTbdHZvDAC2ABi49PZrt8wCQGEb4BDf0R39JYte1ZGDhmdGGRU6QG6K5GZ1lnx3zwH1s9ma2Gm
YUOO3dnMlIazmHy65xDoHEiSdUdmtM8GSxc9V5Qpnc8oljODusGcdm6Qp+ifNfUcZObsePLglBTU
Yen2hTSIHc3JEerP6xpEg9FbKy+5ZSL3t14QF/SCoKaBcgmE5gTTPkw/AzDYkT/1+RutvuDbmDho
13MHL9bJu1wgrXqMSKT0uWxvobWhUo8iXoLsx9GrzL/BmKxQVjSjlumYa4NGG6rSJWpXBjsjv0vX
ZoF/N/JLbPZr5jtF/L8/7XzuILLUtbY0DHYTZ+iXoO9c5ziWtidvmygEA+t+uV4jJseDTd0vF+G1
lVJ66TkzaxjutTc5FGFNqPOvxNvL5WT8l0BktqJIOJpjFuDVJz6jzr7BORBFFuVxIM2CjvlvKLbP
QSNYVvw1cGlSq/G6/ahnusQhJ1DUv+4Fx3GbXBXbpEoBDFjMz6Hm8/msPpcjRkzdkeGAoUetAn+C
cjzm8PF9TGPIRBnWU6kABkm2RSifFnqDgoMsLUPo/SoB6/tuHPtMNYL9D5vkQEmUfFOY+lNfP6Gt
rCgDPvtYXs+fq9mHic4lS3Nys6F8/Y73T/3IKUcVqx8QvU9D5R8dcdPc46nDTfL54cOnulDb53Wl
T4v0ntVwdmkuedE6cfw8q7HexUsAopvNfByZzJqyZAxwTCGnZu1kEWtxgxovwFA9XeO/6HmJXnxe
wy/VlpEnJ2i6OwqkY++vFmpqKHwCU+NfQGn2tetJDvDuZfFje5DawzQOrBlmMwInI+uewfM4k8NQ
07r4hRw4nLDDWxduyMlhBQlW5twmuXtIZhBcBzArsLPt1JoAj6YuW5Jx1w27mJ3YxghCnmQgUjTO
z/+UHw8RjpT2PqgE/Cu0Zte2QFPtjEvZExVTErYRdUxk8r8yqK2teGiz0+0jAXRpTuWIi1syCWDX
Y5l5LeYPzx/LdjaPypmHd0yZfxfj12JJ0TZHSwwMWl4HH6Dye2yLLFouiUaADYJiav/jKdLV5FiL
m9+jSI6UkXMhmvPfqUG9GwV1LN0mkRLVp3X0ZN2ctkPYii1ITKB0qblCul6Df8+fH5Czl8CRlQvF
0PeFssh0yf+uJfJOizTsrAyYvL2ZWTEaq2wCQY2/qs+7smeltdOpTqZdec+oPhd51yoN5iTPgnPo
Fe50+cxmxy61Hb5X4NGCotyC+CXssHR28ASs5x/bGxBOy49QWmYeYtfPoIYfzlom/0E5u7q/fvAu
6eAED1eXbIbqGG5fZa7sAG8GRpUyttfOUaOGyNmEGmqQ2nqlrbLwBrYz4b/UjG86G190zIG8to30
p+teLIehBIN/xUMXaKC0dxGxFKcDTww79gidTFsJNrBF5FArlPYj5InSxzG2YQDVoU9fp7GUwR8X
t5ICUVUBpM4OEkoVs4pFifi/x3yZN9/dSoKJupdrjTZxlj/VhB6rHEC2cPmBxMzPNCpiylKsfFsr
rpegq2zY9gI6K5ejXb4ah/0FBmFcNZtPaL+wnIoOp26TCdHZTrerUCy3AbimioQ5FbRviL8yhw6k
2vafL4/J2pmfvjX+nhCvSowgrTvZ6kl/tj02iNN69p0OqJs5oOldw7XaBaRz6psfB1Ss3TWpb8we
j2rIDHh/+TBjkqiqI+84YkXmFKLs10COj56YnHvYVzDiNOUMDwFzK48IlaenRzlKcKrdKzj/HJKN
1z8A24EQ2dwggj1mj3Z0lA33EBY4bVl0qncu3qiHffMtVwZp+f7M63zzroE/9wLv18yD+fSIWHC7
RIRmHLUVNGuC5S7wvy0G0eRmDJ4TSUbMLAWdW6Umtz1oKKcwwG6MIIUvQ/WN65/V74TmoXGaChje
gQLhgtD8Ugktq58WPhAnUjzVqVdEJ2EAhu1nmQuKIbGAtSnXnb9/2kQmqi4H4qe0PdguIJwnwfBd
9UGn5AAWBt6LEJsMka5IIVWwCEO1Y9qyKuohQWYBTCzCjZgyABxmnziwmWvRD/wMJCvSclIBZ4lh
9q0yqb1UHFidyxLGVzvv5PK5kqKqx0Re2OoBbP7LLH7oIPofQAQfErFnOBbyUuBVPyvxLwT6BL7m
/kSiHfTYtz+5tYb8JYphoiTv2jpVsiLKuhc5szV4673ATnblfJ6K3uQm5yfo/BkgNHYS6wVxnUHS
wI+/gONauWfJZXQ+K2I3434rhqNPb26wpTqQdxaTgsuMmm1iUPtJBUoC653zTbtepP59sJQslg/t
u4KHuanB2vlRPpT9xjhmV0Q2XR2EkWERyLlZPGoXfj5Q4CK4X8fAC/IGzURTJfZlrMp+YEl4lmo3
sRRiX72qpEEQuRLvxQBOQNKg4+w9WIZskwI+TXgp5yqbuhRka9c7GWezS8X8hO4rzApGIraTUep4
DTVCJQuErTeSZCiRENWsITNqK6EK31bR5mPrqHgT6RKpnyDzsol2/25d5CohNhSV3WT/pq+gy5WD
SJTsITkFxBmXI6eSCcbK6wTu7bYNvUkqfRUpV2WRv844LzS9SxKTDMmWjXvKVrqvTW8qd1vnkWis
vnP2oeYgxKnT4RLt1JeH5kZ+w3Y2ZdMWYKGQpxTdQBRfXNSEm/H20xPED3tCPeAoOevckNhp+HbB
EZeuTpd+VEw1NLetAA9VD2GQ7H+lr7T8AYGLMCHPdqhWrmSYdtad7/tvCULbupBGkkK90UrkyYOu
ZoStmt3tkhpszQTsa8rguImBGphb6ZAhG7EaK7Rd75+CqDH0lPnXNdIFIuS7+lqh8F+JaAPGcjHz
zCXOV3Unz6tiOlxnJuLcvOfCuE54nX5S6SiiNEGuHTTnY7azKEPmefwOv6qM70QpM7d2GjuE0a2c
XsZqekRcV2KPQaGyItw4Y5BWs05g+LiN1q+tC9tyYuwKpe1lkwtf6DbyLjGJ5ULRmx34a0FqeXI6
xRkuUaVR078VHUWjjE7J1/AWdhBTwgmfNMBzOlfY68ILhAKnxoNiuRU/oVXLmMCpLaiw/WgRJt1D
qCS/0vD+/znWd8eY3RNetQgxONzyePby831oWzWMUvOMcjrnytq1j9Jmawpxl1SUPpmrQGyUJ+Xq
czK5c5M8Vh0S7nF8dsYRxbNR9vzjwmiRoY1AeZm9ouHEibyfcryw57ftlek6WVxSlkMz4TsK8cv3
KC6IqX1szKPk5dzCTpMgQggVIFj52AhRik6w6lpbR0V5mXdRoZVqA5CjFgbPbJ20FiMv84dFIsdE
Kxh3k3C+zP2pPFGuEtSDhY7DoVqGM/HhHPYX92x0njVTn7lhs8mE0HD1YbfSoucGS709yfym78pn
+6ZYO5dnqk6GXt5MfWLIuzeMtlpXgiEQkCrRWQ5qJ9xcz77Wg/7lGrU8U7T/DML+kPuPgwD3MTx0
tntnNOpJLa96kQTGpjk1F5MlqgqxtPmBKgVA271VbbgcdpiH/YGLL/x2Q+xvEkD8oxXd/+PvlPKa
uyCZ7hHF95S6PxZbr7G7Z+hj5zc44loLJKTfFV441wh1ymKddosKFODb2PcS2rEaPrnxmNEdSkDh
sth8i7qe9ESDeph5eT9BucwOdnIn7eZF+J4iLRavS1oIs6vsUGI5wgDO78f3h8GakzDP9lzw/rSL
NwtzFQdOmMEUnQzUd+fnL1fG5aXut0FnG/xb8mfxmHNEze7PcX7IhkIE7zTwJsFva+B1PBNKJQMI
MNbxEqQe/1o7ADBRP0+HszywEwDUpQIvr7XzdkD2eYY42C1ujWSeWVE9O2hcppFBIGMrlXJ1bmDW
weSfZHmWI//kJdXzoxJcOVRp2/M/M8sovCOx0a82Dv6PN/rL42EuYezem7oWD7ft977B6UEodj4u
y0MkUg5zB0siTurGP+OjWjSDOZvq41LbiN9Lj2mFA+Y1A7L68PniXOtnLyK3FP0yXeMXHABTzNCx
Z3rOamvIEkqM5FWR6l2aXbvWAbPPs+3t0mGiA6KinVpF9n+f2jjSsaqMu9qr67lr8ou7gv+elodh
pjj50qibQ/741DIuldB1T3sy+6TjYhxZuwshoVk+r1L7/T5OYFnndzQTpnCt+fkdL+pIeBwcA/mS
PWNDQUG2X2SiLhqpYWdFKYX9q4MlfdwSjebafkcGyWMzyGzXFJVNED3Vdhg+G1SHIV+u/wcNXAo5
fGa6oMPe74XYLCP/slFObfL83AZEvlTUu0MG1vyMRavpkeIgSNqis9Ltt+6fBv65EfB8rwQqtNm6
GyFQunDfGfj7fHVsykhmDqrwljFUOmiWTxYpHwSXPaOFL3SSKwdT+L4Q+q20di7d9Cy1NdyIUjTs
f6I6bVANBhidEO4RDBTy7QoShl7RBvF23TBntP1pX2TWz527kFUYWJC966AJDE9oRQEqvB+00dNf
33UfyBeLynVZ4t0E4rV9HdxwrN0s6gme1d0hP12oskLnt6t0c3mdTXDe4dT72aAM2pI+Bh7YypMC
564DzuDVevlIaoD6jvEwwa2f/vlqjtRXHjqotPmQ4od8nVQBgLydQam6GOLEn6mdlO+wqDpe5Yvf
EIElttUVUASAm7o7AuKGnmKmMlIK4iO6seV0itMhfP9Z0WFJkROHq3pfIrHa+Xi+Geu1bS2xHDRH
GYPc9FuprXeYaBNOPkhyURt1L7t4BZlB4ETzQaJI9wVs17wuiPIoiE/ylrWBup9FJBoJUgcqEf3I
ACq9eiYP/X9z9+SrCfZ4xN62Nuqf/tONv7ZNPZr0pwI7cJH+uA+4Eq/Di+WMWIjJrY+FVpuFAMIw
UWH2hcKq4cFB1NzrQnvG1KA/diTb2Y6azr6KLwjtfgOMQ0Hj7MkGlGCxNzIgKxPBDaVHbuX3EbDs
0NXOY4C/+tFhL08H8///4/EUi1B32jZ2udoO62Cy0EUqtGbwtf8nzo8cB2Swpsa1269KLYmPztsW
vS2lun9ivNyU9aaC2XstZ2MJLjW9gCNeqzCoNgnqAzTNO6yDHz1DLLKSx1kbaNrNhrtb6KMjjSXH
t4fHadCenXDoyABmULrbnrPGPge9swjHtpC76Anh/LBsrnKFaWweDsAOGKWt1EfSJWgFZ/oUOQCV
pcZVHH3FdeIdTc0y6L86zE55HjiDop4F6FhvAxTE114C2/7W7+3uIfTcKhF9p7SLwkUlBDDPGMeG
sS9TBNHQn63Md6+74Dj5m0uDZpZt/ITx9/WbVXmkCLvnVABjG4pbJR7rNzVfOSZ3l1LBTjoM/whE
hZ++ohOOVfkwX6Ys1FawHrGZ2MaQWlUO6aESlv56qNnfwxvU6xpGXdQdu+fm8QHra+0EMHYtWIPS
i5S+eIrA9SOz/hU7AugxiqGIowFJmCoWSMpie1jPWNRmNRY9ddLSARSnn1dkHB46/Aw1AhG0y1qG
nhH024iclE1yN876fqAtNlly+q+AMr2HOYT3SyFgD9kbC2tUPvUUp3JefHkuH8fedEKZrSrHBb5Y
C2gvwRSAm4obi5tmo2VVWjgvnW82qua1E9NpVAFTsFi8LYLSP+p6KzVSDKSrF5mgccKEuAMtna2Y
2CGJ0P+JPFapiTXBvkOywtR6w221RKHTAj6zv+G+IdXyHG15Va9G/0lD/0H9uX1uhiWdfVwL/J8G
8DFjG8DQQ8Cr4SVoaQEdIZj6H4lcPBuTUBV2ASIFWJ6PWYXRLpk0CcxShjN85uUvidYncR37Ip7K
Y8Kq3dIuLvUsJbxjAm2JvQQyq3uYB9fUw1DPZwzO0Cb5eGtzvEnNX+mJW+yqfjIjh8lJs5hKccLG
5/3mrNHxfVxLUIu4eQKdhHcKNQr3bpHjR5hj5eLulibQRAd4oWrR9yY86G9xmNakKrKk4E5VQt9Z
M9wHP/tf4SEWpfPUnfNJtTQqwqfxJ2SBEa29fIx7IigcKChqGXCBTVcUmj5AIHQ0/joyDBXkvUWt
KUhLQoWEX1ypMP9LAk5MBrOQf7V1uhV498zaRxYYtmz5cS0hqisb9jDf+MCSmXnOwKNihmc8cok9
O0IpejKl6umnPjzFi6Z/pWdA3BuDAHIGCz7TpR9sIA0P8RO+LeG8Vw098wo8SHVFVnNq079ibvPc
ICmakKrVobCvWxuro5fWIMIfeRav+kSlYjDs767RoKnWNVWOQpAieoJjUZszj+Jf9WIy+iVvsf/z
Z/LaZe8PeyP9T5w6pr2fuf/iT0Zqo+tGoMNo9OGnUx7nx9lsDYCC2hOtEgYY2EEDMFovv29kp1oi
GiHVPsbRqaAed2XABuqkssKNsThz3D5fOL2ACIsQxBmzaxcGN+EVjl0dL4LlpRKwSmefSrxx6u2S
Xd7mloN9BcnUJYHSfORQAp8epsm38bNNi6uMEuDY4Qs6phUQzVGH2OEVv35mkuoUuwAREiX+B6pw
LcAmGJGw5JT8ISJoThOd2Jup5oD2hgxbXiJ+U+atJ7mK+zQki49KZllXdowINAHIiVy4tFXTeOZl
jsQb4BJPWxj6bF3yzH+2oMUi+DbtY4xDg1V2Viwzv/0fewgIBisXM6dN3a2LP8LTxcj5K3TNcwjM
C1K3QMfTGquqsrPq5xVLSQwudC+nylnnR8giA5RsB14Xp624PyHtyvnJVysyKXSdvgZa4VxQ46+f
MKB+mOPi9ogWqTKenmd9lfy/V6Lcc5SUsMcD6HOhIx/tcAyzrW3C6w5k1IyPVEaS0TS6KhM04iEj
JPTd7sohInBFSK+9nbPBva9yPpfnsGOnFttwJt1T/mnh0oVijEm0IczVTYqNxuD4FtYPLT3BTPrL
VTHyALDr1JpNJ05n3U22MWbv3JyfwH4Ixa6ZgdAh4SqVRdwIqEo+bdDMZjEgVFMhTHDqFBfmGrm6
ddYJrasoMcO4Lwrjz+o6eL8GcmhD/mg38MXz3N7aV8TGkQo2ybAo0eAOQI9/tUGoE0TlAPJbPT8O
39IHL2YdXoTnTu3rgyxJdmhYUlyH96e0jLAqV7kLGrV9ToLcDjPFrPPXIlCMB7g6MDUIOFPb2Ckc
Igcvd5+25VlilsypMROK9w3dcliwB9f8bnfOvxh4SaJG6YfOe1p025ecG061eQIrYDEWuBIX+Aw0
7LJukMeW8woDRUVyLSTUDG6QxILtohSd34MUXoKAa0kzolGLAjV0sNckzflQmfvWW2OLcZ/WJF0B
tHPzGjc8cNTVD06kX/oWv5J+6FnV1BVKFJrF22E6wc/LXyBZvyR1u44bC+XC9NTIcw4tp0Ubp4P7
Sa48useOBRxog7qodUGdpzHels8PS1tujqk+OW8Em88eFiG78on8qKe+i+OvhA4Lh1m3OKbNHsDn
pHRyMoKrMLr6FNQ0Mge2YcLhyv4isYIrD/QcPs/mDqzGLfPAAy92bYIYkmRV08KM3YjmLu9Pazox
9KQeAVj3cyywmEoBG02feSRhFt+kmwP5k0Sai3riQ5g5e3vqmt2wMrNpV41zLGQa/X/Ef2/XtL16
7V3hGMdQSZIbhvAzoSERTP/FIrW7mnTPWwOLo2fC6kvTH7UU22Ohpt1469OUUStElkNZNR8lSDYM
7sqISRV+xayAvoVBGVgKxRtJMIZ6aHOx0HCFl1vT1VJkh64cCiC1OapKCHSzOJ0+mwWOmlEaG2Bm
TmzP0zDVMsg3jZa16ZWl2S42IahrxIsGUA3Pu7G0UVJTc4ncMHeg9FWjPtKEsCrnaX+TljiDRVhD
uXGEXm7LGWoZcyFK0hk+FJ75tvW2JihomPPo6kRyw5RPSrMKsw9kUeClztmxL2NbWfq+JUt6ibiZ
W96AIC/1WLMJjNRVxcYRF7tKbFTXeDZeE6XoMZumV42uUqOQCEB2sP6hoFIVHYZh9OofLWzmKgIr
oSrit3qXxuu8Rv01pI3oaGLzexc8xWLqzZz1YRy5UczLsX5VwmKIIy7f9XiV3aZ2Sz++cBZ9sA7X
QY/0gan9Wysc3AYe7X9qAuP7L9LACFuYE7fWJkP39qcariQgIEpWeVpUR9zz7baZxkTw5PyWPgL6
mnSnRBlFAuyZcItDzk7gJbjyiPJKzSIYRt+IaoCu6w2igsrkMNZdFs37HVSVHyQGQ5D60+YR1qdd
MxDjePhVd0HEHksLi53fORyKkmair0FEX03et08xqK1YJb2ueC289nRB0CdcIi1Aq3SEZb9JOd33
o0ohXpa1WmjuzyDFmR+XT8eOvo56mcH4f1wxcoKph5467+zUXvWjpu8n9eFwz2gDB8hZzTzON3Xw
y80dRGCG33Cw1CU9r/NazZjcElbP8Nci88MptFoTP4iVCc5IDTOnoom40YAVRm9MHRnRwjxKO8vn
LqDkLpMi9+qT27xKkPRKIBOeiNWKfA3ZmnONiPwHMK6ned3+JCfharGQCh5c1p2Yvvo/ezgQmPEO
qZnN47ywXYV2XlLQ4zPuJ20h5cMr3btwl0hI3C7QZQbIkJVYxRvU+KguSXyk/ElzPZBEPpFsNoEV
YvFtdUnEGO+M5kpOC0DFCYx3Zby4i7UFs11xmnmPUxUkk2Lkvwf1MOBxgzYC61d8IptonhzmEdnr
DD9y1ab8+GrpwJh3AxouVUo0B8sJqnW5YStcXz8HI97ISZBYlLsQI0SKEYr78Znic3RN8I601Aoa
mcsctZ/yrHwFEA8Fn3wmzhzGUOhjSzj2o5/cqGjwTgDicdd3ZzUlBgo5Ysz3lypQ2xeRn9NgAZO1
xuNtYhk125c1rI4iohTdM/tdQ5h7/dZmDHHyMHJKKXjnRfFPCvxyt9focHeGNCEOWGmkstU7Vxkq
W84sBC3TAIIjxDChwJb76TrHZA27p6xUk2HhnENUa7Wbnbfg2l7SxjEF/MS8Yt0vRBQIFyebBSGm
YxL8PvCLWYGaUkmvUfZAaxBS0m/qx8vTOW6+ZIEr1WOYEbh2ztqeQavr8hL/DP6s1aE3nohFg/4w
W5g6OCJa/9tsGPmNsg7Hz30ceJsAZJ16uuW/+l1i3TlbHtsfWax6pUfjYx8h2io7Lnk3+g/nTSiL
RXPAUuIDRSZK5z+PtaMLicKQz9Oftfj/xr1b6Abnlk9njZV/CBp5O3KnrK/HAPP4+tnv1zh7sv5G
N7uJhUE/l19xbMpEC4TrgJCec/FpNA7xL+gGLFOEc/LhkIhAw/XIf37mq+02wkXRZFUfMKaH6fed
lwaqX+mpA/+7ejBkj9df5P3/yFJWGyXD/JqMKh6OMsHXnfQNefr+S5G93DpLOCmHSYhSQsY03CE+
KCDNGjVxi9Msc9PFF2jLPXdlkQlfOfFFHi6mJ37HplrS8pIo6LkeOLdbgxIY0N4/PRfUqtJpXeep
Iozgz106cdcCcJZKcciwxa6IxmVGX6EFN4B6jNP7SD7UQy9bPlK81rJkEivqDUFXAUSswCdrTXUi
R45DPAR60e0HE3NueMJWYEfuoYXfHRMruy2OVqiXAcTAXpnEgSapR7udrp8GLdEY06iPHL99EVLz
5VHzcqEi4f4levGWzYtcLnFGSCe7XRtQHH5zqEhZVjG7IM7kfyulIZcbdxHrfPzPK8HvmnJoRil9
/pNnuP/76XjqSMIWeJzPGvPHAStx0dKHbTGJpYSHpJq+06hlK2VrsS8C8474XZYyt1mhZBe2BO2i
uwDxUSOyN7b34+y809aHSsq9UTn+WCOEc/RcoKClG8YoYYu4WE919fSGdfhg2zykhkmUVeheS4dM
ihSjYoN2GwsdCCox+jjvvYWNgz7dqkpBIyM/bSDcVodAk/UdgiuCaeq9RUcYgn1ejLwypfk6Q3Me
gYRbb5/+UyW5n90qhGfaGx1oxXqc7wTBbMoho49KqjhJA/Rn8kOPVD7HPlWC2b3ESD7Fg+0tmma0
HOSSPuh/Ql/DV4XzZrPKQShV9rK3i1zoCMThqeOoxk+abP7focdREc9mXHfZdWP0NMJ4yekqIh5X
IwMy2qXQvU1WB0N8o3sVmhTWv8jOTOBY7/jGhj8XNkFNIHrtJGocYo8pbTIFJgwVyEkf06m9i3rL
/0OxXDxzDzvGeqpdPeyUP0CwhOmVYj2MQQTSXv7QW6FqD0vl6Gbjq5dV3qZB92RcClqy5qQM2S8m
j5AzQ7/4lfBkzOeo4CgQED/c6n+7kLkCgww/wAyLDPfnsBy0vWCu5/mHAJupNVPQKkAAFOnFOYf/
dGYZYVBU+OMxgw65SHRzwrn6+ajI0AUJcHC9TdwK+o25ponrylPBri0DZvOQgii13hG5XZGD7P3l
jYmrBu/GPu2UYBVDUMN5kJyf4FwX6zGNRXxZ6NIQGuIEP41buZPyb4ZWrCy2bEtYzuthg7cudYsi
osK5TEqKSQhqePhqtBzIuyPWpRqfGBrv47UeXW6AxdGiT1VNcH4/yCa0ztfiAV1VM98Ure9+Pj9G
BFLk0SNVu9jkcNUkW/u7GWSEmlF3JXJZrFh33k8yCqhrIcFfrtR6n4jlBWfyYy+3yAWvJLlFVRwV
nYTpj4pTpYGME7XBclLZ84qYOOQdRU+hPOqE0vCukjBEEds5iNJyDTb0WdkTProElEKTW1ZIAd2Y
tPErpj3r1W9wsOJsvNeElykkm6U7AFNWKYFK3xbOGBrLOAZBkz+x/j0YZOHiTRUZKH4yydFyCatq
USI7QBrN45xCGQHQPHHe8YLYnPAOM5FYWztlDaM1BunrD0JiXztAh6VcSq7A5yfLmHdZeohuPJof
qLrGCd41QSwQnx4ese6PPV5q5Uf6hE2TWP/y+RdpAF0xjGw1j5pWBoXxD+l6Hmv3zdcJXrGOOc8k
Cfm0rmXARGm13TiLrqBfXVff+hzluzDHPp/UevzXBQJNp5T9l+wmEuOX+Qlqq+Ch8WtGnasDdcwo
5epDhW5VItIAL4iB16kLKb+2XVCy5vtMnkzJBmtQzPWCJPuyjqXYxrjMi851i2eswtu98tMh68WM
nOmFDPciowr3IYPM5MfAH895ytwl5b5cfGnpcOlbxmjmGPKKB8Vy4GOauYl4n3OQFyFj+fud9lGF
Ls+rVDmsU0ZfSBpHJ9G9IxYU/5E8NzT3BxKk593JVThqz2iCRRVZhYWAPQbY9hxP9nVwLz/VR5Zn
V6BPhc//WeQKgH8fZ6XiGEZpo6wQG4dlmBF+ZDA+O/7PpfT+Fiap2PhHx0hDq41Weno6UB5tEgOZ
bJYhbB7z/Qn9NfTm6uPt8+1ipBUk+LBdczry/Ys+ILqNXHwdLsfyMjIdiMi5B4zRQWtM0Ogf088z
/5IGDv6gdnJIPwNGCOWR7ZhtheJ7RZodBdCZTH8dEf7PTWVH9ZJDsAkbdurJXLBA84DOMCyrIGZf
OYYivjeIUzFsMGdoI18K8/dnV6frRCE5/ZNBB4buX8qTaj8CJrlHeqdf0PEHBfu0QBw2aXwUGLoi
CPPWX6Q/uYTm/k4ZpcPp0qN3+yuZ1G7MdnzzS3w9Qe4YW9o2v+/75zK0YZkrKnrJfwfai1qIKQnm
kRQaobwU7524L4Bl0WTr9oI9LonZaCplqFg0fyIJvvnId1EgB0X/gV7YvJgXeV2vmYGG4VNU11Yo
+uUnPL2D2Sg109JuCZZvvm932qCgq5aSVv8E6PGHbHpVUjXzHa5F5vCmoVQro5qEjlRFIasL9TIA
5f9GF16UBaR3RBco3UIgToNRuiGS9Edvc1ZyX47wENRc6wwkWihjBXtNywtKTyuZspAVcmn/FBcS
VsZaw5SF/lHAXcUKC48aFYOQoYoUfH2ogJv23jcIsH51DAhEDpNaX03j3pDvuZodajNZ46p5yJZ3
rKekTTWvzv20hucJ6cIUOuETjznyMhDaF0IlaoLIjYP6+JDtAn21kpF1RHvk8gLKAYnU/3yr5b58
2hhOF2ylBiPqra08I34ADSNlFneedQqVrtf4CtksyCGxVP8npnTZ4C57TCD2h8QIkB+QOLa5vU06
Iad6kJke3xRgI4uiXXeV8G+mY/4tfsCDwowZJa62Kvf/FVlDa5uQrDxDqrsJsQ6yllmbCL0hHqVB
UzrmPskgCU6FEjJ1kn79wpm5v/R2Uq+OQAmxLOwL648OmYKciI2+M4AEoJlEne555V9lHXyEnC95
pp3Kf/ubojMUgYEO/RImNlHncrvxoqLZMwM8cqNM+XjtBnTmXqTFhqZLkhFT3iTq2KkIM/Cc+o7D
8Kcxx4+i8X225ubU/pAZmVp4NhhjpS52UXDGV9W+DPA0WM4Ezw6u/6r99NU5JecBzHf/b/x5h2Ov
yfxv74OVkIWhVj9Cwz9CfUlk0YniH1/yW5jplMMkiJxYnP6bt+7xaZctQQDRvjxTvX6CgP2Hp4lv
ZFuoUmxaMNK7w6Nwn7QAmU5AJHEhG8CqS7pWGY4c5ue2rgG43Fy/D6upZPFPPnrWCGEulzF0uIvu
CzOCS76YGLvvk50zQchHrrgY/+Ci9xwrkorxzC0ULcj3f/ixYspA2sIBMitnNO8QE7BcXusXux3p
cezIn5gTs/2aGTXl3LmDiLoshJJp7g1jBlql2RNCUbYyT0EBHkN6rku5K4F2W7fSS66bEIGryp7R
M7nfrwQmoFNoZK5xp7M7Px6mqWKljV6NzZdOCMY/21mjEadiYin4EFYKbcIAxMLVDMmbsqfyXe42
94K4pB4NkQUrJiVqoaQX2umOV+T+hxkMoTdFvAGjg0TqBRfudvDfSUhdpx2gLP1rB92Z0Zqll6Sl
a5BzL4fgeAhliUpgFdbv7eeeiENda4wfkisQBIIZqDBPqCL2c3wTjDF5qrAvlXsWGwpWFDnvwkm4
PcTb5MoENa9xmm+q7Rsg3dNhGKFiBHf6iTbKR9o/F6W9XmT1oKz9O5g62xHiWLWxZrWTvVmliy1U
sMlUBSJ6SznoD5UX23u7TrrjOj0Gq5L36aKggZwUACxRDRjrqhNVVhNZVIgo6hln89TpUx99bFw9
GgLdi1NiM4Y5GYy8OD6qC/DAw47pP/DzALW11afhnNY/Mww1Durx3mArh2qKRwqqlBr+tD7xFnH+
07oEpOj7TqNYoKWq9nwEk+WDjrZeKmRQhdvjZELkG1hVw4I6195HYn4c7qYZTg8w/lw/tv2DyV5O
eWXe1vBbrQi3X+DFKraBXUIjkTaqfAqwUj/D+rEAJbrSyv11boAmby3fGiJuPMfBT2bD016pRrfa
G/rvUBTbVxrVxZ23LrRRFXGv1vg7NB7SIrVsN67rfyt1exykFUnFQjKo+z0Fesle4vAi+Joz+Hom
i82MFwrbxree/komHK4m9dAU+CJ/mUfxfkyjB+e7WhvUq0bAu7ZBgUyLfBhT0SCqWCm/TtbVc8Zn
b/2K056md6HGSqaVV7vS+J8+wZD5gM1F7AGP19q8EhU6pbxIv+B6EDdOfMTo7HMliRirNMJ4uRHD
52p92Ph9+tyIv5ZcK13Q/oZNJUyNGuPmT6XxA2N5lELUpX8VFy3A8ZEKIaabXfdKLl7ELndUxtXG
NtNTFy4ArONLcRu4v851uIqW+24AcKTMbr8SW02OhSEDPByNJ88s42hVGiCBzxO1BQdiCmBtSrDm
nXij2ve/qWIzAw+DkhUiQmlWUr7i+Lq/Z3U4FShbbY09ofKobeT7hFrIkeW9N3xJdSImH2SJNEfm
3HWoQ/0WYjTEcAa3T0YRJgzWz1ePnHZMQJKUviC6lNRh6OcC3PW09TLVVbvS1FSlMyFG5u1v89Ma
SL81xLzZDJf3pQmGyd7zVvEVMUBf3DvFs0DZC7uTP7YgmgcHORA4t5XZmmuRr3G6mdgaKCqh4qZc
ib8ZYtQxhEcekM2GeJhvbAEYOUnIu4AgasI8ftuhxScUJoQv+Es8Hpvfg+W2UI/L+e34Dht2vYGH
3IkkH6swvDKT8vPjkQlJ51mBzXUIvJwAf4TZ6ahMjtK1AxE19w5b+swwvdQEhoOqGQWEfCX9AgEp
2V88If2vvrAb9+Y2GBu65n691MzGVL3eYdIwFMXmb+QYY7NKBRY+yQNQB8pXwfdTBDo3EpCR0Ypd
S5hHggREd8EFAGgtFPp44DK1unfVrnuwGZg5Ec/eXY9zk41cH9N2qqGjc8Gq5F/BU+m3JN0UUyjJ
9D5Q8idm3ORQb8ZGanfWh6zlDemN+soC6VSWUSrsQPIp++ffPDQEV6ZiTl1Y8Oz7MVjducc2Zf7c
jmOXXtHMaHIubkuTvXhmaQLB/GuDinTcNM/qEGEG8ChzxQiDSpS4fUT3VmOfbE+1LBJjsBGTxbrC
aVrn8EHB8irHmG5OUHyJOgiekscaGCrmZCocemzrV1hjgO8G4oSBq0owPJj3Gd/AZglTcKi/9WfP
SjpO78waPg5UAOTdwO21YGrGn6oW7m4CGlyUvjmkTeSNdc8nzIeB+CuXafJVvEqQkOrwvMHEoJwQ
gwTonVOL7PzP/Otwe0G2vxAaAMIpEyqk5CsFFA1BeZu2Z5SrqhtBBz18fYjMdxjjdiRScyHj5Afp
xheJB5n59UrNiVt9RqNB9VYG/IjzLEPumk0qC87PrcjQ8CT78O+dIF87N8R9fAq/ttOEE6px2G+P
7FXyQDIaNX90jDHjJ53n1dQxq6vzNauCjgXCfn80jTfvKEp48SGb+8naggaW1KDIkeFKs/d4YsH9
HLQMiXxF12PQB3IN9HzaU5inT08dWe+aKkHxXpIEFnX6NIIopVK+nQ8r+k1+Te/wg7zozrt6cIW+
gjoKq+pAaUg8+61z0SmrWgDMiQbo27SajBquAC8Y20MfmNXzAmxN6PUoMYaqYSPymDLseNLZ867u
EzZGz1Q3Q8O1mKDrnkCE63B1+y/FC/sZJ8WHQuQdrCoRGSvjMg4Dq3Bxtx+FO9lpu+OYlTVJe2gy
jmzxtgx5hbI31z+7eOLLIu+1sm6PBE73Vt2902qY7T+F2Mj7U+h7EFtYSTn3STLeENcnGcaBtnKQ
XrM9dHKKELguK0MupEcZkZtBNAaD6S/fmgGNDJcLaNvejK/Yeoe8faJEK1ESK8aifky9TQeOiE9D
DDMxAPVgelAqcBJX4FD2eegvokTpaNZaEgsN2ymO7vPNzTzWzjx+UOjsDILt5taVU4UXGv0hSjBz
VjIRwJJLDMyuVOdrmny0kxb9O6Miu/ysGim9ole5FONrfnr2Mg1qsDbrMaVy8lNbZhrVDh5Dni98
4geTLxY9hxPbgC/ui/5PnhJUZsX8DUZ2kem24GergKdKyK5xu+ykdqrmdKRlkZETyd1d2p3jNK/x
pvr+bJYyWpWMsoRo52ZSscVNUeyqLFiZNchwKddR7r6jguKUfiC5XAU9KAsXb3Ejm0quS8vWSUlQ
HVkrbWgEV3CNRP1eSdsh8g5icGsG13RDSBe3uFA05y1Tg2tQkZPOySv230PebZgg9RF11WRgKpvy
4V7kPU28R6ewddTT9M7y+0jhn0qrrWogeJR/zi2n2l0JO7WRNSoke/+7u7PNtubNYDxWV7wH6bJb
QutYdIeK6aRY79LRuHcr//CuUxA9TTnbzuXNNcqyRWM0JXzOrLdeCS1Oo1t9POMWzxu4YOCKMOHi
5Z3YD5UZmKFLymcH1Winc93dTQ+E7/z/mDfgl9OTlQblOkX5/qR0HTM3RzNFi6V2RPL8OzrMnS1e
y4aqBZ+6crSgyzGiTaOJMJ3iffIiNkqU0xk+c1ZvfwLzayIEbRFaCOxToE13EWXaDId51b1yEEtd
gGjioCxRGCoIQzJ9BWBHKBPC6v3Af30Qf7TBCPl/nGd+sS8cvYfzebt/zAFddC3vARv9FEzdx4Ng
zBWjSE+UOSyX6XwEHBPp16Ah9htJrACNrIrHVbGRANThcUfHrb+SpwTnFWz3hHOs9fmOL1U/Ke7v
keaegwjznt9QLmuIvCT6YqcCnWkRtogeRDRDys2Zsuf18J5v1D9D0mIEcZ1mCK4NeUaGD0hy4Bnq
gspGWgwaFqLd47XMjrmd3QSj+2b3u6Z3MY0syjsS1nefQg296fEK5n09C57X84CPlVWudU01QHUm
tdbULMFdZKtsbRKs2ilX/1gbeHMNlxPh1RybeafkVYURbWdCdvj647eXwsRyKTA5hKKm2QFTPROp
H6pf+z7bTbDvUNQxbrWCq6vO7cSFsbN4s2Le/N0XnPBmNFKty7Ln9KHaLPdHrQZIHk1mVh2g5qZZ
bwZIsxelB+gYYwUQ8koxPhR+P7a6dnQTFZi1o5o2q+gkbOlOH3IOxkfgt7XYtXSO/bypAPB/Sd8A
gqAsKXAbQSd/0L9sNDoalY3eByYxhfk0/nBK8X9DlKSCt1+dLsX7LtnKZ2mvcUZxYNm9lXshpC4D
77BuKJBncyhPGwwGPklpTXdyTVnhzkU8opMdDKAFlBYVsNwrHXmFJpNAyP8bHjATiqbb4bH0O8Nl
9kS5y7hbULr/5nNC0PE+Y62ybcxkbzdFq9QFZVA3bNyOWTty5j5ewq1uk4cRWzlLCYMGOAeIbMT8
+GXnzxM0nIVbLeeCjXvFylI7zIx1hT/Lk6+Gp1H1+oIfo+g94c648r33ZBsumSYCHIZIg97gZZiF
s/o5wcX5kmOzrlheHXukAb+fKtmmOjqjcpCaqhXHRa5YJD73a7aBpnHNnilh/7DRqv2kqItqdSSC
fPWXJiamJBQKy4R55lQWIodh91ENNckc7uGbFWb2ujCW17I3RazGfmdXPanVThx7ZeaX/exMXlEC
IygYQRPRexmVffHXU20SyfcULeJcNLwdLU4/VGbkgDd9YORga+19IZZRDmygg101gCLyT2yFGmfH
Wc8+uB2Zy24FkW4NJCPYN65oElTqljyX+giG8VuROwH6FoTuPG++PlgSlUEzTJdsfV4PcXohYp3t
GN5B49GItFujjlzdWihFdmOkTH389csSdxtjAb1r+XN+RAiTG8tKynlDrQYp9xYiqIyXv9jEiKP0
Wz52at3BTBxGHJtidgcDvBIDG4IMNzeVWtRzNAc2BoMegNdRwR3EC/cyVOwWmhmbgHdZmmjG/+Fi
s81OyACqwE/CG3cG26QLOjKIX5/XnX4bL0IHYTl+22B/og1TMwdVTbabVz3m0oFFQ1ibgCUJpXoW
+07d602I+L/S3WZ62NHp/niDKCLd8ZvX7FegpHlaljWmw6mM6Z/S8hVZF74xyB/POuLG60zCmtiB
Obdw7BrGF2oDys/6b579jWe2cN6R5dxyKe8DD3YmIXjoDWly/qZpWOKM40tzW+OXyJD0nBg4zCH5
emvEcw6dZluOfo0VsMn8Q5B5K8cN4bxGgC5lTBHsIO3z5/e57JZYN+MvI5o6NJbAtWbryEzmUK5E
ZyJ98/A2KqpSux72j3BAf6gYKPyfcjU0VRbtTSDCgLkSJ0Bzw3Phs8wHenHK7vTvfPEQ5iKBk4mf
hfOoajOT4nYQZdP/omErH9ppU/UwX2tT13T9CqQg1VQxUBKe94VtrTY3Lc3ntiMdRYu8EfCGLQD9
U9FHQvGDWexYE6OFXUbIbDDqlp1MSzBs4hkk6c8yFK5dC+Rz9k7JcOY0pkdYtt8UK5cWgRSsWdAk
fRjNHyDQhfM7kOmK2yeDDJKwuJTExvw5WL9ds2Zc03BtJ/AiPLeF8X59n+8/jE9+tGto/BRxWeWL
M7enncYSPu6NKcWZyBVr7Qd7OesdUth6eBIJCq+VIwHwKjZB1UYt+0Xc/0BMf0Z7sAcGN4c7api6
mc+8Y2ifizsnrbzBZ+MFTZvk196aNeBLJcT6BFa1D/F4d4CJMb8nscVZ1y1iUL5ojVSK3Lf7o6LT
P8pWMN3AXEIlZJ/D9SOxqTNXNJdu5gbAV1OUsxhxiGiBiOpugZMsW8EPKXyFT7UYJWKZ7AEG3YBG
vHB+qooJZZrqpXfCfk3l9QLglaFDEaVUcDWPzfadEo653qibgbcXLJBmwSb18Jyz75Vy0Jj3e3H2
tg48B4rehGqtQbWMTLywPa9wVhE67Gq34se/qMFalI62tXOeARth0/MYVIRARzHtMFijwpJKvXYV
X9j8AQwRvdXcISHLOaabn2mQuBlOU7E0IeywF69nZRdSbF7y2i0GJ9hduif7WZl7jVGhFi1d7qwG
Fh446K18/bGrwYdJNTFZ2WPym9JlRPsAALzU5jGPQizPwOVxDil9uk8Em2O2bWkrXiTfk9VoGFix
tsdezN1SgtGCdIRYgu6Cv70rr7cfiKhHOXXB84tPh+eeir9VruXSKKKaaoFGZVrd6wrSgsCz78wc
Sr2EeiGDYUzjqh2j3+lcqGElUPKWKqz4AOJd1bJeVL/AgumsWUb5VRBGbLeJF1t2xU2AvfkogQjI
O7OAmVmVf9tGETf3/93T23XPvRh5bAVgH3TTpESCpv11FB32Iej4zEDsZG9JX79xZPvQip9DI5s/
9iwcSOpNpBbCVvGvwat5PrRbz3+viP0dRO8EgJhd8vVhLvVUFfMC3bOlOJTiEUVMO9Axsc9p6Xd1
DMR36nT5VJjA41FESQolHnDyrwmrTQeSbo9oPo0+F3WLWEgdwUEvlhntULktBnzf0f/GGcF5pOuN
J3bXcqBhVSL4Uz5U/vUTV4mYu8iMcfYN/P3pzkbL0mG2YJeITBWL5LLuqLMW4Wr+7yLFXgR7HQfJ
GBz1+NNhTh9fJ2voQIdh7R7B3ppmpNlywTPFDD/kO+6Jx3m7pvXUOFOpUp9oGYELty+2X2abufwf
ybR40yzqn2iZegX1Bxpa51V+j45f+VDFRxan4uafuVqpMyAcpnCoAag9XNUr11oDnQqgyGz7/I90
shZ1Yrz0+qtUJjNmHIT6K/ZOgN84zcX90Y4gPGjgFc4IP16yKpI7bX0p10QFEIAcAyRdsfNjW5cM
jI7wx6SxG8ta4LRIMZc2arT5+HREzkBMYFw20Fa9q0kSOnXV16DWxTj+2zT+t+WWWnY+fMe7tH5t
IrV0GBZCfbuag+Adp8EtSpTF84cdPH7mzUCbrMX1Pc5+Rhv6dLmkidrpV0bwHBY=
`pragma protect end_protected
