// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qurYq840B1gssr2zJb3gJLDfwKyamQFK6OMGyqMNMgqcLoUVZvbyRWHz2VJtbggT4NZvVhtRem3M
aZA9smAdFjLJkz1tGTl9CaZak1wicr5h3Jnmq2u6hkxaG0B28RjlH3C+Rn+y23cqaJWTUjVjuQg2
E8w8sJTN0nhAA7nSHD/EVVTxb11V070mBPyN+FcFNIm3cSqawq33zwpAYO2+LApQTP+ZWIOikA8Q
2IcR5YIIXuRkLqSG7GSA0NnuT24cWjcT+Yo8Lp/PT9rfM2hhagwPgDhYDBdtcBoyl8lSXSgRHn5H
pZmq2gYRIiYCrAg961zlttk3tL4Y2dN8nHx8cA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 28528)
RMtIWf45J5rtfyKYV1RuVkvZLGXjnXBh8m1iViJIrkwSuhJqQOuPyTk4nGplLRWTFlz2y5w8kvGa
F4Ro20Oc2YS0MH0AWkqFF1+JTkiPWhWWVZcXosDsJyCi+y3PwBgGhqPMGp0O4+LbsRwPt7dth9b2
aVnP4PyWglxf6A7kZqGnEjrNCidq6h72ju1MuUqX2kGeSo1XdV42yAbfQkh6UWEjyat3bLCq2Qqd
29XLUgZJgIbbMqkrZs+zdFs9R7FYtjihEW6HHKF9uRbzu/HYUch8EJ2F4ydJUzg6I5FbBh3b5N/v
QJs6nVXv81D7hLnCaZXbHyGXR026aRZY8pkGnZZa5PQ1Ywu6P/ZxXARTCX9Hp5D2soPusRF0ayWu
N+TUGhs3nkJEWmF1QRBC/LkVb0UDVlqmlXUDOU+IdAG0CXDlOIjqCe2JpdVjizaueQvqWaYR1bv6
Lq/8w+OYRlZsxdL+WaRg+VhuVogpidM8CJRQH//Dqot0h+8r7FovYR9T18lFW5AVlkpQ0FcLp9C3
fwieOMNCtr3Y6mkutYfdIvfij8Uckr1K6o2D93ZQzTS2uPANgKp0yGWIbOXeuT6qCxi7ae84feJ5
8IzvWRWP1NOmARKyaJ5KfLyXAvbDVEcpKoYxC4htNEhgXrhADM7FurDRwe2aHnmiAlEBb0/r7jOy
3cjq2nBa4a1rHUaHA9sQ9ouh0a0qUNemR2u3I893K9jQGKTYjlpzxpkqPCvfIei9wB9Jmr7t65VN
QxkI9RiUsdB9ggIBPH8TYdNLHO+T8Qwt4mhPeRr6pkJAEgLzGlRqbQfVwUEuOTc2agLbQfp38PPX
odBjxIINYzh0qDeGbLVYCANyEA2o+c5RuLlrrS8DQpD03VxgwYi1Y8mYWr6xNziVijxmh4UWEqgP
lBi6Z8blW1bbKMOGU5eG6BGzUpDIv49eOK3bjHXMrI67GDkC/BDbVnVCJ1r9F3Vqgm1YC6Ok4czv
Pc9foaNUozd3qsBdlL5sm0GTDo595C10b2OrjSq/fYLvOOiKPSYLkjjHu1OnhWb8/m9ijBxGSX/L
gNWptlTDGO0pmjHlCQUJ7EQmp/V8E2ln9cNecnKBAvgZaAU3gmXCDLpPWgzLlXIucX4jQK+FCeHN
7TGBWPq/ZAyBo+Ubgzpe29wwtb4k+KVHHSiM6efbLUY1Kutx0l/1lU4SgBCy/i9iNpQaNhJm80da
gcdNfxpR22R5ZYrkVlXx7A9khXBgdckrMOdY04045irubn28/noNAStWaQwsmmG9G0COQdYW7sJi
QyiC+mRi2IHDxsKj7F5UXHLVAuQ4v8uxDBrNzBaeeNXTEczq+dxXHg64w0OSsxDPEaknja60JWy4
Z//nGnD4LptbS57Fumx3cPenknCJ4V8dI20eW/L2A8D3fafdUJVMAsGDyR2+Z6EqtoWWqa8FEm/d
23xLY9gumok6sixC0EHIk1vs5UxOqNybZ1SkjfSkmQZwA+3W8onW9q+3GlHJXxYScC6mEm9Ncclp
LcVEWSs5gwxM6GQqImt2arK1PM9zrY2Rdz8FMcMnQdnwrtpcwujph+muBl8hwEQtDCoqSmlX3VXM
bY7aMKOOtyieG2x9I1SZAdCRQpN7NgS0g6KdB/8LhP5rT+qsohCOB21V4hw12fVlNHS36YoCpSyd
Nhr82qLRjr3rCHn4nPRaxldNOCa9xGAYf0x95Tpk70GYn6zv7l0DRGl0p/6rRMn6VUsr3LJchNcd
g9p8/o0fOWHhWWN2f5oJrFC/5cgqQtlC3L7ou9ePGbVBtXOvn5QiMxv6QPt+CrTyl6fs6VUQO2Hq
DCy5j5quE7thzizRU6aNHY8/Bq0BWEC2mEh3mV8bz+on4OhJk8muYnFRz91t2Y/GzC+DxD5pxJkP
rR9lyMw8uo66LMQfgOvMv7MapgzVE2liQYA6C0H70Fc/It3y97SQXg0QIwW0TLcB3YiVaf8H9oYv
OXe8mkmhXCsGR7Mnz4MYGE12Tlh9tQfOKDs4JebKjZ7iEwknwsfArNPlUDL7Fwb/9eaqRDVUlToq
I6aU4E14W1IGwiCi6oePnUB5wAXblDMNrYHeSxWWdg5FD7S7JMWMuGUSQVf3iDOIXnmHHDq4zJoD
l6PSr0at9QF6EiYa9x7bJkngtcJTlymi9h0Jr0xOvAwuOIlVwPdhL3VEYfUQLmwbDI3QayYf9zsb
h6Ivf4WhE7tFpMwcXHtUYlGB7mMlwVL68GmXrtDjw6kE9cSo6EcWA8ijI7Z9Vc3nFT4w/MpPrnNf
KMOqfWuQwbyIYs2q2dHK7VrXat3Zam60AA1dHCAubQnF32RxkapWXr3m3SVQSgkV3LjfBFc3RFs/
kozMf7AJcufREnura4nXr6hzb59QXzEOScAVGtC+gzMcJk2F/cxRMaSZKHoMBQH+wtt17zHP2GVQ
Dw1DmhhXsuLT2Wojp9xafSFEwcO7GMyX5A+JSnOEvi1P35tVulA6H5pCbaLQm7CtrYpVikRpSIf0
72Zie71qn0vBjaYLM8NaPMc6bStNqU+0yErNKznZkb3d/532Ictu7AOzRSoBMRtfZpmTqgNja/P5
Wwt5XfIb/Vs0r6gcuvFecAppHr1E5NNJQtiz4VqMf7TsGmDC8gPiXEYofBe/WHmRFEhkKkLtgeow
LgMyN6QyDUQq339CKFrM5xsbWaRvsFkGInkSZRT7/bol8kgpzkjXiO9W8j+SSXYyAEajeIGzuzVE
dy/9eXLuSNmfbkJ1r4wqV7TBeFjQXnCQCKGZRRujna5yZ2OkUq70sz9Cglbt7vmbA0UDV87meSoB
zVGv6MVcQUJ82bQsXQvfzbKIMFa2iZG9FSrEo55KJJYzzdkY9E4rs2JlmNVR5HOSmCRPA/n1NBt9
rtuBVHlHGQ2dgwU1EpFq393uMUgyneCkG/u/VzDzIKUyfVNxFSa7iF2oQfZQmP65lk28xZQMTsVZ
43tmsX81iTdmXs8GZQgYEmztcaBiLHc8EIsgLMgPExULWrgerIdHHTfUQVRPuuKu+PJW0rdZEtV2
pRxkR7PTG0UCoDKAE24oOH/hOYIB6zd1TUa4QkQcJspDrG85yGsP+9PB5Q/CM3a5rDoP6f/srNjs
wOk/VgcfBLfUtGM2MINs+HzfVQ13N8sFKl7erLQRsT8p77H+/Meh9CG2WQRj8BU6WwQgriYnpxRd
22bCTiXi4u+kNcQtaUgfihR6/B49wq4hbSe8FYPwv/ZbgkXfSO9PLYPZlZ7kVnJEJuF/mySC7oOf
bAcNVReMrE+Zg5hMr86/AXhnlU4orkEyXL7gNptHgawicxNwbkRGylkRRahr4k285XTWXdAlurnv
8tEdQsYc612HduB8tF/Jv0BhTu7qmXhe2q7QZWLWIu7ptkganfDRvnQDcmPSEuvQk22jAQdbPzyJ
DHb1WL/V58yVUE2AcQc6A0vWrYZPwWFKRTgsJsdOrVvEanPylkN91A8NAPBLEz7dBo5TUf2e/zpB
HoVjOGX6ZWRMTVTX2D9wTTMbSKQOFk/j35hs6Qle/fYaFAmorctj8jiKNzzi+8IkDIGr0vQYr0w/
S40gVr5BkZlcLqRptb4iT9h00M9HVAdzSGYMAFXxQRTioSZHyMC3Q+lsfAo1QbxTJq2SD3ZRJn4G
2spuSbChDn0kQrp+Wzx8tvRfjOVmmzYSZZxlT9ZmIbN0B2di6RDrf/mfaJt+KnLKmDZSW9LZCUDD
SHFXZxzRk2ftK8COSEazPydS0N5d6tF+8JhKW7AN+niIkM0Ab0KgdofknSRfwWmk10YZdDOy4/s6
UigJ+aV0btRQ0FLoH6UPGVK8emZXfEIvdJIH7S+L8LOsq3QsnfG+1k4FRsLECeIr/CGxNS1Z0otR
QsKraa5VFZnj2/8veiiZSkSofq3iQfYgjFHZnuFEltKX33QHMrbgwWYFdP9RbegUiGbpUiwMZdKW
MS/Q1op2+qBohqSjo1jtbuRjU2FxWH6PMfUb2qGuvMwZANkk/67q/yCe9o63+2TvITEIyPwbEgBJ
U8lC/R6koRcGPajX47CREbLgoFZsildI4rzhdIi050BdlsSpy1oL2tWKjyy0MpSAQROKHSTUWyiJ
8c10fIxrWr9/x5sOLI0D3eAf55QO37HXUTVno03nLl/bqvsq+ZGzjC24U2Zn1WB2ufXSm7+7DXjU
6Hg9bFB/rQTDfKJz3i28otQATD2WoJCVgYPg03eSWETmEWqAzB/daVbg3aEGHFpLNrSSiO6H17cY
qll4Ujx/PcTzzztNNPe2a5Qdta2dXujPtBDqQM6Ms8SzxowDYTBS29K6b7MXIbJWAqYM/UMQy8Bp
njsyZY8mRWKA7RsyEiu0nmbiy7vxihYy+chCUakqd1styCsqs8F9xLnZaWsUJcTP988S04MH/0Wq
k2LEZBFTblw3ocr+pZOQk5nmAPExWMGxk8gP+8NSEC779nuR+6AuaMidcuYkGzcC/Sur1awjCEbU
LwdZgwzp06dBsFdR65MdHS7dH0CZQhUFUVj1pdbaglgf+X4CTN351XWr0m7lb/eLaIrK1prnJX35
7zQtNQm/z4WvnAoGr/jF0Hqkais3oydjp/H/H9SGKLkIELhS3BfFiV/JOW4dn55GLy/W5meqv+Iv
0uQOSFB7b8jfnKrarQjkzOsb44mrVEzux+8rUaIk0tFfg0A1yqD67kNskIgQb6vNT0Eg9rhY3+CE
7dSxhWQdr8uQfPF1SL2yZ2seoe3Bi7tO2VkauxsbQ4Og87v/rt6C27GZGtsOk3PhaGk3ouJ2zYCN
skkpbwGbKDuWs88qDB51lDNt1BEKfCShl4q7uaJQWLVVL0mjL5Ol86xnIWD9a32DEoPTj12dLeyZ
fNQRZkq4IPZghfDQfF9/OOuHFln97w7wGYDo8LesgQRrsx45K7tKj+0kwYZ42GgbwTg/mZQjdWrT
tCh1gtpWf9oInct+rITshwU/Pfz6jrYlxUiQR7y84nERqEFtwdLh1x75z+LL4A+pus3SjtBpl5oM
h6e4Mm9s7Fnj/PF+pM3RtF4BXnfmCPHSUrU7uU4LuP8esjR8j7GtECnRpLCa/M1pbM6puVkpu1xn
G4JCeBprscfosHb+rsdgmPqwiOZaZN84+ei7SQV+U945f4Eaneq4kMo8Pt4OBo+Qzr3OdpfTUthD
B9pyTjxOL9Dvu4qiofefUZofXnPPuRgbItERd1rr2Tqr8Kk62SpBS/ORADD7eN7Od+mc4M8BNiWU
tPppTZOicJHfL3RcSjYpxEuSiOY9kJOTEO/pSbQU1EHFiZn+Sc3N+L9VokqzC6PgUVlrsPJN93gf
pfOUxxyNK5dCWh2mSpRg+SBmnYw0Vh+9nniluSIemPARJCHGsT9tEiawz/vG/XN364FY+WoE1fHu
yfBPnNb1665lUmwajsYQz9fs7fMyIWQmyKCt2JcVkTwOaMtwMjtiBH6ebW1cu3Qr+f9g83Tj4kGh
7moNFl4K8Eoxmtpauyxb1gRkUJkqrKq/qCa+JcWvcgJRS96FIWR173XLXh8ZK8IiDCAw/SVVIVey
0ZudrOAU5ZDoGO93hOH4J1k5Y/7Irpbi8RubCKyjnA7ti2CozpTh6wtQXQOrerw+8783H7G+D7Al
bnFHkxO3Ck/lsn134hkm7Ob4kScAzyk76l+H+JeZhvHL4JJErtkiVZAyIR1G+34cO5tFL8Y2D+ZK
xywyw21+VN/Bf2AdX9a4jkbTo+LDYNqrjII/l2o5xKr/G4D3JtE/Q1euiv+0rh2JD6HshAv31+4z
TWK2ywwtXZd1k1b/d7wP8qvcNhbM5QzEAajIo0w57uN1XknSdEBz+Ed7GV1JMyOycj4RCU2QjKbP
OZxkX9oRXrCSaW/9wQn7wAHEODJKMCqP2RzMg1ReVBYnFv6oa/cITB8nYd92LJ07ZCMHDJmaLJe/
I3JO7AEJV/3QAVg7WKI8b/F5FSQS4PTE5KS+GXojneFZdbxuJC+IzLbfiscX+XjVTcWurXF0pfgz
dxHog49QrBZ7kDLuAyFEFlHzjzLyOtKLYnZAsNINee4rll8T6MMo/+2eaejIMMnpTuXWAjM5Y66V
0wX4nIBp3rqXBrvv3Z9mzusXZ8gIQBWlhyuAtXgi1pS+cJHRaYMNBnBvnzqG2UCTYvoAF7/BzWnq
X/kQXfy8ISIgkbaaMmArAR0GiwKLQjD0/rIPQf3ShZULTskGO0InfI/KbkyIK0Gu06sxe3Skc0nI
xmlNwE9Ivx6AwplhhQBtmEOgnP8+km7Iib0Q4yMnNbN42wlkIWm4/GKWt8ZbFvjwQUixAwbt0e+1
89QCST8MtzYHYpEbkHG8NOR4QBO+2tnNloUy60Erl7sBIuEiAD8QRR3Bl1jRhydehQiYgJJFCv1i
SbZvOXjZ/mn37xwzNkAdzTHxd2lyxhfen7mmgGy8Ixz5CUNNIAjd1AijO8HBKCnwtuzQBv2N6Oo1
QI26DaWy3wKRn2QiNIha8bwdKsKNgMfKqGAxxbTZ8GKc/6Ap2e2QRdULp6sjjrDQTzfiyllq6mhb
8MuBdNOZx9y60wTM0U0sgWPEyMG6+a+LjfF3eDY4iGqfTzBBfE0nOGB8jdumdGJNp+GDBxAZgBby
jE4Fg+S7enPRzVLyHO5Wt1Ri6VrpDG1PN/kIH8+Jmr18hG73mJMx5PPaTC4L4FwxYsnqttFDiiKN
qGWMJFx8j1VWYs2AKxtMScgEwpMvrQbqih3yGKLXltXnilMxsWn59Veh4vaD4pMAC3gSh4JSywNB
A77BPRn1a4+6XvCeKPX8rjvzCaeTAE5Q/ow+aGnBqwY/YMQ8i3bsrPfTOOjuSwyD5I2LVsyk2pFm
kVHuAgDP8rOEbfW8VIh7reKMt/XxGpKi9k+M9NUqIO/fTD0Kvqc5kzMqaf5sfzlozTzF4C2qvmeM
Ww/Pyfo4CsQCFQAPPSKG69Aq0abaXsRXVW21RIyq7wMV5rOr+dJ/zDLduUhajPWlNcPaZT7KSRID
/O/jyVTPdCOG0zE2VLEy8/Q/hnzQxEwe09bBX3bzs1djD6tRbwtngbCqhXoS9MLnol2TZidyPA9V
7Quo9NDC3DxmOqAcs4SLGDJMX6ftH1/fQBE5+9p1187oyemQqNQp3O4Fd5YN641y3IVwAS18qeB6
zLRnT/eqNFNWJcBG6OuYgjNgjKS/17ZhjRWO7hJI8F7D1CSHUTsDSYWknnmQVftLtxKlE0VKhmTn
SR2Vuq2MBnhu0Iyky0PmyAiC2nyvb5SYYZkux/mWvAkj2yq7yIT+w+ROdrfd/BuAHjQdVuyryAQO
KUH6cciyzl/YQvr7jmQmnxnKrdTvM5xOwU7hJyw9mCTAvQ4rScKymOmSfiDc/VLG7Pb6C2VTBuZS
x4+rNlX/iUXd6UqODA1wXPjFeWJYWEq5OSUtNwiJTOVDSCs2t6R7P2IhdqG8BgMuIzUObB25bbNe
bwIE/fObUtAYBJiIfrA6bWk6zoKstfTXMBwKbjQJQsuLkJRFnj+zEWEkvIHizyXXPPQu1PmTbXIR
jmWnXgFP0/ufvI2/CIlmXIdHj+9R4Spq48l6l1yVa2WnqVta5OSA2DpV1O0KWsEZT+CE74koTqp9
B4X3vPZdqbKkozegoBDCBvmsFG1eehmbK7aEv3QQuJE2QlA25FiZuvkrJTYnGclbF8FmrMoYQ6/c
B8nzioGpWOaSbV+mMArnHyCY2jOzierwn8Dy0+vWZ9SiO+0MMLRGGdfayjc9WS/mpCy3ad1fRX7S
sUBn5kTx8cFLeI/fFv4QVP038qXI1aHQAxpIoanAiyTgTiGgqJGxfZZkgW2vLOFp8qgX8UQv1zoS
pDEWYl/oy5XEM7wA3nu7saw4PzDYCfziP5EwlUmQMvVZtZy+GfODdDrJGR3Tu2BifCTivCjFB5nd
vkpTaqF9nigEnOQmfqxHvUqW1Whbl7EmbUfS358T7tLO4CeJZwCghH4BpXneZinlF3182ZpLYy+h
wzjyPE5xzv3jhj8NhrD4+3UasxoCnHJaeMmM42IrGtCwQlCpIC49RfattGuMFO82vqsek2pglIyq
ZNCP3LrwVIZ1f+MN3tU0+sKCpMMxHswyDeCxLoPiK3xnaytogon+pcqWJo892E0k0rpvPRv+x70Y
NcXJAhyVssrUcm7OqbOWZHVBieO/mpR9pvjC2syzfNE7yg5lEXG4hiu6ZatUZqslgoNo1JFu1BbJ
eJWIKxVRbeSX2UA0S71hcZklcMxDWjdHtDngP+JJm7vlefFqLEgxjskshJG9GemUj80jBvFRq9y1
WX8q9iNqmMDCu/Z24paAVYj4qkwq1OoSIJl0m9AFBvy34YlPn7bInbo0QmStIFNoOm8XhSA8NJzI
gKD9c+3ouuRPGtrR8XCLCWUO9ludt3qgcfZyYmaZCEO0BiUMafhLwuQDady5+fbnarR5/IQmJEqx
ILw9dWh+QE+3KFvGUEpCYLeCBLzXRN3NZEpuMLUH6zxgqNSf5UL/WJkf79YiuQ8lQ2YRmlJZwTF4
9Qln63AY8FvsM6+Nk+Dc8aQT5GWB+lblGFdRfpJGBx0QKnkwLAQzYKE5KYsaa37ArRiiyqMFITHG
tzXZIZ/yLZP9UftcTjTlH0Yw/nbF1j9hcTCHjMCVPUUW/AgaCP7BVQudPSBOwoVBNulChoVc1k3R
O1rHvUs/HOFqH+UQ91EqwKGm/qtjEVV4Buh7gHYc0zLSuuabx4dKNtGQ7kVK/s1IvQ6pwDOpPy7l
nBI05hevD0V0c4ft4KiCXaCZLu14XDdWIDlxkbzKgqAYAHm2gcu9ESGgtJTTU4IWkCEdy+DgsHlr
LdF0TkIoQnqOIFjQW+V5qo4HQxmssx0tpswZa3anjXkKkWzrSgiMsNl/Fd5qYN2WDUZ7emcm7OYX
QJmUpRepUtBfSq9hdujyPsAmDYwdPs4srivDp9dljMWz1wwvGXZtOs2SsNEvIdLFMqC0D6meR9Hy
/tXdbHi9sRqKh890BVMG4cTQ8bSca6TB4O4b1dlVQ83+zYtVtjQc6qSxHIPBl4ACxhvqJY/RwlkM
cxPMBe7YiUPWRPF3wl3lMBtDcOaf6bHzKriaz0zu4vqmOkkAl+fLLJB7Ya0xXyWeb4Hoe4Y1p4o7
4/3sgR9EwIbjmWWj9eJUe6oyZXdMs5FSOMl2vdwMXiP4LYJRgbi67Q1nWRUwZhwVHcmCTgOZUu7K
RDGLbTcKSurBwCpjiKICd6716oA4otBM+T0SY4+pduXlzab19IdXaPFaAURSfDghTgnwd3a0WTVs
XrUu7g1ZcbP637hz9d2kvqLR6wVGHDrWXhwG5H4g6neYVkPw86Lf+plaPhmtzQBuUSamzw2SO92t
eWaqU2izjgPFUeIb8uhYnD5hlonEUpJxoA3XLqfHZQPHccs80Bn7Dl/bdP+Avkjj0uMGcMq16W7g
y3s7lu4xSOB6eo9vrRBzzU2QTJFqkypD2pHgh4K991dbcL/T57v3JiMsVm+2yqXbnKysHOA5KJEY
llXcZodAJNaTF6dh/eLRzDcZB7a6MtzFCc/1jptDMGYUYJH34U2VaMh+ee2EzvemZdcYWMW3aUuF
QQrXRp/+5r8vQ+3cpeYjXyWAAdBQ1fnh8tupfX0kggtS6b+od6F6VkMvqH2j2dybBsoVyMGqfZbu
kCa+hyeS7RRqy+RllQvPLhbl9Yw6u4V3FMVbUjvWQSID25OmBm/cet7yLcmoxkzekmil8YS7dmoR
gz+dwM3mvmAbCFsxMJupD3QqH15rpGhi+NNt2hreI6WG4TWxT6VqKaCc6DAtpKqq1kAVYOxcFkJe
id46LEMTVllz5xP1wiRDA3CXBzoyKH0XrASE2zBq3Ds4KUuy3EaJ4v/aZaKsYB/Z1g5nLIwzO13J
fvscdJF4/UnfEeYNUB3A5u7oyzTHba1hjp8xvUfqXLoDyc4oS0MtFNxuYOCs4HZ9wijqdyOqRi7O
NQhcERgYEC5LJLmdtb3ro5xWbyOmq2LKoLsY/7xLnZNV8HwAUUJ7nJNP5iBLWLXyCMYAH1A9pIIV
rxLTAEKOF+BB06k8yo2MbshhWHXB1IGUnBk56Xj7WEvEj+3vGYqupHZu5uw+Vd4OCu+0mdpl/68U
kcdEfwrVkGQSfvJhTs3zNPbO05Kn17IL/L4acN+bVX+M2D7JSDHf576fngByIAhOqgMKcVxPz3Pv
Ffx+DANyA8ZGpFFuXpGI6Ua/n8sKZI5ffqo2VC6mscJJ5oFDse+BYK66VDj7EwMgChesD8NBmkyM
PbJ/0lZTfay9RLmPnex4cyFwOPuJfbmlXDdnBD1zHNYgUwiajuZiGlv4fMD2Cw6CoDkEhvoai6Qf
zcsWpN4O27yF9h2wUDlHGzW2MdqIt/p5dGHpgVxlwrJTLz/7jEeJSIJsiT0jHauVCUDSE/XEKOUp
MA+nwnjOQrSxDHhf9eyhJYbGQzYP6eRKtSWJO6TGQ8Wd3YnwRA4dG9fmnvnFMkmYIs0v0nCsqt9H
Kwc0Emg5I1gPS/wmwF0VcL9TsjyO7hjFHMEBPrR2icvJgEJelMsLq69ZBT9I0BTgO6RVoJ5+dMIF
iy5ulMFTV16f1fWRGbTaAjisTHFGihgJHadsyLiTBnB76MPzdd0MeyKyO4vGwMMYMWIFGX8sdEYU
N4VaNHaZgLDfG7p6epsbvteIyZbpvlG9yFia7J3WSShQ9CU5CCMevKRmmt4ZHcFTidO7YtR8094R
LTc3aVbQp7+hTx6GG0fiFugLj0fuT3A/MzA8//uifjntq4BdCqeimpmSY74WEGC6h+5kcw2o+4+g
Vl9yK5LXbGWWMzynDD6xrZ2sq92x1jSeCJpsJXLnrTB1VZKZU2vPyhUGn99KG3xAs7vbOeZFu8HV
xd+2WGbFUoRRm4nGDQAcAtEMerZV7MpsgIiWSSlWDu6+KeUNs1NuWunG9638aXDxUZtZNJ+aurrJ
mICJwG/Igf4y0eKDqfRSP1brEyQoKzvmoJIUR54zTBzmDbru+Lsdq1OWCAZfYqPxAzb+DifwoHX8
mIWitQH5fwqMI00RNSllzRf+2fhOBoL3UANvRbftGbZDjPt0OVuD9TGUp418JGJGWdFeCxA5aRni
gbAaXoIVnO85tAMt/AqMzOdnjNpJOazmDWLKDUqRyKWuCBgPNL843TtdZ1SJLcvU3aLPzpJKTGcO
Yu85xrjuFbNOKwqwN1kYn7CgrGgyXp+uEWMuPDvfUnMhnzvXuSGutrFTufZEtgb2M7zevQJsSxFi
+3nJ0xR4Qr4+QayUzcmNc8B0/Q1V2kXDVewwl+dbyHfFw7oHGGGLazw2H6egTmALClJKZvIQlhz3
U9tlyIKgf3Z2AHfqDoDcG0ntZd9jFuL2LTGuOXtIZidppe1dUfRu8JJPd2l20CC53r7teV1TmwEq
5inD6bVwc6skN3U6T9NX+gKIdjeKR52d/WO08v+MsAWy3O0noa3Qlg1rpM27Qr8I2smpM+NJzkMN
SoFxiAY7tHTvw/kdJhApzwHbgpA00jE7BRPdyxQ0qrm4QOkzIFaC5xM1Nss+ntQ+kp+0qdBnKle4
hZj9+Eiv5YQSNrw6Hxy9pEccdHGyqqN/ocnd/nQXmjhru8SNweGFxCYXERxs1wzdf9CCsqEgjndW
2mCY387/6r1VPrr+fT2VTUAfyzPslAP6U2Csvs1iNGdlgysihf/gYtW2ZXemz+Dx5yK95lR4tvBO
M500sw87X0HRVCYdHpKivw99m2lOj8N9bEnsihaOULBu4+CZXnwa58DXoqtaqMPpP7B1d7dySrla
bO33BF4OmxKIoKbQrTP9mBUWd/KZIRznbASRzSZ1qi4+lH52O3YXBBy8Rf7b8ghrBLB4k1LPd3/6
LE/mt237UYJKdymYAo/nR6UrunMNbFbRbRR7XhWpqeKf5iwoRu5tjK3QhTUz2dNaWb/M9dJ17Qfu
82JDkhPZikSAl5ZDpL0Fun7h2l0yZZuLnCBi8D67i0tp1Za48dKlWNX1insfrVSZmV3N7pEPADWE
9jfqEh7Tz/sHh6VrcQIGYuEpYTcwtOD2oeYAtL2MAkiJXYtxhsbZOVZvpISqu80ZGBtq1sxAiOVg
b2rcDMa2lEvPzsLCuFtSgy/sTzrLcDpoojiFKia730zVVKnnm484SZDF/3reZCqHpzzB4xfIrocl
0GXDQnBADAdMFiUd7FgTm3iwH7pTh9Aox1/2+xAnVaHwTItx5roRF/WU5P1Mk5wFKBStr3RdG06f
ht4EMJBZF4GWO9zGs41M/uH7g8c9Y+4uNKIF2nmofxVqnb4QkHNu4TMCBj8zEyWOnaKa+t3UGTwz
j+FSJHB6emw6n/fN0FTd66YxLyAYoZ010e5hGdC95U4Wtmg5JHbwDvOlp9BZACT05Tflr0J75t/Q
0LfsOmPuVisUESRdGqSswEd8+LM7CVuYuzom8jElCTkiVNdxyczfA7m+QNK7c6D13vxXPaDL7xv5
QILq6oWzdrnsT/4MN59gkHWEqxhvCjS+QRjRr+FlrC1dKUfc+BeaID+2JYXjGEFvrXegmiJI1mvm
yMPALRUHLIYE5GvMM5Be0qJWt7bSldryV6EHmDfAwKKOE+iasEeLkSsmVXXrQwT+6HdgSDjEPLHJ
xdqM7E1k05DDoODjI4WHtWF473X2hEJrLE4Q2pR40pg5Ppy75dfxF/ib9e4MzZwdE4acwyMT+qDn
69JvbPEaZPdSuuWko9AZHwkbI3jG50ROIqiMKAkse37K0rkbS86N9h6ZVisLgUG6sG0CflsD6543
hcw1XhPM7nhwSW1L2zK7mq2QxzjWst36t+37LwBNZVsQRKvC4jqfyiS+5EgC8AOBo3tnvg6L8mxw
Lwfl73TXz7TmNUJTtTnMguBscMGVqHrCIgnOX32B8klXnSu6b0EF+Ah2sUrvtf87LDFlnsQWkzOM
oO8b5XCvpeG4RgWSUEW/yWOabYxA/oXUZZHZw0WYIo/53ULlE6Bgdwu3+vfz0/VYqfSj/MuvIeJJ
KBp6ubTwGtBOetgSQHZZQd95+JfH7W2aaE0x8zzm50/Nm9o+IqadgFl2MSCUbY11p1iBUBy99MU8
1QKchyvNkK7XrXEJF4YcrvLI4UM6mxCxubvGEMWx9x016hM0i/ZUlLPvhgLtdlQ+ZBw5uCuU4C8T
CyDRNxo4QJ5r1MGf48O8Pb4JSMiyWiNAm1r5J0FCEqLrOwQENzQG71TB1Sve0B+gCifPSeTHJxBZ
svyy5C7NFuNeO5vk2fSkav/Q8XNW9mm9Kn4JpJJHpAhFwXRTDxpverMcWxFO6VvP6ELr8jPrOulM
KD8MI9EEL3G5gR4eY2FiIxnNKbLkJoJkyv1dcYq4OkEmnwlmTnuh4ho5sVqf4A0IEMS3+KxBlYrI
gvtBvgC9TRZLSoyhTBE5WCnD3oZarKth6xH+dmQLMgactAcDOFLXyCRf938oE/X+7Yt9ESuXJjoP
Yt4c8ebYmVUIzvU/77rPSSYpq0gMPMMllcML/QH66i2MmSQ1ZG7EO7mE8tOdee3f/qT7VqWnjCmA
EaFUKbnLs9swWkyUgFYQ6bHsYF4ki0XRV87QQD+AvPQv5sndijqd6WSn192xECIvSD+T1NqjHsxA
po0sgHWMkjevM9OeLmx1HjlhL6krAq9QJ7XTwbeAsv5VzNCALEeTgW9ZN0GtBZ5fM0rF+M4n7ta7
H9bOMnPy4KWcJWuhA5KCcOE7e6xppnQ9T12l053dP2qpS4MzKlOAkS0QL73Z2pKRRo1I+XctJTUT
vPCxodhywBfzU0kB+4kZBXp4mlKFio/qmgHqNvTYoUgcZOVl/9+/K15O9UbXj3tCF5iyjg46Icmb
h/pzf2XHbVFJJ/HuJG9noyfINKdmSDtA/3zim+uiXraR/BV6MmQy2v9lzAizSwzx/0zHzgY/20sr
/yOMJFa22LyLhbA749tIioE8apeT4PRe8iJ1s7V+OrMlybxfpoHsE2j6Gamurs90EMzkAU7EXCOa
R6aCPWyfLXg23f2/8oFiIAB/9bV0/vxNynsWbVxwK7T52Sf9xhH/jI8WKoLL5d4nF6arV4ID79OA
QqD5mlJsUHsp80HppchhVEMMVo+3jmuxw/ccl/9QaWXcDqIrWChDV0+G+Y+Qyul8q9Zqc5h5wo5q
H9Qj3RPKRwENTxrGc5zdxVcnlnEBSXSQXGCnoenwfnEmfLNuALjC4kxDTGgSQDhC472qcrW951CI
ftw2bnPm9nIfFi5NHDsPh+0l3RA7/MUykeAMLQtFIg+bgGJEtD7xo/AxsL1dhBJU1QAu5PqCEW9I
sNuRDHJZxYoJThPHWRUsVm0QHUVfl1EWCBUIEkPOo8tPkagKqgvBfHgLITinzDvIXJeOeg/8fifb
hBycQjwDO1wTUbFiS0+TrU+Zso63H0neqwubC4SOBLvty93fh2xa9Luu8c7HseeMKJkmIBJvwtMH
7R5CQg8m5mT0KOY24q7jcaoTvKzDkMPILjYKuvEVyPWVPpSJMcEr2S50psCHV9kTKq1QO40bKSqu
vQBEtBl0aNooXjHh0C7mv0QbycpGSvg8/tMXpCpmnldkHzhz6cc8Zj7jcbwWdJxs1OcKEseU7Rld
t/Fcf1wguwp27QiM2O4JZu59VLeJQT8wBr+Szdks7qmiHWOBYDaXPnA4WpRu+Or/xwu0yfQqpbtr
gMN/ItFWvPVvwDXMUgaHGJJF6WRteiXRp0hm729lausZNSlt1DGRMy7cYlGU+Di8ZXJZx60XWJTq
S1ZTCViGyxqOTXGz4ycV1KnLm8Vs7OinrCSmpQXISzvttmgPfJiApoPDxIRIXg0jExABrRG5HTuI
yAJB670IOWmGOc7LV4kEUuF3c2y/sOJe2ugDruF+oTFFuR+m0LDNPq9Y6fEUNXSpcH81BNimprj7
21lHfZ/HZqeuXc/l04z8494a5iWVD9C1VssjIQMA6vJxFfYoDqYRV6AqVOVo2xcAhgXOKPVIfuwY
rS3QKdMEFxN2PzZ7VoaV0LcR8W5dE95I9i+Iu82qRKBOU8tpA7b9iJLMQGgOGhoxX03OgqK5nvIF
Lz016er+avrSmhqVMsTOOIfXk6H9cDw08L+OBwcR/NGj1pLTee6QbVozxnSZlzTA9i1K/hyOwvYB
BILfA4wRDm2AP+5v7DoLd70WecJUCZ8QcDMHyUDrwW3YNUq4gLVXVtMJXFqqzWE/EOOfsytJ5A1/
gnZ5OZuOuidl3i/7mKxk6B23I585rH2wvpuxvbWB+ljVUjNn6IlJnPgio1oCwPEWKz38gJgf0mPE
8tKaLEDIdxel/GMoaGw3PsKEAcrPNl4m1F2UYJC262gudcvdzAEGio4AuWAWhn8vjksIO7G+YYBN
ruocuejFf1ANtjBHnw//zGIh7a86M97jVh2XJRUmwLG7qsJ5rk0AQQ8ADSXXG464LT7I50nvVuxW
jCT1KnZq5Q0Gy4U5Rr0E2b+WcSyaOSgYu/Yjiikt0tW4191s/GxCucHqxjT+i/9CQvehxYwjL8uZ
FADutVgS0qgd2P4wYn7qbDgRIrGQgfNmGxUfD+srjPhjtZVhw4wUXiGHoioJpuAVNgTcRkXror63
RZ4/CEtwGY2m7C2P23AX2oSM8g5V7t03JqLykCHRX5SiC6t3EcvnsE+9cDykw+SbNpRS+dcuEziI
aMvX9ruLWoi5WX594Auvb5QiseONkVRwHF1aB4anL7aZe823tJjpbYAS7jnb+AJQdLtAN36eZDpu
2TEDnOsLP0AOSOPKwlynk8PKwtf/BY7635ilLhzzi8uvayD4bayoWSHewr/T6ufO4qjk7/Oz8qhq
Ac3EXBwvp/bD8viTiwxrzZp1V4lr1y9PgzNPBLPIa4wFfGO1aPNDzt+0dhg6DDZHxGpLsn4Kb3Uw
KSFycFmfbov7Za1cl7coYByyAkRyk9XcLdevu62Kc8Kwh6hR+IfXZLAo00zlPaAxjCuoRf+RrbZl
8fsl49diXHQBBUcZF89U30UqNc1r1mESsmpoMTAaI0ip5OCfjLzarSsO8gu5jfHSFIalVhAwdWvt
ilw/p1EEr6kUURptiUc0pTWsQKxJjO1ZHchKn17iQWXGxKIZBZ56x26QeGX/oVj62NJ9yjwBt8Ev
8neUzgeoEYWLy1S6rzPbS//yO30z9ilNjH+YHlgl5h1cz9dcSLZfpQ/RbRX4i5FK61u/4Ohruo4S
t05X+5SycipvxPnfh1fPJb7fZ+CRh9mIhGeSzeGG4znXQRkS5ycGGC1VY6YnTrOGflNX7Gpr/KDk
zLkAoxIFB0IXDt9njoZbu+GbN2JhnwWge3Ad3gPdtyLdaisdKLddsDM9gVD5WMoGiPGPbn0Hlv3K
yfIVbqG7knrrjWi2wZ8LQRKSR1m4+QvQEhXmdritbt7d+loAhgfrZypWP2WIt9er1BrRdRj91iKL
2KhDS6cblRFSYw2YhEAbobeuN2PiYYAucGaZwZTrn6OvUJsJp3KS4LVnwUTNgpp4jKUTE21tUrYs
0YKaw4ofUV1n9v07xczv96r92/qMQqPKMIvibdQQm4WwEhN2M7BgGCecgYjBCfhJz+LhbHeGiqVV
yK8cLutqg0601ewq0YOxDycpkv6B7wHVWNdVSd4AtzpAWCrsm3g148Yo+G/6R7+jCYxZHqsUuOTw
0DFEzYbJUKvHTIt5Ta7tg2cSRVKXplceRjudUNLyL7j6FJZnpANqEcVSrCpAWxylg70owlu5QAFf
Y4Ta7tvb63RkTOfffLIBD3I0PjoI8NPxoU3M2Jf+OwT3iNLDl/xVypJGFm4C83jfY+As4FYv6LMG
74ALVZQatVRbcXb3UCIJE3aHUCrA2f6VCa+phKUPosgvnZC5DJo3UjWNB/9FBqQcwaZ5CtKFvhfq
OJsXlTdfUQ5nIjY5C2KDEKAfTH8d6rHnTZZitxPi1ik05wVkH3eSmmJkjMYf5/CYtyFKpCcZagXg
Om0XUaCT3YalXvdNl/jOkndcyUKRdFNNH02TtHT5YS2L7t9dbJQ+R0PABMQyBOpFHtJzHJaLxp64
7VJsYI7wpEwrWcXf+lJ5YbastXAwL8mddumUCYEYl/2Hizs8FIl1f2hF8tihxSjEY8rXCz+BY1Vt
9+jdRayZAbsoNFF917YqGz8egiAbseIO77w9ggXhVd5MYLG0SaN8YS6OA9PPluIJcvVxJI58QWEI
JeEi7DX01q9hUcrP8UmpH4bAC4EV3YpFIGNvauNRupK6p5MKxmxSvxt0XyYGXNRs03MN459SSyHR
JCMotoH6906wDAEUpGZvHlZuhKEjmojdWFZbynXvzmrYYAc/6ZZ9u/MHsGthfPN/ge4pfC9twmTG
NJnHOnziESEI9/VjRvHvTqfYhNrACJ28+33Yub4bxNM2OyYv64F5FaiUGVTXcC2L3VUbxJq4E+wZ
9Ak3yl71z+fF+wx4i+DUCORBCfyczpjgwQwS3tvgZP8uNzykquktXvkteK6nJDUTmv170yfc2Mr9
TmVxyrERriS3seE4h1WbXL9OJS+CaXJw7BUCO5WORm2awVDwLajCgZRGCbIXZZrclNf1vC11aOHL
pdTHE/jTLVityb2FhksVVJtU+9ErbiMOQMMd/I/RIniKfsaoEkwmaKaW7RPgI/7eJuhl9UUHGe+o
D9i6mVwx+omytt9KIOWMIlWZoxdOr5W7bkRd+zYxKFGTxK4DBLTIRShCQ76B2RWc64rJqQsOlC+5
Rrk2yQYFJ9+qW2OsijA7IRCozJTZ3r33agDkv0e/O2L1LqUiWbUdwMjUpMg9rR0n9WjXzBhrR7aw
m3sUatq+veKc13WYGuKHHMW8kijdv7s1hzlzOpBPpT++LBh50scWU8NInagSz6jFGG5/hDVR7XwN
Ma6kiHceSgKFnK4+zR+w3nEZs34W4vb14eXR6PIN7Xi4NBbKyECeMOGx951kR9umoq15DbO0vkWc
6nAmuT9DuPkXvw47lll4t0ns7goP8aBk7RN2TS9OTSULcmBSbKepvAuCCXoSw0eJgVlULREvZBFk
uqQnlzelha7SvBrHehoblgb9wH+ozmah+Xx3j2V7QG3zVyk3AjYMDvqT29lPGkjv9A2e286c5cbp
Dx76uTTWaNzvqtSrvMmVPqtpSPLq0H1PmWvwE1Qs/edWQYsU5cB5zbZCAEZ3CrQr9GlkqPXSwJA4
AvnmLLsTwLBuBVr42ESTiY9rI9xcJ+j0kc2kz99MmqLcWcKqLTq8xMikXqkyeB1YTHZP0jcBcD0b
efOzP6yHt/oB5mO0K0NLMEaPHkpc6MqnKE6CniIMMDvHMmOt/DWgK5zwTwPch6d7OlKH6NpZX7BA
oftzQ3CEVeW6Y9W8TrGaDSkxyQ6g9JPL/WSsUylHLIzgva+x9zYoy4wjD+8b7NuVjHohFMYWNYLO
ZtnQPN97MT5O75trpNQf1yp6mw72Qmf6YiwKVCIRrcrpVGYDNM1Hl1gDLjRW6PYSL3gpwDlqFxhj
5N6L8N5W0YH/P+bm67upadouSBgAcGackrFhDLEsJ4+Z8fBWqzpvIh28rOo3j3rNyEE1k5HTt5tI
SfVEdhujZuF2TlXqHZR2br1fdHZHpZWaUid1QRo/rxiRmEBq6ZFSq/Dws1U/BAenurJu4kVAR/Wj
VQveMh/UIWm7L1zisiB7uHgbT3o+K3V23rmticthaOCx/Z+6PznaP4H015XeOsrSFyv2vMMXM1gy
lKZgHXHWtXxr8K5venIjtzu1FSv7/svo6morCL76b9qWAGXL3g4FdSx32HHg/k6F5o0vj5IWdeXS
g4L5DTVPzNQCgYicDxJHD606ae2H3uU9DWO12VbgGVC8rYcVMNSIX8+zyYuJ5Xfc3z7KTvK8agpV
037hHdHgUHlyWZuXir5KXtQiNKYjEctggmEly1cZRuMTuktcoNMn+gZo1s2pObkM4E4XvncwU6T0
eAfhdWLfYZem6HGEl/ua2xVfKdybQ3UTdScG8FTvHRYl3pNR7rh8c83l5DWkOxQANl9WCwfrGORN
6DSpxjmN9Fwz/Fw71fiv14AHa6nQevG3YYv8jbO4FdfE6H7TwfFVufXliXo++znvmXpF8H5P+KjE
RF4i0Dgz3atzM5z5fy9ZOnmz48H+lPGViN2oAh1BQN9QFHU/3kSJHkN+1UrreXc/LhUp4Mpn7XMe
mrL6lC3fDJHa8DNRjUCXz5+1KIJ0ueBwuGgxZhYiURYlSBbyll57zLQWMG7bEN+YCY+yK6Fzuvb3
ZkRY0i7TIEKLXOMBWcrHjMG6qY6xsn5OFUK0QbtEMU5MKLgDvIqH4YMi2SGxvhA5MXzeuV4t9Av8
7TGjFUZ2DpzsUe2JYKGKbNstu9BCX91HcALd+DO5Mh6Klr77DTcA6UIUyMkWrjdkZDvx+niIvO9t
0ooxwnL3rvP5SLb15kvSfyf01hsTbq1rUm5AGS/3BhV4VvxDL4xAR3pFM0BCWYs/wLxmLmM5ridl
qGPKVv9Ceo1WbTbN/17VE0xt5vlTqG/uWPVbKyoOlDCU1dUoI8713mY2WI2g8Ict3GN1o0VFAeBj
CPgfprpdYPUUQgIBFqyPT1/nJm4Wl0+S2Eluclkz9SyBzqeEdA4dZprHFtUviDF+3FVvk+HUVOtF
g06+il9RYyRUNflPm7xkmcTL32OqarHH2oZz5h4ds3noHfcgmHwu/tsXtWgL/u3yTBQ/0Gk/IJb3
X1OV30Wn7RzxWuIhwy2sA1g7znBrTf8BaR4sneXX4YdNeMA/TT5p7jkl717IT2vTyz5HIjIg1Xi8
Uf/XSxzlQIFs75I522JuU1Fn19gzKKuSw4GfXhK/7nU7pQNnxrDbqbhpj9mDhuWW7tN9vpWq93a9
qsuP1M8prjrjv9D21L78YOKm0E66KpxG3zLZBLhoYRXV5EsuNR6f/nbIotf9RlwqFmDBcCXh0UbY
4Yl+cL9oQko6jhkcOtwCD5/JjNSVy3djamdJi+vbcy13nubnbgBr3NDFQwxzyx86Pmw6HCUtk6+Z
AP+mpbEgyUP88W8Yn0nuT6Qz959tuOKk66YOSZPsExkrb2rq1rdK2NRuwXctIi5JVoLw++hqfrxp
wDHGlrjuEB7PjEWhEjDy6ovQjGrin28BkBcylANTouImjg1Jcd2/1f/Sn56LHleNkktxjxAWt9/S
9sEBW+32JecmXzRgbvEGNLMc30PKEzj3dXURgDj8skgdL6ZOe9mCTIuyp6ElUMKCGpsfVu28lNGw
qaWuZufsClUpfsr8p0Qz7K5IlbRxGH5Gr4SpwBCTrpjqCKCy2ghi3SS+cYY1n96xs41FP1la0cr2
pZwK03edWTqrprRYAppDwSfmidM/SzRxf7/vOpprA5Q1O0hn41ybzhdYpKJVBWgCB0U+nbltTxRO
afcsZvgsG5lblGCjeFM8NXZLpErD7GmGyYUSsqbf4WcB4MKAZJ6sYOLapSxbrwr4AWjxqE1IDrxC
PsyELVhEbdWDye54lzJQD8Pdykw+QX8th1AAI6sPKrF1JFPe1kYVKIg2QPUHdGAT/be6y6sk8mAL
yL3hmxgolMj+eyGYqz5GKhBpgXUEQ0xJxpOuMK6zNYYXzgglFrCQqA8STIw1OWuMRpfBsC4qIkwQ
RaHu0TkCrM+UDxN1AMo84Fj+LIzMRytdH/TleyCcD2X5qVCUM0WRFJVcfCmEaGMw9dIQb+dH2lZk
+gHn4w6UH6IeiEr0gZyAtDQ+X/ybMq7EheTQfRuYHrXuVjL/jh7l5nOzloFV6KnntUg5Geb0zOKH
XCu05SeRw8vcpG3jnMIcLWJFU3Wu8VwJsjOn5DRfWKkLKiFwtmLJIE00opfN4FxewFg5egzoWl9y
DIflxkR0oOy8eIqkvpZxE2hHFZygLaniUiWMWED1w5atfuFhRSxPArbvHoyA+vcZ/jiVKjddEvdd
7HX0CNAsfk4jN3S6sL3JTPgAYgZ1yjt1LF/HTYkvdxilFKD5Jtj5GWYMUS3qaUiHH51GYTOH+mNB
R6FmdCCLsSJs5UfVjf23QuB+jV+vxtX9Z+S47cTVCg0T5owhC73EUkFmPiIxtOMBy4PVlg4Ll0Sa
Ip1rTm9dQv49nf3pU9jA7mb5nrf0TZUJYM1jhixQLdH5OLI0aWo1CW7ebpzI1IJtUM697hoFjBOP
q7EZpL7G3OJ38VZCByTRTm2sM3/48rmbTym5oQIFHcEkgh7Sd57ppeAEFvVY6nczmHVgHe88oUnG
iVRCor4yHAFCLCj5aI9l0Ir4getJ5H5wzca/5qvi8+mZYx9JWO8OxmTeGH7MPxeq7WjDDg02Wla1
IMUa1w6dgpWKbB/iWPUvDnBnvnB8E9pObjCRyJsc9Uf50WrtWQME8/s1V/oJE4N0RSpZZSn32UDC
FXugWlc5ESamVOuwRcxmzbYQ0PHdEFZoWS6hAp8hPG6BMiC67a0XLGpvoFw8rfWKp90Pzcls18/d
A2XqKTWz5khs5VBgP50dXMtGIimUTkqlj4OuWv/G08yr6HzejeLHN5LfJLto0k4PwZshjIXidXoU
kojQlqFaHaUEwOQ+wr3MvawNC5tSKsbWdsflRO1zLo93uMrA+IW+RxfbkTW4BoD1lqmeIwxx+4eA
3qTnWX4IppVzhnaVqFwsEey7uKhxBk1/8XUACwtDeLBwXJNj+QtiQVOS9v5Q3/XHTLcS+A7oXPYn
j9WvH9kLZzyUOQBK174uhg10cqjpkQak7x41RBN91jD80pvlDHWYok340DDGhGmoU57tdRPjAhPZ
5G6ekQqXA8IrMDAoU7b6XuCRSSHhQZq4xc4nT2wJWSAjupjAP79LvgTha0T2CAFQFYRZOHqyDWtO
46LhcOoGDZONAadNT48wLbXIl/IikP9PU2cuMcxSzYjT2eDMm+Dc7HUFnioYoMphPgJAi6W0AK5y
AMRW7rjLRcTKknbmR6tgG3+S9kxa3v7DuoLsqrQHsTAJvgTmu0YK+87v91SF24ctvEZ0oFcBELey
7k6hB9abw4AX4yaw+oXBwM+jKO71qSAqhZO9uuHoWPjMDECze9DQqNUQexzAuH9oOP9OGSd68+JY
iXbvqL/nfRoUzcrOCowmJltgsl21IksC2cr0kQQk+GTNNbSbCotsNcHllMJ2ZyBQTRP9NcuuyJ9d
JTUDj/l5GfZ/3F1pXSRjZL/jLw8GV6n7gc+1XJrw/fIQgsZqcIbhpxx9VagODpsthrm0Ewa6taqn
BbzCZvlhDu6+TVwapGyEfntJDpUapZV6Vjo/UXDVjAKYUCeS9x+ej0qzrIPzVHFlA2AwJMilNMSX
4AhCmJNTiClj0o1i0HeyyoGnsJssGb2SdTvIfBF6MwK1ej4lyJDx/f3OObrcABfsbCk2ccAv1+jZ
PZkmWuuk2MKzSYHVf6KTEF/b1XmzLxmVHuKr87Fg7dSvct65fjwEHmRqHtVi5rYnfSCzrjQFPIms
oj1x4siAaLc+Ss8IrXc/CdiCT4HA23YlTX/5S5NEivxEYU4lyQC0LnY4LfPTvgG6gMNYyzi9Z5XA
Zx+k1CCuVze+wU1AOAHmcOqvltc5n4op8W/+sfwb/eZnZOinSkmrn+/CafJECo2aJWvNdvv3UZTU
VsIKDN1ad7GDFkT8fsQmOc+jC1IG9jndISh8oyC5hT/8xatnYzjffd/q33Si7rfzcG+hLdDJct+I
hR9EYGACCiG/pO8VLOrGNkslJpx7lNOAW7K5rN9QeJUeQ8MzrtHHMoQZz8xem8gniUZmL/POtZGu
l/c+WrukeEgHHvMKBIHVUi1RopO0lH9yuL37kVncawZEwYAi89xNUDQPPgJo2IxEARMiBjaFG6GQ
giMlgeNGJhDUKPMZY9cvxMFUHKGj90mT04bdKrU/NmVPhgUzuk03Wk+QR9cbllGpq/YBgLzmyq2V
xcKVYpAz91SdckzGcomUeiAtxjbgZesW24U+/KnRMuaPZiHOeJSllkphrryA1h22iqWwxIajptB2
WbU/pBrUVIbhouCnMCU6YGdMN5eCorCCCu0u2sx3DFYToC7MYd5yEwRgcTDeZ3IFwIiDX0gj40sO
JyqoYNkt/w6Sndo/2hQe2vr+4InUZ9SyN4S2Len76PGbyJQ5ahECU1yYfmo5e87F9JNUCRp6l4mH
zGQWfenhoBHK+I3AA3/d55wrqgfWz5YEvazIuhPNRNl9I4yrf4VXoODVJErYdlPqdL2LxmV1U/8Y
4DfHyIKi1gKdrT1/RknjoNL1Z/K5DD9+bHgLSdumKmfqD3ooYHvydpb7r5WuSuSUGjhqbJfFysj8
WVEOpgqYjXv/X/5S9O1La6l+LcrNKJwwi28xP7KcfHePiIFAgYaNtk5/OreWvDaHCHv4cfSbs4bl
CLgmYj0Xw0MGI2EC0MQSC3Tc39njvsi4wIjjIg+UNAdxY0xAhHQmVcMyIJ9qSMGFpAK6+E58daFp
XE4KxWcxTJxrlxUJqi0GmeahfPah0dLfQ29E4HcXsXh4QSJoDSodz/E2raaHDphJRN1/4fdqredB
Xl6+DWrfwig5GZBsn82VGq5NbpVdQ4jbixGeiwsFng5W02DaIk2W20M51se+z+pF2gxeyYgCnNG9
CC+6qVgSLaFfewnaqCqzYGxR+j1H8t+dCcsR+XqdHNBpjZHXd4nm+7tghFez4ziChFUVx1r1fKug
0aepenVXI/o3B0LCfgXBUnE173QML7yjqxPUzRTk83qLLiZZsbLnb1EHef01dyVBG4sXXZCy7V6Y
8ug3ifVoKmiQEydPYwWf4NBDi2q8IUA4Kcq5nOhoYEUsqisnadHO/YTcbJtgAlm9EnNkanvI/ghv
W3DEB+4y+gJc3x1GLS9UNlk1n+V3KH0fqHE8rPe7N/QRh4bnnpuQXpaBfGfhcPOiiXIE9xRcL8Yl
iKwnD3zA+UXOQqqU8gSkqxe1y/g8tnRRJkxEM/ILqD2uxe6tyCWeOAP3dsfZFG2jSFFQgH/CYmZm
wP6FeZeNPxeWE4rMj4IHmWPh0ejeaebrM4Rr2MS0Dl27YYjtwprZpBbT+GWP4wXCHMn9gL9MlXen
uUYpLWLhriZp92r2sp5VhJzym9qrPOINhYl5KzmOjH+xiROpZEcgll/86LED65Dv/OgkDh4Q/3cZ
TJXGCoLsaYRdf8NQgnmKV5UPs9EDYHg8PF0FefbdNKjT/1xG3XtpIMxBLLHOXv1q1WDP4tDusQvn
y+aQhywtwFII2gtCITR51mqkvW6kBibtOGUSScQ0d/NEyb4/Zezut5qQ/D3iRa6y22+kW7/DhpAQ
QO6VdraRjuZtF3VfDeTNZd/WTGlm/alPf56bJ1FD2C2NP5ZiNERhkylacxGL9/BdaEvYO+xjBt5E
81Kk/iZ/eur/uUKXbwGzr/21BM/eUIKL+BIHn6sleoE7bqBBBIXAbc2ai2kWvcIDStMvkd05LpTR
xds8jEFyijyydwGnIJoFx9xoeLT1FjToCC9QGBHttfwjZirt1u56eu5uU6CkA3H8+QjNbo+9Lxtz
HVQ9euhz5JhnoKqNkYyTtKq3udiHymFnP5FQd0HuKCeMwv45+uZpWLT56Du9zixdkZaWWp4LqhY+
F6vZh5xSfSD+JmTCmjxLC/DrKKg6DvAEG4uJalFzzqn0w+4/s9BbO5KciqIuBuFyGMt2EV4kQFW0
gcgqlciwOdQbLzBTPkRq+QY5ePWXR6wlaLrLdIBtQ51zStcXjMwS+PF77Vp1YmI2yUHyaKArov4h
50+4i769cnjerjsLb0NRkw00O93WFCmedW7+Dg+/F5RbiKdKrLlK4RhaTZ/zqRWFOErbiAXY0lUO
6ZWuiwPt5d+c6XzrIbrs96pwFpshbTXyiMWdrqBI4FAE4J6dVgyOENoQDMKJdzOOwojertnvppyc
5Io6DCKqSpAeR4LFt0t6YgZovEJCDCt1WLvG9t3ixO1peDq4xliMJsainmbZKrFHziCPXvnNqw+z
qzPK9EzOiofs7AKCD95rkzKutV+5YaVdZpws9QgbjckyYKTap9npRz8wxrRMrDNDlNi30XALGrzu
1QyMA8oHGqIsT+BI3FWKAx+uUwPpDNQixXQLoYsQpcGJ24+C4QyH5F1VR4dvwnRd+qFDveDo2TpM
dFNqq1VDDkE/td0OfpNEfYjn2COswiZOmk4pMgj7nKRDqPchBi4ynsKXcK+7q3WryTWlja2vBtkh
8lhrDCzX38UqmEudNcDwcorwDqy5+chPTz0ukisH5+WQzpqQY1uMfQ/Yqsh1cJ16D4lbzZafxEFe
wM01yqFtquc1UkxQYNZ0Zxg/0NPivbkZz/c/L3jqGbX1PRhFtwXzP8msCp7gb7LNJ7GYhVNhpevL
4mPfxNFPOL3sYJ2FscVWGZvmNhps0t+tmKydGVSvwoKcgJOaoxqTWXhnNS9bwieMt9ZKpjucVmNr
lc+OSaTcYHaBDuryDVCZE1f/tWNqG6/a59J0XwOmQ0zj5QAnqhJaWNAMkhdSSs+b71sUbAykch9+
hCkrvRw8jdg31zl3dRujCRAbDMcNc9jSe1mkk/IfLqIA98VAdLl1NXkgpLYnI8fG1HJjnUwhHeK1
txAU/1CgkgwVBtwUwCAHBPkewfZGt0POeBTfv1IpL0geuPziIGnbzhh4bSo5X7I2Vf6bl8L3deY6
xev8p0HQ6QONht5ORNcA/iglADH33Ik1iJFAQKBYSHO++pfh3D7PyK/cz45xqgdjOh79bsFNU8e6
/MUH8O5TLAMycN+uHF83Q01cMMYDOEVfkAoQx+VbUJaqpgxYKaZY+1jjMj9i4qgmJv+cKqRX5AlL
7+bcevYbuJtGsavyZEVz4EzxRpo/TgTDCSEsDI8VgqDu7D5JrtQITKLwdvCwub3W0nq2NZWyXSUL
W5e85TdqTQxSdGTahEn1K+7MPmxUgDIFve+eGW5qM2XA58R/ZnkMs469BanZwtGwKeySgaUOfsht
9ELf6uERGNUvrNsx/7QO91BHyGK7bV+P4h42+K5rJH+5mMWY993e8ZlfOb0PAyIFj16lxLIBSHn0
75H+MzrZB+cI7OMEJdPx+gUvB2BjC2XjfBqKi98qCMkKwnciM+KOSQYJkgixcYuZV/XHyGEdizcb
3Yyklqv7+oj7BCRa62gsucWKMCM1bV93fVmzEKqwOVvykQrDBbvvBz/J0wtRhikHPm+MHEvjxOJe
wGmoqq/OTFcBWzq4suKUgqjDXZ9sY8vkOSbIGz7nd0Wbad8wn1hPKDc3w4PDe4CBGNlQWt1TI5gW
ZwZLmZjAY7zwSud3cFeK8Q3CtVmWHLUGFUyxZSnzDZACZ3PWyRa4xH78KSv/ko1+LPAXvIRUarAz
PIsJec/BohCItinI8qV0FwQML/a8W7zTT+MFFzT0dkjczN8lMWfekzJ292yuSejYIC7rQeeIv/Zy
cVYlF9FA9b6gnKOUSsecsgnhyM5nHyum9Pp8sPal/YpttnZxLKhoSHxmsWf4Iy8gmrpctRHtjzel
WPigEExrCKuyxx6oBxcksyoEk5FBNAmEQnx/GRyDQRLALQRe7Lsd9/p8nDa98ls1qYmSQ6RxDoIo
hKJ1/2++9OfnmW5Kd+RsuwAwq5mW3OQQdi/pexRCJ6mOKnEhjth+elXarGtNhH329taEAY6AO3Nz
BQE6hbWE20MWaI7ig6NlhkcPrYynz3MmQCkRh46BOehbeS9AHxX8lqspAOF7zztW+jK/LCZNiAty
uZ1FgseHPBRq2PhbRURxSawvlRNcXwCpox1XxviyE3qqDA8l6EdV2//sXXHEYQl4PX78Wo8Bxk8g
DF7yFXRrCVbA9uG4PseB/gbOAOdcGdkPl5cRu7oJfnBoNiUTcNfaRrzL6c0PnFBGrGZfv5nntXL4
oJUi8nOQoSUq+BY+rpulcDSVy5ZHb3oBLdp5+NGLXbtUkxnqW6Hp3xGilNS+cmJtX4FQCf6kzvXx
IWWPq9/UZ2r4Ajji+Y+TLtTeGNzix1DiwuBmUukMBkyT7KfmHL/FP82E+a5ygsMEw7SffHQvUU88
Sa9NO2pOVe1TrqYC+FZVihC33yZs0LLCNPdwTk3t+1OV3FayRgjNpo42B6RD/PkcwrRtNDWyq9Qv
FeIw0q9pbrAWT81LAiGU0Pz0fYIZgNDxsliPTbfcMEhKRsOvcAoz7r8vWjVWcluiMvcjPbvu1Zkb
lVV1CQN68q9sJqsI9tNPPb1llXEqdOdI3+XE4WXW34mAQfC34w3dLuvRmAy7Ha2tufFAaXhXm5c4
iPDGNtQ4AXN8A54aB34Ulj8BuZhAZqB99NtMNn4AZd+saC57D8vOiMvRxSlyHTQdgQk3So0m2SZG
0AO3/vj4gnwGHVpezkky5fLyXJLvn/hj9hmsURpioEoP835xAyESqtJInE5ZPopsq4y0C6tg32JS
0dKZsAFUWbXwwfo0fOwhfbrTcE1vNhc4NKbzt9uDjRxNo+xWBqYU0GIFtWJ/SNv1CNyRWt/4Zva4
uPGzePiSzIgHWoeXq3PinZXbLPuutJyWH5XtPxbk67jbi16lC1SuHHIPoJ33wmnM94UPSdFBuPIq
jo5n0T5rCemoHWKMAWrwR2iPUdXxrm25gYMV07AFerPtb9R+VubQ1nyqoRa+rxthXTYD+XbFksfJ
tiBtEfX8xvblPQCHI246PPs4QgPARCLWH6nL/Ajkb9iauenIk1VMcw4IzS3ubfT4ugIB3H+BA4VV
hevTajk6Q9ekabpcAqvC8GN1I+0eaQI3Jd8P7MSRft32CjvnVAdloQ6bOe9YcmTVi6jX+rdG6jkM
HIXO73McoVt6XBEqX769t7MEz+DPws4TlQRTPPeMGgB7MtSuTD14FmaeKVBzMb8fjym5bYOIn0pC
mVWNhjomloKG2xBRi8nXFhgaelGX36yxxgAeWDY3mN6K7g5QuvJhTM6zc4ImFwjjgdfPMGr4f8Qi
P/zeEuqhEGfkkWBM7EHkzapzjA1XsE241rKxjaal9i5HM6l4ddk2HQO4INbeJryKDHk0Wvu0tZPT
oOC7okD/smYxVA6gblX7/EMO3ezWFLytEMs/4d3Q9FSOBq87HumqJJrrhXpPchmbd/dW17QYGLcy
srDEuryfdQ2dNXD+noUmUfhtoXL17o6W79m6BIQYtGaat4Ji4GKC+MrZkr8wWtfkp5foYePQTwvS
DxbRwp+sLNvD9OL9LJ5w/cXmxqghTskucXMADNdQYBpm9rPyN4IGmaxGW0vbMXKBZeEmgK4IgUwa
uEt3iSNoeVJ9IoycYJrzT6YTWcv4x6P3RyA0QHLMpeIs8HIQZYGIErIFDiltYzOF7jChTekmUZAu
JwuUZWjfK0beeV+lhTrsIEf4vWhzW+jDcVyPWYoRJt3yeLlbJNDJrVmZEa3VlVPVu43jOUf5w+xI
e0LRHuBdAo+MClKMz1lhsz3kTshOhEF2Wm7LJi750zbx4Vl/6QDIxOzsAbCij65p8ib6WDrEGwFX
Rrejri2euL7hjXVdq4mxaHLWx0YJgpUr7HjhxjJq/fctr8DCBPtQo9fH9RlGK4AC09a+r2RVSUua
JaWRgj3gvKDRiChb7NLSfbMCxV8HZkEPnnDHU/I4V0w6QSU6oOsse7N71EQ1G39OgHHzhM0472uf
HQ5D/ZcrpEchXEgGUsz5h/7KVRmkKfpSe8DogvpA84/iTZKhY7cZqCKIAqGNkjP9TBcFenHb99cw
u+A2GuhESlrMxOfgOCU5pShqtW29+FEb07b0G8B8bAZpID8oJvzFwmzNLYlc5q8LqlrkAJ2NVpke
LuVK2+V54KKgqpv3Dv7gSpam0jMkN6FaAp9DSdLQDLakn5HoSw1fWOOsmJerc5+Hg+zY9WKmv881
vaiYjhLzjncMxXmwp9h88e01CQd6Yp36m4gq2Xu+mvjjYQjbdKqawxBdLFZR81dSxTvsuUoIEzTf
fA25peQRQGuVgxqmujccqmMRrcH+Ze64hBRlZEq5LEQicVf/bbH9ZDDLNTU+qlMN79Zxu0RvxydV
BzZtgmjNT3eDLbLds+LoVNzapK7DeCXQUeMdXJ002HLN/ryIWTf2d9Y5aWciclBm2zTpifgrTcoj
4J0h0kX6pnMOGTpDmkBIkFmfCMgpP1lcEaaqZb/zIEJEfvvCfhhOp8chVmI2Tqruwx7sSy9Oy8WO
e6vqGfbWzken5x76m/NmNnnkqAfSy3bYW52oenjMWzFeQwHgyfEV2IQ+X3M4Yf2GCgGQCdm4h4rz
vfy0FmlEAbHTx3gD91yMJToeWHQpUOUJWRKTYW7DpMI5Q8K/slil3/ZjWTmp5drkW2zDkqpeEY28
BaIa54SZzxgervTE7ms12JrcLEysqrbRDyH4EBkOsIOV7DzPBboc9OpBiY/bo7fIZjDNpL3ovp1N
soEd1IyRi7myZE16a/TWxSFZwXvbqpyWyDylgTiJQo+f3LvrCU0tZUUOvliKjNrEWEIOq6XBwQbF
SSyG9nc1xbu+Ef7Sn+rU2hfHeGqLtnKOesY2ksJ5scS5sW0zKpzXqEecWp/5BZNg3QDLiFTZOFv4
7rbutAxY2E4bOlmju1qLTXu8pbbl6fPdkdJXSsu0PtFt+yh+iYg6qNpc3SqYDT9h8cNkRMPYoH1V
Ov9QFs2D2+fVUteuGQaF4ITfeO8DKG5C2tDtP4r1f6Z+dcjKkD9acA5RCcZxF/uX31qP8oRFMs8c
EPNNzhF0kpHIxzQ+mTS7k1V44y7KFsdyxP+HEiWB6/a/Zri9lmk87ezcqxwTVfsVT9ZoM2Yj7u3G
rcX9CwKMOUJkM6jTD9G5dmLLV2Q5JFJCASSRinvxK/xPv/Qmg/RK7mZdLHg/r1mEgRrdSGZaAIpQ
Y2mE/AjLLtXtocIjd7VAA5p8KywyxDORrVdqbtSRkA8ESRnYAF+apKJ1vb30dEucFRhEiweISG8M
Ux+VA1neRdtTqSEzDnP2juYI7mul2BleYCPYV+GLMLnmi6aViSl57kE29FdKeWOktAWCHctlhi44
zgBmgG2oTeRhVreDCnuXGvEnWUrz8HHJ2jd6PjTkii5Wm6oZnhQWsOPZ6GTSCELBPzapccy4pdHM
nof+ICBF38aYwr2Un7E3U469QC1RdKofJDSXsRYDbpaXM62gB7sPMgpsJhjbHwhYbWafSRO1S7SI
aoFhpoqD60PZuyChH7xH39FtllxnChHLbZNTl3+dpEA4hHVKz1Xb/DFid3IHBQru66dYATre/KYH
qXWv5TbLeGGtw+rI2Fkv1fCRaWp3Mmtnp5YwBOxv5fIQiZo9gIrzVzGnaQPyFWFhAfEBVfXFG/4f
lSptYSnPU0kv1c8WwbmSdJxpr1MWehIizoSNDEP57F9g2h2bzTEZPcMJg6/zIftdZhl58jUHFZXR
uNXZZj3Xj3N4unirTBvmhQJWpQ+UM78NdeOqVYp7a7YvSo43nctbI8loipYEpvJpRaFQe/mwpnKJ
Bb9QTWw3nuHvSjLHmhaDtCBaLOL5vurAZFpW64zbQLJd0TBq2zmmIJ8hFOvlm7qA3CD4jTzlsqX0
86Mu/7RtF/5X4YJbrOvD7LXukGy4JR40c1s496za3MALOyJfjyGVEoKgwVc7YGQRYSYiau3H0Gfx
VizeisjvLah/pTr8biL1KVICbMbn6V7LGyzYYJPW7Zo67SWP5T5n0McYyAc3tX9bT86X6smmK8e2
ktZdTNDIvxahv8EifKqq4zvLNI7GL8YvolIagrJ/G/ZhSO4SSWDz0bmeRZALPovwWBm3PBu40CWR
MtPPij/MBRlPfe6HPIWZJl/mvJmPJTQ4COTOC09qwhEzsuYaaBqKpgKgC+CoaZF9xc4TQAlOzr5/
YwLymsQLfetFGItwDZvEWzmNd4onPMBH7uXyM98L34ZvV7XoQsG3QQlPdPd3zlWNHEV7UU1C5GXF
4z76adLTQcKikR8pBlHNYEB/dFSpHIynMJOqc0kwtJvIf1CJEQklKo6PSa14AyUh8iOfVlOuMqDH
Wli1h1PYGeAD1oscNeIYJFAr/RMH13EXgV27JDPEP5NLCUDhWrqArI75j7UYFZg1ip8zby5rTW0b
KhqzJhMBUo5Q8yhwMfYBgwBcz6Nx22dMCAzz5XhIiofVzpByv9+f5St964qiN2QalNw0oJZfOQVK
zu9gwcWVVVJsGmtr2qOxI79UTlW/GdgQuHa3dv4T4OoRJNrcnm40Y5SYhfZfZgZnFgGgtQUxeV/9
FVFXWpJKZUJ9Ybe3ao1zFVMwD6Lo2JREmjhBs5asdVnmN6yI0pxCzi9DG9nJEZjVUDHVP9OWOwXt
Bio/DSvaE65DTi5klRMODvRvp1gdmP7al9deaF5TWKHNJejZnP32lkJB8ulcfDCuDJydyLSki+jX
2Xe531UxjQ9KIWWWgHTZJkMYZJOWmDRZE3L121D7ZfdZ86GCE4Ak2jP50LGoHf9vAk015NKwG6gJ
VNe6pxQdThgh1m+xmfGwALS7OUNiNRuwfWQI5uugDZCn1292k6A2Ocare3Cm4KVOYIreFFMBa3qt
5fP4D/t3U82+HqcuFpF2o2jRWAiKmTTUCBbGf9wGtyfXfy3tdgwI5ZZ2xM7nPNWfcPjikXeuc38o
abDhskiTR5k4vEVmmJhI0qNTavMH/xCFWw+sU/W5QeFSeF4uvpE3SXd/hWeVRPmBRf3mEC3N7Cs7
xnwdEQdCANlvOca8ZahE76r02XzhxGP1G8RUZ+M4g9hgZYLwiFUfD5MMF+O49PDo+48dP5Oj4UBi
bgUXetAzNOiyyI51kIduVsC/NA7dYQhvjp7nt6E6HyugKIHUgD2Bp9E0Ra0epTVUYFr4l3C17hS8
X5BnSAHzLtNTkZURhFFq2bKtybBQ5vZ1h7NSZkPiLKSfobibU0zieH+oMUaSOnzsoaSkhnu/9klI
mudtkCyUsIlL6WRy6k+Z61ahROJ3alF8Zd8YDBHcbabS26ceMUNyqPaNRhUcKZpdsuDXvZkxTsf5
dJZq3i6KDqsopzvkyRMtO0YKXo6VQAHb+7FKT0u7FveK58Ed/FkX/toEBmFjYKyUFSEG9nWWUaG0
JnzCOBMnmkm+p1chLcfRzec09UpBxwvI2pgwhu5KK/1M9t/gR5LMJfcFQ+PrFHxF+Fyiv5k4huGq
1nUGo7PbF1tYIrke03PoGxhvpF8ZoRbWDpCyZmkbZiwRFKw/hpjBUf7cmpFMGk+Nl2MoatWJeBio
7lEDmx72lOwHNrSvMf1xG2v2QxqTikbm7kdpcHSYSiJdYsmQRBjW+Dl8RK6H6B5LM+mVX5Qwt3Zt
7EM9mnR3ghBckp/JYMkZ/gvd73boHuagKfmEIMqD6nlMR5fpX3CpN7KWm6TVt10fRb80JlHYVoDH
dqGggvs5rJxjy6eJ0hDNWWeYn+nmdkRG2dYm5PL7yh6s4VMpOYkpA7KG+be7tiB3bClAwYrPobmT
z4uRVDmrXyhWo3gM9SMbTj59ajFpFG0EzIhYjkobrBjQN/+fkuwCsoWoUGJee3BRhvFyIJC35d+R
Wqtfo7KzuJ91l9IVozGDDuJXIjy2tgUUjVF+PwJEoB+9NNxMYdVq2SFlOgPjutI01367hI3GPJP7
rEOH17g5F6TwMNDrGEwvFWsCTVjzD6RhPCHtJZ3pTHbBvRpA6g5tbm/i/OZQKHfNFQH2/9C6JmG+
1vdPr7JqS1q9oqcnRgmvYyAlTfh1Ck/PTWBo11PNySAqbKHMSss0mo4S/wAQuYUk1GGP6Gh52kUr
6CwQ52hrgRDNPDuthEqV0qhb3olIvF6Tcczbyy46OIR+HEIctWSkNVm6Q/eOwGLB1CHYmZVrCHxn
AkPX55Rh8RejV/TAAMWXTqe6QzZbbt6pvs1XUCNJ2oalgrBAtWhjZZmo5z2CeJBZd33LuEx7DDI3
Ds+A4PxxpERsm+mJwy0lLOWo3vE3p1hu4KkpeqHvTGikBs9A7187KXjbX7NdJ/OaXN4mb1OD48mw
7U4T3f/FMz0QXQkBEU3NypfUU//FaMQPHppSNlSy/h3vgNGoAF1H5GwF8ZmKzdzDSbhFj3et8BaK
WcToSQpLcUtjgiitShg9bTnoXAW4ORyl6blssobVcoXxES4kuehzRVIkdkdGV1GPEdwUBEbarf74
XRet8ZIfSgFOxGliATdMsCYlOEf/iulCfz2M0Uq8fCfeX3/WmEYMXa3K9BgllCMtzTu49sKoFoZh
zMtVURUYUvAknx89i2dH+nUbWb/kbVrmuL27U99WlGe+Pc8aZlUUJr+Sutda7bg0sSBThB4H1FjE
UohZg3WSowop6jBbaUniVlKGWwOhUZZhQdbVQhmmBuSaCFtEFwxwegGYNcVlocZXlV09lL/Gh2ip
yp8nU070M1aaf/ODwI/6ejNQxnrINjYd4+kmreJHqGIF6KjQ3CPNk6v5Nj2ZlmN8f1fBk5PHrIy/
bj4XEIn5StAYfLMrrH11ZWEfj1U3mCxsHgh2NhNld89+jbLf2r2/VH7H0+aq4qlT5R6UkTG05arQ
+ZD8GBFLgjxisv/ZZ/n2sK3mm9s1OnpK2lMU6yIyfceb19AgQmtHAObyeqLHAGJ90atbn2kb/R3e
7utKLBeOYlJgWU4tHIWXGF87xPcO/bAvzNHzqMqlGwrvWot69W0fIlKzmUlRLyd++roM/QpZTukW
hBbimoyYhnqRs97aWXB7L1gdoRHAQvzl8G+0UcPlJVCrvhLJA64Vm1C9dHbv/atciNT1H06+4bdU
E+tc5yyIdLJqefWWIznmiACFDgBR+Ry4rYOO14CNtjp2KvuG/9e34juE7ftxY/KG4xtqDkRG6g/0
y/OEpl9nASlE6WpeIkPJjzxEomqoO/FlE0FWH0NQjiEhNGyjVxMbDeKyEmV4Qt9mhdqnLP+haRTE
x+1umpnnIt3wYUNIK5K/8xKZ+oNsTAe9WnW65vtKc69KI/tkK0cIJSrW6b7ZG4Pha+2ikDmsxsMY
kz9VljitaBRe3398LzmRkduzQBoiPM43zPfdog1MmUztDOYfWrtkLTX+ufRJc13MwLDly6J6y+N2
3F06JQcTcbRxuqsEdBPAxnhWH/iW4aHbuXRXi1J96KRxVtS3sQAO+HSPrTiOGj2bZ9l1/SM/V/2T
y95REamX5Br7yFEglQvFeOK2pSukOuxz2gMyEuicXgQPcopWPssWMB/8zw1mjdBYgFZdGkU3KP24
+vRQX1kErIMxPPDaLZPoRBNTkla2Oz+Ug2lv4gfG48r8eygO52bACzVCGMtCyMrnzOVxXqkbq9MZ
hIR47gmUApvgdHlIVkNXJKgvWrYPykAzMGpau+yWfbERhhghwtK5AJUvksXv2PaPL9tGpzK/8ayy
D1hYBBVv76SLN0ngjwXnJDzBQcL6YuhIfWy5Sg7cw9ZIynDG7dw9mXeq5n987f660NBN1ZehiwUk
deTAxbhAA2+4reJRMra2lxGQmPIJwBbdY47G4MxQIY2poQfcwWMgqONzUEZ8lZnJEKUxN9mnbIvc
BIalj5gbv00yHjsIZOWrsUqO2jVprgi87R+9TffBFXbePAN/D8M5myErtPD1c7RQIyBoazNIIQUw
XkIO493y1pqtcU9duE0BFG55baM+AKHB+XqhpDxZ5Khc6GnJgrIMPgSEroGzFpIa08MPIwT+nzR4
Q4bG2m749l1ucHfa5S+lxwItTbKXn3m2WrR6taS6pCrFNlBrh6lflTftEIt6u8An7xxO7pgDsflg
BtnmrcfUGwqvQYDfnIdIBWNqP1Sl/QX6xUSmMo+qXi/1A7V3cBYtmy5uBWhXmEwv6iL+GT4Dt09L
xBtotYQBy0HZR5oJwuEl23I6TDwWy6Pn2uFQAGutqLxachc/biiTJeyzpJIJlMFUrNS9tCLHCTzt
8Qcr5oCqhPfCIDodiC2XW+99exLiUTnJyLszXTQ68V4krAuvdPwgUTmwe5wHH+DG5+ZHzLMlzxxY
bQ3WxgphNBqhyAT7SyXliIfZAJx7msfc1s19pyL69sFifLS8A00Rg0Xio/LCzXoJzQ/tkXe7nB9n
zS/AxEUx+CJj0+2Ty+9uZklpT5/mnsl73jJRIXNJY0Xq5cuIB3hw2IgziMW/XKRjRj6QyI83H/G8
j0xWMUqdz1u2qIjTmPx9MndOEVz92wMsIMU21N5CWVCLQ+4hQgl6Y7QWarUdndKs/omAVJskMJXJ
ntBJTexXL691mj2PxZhjdwOy6buuXWdnzIX7b21/n05QtOpL5BDCvJRY1fzAZa6tyn1Bxw3lSsJH
ExP7wrKZLwSgWAWQaYhStW9d5HbCLODur7szSJUoPtl3RAViZgbMb2A5YrLKXzSiRoWaV+FIbQs5
RrmKzOTk23yp8r966w0B2Eq91kfMG6eQu40dJogFTQ0SsCXVOIQE6q2lDuOV9Y0725X77gfIwfLq
ihztgKh/lU03W5fOLiHRqyqeX/elTQiU1yOVbvQNrgwjWJhcPD7PJHjKI21ELo7nMBPz5lsJi26x
Pnzwqd6u31Ti5SZUYQcqtPB0ybRfWVkMtjN3/pcDYlnXCTEYb2W+IDCxPhluSwz3EmAco6XF5p9p
r9O+dgseJO9brEmUC+9ApR+R5CQ3Bcr3+jQi2t8fYeyuIBtVdFc3lj+geRfgalozCU6GvR2wkc9K
rCO1DmCLuJ0wKrZQlTEAYjkZGUmhA5S3PFscQJP6o+IlI0o+DrgoSFb10mr3B/Ao9xZpBnmJRQlZ
cSDRJkSJv8h+xDHSf4eP7Q9bWjlMpddCZpckUYjZW3RNaGjIqi61KT32CXCpsNqxNiuonqLOVRRO
cfw/qqGe+Ev9III/DiqlwItYJMOpD2HWVk5GbCgTu2fZ/aJVtA6O/W2o7MhvOmIYjHCD4bIbcKTe
xLAqcd3DUk6Lkkg8yRLbwjPJyRpnxMbxq8HLJ7Vdp1FV43u6tki+ATK15iR+iKLgy592UXnnvwRw
QbxFT6HH9YdlaHbuGjp/1imV2uUT/5i6XaeIXJH8Mx9bh0i6BJBBXsgMqSRHtLdSbqADM/yU3h09
7y1Dzf3cbt20wVMOO2FpyIXE8yC9Kn1aWx8BaHgfu3X6l8i/H8atvDUpscw6kx2cA9ccBz6Ot4bS
vr9k7/Pr6JhqSvrUZTqhghmJuHBf63m80hB8W6k6KGbCyWW+jXGuIx8cBCDom8MaFG7GVSmJFbuQ
7snevGmhDMoDYrM5YA6IDCF53Gec7O/7YkKTZln2J17QiowH535eAmOttWUoV3nskk6G8S12hfS3
6IKNr4KLe65WgueKZxl0Zdlb65jVFW/4UCs2GIX/iALiC7NF+pZHbz24BcrutKHae3sGXfllIJLd
sN8tO4E7QmYtDhL/fMeCt0DN/rUfAaG4McbaTvKAuOn+pUCVruUj3LlVB20OQVntN6mQS1lVLMY+
640XH43FnndFsgKpeFF+RDIuCTgBjyPn0aExA9CcVw+r4V0tj14fRVWhEs0IIG2mv/jNxDnpqzkC
gGTAlhdQLcshAyv4GWmT8lqkqfaEOx06uOcn7X3uWASNc7r7dK+OqU5CZx3V+mr5XLqGE0dbXV80
TXY+2k1r54LNO7RkZzE805eDf9mOT1ANmJtbaG1SReKGt4gnDHKKwgqEswiY1GkY8wO/B+BKJv7L
5mkBDaF46/CgyZBYS/FGgz3UzV8inCyH9Qn2lXpQ/HYDAfmjDMXfONcGUf1fO/0Ul7y0e5qiDZwv
G3rGyp/51sKNVvB+Vfuj1jjGUZ3E5xht2DTP7DsDsjg/kAvDOw4+VeQuuaA3/A+PGh7TayR7ukxM
vBr45yPj36MEEVWRD8XXhIzD27rnHSOBoZSihVEZu/gfxtnTGycUttIiRoLyPZFQ3ZpHOO95bFnA
qHvJNSgQ6cO/Ed59h6D0I8lxig5DZRNp90wCa9uzXS/1roIXB1Y3BWpX9ybj+KFibiQWHhhxonEj
7MyvjeYyXtDFcX8KpA2LLQc0bgbMHv+8fk6S/obZpUQlQFh8Qort7/cp4tL/3gCvrpYXVGdI7aWN
AitejihJw8I+3Cy/KGuxDN9XOmwwMRvyFHaGHLcqLkcscHKblks9udLcjvO4KEHkOCWM5XoNmuef
V0dDsau1E+VWt5lyaMrkzWkIet1SdXiPBxsZYGdS5nPy9ozSR6bZigvmzw0ExZz9O+Qv9u+vd9rD
e/MnKLzlwZKJoEFjbFC6qqY5i2Jn9g9SrjAVpyXtYTfWHBSGXnsBDXKKpgHEN2zjAEpcA2qDLqPw
TAQ9JR2fKD8ui3i/rP+3DeR4CohapJLEdxumjj1wHTQy9Fu9QhJKuHR4ajEv+bKEZdQkLnRNaH5R
eH5rMYo5PNcGbfeol7t/k6/70eKDxfB7DwZN8T0IOAsaXgYP5RSq6RHlVErLtyve2DRdRi9FOBBz
1ZAZUKPhuNwCSk8S5iNscGPId0X+8eI030wdjHfd+m/ri//cCsqeG+15+uzrhNiw9i49gqocSLdE
np91wZHc9RPpZnzaIQcZ9DZVeUF3uY8vX1jTdkiwmlo0+2uVUyTDQkgckBK0886qWIcHZP/Znq1X
6Royhu0zwat74jqiiLocyY5yqEJyXiLzzjlmXBqsuajPK+NfkiJyr8ft0FO9TmA6l3+TnmdOQtPR
rwTZXETL992BsyHpnOWcosenEWrbJMdtb5Lb/ERbU7fQtXMt0g/k/z55vEwLwZcUfzKBGv05oeQx
uylVaG1sOFsUTEWcVwlfGWD1ahdM8eYNOkPlzJcY5fCKNU9g47f7P9rcLWjkZrS/oX3+DZhfeHGp
hPEQz9jwi+HvQlf2E1SRjoGzBA7KzhYrRjHNXrRDP2y/7lwu+J80A9nj6wCMWMTzOODT2CCwvk0s
7dSHp//Y9Ry8nHpfZaoQEOXt05LYOiZMKoyH/cVRgYQy0p0tHQ6Bgidf2iMNyMe/kemcMkMrq3nE
zTrPgCowXjkC9d+zS2lo4acJ2Ojsa5iO0AzBqtJWGGoN7xx3h1FHfS6SCcbqj5VtvZXpu+iDdDdz
p82g2EkeBGYpsTrv2GzVpwNezxj6civ7yoEyGX3mHqiQlYFjeSGu/e2Sh3dKGfWqR5sqzFVxCdGS
1v5983Ams+dZ6lXBFCYptcMSlWrS3D3kPbDAzQ==
`pragma protect end_protected
