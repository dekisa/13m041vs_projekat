-- system.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		clk_clk       : in    std_logic                     := '0';             --       clk.clk
		reset_reset_n : in    std_logic                     := '0';             --     reset.reset_n
		sdram_clk_clk : out   std_logic;                                        -- sdram_clk.clk
		wire_addr     : out   std_logic_vector(12 downto 0);                    --      wire.addr
		wire_ba       : out   std_logic_vector(1 downto 0);                     --          .ba
		wire_cas_n    : out   std_logic;                                        --          .cas_n
		wire_cke      : out   std_logic;                                        --          .cke
		wire_cs_n     : out   std_logic;                                        --          .cs_n
		wire_dq       : inout std_logic_vector(15 downto 0) := (others => '0'); --          .dq
		wire_dqm      : out   std_logic_vector(1 downto 0);                     --          .dqm
		wire_ras_n    : out   std_logic;                                        --          .ras_n
		wire_we_n     : out   std_logic                                         --          .we_n
	);
end entity system;

architecture rtl of system is
	component system_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component system_altpll_0;

	component system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_jtag_uart_0;

	component system_manager is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(29 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(29 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_manager;

	component altera_avalon_mailbox is
		generic (
			DWIDTH : integer := 32;
			AWIDTH : integer := 2
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			rst_n                : in  std_logic                     := 'X';             -- reset_n
			avmm_snd_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avmm_snd_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_snd_write       : in  std_logic                     := 'X';             -- write
			avmm_snd_read        : in  std_logic                     := 'X';             -- read
			avmm_snd_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_snd_waitrequest : out std_logic;                                        -- waitrequest
			avmm_rcv_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avmm_rcv_read        : in  std_logic                     := 'X';             -- read
			avmm_rcv_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_rcv_write       : in  std_logic                     := 'X';             -- write
			avmm_rcv_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq_space            : out std_logic;                                        -- irq
			irq_msg              : out std_logic                                         -- irq
		);
	end component altera_avalon_mailbox;

	component system_performance_counter_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component system_performance_counter_0;

	component system_req_fifo is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			wrreset_n                        : in  std_logic                     := 'X';             -- reset_n
			rdclock                          : in  std_logic                     := 'X';             -- clk
			rdreset_n                        : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonmm_read_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read         : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_waitrequest  : out std_logic;                                        -- waitrequest
			rdclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			rdclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			rdclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			rdclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			rdclk_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			wrclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata     : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component system_req_fifo;

	component system_sdram_0 is
		port (
			clk_clk             : in    std_logic                     := 'X';             -- clk
			reset_reset_n       : in    std_logic                     := 'X';             -- reset_n
			sdout_waitrequest   : out   std_logic;                                        -- waitrequest
			sdout_readdata      : out   std_logic_vector(31 downto 0);                    -- readdata
			sdout_readdatavalid : out   std_logic;                                        -- readdatavalid
			sdout_burstcount    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			sdout_writedata     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sdout_address       : in    std_logic_vector(29 downto 0) := (others => 'X'); -- address
			sdout_write         : in    std_logic                     := 'X';             -- write
			sdout_read          : in    std_logic                     := 'X';             -- read
			sdout_byteenable    : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			sdout_debugaccess   : in    std_logic                     := 'X';             -- debugaccess
			sdram_addr          : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_ba            : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_cas_n         : out   std_logic;                                        -- cas_n
			sdram_cke           : out   std_logic;                                        -- cke
			sdram_cs_n          : out   std_logic;                                        -- cs_n
			sdram_dq            : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_dqm           : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_ras_n         : out   std_logic;                                        -- ras_n
			sdram_we_n          : out   std_logic                                         -- we_n
		);
	end component system_sdram_0;

	component system_shared_ocm is
		port (
			address     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component system_shared_ocm;

	component system_worker0 is
		port (
			clk_clk            : in  std_logic                     := 'X';             -- clk
			reset_reset_n      : in  std_logic                     := 'X';             -- reset_n
			wout_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			wout_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			wout_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			wout_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			wout_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			wout_address       : out std_logic_vector(27 downto 0);                    -- address
			wout_write         : out std_logic;                                        -- write
			wout_read          : out std_logic;                                        -- read
			wout_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			wout_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component system_worker0;

	component system_worker1 is
		port (
			clk_clk            : in  std_logic                     := 'X';             -- clk
			reset_reset_n      : in  std_logic                     := 'X';             -- reset_n
			wout_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			wout_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			wout_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			wout_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			wout_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			wout_address       : out std_logic_vector(27 downto 0);                    -- address
			wout_write         : out std_logic;                                        -- write
			wout_read          : out std_logic;                                        -- read
			wout_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			wout_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component system_worker1;

	component system_worker2 is
		port (
			clk_clk            : in  std_logic                     := 'X';             -- clk
			reset_reset_n      : in  std_logic                     := 'X';             -- reset_n
			wout_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			wout_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			wout_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			wout_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			wout_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			wout_address       : out std_logic_vector(27 downto 0);                    -- address
			wout_write         : out std_logic;                                        -- write
			wout_read          : out std_logic;                                        -- read
			wout_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			wout_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component system_worker2;

	component system_worker3 is
		port (
			clk_clk            : in  std_logic                     := 'X';             -- clk
			reset_reset_n      : in  std_logic                     := 'X';             -- reset_n
			wout_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			wout_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			wout_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			wout_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			wout_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			wout_address       : out std_logic_vector(27 downto 0);                    -- address
			wout_write         : out std_logic;                                        -- write
			wout_read          : out std_logic;                                        -- read
			wout_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			wout_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component system_worker3;

	component system_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                              : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			manager_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			sdram_0_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			worker3_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			manager_data_master_address                                : in  std_logic_vector(29 downto 0) := (others => 'X'); -- address
			manager_data_master_waitrequest                            : out std_logic;                                        -- waitrequest
			manager_data_master_byteenable                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			manager_data_master_read                                   : in  std_logic                     := 'X';             -- read
			manager_data_master_readdata                               : out std_logic_vector(31 downto 0);                    -- readdata
			manager_data_master_readdatavalid                          : out std_logic;                                        -- readdatavalid
			manager_data_master_write                                  : in  std_logic                     := 'X';             -- write
			manager_data_master_writedata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			manager_data_master_debugaccess                            : in  std_logic                     := 'X';             -- debugaccess
			manager_instruction_master_address                         : in  std_logic_vector(29 downto 0) := (others => 'X'); -- address
			manager_instruction_master_waitrequest                     : out std_logic;                                        -- waitrequest
			manager_instruction_master_read                            : in  std_logic                     := 'X';             -- read
			manager_instruction_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			manager_instruction_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			worker0_wout_address                                       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			worker0_wout_waitrequest                                   : out std_logic;                                        -- waitrequest
			worker0_wout_burstcount                                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			worker0_wout_byteenable                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			worker0_wout_read                                          : in  std_logic                     := 'X';             -- read
			worker0_wout_readdata                                      : out std_logic_vector(31 downto 0);                    -- readdata
			worker0_wout_readdatavalid                                 : out std_logic;                                        -- readdatavalid
			worker0_wout_write                                         : in  std_logic                     := 'X';             -- write
			worker0_wout_writedata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			worker0_wout_debugaccess                                   : in  std_logic                     := 'X';             -- debugaccess
			worker1_wout_address                                       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			worker1_wout_waitrequest                                   : out std_logic;                                        -- waitrequest
			worker1_wout_burstcount                                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			worker1_wout_byteenable                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			worker1_wout_read                                          : in  std_logic                     := 'X';             -- read
			worker1_wout_readdata                                      : out std_logic_vector(31 downto 0);                    -- readdata
			worker1_wout_readdatavalid                                 : out std_logic;                                        -- readdatavalid
			worker1_wout_write                                         : in  std_logic                     := 'X';             -- write
			worker1_wout_writedata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			worker1_wout_debugaccess                                   : in  std_logic                     := 'X';             -- debugaccess
			worker2_wout_address                                       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			worker2_wout_waitrequest                                   : out std_logic;                                        -- waitrequest
			worker2_wout_burstcount                                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			worker2_wout_byteenable                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			worker2_wout_read                                          : in  std_logic                     := 'X';             -- read
			worker2_wout_readdata                                      : out std_logic_vector(31 downto 0);                    -- readdata
			worker2_wout_readdatavalid                                 : out std_logic;                                        -- readdatavalid
			worker2_wout_write                                         : in  std_logic                     := 'X';             -- write
			worker2_wout_writedata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			worker2_wout_debugaccess                                   : in  std_logic                     := 'X';             -- debugaccess
			worker3_wout_address                                       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			worker3_wout_waitrequest                                   : out std_logic;                                        -- waitrequest
			worker3_wout_burstcount                                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			worker3_wout_byteenable                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			worker3_wout_read                                          : in  std_logic                     := 'X';             -- read
			worker3_wout_readdata                                      : out std_logic_vector(31 downto 0);                    -- readdata
			worker3_wout_readdatavalid                                 : out std_logic;                                        -- readdatavalid
			worker3_wout_write                                         : in  std_logic                     := 'X';             -- write
			worker3_wout_writedata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			worker3_wout_debugaccess                                   : in  std_logic                     := 'X';             -- debugaccess
			altpll_0_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                        : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                         : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                   : out std_logic;                                        -- chipselect
			manager_debug_mem_slave_address                            : out std_logic_vector(8 downto 0);                     -- address
			manager_debug_mem_slave_write                              : out std_logic;                                        -- write
			manager_debug_mem_slave_read                               : out std_logic;                                        -- read
			manager_debug_mem_slave_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			manager_debug_mem_slave_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			manager_debug_mem_slave_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			manager_debug_mem_slave_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			manager_debug_mem_slave_debugaccess                        : out std_logic;                                        -- debugaccess
			mbox_m_w0_avmm_msg_receiver_address                        : out std_logic_vector(1 downto 0);                     -- address
			mbox_m_w0_avmm_msg_receiver_write                          : out std_logic;                                        -- write
			mbox_m_w0_avmm_msg_receiver_read                           : out std_logic;                                        -- read
			mbox_m_w0_avmm_msg_receiver_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_m_w0_avmm_msg_receiver_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_m_w0_avmm_msg_sender_address                          : out std_logic_vector(1 downto 0);                     -- address
			mbox_m_w0_avmm_msg_sender_write                            : out std_logic;                                        -- write
			mbox_m_w0_avmm_msg_sender_read                             : out std_logic;                                        -- read
			mbox_m_w0_avmm_msg_sender_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_m_w0_avmm_msg_sender_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_m_w0_avmm_msg_sender_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			mbox_m_w1_avmm_msg_receiver_address                        : out std_logic_vector(1 downto 0);                     -- address
			mbox_m_w1_avmm_msg_receiver_write                          : out std_logic;                                        -- write
			mbox_m_w1_avmm_msg_receiver_read                           : out std_logic;                                        -- read
			mbox_m_w1_avmm_msg_receiver_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_m_w1_avmm_msg_receiver_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_m_w1_avmm_msg_sender_address                          : out std_logic_vector(1 downto 0);                     -- address
			mbox_m_w1_avmm_msg_sender_write                            : out std_logic;                                        -- write
			mbox_m_w1_avmm_msg_sender_read                             : out std_logic;                                        -- read
			mbox_m_w1_avmm_msg_sender_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_m_w1_avmm_msg_sender_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_m_w1_avmm_msg_sender_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			mbox_m_w2_avmm_msg_receiver_address                        : out std_logic_vector(1 downto 0);                     -- address
			mbox_m_w2_avmm_msg_receiver_write                          : out std_logic;                                        -- write
			mbox_m_w2_avmm_msg_receiver_read                           : out std_logic;                                        -- read
			mbox_m_w2_avmm_msg_receiver_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_m_w2_avmm_msg_receiver_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_m_w2_avmm_msg_sender_address                          : out std_logic_vector(1 downto 0);                     -- address
			mbox_m_w2_avmm_msg_sender_write                            : out std_logic;                                        -- write
			mbox_m_w2_avmm_msg_sender_read                             : out std_logic;                                        -- read
			mbox_m_w2_avmm_msg_sender_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_m_w2_avmm_msg_sender_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_m_w2_avmm_msg_sender_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			mbox_m_w3_avmm_msg_receiver_address                        : out std_logic_vector(1 downto 0);                     -- address
			mbox_m_w3_avmm_msg_receiver_write                          : out std_logic;                                        -- write
			mbox_m_w3_avmm_msg_receiver_read                           : out std_logic;                                        -- read
			mbox_m_w3_avmm_msg_receiver_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_m_w3_avmm_msg_receiver_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_m_w3_avmm_msg_sender_address                          : out std_logic_vector(1 downto 0);                     -- address
			mbox_m_w3_avmm_msg_sender_write                            : out std_logic;                                        -- write
			mbox_m_w3_avmm_msg_sender_read                             : out std_logic;                                        -- read
			mbox_m_w3_avmm_msg_sender_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mbox_m_w3_avmm_msg_sender_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			mbox_m_w3_avmm_msg_sender_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			performance_counter_0_control_slave_address                : out std_logic_vector(2 downto 0);                     -- address
			performance_counter_0_control_slave_write                  : out std_logic;                                        -- write
			performance_counter_0_control_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			performance_counter_0_control_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			performance_counter_0_control_slave_begintransfer          : out std_logic;                                        -- begintransfer
			req_fifo_in_write                                          : out std_logic;                                        -- write
			req_fifo_in_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			req_fifo_in_waitrequest                                    : in  std_logic                     := 'X';             -- waitrequest
			req_fifo_in_csr_address                                    : out std_logic_vector(2 downto 0);                     -- address
			req_fifo_in_csr_write                                      : out std_logic;                                        -- write
			req_fifo_in_csr_read                                       : out std_logic;                                        -- read
			req_fifo_in_csr_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			req_fifo_in_csr_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			req_fifo_out_read                                          : out std_logic;                                        -- read
			req_fifo_out_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			req_fifo_out_waitrequest                                   : in  std_logic                     := 'X';             -- waitrequest
			req_fifo_out_csr_address                                   : out std_logic_vector(2 downto 0);                     -- address
			req_fifo_out_csr_write                                     : out std_logic;                                        -- write
			req_fifo_out_csr_read                                      : out std_logic;                                        -- read
			req_fifo_out_csr_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			req_fifo_out_csr_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_0_sdout_address                                      : out std_logic_vector(29 downto 0);                    -- address
			sdram_0_sdout_write                                        : out std_logic;                                        -- write
			sdram_0_sdout_read                                         : out std_logic;                                        -- read
			sdram_0_sdout_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_0_sdout_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_0_sdout_burstcount                                   : out std_logic_vector(0 downto 0);                     -- burstcount
			sdram_0_sdout_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_0_sdout_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			sdram_0_sdout_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			sdram_0_sdout_debugaccess                                  : out std_logic;                                        -- debugaccess
			shared_ocm_s1_address                                      : out std_logic_vector(7 downto 0);                     -- address
			shared_ocm_s1_write                                        : out std_logic;                                        -- write
			shared_ocm_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			shared_ocm_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			shared_ocm_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			shared_ocm_s1_chipselect                                   : out std_logic;                                        -- chipselect
			shared_ocm_s1_clken                                        : out std_logic;                                        -- clken
			shared_ocm_s2_address                                      : out std_logic_vector(7 downto 0);                     -- address
			shared_ocm_s2_write                                        : out std_logic;                                        -- write
			shared_ocm_s2_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			shared_ocm_s2_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			shared_ocm_s2_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			shared_ocm_s2_chipselect                                   : out std_logic;                                        -- chipselect
			shared_ocm_s2_clken                                        : out std_logic                                         -- clken
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_001;

	component system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_002;

	signal altpll_0_c0_clk                                                     : std_logic;                     -- altpll_0:c0 -> [irq_mapper:clk, jtag_uart_0:clk, manager:clk, mbox_m_w0:clk, mbox_m_w1:clk, mbox_m_w2:clk, mbox_m_w3:clk, mm_interconnect_0:altpll_0_c0_clk, performance_counter_0:clk, req_fifo:rdclock, req_fifo:wrclock, rst_controller_001:clk, rst_controller_002:clk, sdram_0:clk_clk, shared_ocm:clk, worker0:clk_clk, worker1:clk_clk, worker2:clk_clk, worker3:clk_clk]
	signal manager_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:manager_data_master_readdata -> manager:d_readdata
	signal manager_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:manager_data_master_waitrequest -> manager:d_waitrequest
	signal manager_data_master_debugaccess                                     : std_logic;                     -- manager:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:manager_data_master_debugaccess
	signal manager_data_master_address                                         : std_logic_vector(29 downto 0); -- manager:d_address -> mm_interconnect_0:manager_data_master_address
	signal manager_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- manager:d_byteenable -> mm_interconnect_0:manager_data_master_byteenable
	signal manager_data_master_read                                            : std_logic;                     -- manager:d_read -> mm_interconnect_0:manager_data_master_read
	signal manager_data_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:manager_data_master_readdatavalid -> manager:d_readdatavalid
	signal manager_data_master_write                                           : std_logic;                     -- manager:d_write -> mm_interconnect_0:manager_data_master_write
	signal manager_data_master_writedata                                       : std_logic_vector(31 downto 0); -- manager:d_writedata -> mm_interconnect_0:manager_data_master_writedata
	signal manager_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:manager_instruction_master_readdata -> manager:i_readdata
	signal manager_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:manager_instruction_master_waitrequest -> manager:i_waitrequest
	signal manager_instruction_master_address                                  : std_logic_vector(29 downto 0); -- manager:i_address -> mm_interconnect_0:manager_instruction_master_address
	signal manager_instruction_master_read                                     : std_logic;                     -- manager:i_read -> mm_interconnect_0:manager_instruction_master_read
	signal manager_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:manager_instruction_master_readdatavalid -> manager:i_readdatavalid
	signal worker3_wout_waitrequest                                            : std_logic;                     -- mm_interconnect_0:worker3_wout_waitrequest -> worker3:wout_waitrequest
	signal worker3_wout_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:worker3_wout_readdata -> worker3:wout_readdata
	signal worker3_wout_debugaccess                                            : std_logic;                     -- worker3:wout_debugaccess -> mm_interconnect_0:worker3_wout_debugaccess
	signal worker3_wout_address                                                : std_logic_vector(27 downto 0); -- worker3:wout_address -> mm_interconnect_0:worker3_wout_address
	signal worker3_wout_read                                                   : std_logic;                     -- worker3:wout_read -> mm_interconnect_0:worker3_wout_read
	signal worker3_wout_byteenable                                             : std_logic_vector(3 downto 0);  -- worker3:wout_byteenable -> mm_interconnect_0:worker3_wout_byteenable
	signal worker3_wout_readdatavalid                                          : std_logic;                     -- mm_interconnect_0:worker3_wout_readdatavalid -> worker3:wout_readdatavalid
	signal worker3_wout_writedata                                              : std_logic_vector(31 downto 0); -- worker3:wout_writedata -> mm_interconnect_0:worker3_wout_writedata
	signal worker3_wout_write                                                  : std_logic;                     -- worker3:wout_write -> mm_interconnect_0:worker3_wout_write
	signal worker3_wout_burstcount                                             : std_logic_vector(0 downto 0);  -- worker3:wout_burstcount -> mm_interconnect_0:worker3_wout_burstcount
	signal worker2_wout_waitrequest                                            : std_logic;                     -- mm_interconnect_0:worker2_wout_waitrequest -> worker2:wout_waitrequest
	signal worker2_wout_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:worker2_wout_readdata -> worker2:wout_readdata
	signal worker2_wout_debugaccess                                            : std_logic;                     -- worker2:wout_debugaccess -> mm_interconnect_0:worker2_wout_debugaccess
	signal worker2_wout_address                                                : std_logic_vector(27 downto 0); -- worker2:wout_address -> mm_interconnect_0:worker2_wout_address
	signal worker2_wout_read                                                   : std_logic;                     -- worker2:wout_read -> mm_interconnect_0:worker2_wout_read
	signal worker2_wout_byteenable                                             : std_logic_vector(3 downto 0);  -- worker2:wout_byteenable -> mm_interconnect_0:worker2_wout_byteenable
	signal worker2_wout_readdatavalid                                          : std_logic;                     -- mm_interconnect_0:worker2_wout_readdatavalid -> worker2:wout_readdatavalid
	signal worker2_wout_writedata                                              : std_logic_vector(31 downto 0); -- worker2:wout_writedata -> mm_interconnect_0:worker2_wout_writedata
	signal worker2_wout_write                                                  : std_logic;                     -- worker2:wout_write -> mm_interconnect_0:worker2_wout_write
	signal worker2_wout_burstcount                                             : std_logic_vector(0 downto 0);  -- worker2:wout_burstcount -> mm_interconnect_0:worker2_wout_burstcount
	signal worker1_wout_waitrequest                                            : std_logic;                     -- mm_interconnect_0:worker1_wout_waitrequest -> worker1:wout_waitrequest
	signal worker1_wout_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:worker1_wout_readdata -> worker1:wout_readdata
	signal worker1_wout_debugaccess                                            : std_logic;                     -- worker1:wout_debugaccess -> mm_interconnect_0:worker1_wout_debugaccess
	signal worker1_wout_address                                                : std_logic_vector(27 downto 0); -- worker1:wout_address -> mm_interconnect_0:worker1_wout_address
	signal worker1_wout_read                                                   : std_logic;                     -- worker1:wout_read -> mm_interconnect_0:worker1_wout_read
	signal worker1_wout_byteenable                                             : std_logic_vector(3 downto 0);  -- worker1:wout_byteenable -> mm_interconnect_0:worker1_wout_byteenable
	signal worker1_wout_readdatavalid                                          : std_logic;                     -- mm_interconnect_0:worker1_wout_readdatavalid -> worker1:wout_readdatavalid
	signal worker1_wout_writedata                                              : std_logic_vector(31 downto 0); -- worker1:wout_writedata -> mm_interconnect_0:worker1_wout_writedata
	signal worker1_wout_write                                                  : std_logic;                     -- worker1:wout_write -> mm_interconnect_0:worker1_wout_write
	signal worker1_wout_burstcount                                             : std_logic_vector(0 downto 0);  -- worker1:wout_burstcount -> mm_interconnect_0:worker1_wout_burstcount
	signal worker0_wout_waitrequest                                            : std_logic;                     -- mm_interconnect_0:worker0_wout_waitrequest -> worker0:wout_waitrequest
	signal worker0_wout_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:worker0_wout_readdata -> worker0:wout_readdata
	signal worker0_wout_debugaccess                                            : std_logic;                     -- worker0:wout_debugaccess -> mm_interconnect_0:worker0_wout_debugaccess
	signal worker0_wout_address                                                : std_logic_vector(27 downto 0); -- worker0:wout_address -> mm_interconnect_0:worker0_wout_address
	signal worker0_wout_read                                                   : std_logic;                     -- worker0:wout_read -> mm_interconnect_0:worker0_wout_read
	signal worker0_wout_byteenable                                             : std_logic_vector(3 downto 0);  -- worker0:wout_byteenable -> mm_interconnect_0:worker0_wout_byteenable
	signal worker0_wout_readdatavalid                                          : std_logic;                     -- mm_interconnect_0:worker0_wout_readdatavalid -> worker0:wout_readdatavalid
	signal worker0_wout_writedata                                              : std_logic_vector(31 downto 0); -- worker0:wout_writedata -> mm_interconnect_0:worker0_wout_writedata
	signal worker0_wout_write                                                  : std_logic;                     -- worker0:wout_write -> mm_interconnect_0:worker0_wout_write
	signal worker0_wout_burstcount                                             : std_logic_vector(0 downto 0);  -- worker0:wout_burstcount -> mm_interconnect_0:worker0_wout_burstcount
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect          : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata            : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest         : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write               : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_sender_readdata                : std_logic_vector(31 downto 0); -- mbox_m_w0:avmm_snd_readdata -> mm_interconnect_0:mbox_m_w0_avmm_msg_sender_readdata
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_sender_waitrequest             : std_logic;                     -- mbox_m_w0:avmm_snd_waitrequest -> mm_interconnect_0:mbox_m_w0_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_sender_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_m_w0_avmm_msg_sender_address -> mbox_m_w0:avmm_snd_address
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_sender_read                    : std_logic;                     -- mm_interconnect_0:mbox_m_w0_avmm_msg_sender_read -> mbox_m_w0:avmm_snd_read
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_sender_write                   : std_logic;                     -- mm_interconnect_0:mbox_m_w0_avmm_msg_sender_write -> mbox_m_w0:avmm_snd_write
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_sender_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_m_w0_avmm_msg_sender_writedata -> mbox_m_w0:avmm_snd_writedata
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_sender_readdata                : std_logic_vector(31 downto 0); -- mbox_m_w1:avmm_snd_readdata -> mm_interconnect_0:mbox_m_w1_avmm_msg_sender_readdata
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_sender_waitrequest             : std_logic;                     -- mbox_m_w1:avmm_snd_waitrequest -> mm_interconnect_0:mbox_m_w1_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_sender_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_m_w1_avmm_msg_sender_address -> mbox_m_w1:avmm_snd_address
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_sender_read                    : std_logic;                     -- mm_interconnect_0:mbox_m_w1_avmm_msg_sender_read -> mbox_m_w1:avmm_snd_read
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_sender_write                   : std_logic;                     -- mm_interconnect_0:mbox_m_w1_avmm_msg_sender_write -> mbox_m_w1:avmm_snd_write
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_sender_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_m_w1_avmm_msg_sender_writedata -> mbox_m_w1:avmm_snd_writedata
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_sender_readdata                : std_logic_vector(31 downto 0); -- mbox_m_w2:avmm_snd_readdata -> mm_interconnect_0:mbox_m_w2_avmm_msg_sender_readdata
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_sender_waitrequest             : std_logic;                     -- mbox_m_w2:avmm_snd_waitrequest -> mm_interconnect_0:mbox_m_w2_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_sender_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_m_w2_avmm_msg_sender_address -> mbox_m_w2:avmm_snd_address
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_sender_read                    : std_logic;                     -- mm_interconnect_0:mbox_m_w2_avmm_msg_sender_read -> mbox_m_w2:avmm_snd_read
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_sender_write                   : std_logic;                     -- mm_interconnect_0:mbox_m_w2_avmm_msg_sender_write -> mbox_m_w2:avmm_snd_write
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_sender_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_m_w2_avmm_msg_sender_writedata -> mbox_m_w2:avmm_snd_writedata
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_sender_readdata                : std_logic_vector(31 downto 0); -- mbox_m_w3:avmm_snd_readdata -> mm_interconnect_0:mbox_m_w3_avmm_msg_sender_readdata
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_sender_waitrequest             : std_logic;                     -- mbox_m_w3:avmm_snd_waitrequest -> mm_interconnect_0:mbox_m_w3_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_sender_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_m_w3_avmm_msg_sender_address -> mbox_m_w3:avmm_snd_address
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_sender_read                    : std_logic;                     -- mm_interconnect_0:mbox_m_w3_avmm_msg_sender_read -> mbox_m_w3:avmm_snd_read
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_sender_write                   : std_logic;                     -- mm_interconnect_0:mbox_m_w3_avmm_msg_sender_write -> mbox_m_w3:avmm_snd_write
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_sender_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_m_w3_avmm_msg_sender_writedata -> mbox_m_w3:avmm_snd_writedata
	signal mm_interconnect_0_performance_counter_0_control_slave_readdata      : std_logic_vector(31 downto 0); -- performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	signal mm_interconnect_0_performance_counter_0_control_slave_address       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	signal mm_interconnect_0_performance_counter_0_control_slave_begintransfer : std_logic;                     -- mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	signal mm_interconnect_0_performance_counter_0_control_slave_write         : std_logic;                     -- mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	signal mm_interconnect_0_performance_counter_0_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	signal mm_interconnect_0_manager_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- manager:debug_mem_slave_readdata -> mm_interconnect_0:manager_debug_mem_slave_readdata
	signal mm_interconnect_0_manager_debug_mem_slave_waitrequest               : std_logic;                     -- manager:debug_mem_slave_waitrequest -> mm_interconnect_0:manager_debug_mem_slave_waitrequest
	signal mm_interconnect_0_manager_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:manager_debug_mem_slave_debugaccess -> manager:debug_mem_slave_debugaccess
	signal mm_interconnect_0_manager_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:manager_debug_mem_slave_address -> manager:debug_mem_slave_address
	signal mm_interconnect_0_manager_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:manager_debug_mem_slave_read -> manager:debug_mem_slave_read
	signal mm_interconnect_0_manager_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:manager_debug_mem_slave_byteenable -> manager:debug_mem_slave_byteenable
	signal mm_interconnect_0_manager_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:manager_debug_mem_slave_write -> manager:debug_mem_slave_write
	signal mm_interconnect_0_manager_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:manager_debug_mem_slave_writedata -> manager:debug_mem_slave_writedata
	signal mm_interconnect_0_req_fifo_out_readdata                             : std_logic_vector(31 downto 0); -- req_fifo:avalonmm_read_slave_readdata -> mm_interconnect_0:req_fifo_out_readdata
	signal mm_interconnect_0_req_fifo_out_waitrequest                          : std_logic;                     -- req_fifo:avalonmm_read_slave_waitrequest -> mm_interconnect_0:req_fifo_out_waitrequest
	signal mm_interconnect_0_req_fifo_out_read                                 : std_logic;                     -- mm_interconnect_0:req_fifo_out_read -> req_fifo:avalonmm_read_slave_read
	signal mm_interconnect_0_req_fifo_out_csr_readdata                         : std_logic_vector(31 downto 0); -- req_fifo:rdclk_control_slave_readdata -> mm_interconnect_0:req_fifo_out_csr_readdata
	signal mm_interconnect_0_req_fifo_out_csr_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:req_fifo_out_csr_address -> req_fifo:rdclk_control_slave_address
	signal mm_interconnect_0_req_fifo_out_csr_read                             : std_logic;                     -- mm_interconnect_0:req_fifo_out_csr_read -> req_fifo:rdclk_control_slave_read
	signal mm_interconnect_0_req_fifo_out_csr_write                            : std_logic;                     -- mm_interconnect_0:req_fifo_out_csr_write -> req_fifo:rdclk_control_slave_write
	signal mm_interconnect_0_req_fifo_out_csr_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:req_fifo_out_csr_writedata -> req_fifo:rdclk_control_slave_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                       : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                           : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                          : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_shared_ocm_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:shared_ocm_s1_chipselect -> shared_ocm:chipselect
	signal mm_interconnect_0_shared_ocm_s1_readdata                            : std_logic_vector(31 downto 0); -- shared_ocm:readdata -> mm_interconnect_0:shared_ocm_s1_readdata
	signal mm_interconnect_0_shared_ocm_s1_address                             : std_logic_vector(7 downto 0);  -- mm_interconnect_0:shared_ocm_s1_address -> shared_ocm:address
	signal mm_interconnect_0_shared_ocm_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:shared_ocm_s1_byteenable -> shared_ocm:byteenable
	signal mm_interconnect_0_shared_ocm_s1_write                               : std_logic;                     -- mm_interconnect_0:shared_ocm_s1_write -> shared_ocm:write
	signal mm_interconnect_0_shared_ocm_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:shared_ocm_s1_writedata -> shared_ocm:writedata
	signal mm_interconnect_0_shared_ocm_s1_clken                               : std_logic;                     -- mm_interconnect_0:shared_ocm_s1_clken -> shared_ocm:clken
	signal mm_interconnect_0_sdram_0_sdout_readdata                            : std_logic_vector(31 downto 0); -- sdram_0:sdout_readdata -> mm_interconnect_0:sdram_0_sdout_readdata
	signal mm_interconnect_0_sdram_0_sdout_waitrequest                         : std_logic;                     -- sdram_0:sdout_waitrequest -> mm_interconnect_0:sdram_0_sdout_waitrequest
	signal mm_interconnect_0_sdram_0_sdout_debugaccess                         : std_logic;                     -- mm_interconnect_0:sdram_0_sdout_debugaccess -> sdram_0:sdout_debugaccess
	signal mm_interconnect_0_sdram_0_sdout_address                             : std_logic_vector(29 downto 0); -- mm_interconnect_0:sdram_0_sdout_address -> sdram_0:sdout_address
	signal mm_interconnect_0_sdram_0_sdout_read                                : std_logic;                     -- mm_interconnect_0:sdram_0_sdout_read -> sdram_0:sdout_read
	signal mm_interconnect_0_sdram_0_sdout_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sdram_0_sdout_byteenable -> sdram_0:sdout_byteenable
	signal mm_interconnect_0_sdram_0_sdout_readdatavalid                       : std_logic;                     -- sdram_0:sdout_readdatavalid -> mm_interconnect_0:sdram_0_sdout_readdatavalid
	signal mm_interconnect_0_sdram_0_sdout_write                               : std_logic;                     -- mm_interconnect_0:sdram_0_sdout_write -> sdram_0:sdout_write
	signal mm_interconnect_0_sdram_0_sdout_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_0_sdout_writedata -> sdram_0:sdout_writedata
	signal mm_interconnect_0_sdram_0_sdout_burstcount                          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sdram_0_sdout_burstcount -> sdram_0:sdout_burstcount
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_readdata              : std_logic_vector(31 downto 0); -- mbox_m_w0:avmm_rcv_readdata -> mm_interconnect_0:mbox_m_w0_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_m_w0_avmm_msg_receiver_address -> mbox_m_w0:avmm_rcv_address
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_read                  : std_logic;                     -- mm_interconnect_0:mbox_m_w0_avmm_msg_receiver_read -> mbox_m_w0:avmm_rcv_read
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_write                 : std_logic;                     -- mm_interconnect_0:mbox_m_w0_avmm_msg_receiver_write -> mbox_m_w0:avmm_rcv_write
	signal mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_m_w0_avmm_msg_receiver_writedata -> mbox_m_w0:avmm_rcv_writedata
	signal mm_interconnect_0_req_fifo_in_waitrequest                           : std_logic;                     -- req_fifo:avalonmm_write_slave_waitrequest -> mm_interconnect_0:req_fifo_in_waitrequest
	signal mm_interconnect_0_req_fifo_in_write                                 : std_logic;                     -- mm_interconnect_0:req_fifo_in_write -> req_fifo:avalonmm_write_slave_write
	signal mm_interconnect_0_req_fifo_in_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:req_fifo_in_writedata -> req_fifo:avalonmm_write_slave_writedata
	signal mm_interconnect_0_req_fifo_in_csr_readdata                          : std_logic_vector(31 downto 0); -- req_fifo:wrclk_control_slave_readdata -> mm_interconnect_0:req_fifo_in_csr_readdata
	signal mm_interconnect_0_req_fifo_in_csr_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:req_fifo_in_csr_address -> req_fifo:wrclk_control_slave_address
	signal mm_interconnect_0_req_fifo_in_csr_read                              : std_logic;                     -- mm_interconnect_0:req_fifo_in_csr_read -> req_fifo:wrclk_control_slave_read
	signal mm_interconnect_0_req_fifo_in_csr_write                             : std_logic;                     -- mm_interconnect_0:req_fifo_in_csr_write -> req_fifo:wrclk_control_slave_write
	signal mm_interconnect_0_req_fifo_in_csr_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:req_fifo_in_csr_writedata -> req_fifo:wrclk_control_slave_writedata
	signal mm_interconnect_0_shared_ocm_s2_chipselect                          : std_logic;                     -- mm_interconnect_0:shared_ocm_s2_chipselect -> shared_ocm:chipselect2
	signal mm_interconnect_0_shared_ocm_s2_readdata                            : std_logic_vector(31 downto 0); -- shared_ocm:readdata2 -> mm_interconnect_0:shared_ocm_s2_readdata
	signal mm_interconnect_0_shared_ocm_s2_address                             : std_logic_vector(7 downto 0);  -- mm_interconnect_0:shared_ocm_s2_address -> shared_ocm:address2
	signal mm_interconnect_0_shared_ocm_s2_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:shared_ocm_s2_byteenable -> shared_ocm:byteenable2
	signal mm_interconnect_0_shared_ocm_s2_write                               : std_logic;                     -- mm_interconnect_0:shared_ocm_s2_write -> shared_ocm:write2
	signal mm_interconnect_0_shared_ocm_s2_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:shared_ocm_s2_writedata -> shared_ocm:writedata2
	signal mm_interconnect_0_shared_ocm_s2_clken                               : std_logic;                     -- mm_interconnect_0:shared_ocm_s2_clken -> shared_ocm:clken2
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_readdata              : std_logic_vector(31 downto 0); -- mbox_m_w2:avmm_rcv_readdata -> mm_interconnect_0:mbox_m_w2_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_m_w2_avmm_msg_receiver_address -> mbox_m_w2:avmm_rcv_address
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_read                  : std_logic;                     -- mm_interconnect_0:mbox_m_w2_avmm_msg_receiver_read -> mbox_m_w2:avmm_rcv_read
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_write                 : std_logic;                     -- mm_interconnect_0:mbox_m_w2_avmm_msg_receiver_write -> mbox_m_w2:avmm_rcv_write
	signal mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_m_w2_avmm_msg_receiver_writedata -> mbox_m_w2:avmm_rcv_writedata
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_readdata              : std_logic_vector(31 downto 0); -- mbox_m_w1:avmm_rcv_readdata -> mm_interconnect_0:mbox_m_w1_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_m_w1_avmm_msg_receiver_address -> mbox_m_w1:avmm_rcv_address
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_read                  : std_logic;                     -- mm_interconnect_0:mbox_m_w1_avmm_msg_receiver_read -> mbox_m_w1:avmm_rcv_read
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_write                 : std_logic;                     -- mm_interconnect_0:mbox_m_w1_avmm_msg_receiver_write -> mbox_m_w1:avmm_rcv_write
	signal mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_m_w1_avmm_msg_receiver_writedata -> mbox_m_w1:avmm_rcv_writedata
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_readdata              : std_logic_vector(31 downto 0); -- mbox_m_w3:avmm_rcv_readdata -> mm_interconnect_0:mbox_m_w3_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mbox_m_w3_avmm_msg_receiver_address -> mbox_m_w3:avmm_rcv_address
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_read                  : std_logic;                     -- mm_interconnect_0:mbox_m_w3_avmm_msg_receiver_read -> mbox_m_w3:avmm_rcv_read
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_write                 : std_logic;                     -- mm_interconnect_0:mbox_m_w3_avmm_msg_receiver_write -> mbox_m_w3:avmm_rcv_write
	signal mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:mbox_m_w3_avmm_msg_receiver_writedata -> mbox_m_w3:avmm_rcv_writedata
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal manager_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> manager:irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:worker3_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal manager_debug_reset_request_reset                                   : std_logic;                     -- manager:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in1, rst_controller_006:reset_in1]
	signal rst_controller_002_reset_out_reset                                  : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:manager_reset_reset_bridge_in_reset_reset, mm_interconnect_0:sdram_0_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in, rst_translator:in_reset, shared_ocm:reset]
	signal rst_controller_002_reset_out_reset_req                              : std_logic;                     -- rst_controller_002:reset_req -> [manager:reset_req, rst_translator:reset_req_in, shared_ocm:reset_req]
	signal rst_controller_003_reset_out_reset                                  : std_logic;                     -- rst_controller_003:reset_out -> rst_controller_003_reset_out_reset:in
	signal rst_controller_004_reset_out_reset                                  : std_logic;                     -- rst_controller_004:reset_out -> rst_controller_004_reset_out_reset:in
	signal rst_controller_005_reset_out_reset                                  : std_logic;                     -- rst_controller_005:reset_out -> rst_controller_005_reset_out_reset:in
	signal rst_controller_006_reset_out_reset                                  : std_logic;                     -- rst_controller_006:reset_out -> rst_controller_006_reset_out_reset:in
	signal reset_reset_n_ports_inv                                             : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv     : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal rst_controller_001_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [jtag_uart_0:rst_n, mbox_m_w0:rst_n, mbox_m_w1:rst_n, mbox_m_w2:rst_n, mbox_m_w3:rst_n, performance_counter_0:reset_n, req_fifo:rdreset_n, req_fifo:wrreset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> manager:reset_n
	signal rst_controller_003_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> worker0:reset_reset_n
	signal rst_controller_004_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_004_reset_out_reset:inv -> worker1:reset_reset_n
	signal rst_controller_005_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_005_reset_out_reset:inv -> worker2:reset_reset_n
	signal rst_controller_006_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_006_reset_out_reset:inv -> worker3:reset_reset_n

begin

	altpll_0 : component system_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                 -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => altpll_0_c0_clk,                                --                    c0.clk
			c1                 => sdram_clk_clk,                                  --                    c1.clk
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			areset             => '0',                                            --           (terminated)
			locked             => open,                                           --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "0000",                                         --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	jtag_uart_0 : component system_jtag_uart_0
		port map (
			clk            => altpll_0_c0_clk,                                                 --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	manager : component system_manager
		port map (
			clk                                 => altpll_0_c0_clk,                                       --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,                --                          .reset_req
			d_address                           => manager_data_master_address,                           --               data_master.address
			d_byteenable                        => manager_data_master_byteenable,                        --                          .byteenable
			d_read                              => manager_data_master_read,                              --                          .read
			d_readdata                          => manager_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => manager_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => manager_data_master_write,                             --                          .write
			d_writedata                         => manager_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => manager_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => manager_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => manager_instruction_master_address,                    --        instruction_master.address
			i_read                              => manager_instruction_master_read,                       --                          .read
			i_readdata                          => manager_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => manager_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => manager_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => manager_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => manager_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_manager_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_manager_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_manager_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_manager_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_manager_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_manager_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_manager_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_manager_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	mbox_m_w0 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => altpll_0_c0_clk,                                         --               clk.clk
			rst_n                => rst_controller_001_reset_out_reset_ports_inv,            --             rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_address,     --   avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_writedata,   --                  .writedata
			avmm_snd_write       => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_write,       --                  .write
			avmm_snd_read        => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_read,        --                  .read
			avmm_snd_readdata    => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_readdata,    --                  .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_waitrequest, --                  .waitrequest
			avmm_rcv_address     => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_address,   -- avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_read,      --                  .read
			avmm_rcv_writedata   => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_writedata, --                  .writedata
			avmm_rcv_write       => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_write,     --                  .write
			avmm_rcv_readdata    => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_readdata,  --                  .readdata
			irq_space            => open,                                                    --       (terminated)
			irq_msg              => open                                                     --       (terminated)
		);

	mbox_m_w1 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => altpll_0_c0_clk,                                         --               clk.clk
			rst_n                => rst_controller_001_reset_out_reset_ports_inv,            --             rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_address,     --   avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_writedata,   --                  .writedata
			avmm_snd_write       => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_write,       --                  .write
			avmm_snd_read        => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_read,        --                  .read
			avmm_snd_readdata    => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_readdata,    --                  .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_waitrequest, --                  .waitrequest
			avmm_rcv_address     => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_address,   -- avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_read,      --                  .read
			avmm_rcv_writedata   => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_writedata, --                  .writedata
			avmm_rcv_write       => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_write,     --                  .write
			avmm_rcv_readdata    => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_readdata,  --                  .readdata
			irq_space            => open,                                                    --       (terminated)
			irq_msg              => open                                                     --       (terminated)
		);

	mbox_m_w2 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => altpll_0_c0_clk,                                         --               clk.clk
			rst_n                => rst_controller_001_reset_out_reset_ports_inv,            --             rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_address,     --   avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_writedata,   --                  .writedata
			avmm_snd_write       => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_write,       --                  .write
			avmm_snd_read        => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_read,        --                  .read
			avmm_snd_readdata    => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_readdata,    --                  .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_waitrequest, --                  .waitrequest
			avmm_rcv_address     => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_address,   -- avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_read,      --                  .read
			avmm_rcv_writedata   => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_writedata, --                  .writedata
			avmm_rcv_write       => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_write,     --                  .write
			avmm_rcv_readdata    => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_readdata,  --                  .readdata
			irq_space            => open,                                                    --       (terminated)
			irq_msg              => open                                                     --       (terminated)
		);

	mbox_m_w3 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => altpll_0_c0_clk,                                         --               clk.clk
			rst_n                => rst_controller_001_reset_out_reset_ports_inv,            --             rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_address,     --   avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_writedata,   --                  .writedata
			avmm_snd_write       => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_write,       --                  .write
			avmm_snd_read        => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_read,        --                  .read
			avmm_snd_readdata    => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_readdata,    --                  .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_waitrequest, --                  .waitrequest
			avmm_rcv_address     => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_address,   -- avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_read,      --                  .read
			avmm_rcv_writedata   => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_writedata, --                  .writedata
			avmm_rcv_write       => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_write,     --                  .write
			avmm_rcv_readdata    => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_readdata,  --                  .readdata
			irq_space            => open,                                                    --       (terminated)
			irq_msg              => open                                                     --       (terminated)
		);

	performance_counter_0 : component system_performance_counter_0
		port map (
			clk           => altpll_0_c0_clk,                                                     --           clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,                        --         reset.reset_n
			address       => mm_interconnect_0_performance_counter_0_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_performance_counter_0_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_performance_counter_0_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_performance_counter_0_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_performance_counter_0_control_slave_writedata      --              .writedata
		);

	req_fifo : component system_req_fifo
		port map (
			wrclock                          => altpll_0_c0_clk,                              --    clk_in.clk
			wrreset_n                        => rst_controller_001_reset_out_reset_ports_inv, --  reset_in.reset_n
			rdclock                          => altpll_0_c0_clk,                              --   clk_out.clk
			rdreset_n                        => rst_controller_001_reset_out_reset_ports_inv, -- reset_out.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_0_req_fifo_in_writedata,      --        in.writedata
			avalonmm_write_slave_write       => mm_interconnect_0_req_fifo_in_write,          --          .write
			avalonmm_write_slave_waitrequest => mm_interconnect_0_req_fifo_in_waitrequest,    --          .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_0_req_fifo_out_readdata,      --       out.readdata
			avalonmm_read_slave_read         => mm_interconnect_0_req_fifo_out_read,          --          .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_0_req_fifo_out_waitrequest,   --          .waitrequest
			rdclk_control_slave_address      => mm_interconnect_0_req_fifo_out_csr_address,   --   out_csr.address
			rdclk_control_slave_read         => mm_interconnect_0_req_fifo_out_csr_read,      --          .read
			rdclk_control_slave_writedata    => mm_interconnect_0_req_fifo_out_csr_writedata, --          .writedata
			rdclk_control_slave_write        => mm_interconnect_0_req_fifo_out_csr_write,     --          .write
			rdclk_control_slave_readdata     => mm_interconnect_0_req_fifo_out_csr_readdata,  --          .readdata
			wrclk_control_slave_address      => mm_interconnect_0_req_fifo_in_csr_address,    --    in_csr.address
			wrclk_control_slave_read         => mm_interconnect_0_req_fifo_in_csr_read,       --          .read
			wrclk_control_slave_writedata    => mm_interconnect_0_req_fifo_in_csr_writedata,  --          .writedata
			wrclk_control_slave_write        => mm_interconnect_0_req_fifo_in_csr_write,      --          .write
			wrclk_control_slave_readdata     => mm_interconnect_0_req_fifo_in_csr_readdata    --          .readdata
		);

	sdram_0 : component system_sdram_0
		port map (
			clk_clk             => altpll_0_c0_clk,                               --   clk.clk
			reset_reset_n       => reset_reset_n,                                 -- reset.reset_n
			sdout_waitrequest   => mm_interconnect_0_sdram_0_sdout_waitrequest,   -- sdout.waitrequest
			sdout_readdata      => mm_interconnect_0_sdram_0_sdout_readdata,      --      .readdata
			sdout_readdatavalid => mm_interconnect_0_sdram_0_sdout_readdatavalid, --      .readdatavalid
			sdout_burstcount    => mm_interconnect_0_sdram_0_sdout_burstcount,    --      .burstcount
			sdout_writedata     => mm_interconnect_0_sdram_0_sdout_writedata,     --      .writedata
			sdout_address       => mm_interconnect_0_sdram_0_sdout_address,       --      .address
			sdout_write         => mm_interconnect_0_sdram_0_sdout_write,         --      .write
			sdout_read          => mm_interconnect_0_sdram_0_sdout_read,          --      .read
			sdout_byteenable    => mm_interconnect_0_sdram_0_sdout_byteenable,    --      .byteenable
			sdout_debugaccess   => mm_interconnect_0_sdram_0_sdout_debugaccess,   --      .debugaccess
			sdram_addr          => wire_addr,                                     -- sdram.addr
			sdram_ba            => wire_ba,                                       --      .ba
			sdram_cas_n         => wire_cas_n,                                    --      .cas_n
			sdram_cke           => wire_cke,                                      --      .cke
			sdram_cs_n          => wire_cs_n,                                     --      .cs_n
			sdram_dq            => wire_dq,                                       --      .dq
			sdram_dqm           => wire_dqm,                                      --      .dqm
			sdram_ras_n         => wire_ras_n,                                    --      .ras_n
			sdram_we_n          => wire_we_n                                      --      .we_n
		);

	shared_ocm : component system_shared_ocm
		port map (
			address     => mm_interconnect_0_shared_ocm_s1_address,    --     s1.address
			clken       => mm_interconnect_0_shared_ocm_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_shared_ocm_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_shared_ocm_s1_write,      --       .write
			readdata    => mm_interconnect_0_shared_ocm_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_shared_ocm_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_shared_ocm_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_0_shared_ocm_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_shared_ocm_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_shared_ocm_s2_clken,      --       .clken
			write2      => mm_interconnect_0_shared_ocm_s2_write,      --       .write
			readdata2   => mm_interconnect_0_shared_ocm_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_shared_ocm_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_shared_ocm_s2_byteenable, --       .byteenable
			clk         => altpll_0_c0_clk,                            --   clk1.clk
			reset       => rst_controller_002_reset_out_reset,         -- reset1.reset
			reset_req   => rst_controller_002_reset_out_reset_req,     --       .reset_req
			freeze      => '0'                                         -- (terminated)
		);

	worker0 : component system_worker0
		port map (
			clk_clk            => altpll_0_c0_clk,                              --   clk.clk
			reset_reset_n      => rst_controller_003_reset_out_reset_ports_inv, -- reset.reset_n
			wout_waitrequest   => worker0_wout_waitrequest,                     --  wout.waitrequest
			wout_readdata      => worker0_wout_readdata,                        --      .readdata
			wout_readdatavalid => worker0_wout_readdatavalid,                   --      .readdatavalid
			wout_burstcount    => worker0_wout_burstcount,                      --      .burstcount
			wout_writedata     => worker0_wout_writedata,                       --      .writedata
			wout_address       => worker0_wout_address,                         --      .address
			wout_write         => worker0_wout_write,                           --      .write
			wout_read          => worker0_wout_read,                            --      .read
			wout_byteenable    => worker0_wout_byteenable,                      --      .byteenable
			wout_debugaccess   => worker0_wout_debugaccess                      --      .debugaccess
		);

	worker1 : component system_worker1
		port map (
			clk_clk            => altpll_0_c0_clk,                              --   clk.clk
			reset_reset_n      => rst_controller_004_reset_out_reset_ports_inv, -- reset.reset_n
			wout_waitrequest   => worker1_wout_waitrequest,                     --  wout.waitrequest
			wout_readdata      => worker1_wout_readdata,                        --      .readdata
			wout_readdatavalid => worker1_wout_readdatavalid,                   --      .readdatavalid
			wout_burstcount    => worker1_wout_burstcount,                      --      .burstcount
			wout_writedata     => worker1_wout_writedata,                       --      .writedata
			wout_address       => worker1_wout_address,                         --      .address
			wout_write         => worker1_wout_write,                           --      .write
			wout_read          => worker1_wout_read,                            --      .read
			wout_byteenable    => worker1_wout_byteenable,                      --      .byteenable
			wout_debugaccess   => worker1_wout_debugaccess                      --      .debugaccess
		);

	worker2 : component system_worker2
		port map (
			clk_clk            => altpll_0_c0_clk,                              --   clk.clk
			reset_reset_n      => rst_controller_005_reset_out_reset_ports_inv, -- reset.reset_n
			wout_waitrequest   => worker2_wout_waitrequest,                     --  wout.waitrequest
			wout_readdata      => worker2_wout_readdata,                        --      .readdata
			wout_readdatavalid => worker2_wout_readdatavalid,                   --      .readdatavalid
			wout_burstcount    => worker2_wout_burstcount,                      --      .burstcount
			wout_writedata     => worker2_wout_writedata,                       --      .writedata
			wout_address       => worker2_wout_address,                         --      .address
			wout_write         => worker2_wout_write,                           --      .write
			wout_read          => worker2_wout_read,                            --      .read
			wout_byteenable    => worker2_wout_byteenable,                      --      .byteenable
			wout_debugaccess   => worker2_wout_debugaccess                      --      .debugaccess
		);

	worker3 : component system_worker3
		port map (
			clk_clk            => altpll_0_c0_clk,                              --   clk.clk
			reset_reset_n      => rst_controller_006_reset_out_reset_ports_inv, -- reset.reset_n
			wout_waitrequest   => worker3_wout_waitrequest,                     --  wout.waitrequest
			wout_readdata      => worker3_wout_readdata,                        --      .readdata
			wout_readdatavalid => worker3_wout_readdatavalid,                   --      .readdatavalid
			wout_burstcount    => worker3_wout_burstcount,                      --      .burstcount
			wout_writedata     => worker3_wout_writedata,                       --      .writedata
			wout_address       => worker3_wout_address,                         --      .address
			wout_write         => worker3_wout_write,                           --      .write
			wout_read          => worker3_wout_read,                            --      .read
			wout_byteenable    => worker3_wout_byteenable,                      --      .byteenable
			wout_debugaccess   => worker3_wout_debugaccess                      --      .debugaccess
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                            => altpll_0_c0_clk,                                                     --                                          altpll_0_c0.clk
			clk_0_clk_clk                                              => clk_clk,                                                             --                                            clk_0_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                      -- altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset              => rst_controller_001_reset_out_reset,                                  --              jtag_uart_0_reset_reset_bridge_in_reset.reset
			manager_reset_reset_bridge_in_reset_reset                  => rst_controller_002_reset_out_reset,                                  --                  manager_reset_reset_bridge_in_reset.reset
			sdram_0_reset_reset_bridge_in_reset_reset                  => rst_controller_002_reset_out_reset,                                  --                  sdram_0_reset_reset_bridge_in_reset.reset
			worker3_reset_reset_bridge_in_reset_reset                  => rst_controller_001_reset_out_reset,                                  --                  worker3_reset_reset_bridge_in_reset.reset
			manager_data_master_address                                => manager_data_master_address,                                         --                                  manager_data_master.address
			manager_data_master_waitrequest                            => manager_data_master_waitrequest,                                     --                                                     .waitrequest
			manager_data_master_byteenable                             => manager_data_master_byteenable,                                      --                                                     .byteenable
			manager_data_master_read                                   => manager_data_master_read,                                            --                                                     .read
			manager_data_master_readdata                               => manager_data_master_readdata,                                        --                                                     .readdata
			manager_data_master_readdatavalid                          => manager_data_master_readdatavalid,                                   --                                                     .readdatavalid
			manager_data_master_write                                  => manager_data_master_write,                                           --                                                     .write
			manager_data_master_writedata                              => manager_data_master_writedata,                                       --                                                     .writedata
			manager_data_master_debugaccess                            => manager_data_master_debugaccess,                                     --                                                     .debugaccess
			manager_instruction_master_address                         => manager_instruction_master_address,                                  --                           manager_instruction_master.address
			manager_instruction_master_waitrequest                     => manager_instruction_master_waitrequest,                              --                                                     .waitrequest
			manager_instruction_master_read                            => manager_instruction_master_read,                                     --                                                     .read
			manager_instruction_master_readdata                        => manager_instruction_master_readdata,                                 --                                                     .readdata
			manager_instruction_master_readdatavalid                   => manager_instruction_master_readdatavalid,                            --                                                     .readdatavalid
			worker0_wout_address                                       => worker0_wout_address,                                                --                                         worker0_wout.address
			worker0_wout_waitrequest                                   => worker0_wout_waitrequest,                                            --                                                     .waitrequest
			worker0_wout_burstcount                                    => worker0_wout_burstcount,                                             --                                                     .burstcount
			worker0_wout_byteenable                                    => worker0_wout_byteenable,                                             --                                                     .byteenable
			worker0_wout_read                                          => worker0_wout_read,                                                   --                                                     .read
			worker0_wout_readdata                                      => worker0_wout_readdata,                                               --                                                     .readdata
			worker0_wout_readdatavalid                                 => worker0_wout_readdatavalid,                                          --                                                     .readdatavalid
			worker0_wout_write                                         => worker0_wout_write,                                                  --                                                     .write
			worker0_wout_writedata                                     => worker0_wout_writedata,                                              --                                                     .writedata
			worker0_wout_debugaccess                                   => worker0_wout_debugaccess,                                            --                                                     .debugaccess
			worker1_wout_address                                       => worker1_wout_address,                                                --                                         worker1_wout.address
			worker1_wout_waitrequest                                   => worker1_wout_waitrequest,                                            --                                                     .waitrequest
			worker1_wout_burstcount                                    => worker1_wout_burstcount,                                             --                                                     .burstcount
			worker1_wout_byteenable                                    => worker1_wout_byteenable,                                             --                                                     .byteenable
			worker1_wout_read                                          => worker1_wout_read,                                                   --                                                     .read
			worker1_wout_readdata                                      => worker1_wout_readdata,                                               --                                                     .readdata
			worker1_wout_readdatavalid                                 => worker1_wout_readdatavalid,                                          --                                                     .readdatavalid
			worker1_wout_write                                         => worker1_wout_write,                                                  --                                                     .write
			worker1_wout_writedata                                     => worker1_wout_writedata,                                              --                                                     .writedata
			worker1_wout_debugaccess                                   => worker1_wout_debugaccess,                                            --                                                     .debugaccess
			worker2_wout_address                                       => worker2_wout_address,                                                --                                         worker2_wout.address
			worker2_wout_waitrequest                                   => worker2_wout_waitrequest,                                            --                                                     .waitrequest
			worker2_wout_burstcount                                    => worker2_wout_burstcount,                                             --                                                     .burstcount
			worker2_wout_byteenable                                    => worker2_wout_byteenable,                                             --                                                     .byteenable
			worker2_wout_read                                          => worker2_wout_read,                                                   --                                                     .read
			worker2_wout_readdata                                      => worker2_wout_readdata,                                               --                                                     .readdata
			worker2_wout_readdatavalid                                 => worker2_wout_readdatavalid,                                          --                                                     .readdatavalid
			worker2_wout_write                                         => worker2_wout_write,                                                  --                                                     .write
			worker2_wout_writedata                                     => worker2_wout_writedata,                                              --                                                     .writedata
			worker2_wout_debugaccess                                   => worker2_wout_debugaccess,                                            --                                                     .debugaccess
			worker3_wout_address                                       => worker3_wout_address,                                                --                                         worker3_wout.address
			worker3_wout_waitrequest                                   => worker3_wout_waitrequest,                                            --                                                     .waitrequest
			worker3_wout_burstcount                                    => worker3_wout_burstcount,                                             --                                                     .burstcount
			worker3_wout_byteenable                                    => worker3_wout_byteenable,                                             --                                                     .byteenable
			worker3_wout_read                                          => worker3_wout_read,                                                   --                                                     .read
			worker3_wout_readdata                                      => worker3_wout_readdata,                                               --                                                     .readdata
			worker3_wout_readdatavalid                                 => worker3_wout_readdatavalid,                                          --                                                     .readdatavalid
			worker3_wout_write                                         => worker3_wout_write,                                                  --                                                     .write
			worker3_wout_writedata                                     => worker3_wout_writedata,                                              --                                                     .writedata
			worker3_wout_debugaccess                                   => worker3_wout_debugaccess,                                            --                                                     .debugaccess
			altpll_0_pll_slave_address                                 => mm_interconnect_0_altpll_0_pll_slave_address,                        --                                   altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                   => mm_interconnect_0_altpll_0_pll_slave_write,                          --                                                     .write
			altpll_0_pll_slave_read                                    => mm_interconnect_0_altpll_0_pll_slave_read,                           --                                                     .read
			altpll_0_pll_slave_readdata                                => mm_interconnect_0_altpll_0_pll_slave_readdata,                       --                                                     .readdata
			altpll_0_pll_slave_writedata                               => mm_interconnect_0_altpll_0_pll_slave_writedata,                      --                                                     .writedata
			jtag_uart_0_avalon_jtag_slave_address                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,             --                        jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,               --                                                     .write
			jtag_uart_0_avalon_jtag_slave_read                         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                --                                                     .read
			jtag_uart_0_avalon_jtag_slave_readdata                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,            --                                                     .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,           --                                                     .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,         --                                                     .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,          --                                                     .chipselect
			manager_debug_mem_slave_address                            => mm_interconnect_0_manager_debug_mem_slave_address,                   --                              manager_debug_mem_slave.address
			manager_debug_mem_slave_write                              => mm_interconnect_0_manager_debug_mem_slave_write,                     --                                                     .write
			manager_debug_mem_slave_read                               => mm_interconnect_0_manager_debug_mem_slave_read,                      --                                                     .read
			manager_debug_mem_slave_readdata                           => mm_interconnect_0_manager_debug_mem_slave_readdata,                  --                                                     .readdata
			manager_debug_mem_slave_writedata                          => mm_interconnect_0_manager_debug_mem_slave_writedata,                 --                                                     .writedata
			manager_debug_mem_slave_byteenable                         => mm_interconnect_0_manager_debug_mem_slave_byteenable,                --                                                     .byteenable
			manager_debug_mem_slave_waitrequest                        => mm_interconnect_0_manager_debug_mem_slave_waitrequest,               --                                                     .waitrequest
			manager_debug_mem_slave_debugaccess                        => mm_interconnect_0_manager_debug_mem_slave_debugaccess,               --                                                     .debugaccess
			mbox_m_w0_avmm_msg_receiver_address                        => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_address,               --                          mbox_m_w0_avmm_msg_receiver.address
			mbox_m_w0_avmm_msg_receiver_write                          => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_write,                 --                                                     .write
			mbox_m_w0_avmm_msg_receiver_read                           => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_read,                  --                                                     .read
			mbox_m_w0_avmm_msg_receiver_readdata                       => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_readdata,              --                                                     .readdata
			mbox_m_w0_avmm_msg_receiver_writedata                      => mm_interconnect_0_mbox_m_w0_avmm_msg_receiver_writedata,             --                                                     .writedata
			mbox_m_w0_avmm_msg_sender_address                          => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_address,                 --                            mbox_m_w0_avmm_msg_sender.address
			mbox_m_w0_avmm_msg_sender_write                            => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_write,                   --                                                     .write
			mbox_m_w0_avmm_msg_sender_read                             => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_read,                    --                                                     .read
			mbox_m_w0_avmm_msg_sender_readdata                         => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_readdata,                --                                                     .readdata
			mbox_m_w0_avmm_msg_sender_writedata                        => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_writedata,               --                                                     .writedata
			mbox_m_w0_avmm_msg_sender_waitrequest                      => mm_interconnect_0_mbox_m_w0_avmm_msg_sender_waitrequest,             --                                                     .waitrequest
			mbox_m_w1_avmm_msg_receiver_address                        => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_address,               --                          mbox_m_w1_avmm_msg_receiver.address
			mbox_m_w1_avmm_msg_receiver_write                          => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_write,                 --                                                     .write
			mbox_m_w1_avmm_msg_receiver_read                           => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_read,                  --                                                     .read
			mbox_m_w1_avmm_msg_receiver_readdata                       => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_readdata,              --                                                     .readdata
			mbox_m_w1_avmm_msg_receiver_writedata                      => mm_interconnect_0_mbox_m_w1_avmm_msg_receiver_writedata,             --                                                     .writedata
			mbox_m_w1_avmm_msg_sender_address                          => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_address,                 --                            mbox_m_w1_avmm_msg_sender.address
			mbox_m_w1_avmm_msg_sender_write                            => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_write,                   --                                                     .write
			mbox_m_w1_avmm_msg_sender_read                             => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_read,                    --                                                     .read
			mbox_m_w1_avmm_msg_sender_readdata                         => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_readdata,                --                                                     .readdata
			mbox_m_w1_avmm_msg_sender_writedata                        => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_writedata,               --                                                     .writedata
			mbox_m_w1_avmm_msg_sender_waitrequest                      => mm_interconnect_0_mbox_m_w1_avmm_msg_sender_waitrequest,             --                                                     .waitrequest
			mbox_m_w2_avmm_msg_receiver_address                        => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_address,               --                          mbox_m_w2_avmm_msg_receiver.address
			mbox_m_w2_avmm_msg_receiver_write                          => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_write,                 --                                                     .write
			mbox_m_w2_avmm_msg_receiver_read                           => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_read,                  --                                                     .read
			mbox_m_w2_avmm_msg_receiver_readdata                       => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_readdata,              --                                                     .readdata
			mbox_m_w2_avmm_msg_receiver_writedata                      => mm_interconnect_0_mbox_m_w2_avmm_msg_receiver_writedata,             --                                                     .writedata
			mbox_m_w2_avmm_msg_sender_address                          => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_address,                 --                            mbox_m_w2_avmm_msg_sender.address
			mbox_m_w2_avmm_msg_sender_write                            => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_write,                   --                                                     .write
			mbox_m_w2_avmm_msg_sender_read                             => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_read,                    --                                                     .read
			mbox_m_w2_avmm_msg_sender_readdata                         => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_readdata,                --                                                     .readdata
			mbox_m_w2_avmm_msg_sender_writedata                        => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_writedata,               --                                                     .writedata
			mbox_m_w2_avmm_msg_sender_waitrequest                      => mm_interconnect_0_mbox_m_w2_avmm_msg_sender_waitrequest,             --                                                     .waitrequest
			mbox_m_w3_avmm_msg_receiver_address                        => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_address,               --                          mbox_m_w3_avmm_msg_receiver.address
			mbox_m_w3_avmm_msg_receiver_write                          => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_write,                 --                                                     .write
			mbox_m_w3_avmm_msg_receiver_read                           => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_read,                  --                                                     .read
			mbox_m_w3_avmm_msg_receiver_readdata                       => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_readdata,              --                                                     .readdata
			mbox_m_w3_avmm_msg_receiver_writedata                      => mm_interconnect_0_mbox_m_w3_avmm_msg_receiver_writedata,             --                                                     .writedata
			mbox_m_w3_avmm_msg_sender_address                          => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_address,                 --                            mbox_m_w3_avmm_msg_sender.address
			mbox_m_w3_avmm_msg_sender_write                            => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_write,                   --                                                     .write
			mbox_m_w3_avmm_msg_sender_read                             => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_read,                    --                                                     .read
			mbox_m_w3_avmm_msg_sender_readdata                         => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_readdata,                --                                                     .readdata
			mbox_m_w3_avmm_msg_sender_writedata                        => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_writedata,               --                                                     .writedata
			mbox_m_w3_avmm_msg_sender_waitrequest                      => mm_interconnect_0_mbox_m_w3_avmm_msg_sender_waitrequest,             --                                                     .waitrequest
			performance_counter_0_control_slave_address                => mm_interconnect_0_performance_counter_0_control_slave_address,       --                  performance_counter_0_control_slave.address
			performance_counter_0_control_slave_write                  => mm_interconnect_0_performance_counter_0_control_slave_write,         --                                                     .write
			performance_counter_0_control_slave_readdata               => mm_interconnect_0_performance_counter_0_control_slave_readdata,      --                                                     .readdata
			performance_counter_0_control_slave_writedata              => mm_interconnect_0_performance_counter_0_control_slave_writedata,     --                                                     .writedata
			performance_counter_0_control_slave_begintransfer          => mm_interconnect_0_performance_counter_0_control_slave_begintransfer, --                                                     .begintransfer
			req_fifo_in_write                                          => mm_interconnect_0_req_fifo_in_write,                                 --                                          req_fifo_in.write
			req_fifo_in_writedata                                      => mm_interconnect_0_req_fifo_in_writedata,                             --                                                     .writedata
			req_fifo_in_waitrequest                                    => mm_interconnect_0_req_fifo_in_waitrequest,                           --                                                     .waitrequest
			req_fifo_in_csr_address                                    => mm_interconnect_0_req_fifo_in_csr_address,                           --                                      req_fifo_in_csr.address
			req_fifo_in_csr_write                                      => mm_interconnect_0_req_fifo_in_csr_write,                             --                                                     .write
			req_fifo_in_csr_read                                       => mm_interconnect_0_req_fifo_in_csr_read,                              --                                                     .read
			req_fifo_in_csr_readdata                                   => mm_interconnect_0_req_fifo_in_csr_readdata,                          --                                                     .readdata
			req_fifo_in_csr_writedata                                  => mm_interconnect_0_req_fifo_in_csr_writedata,                         --                                                     .writedata
			req_fifo_out_read                                          => mm_interconnect_0_req_fifo_out_read,                                 --                                         req_fifo_out.read
			req_fifo_out_readdata                                      => mm_interconnect_0_req_fifo_out_readdata,                             --                                                     .readdata
			req_fifo_out_waitrequest                                   => mm_interconnect_0_req_fifo_out_waitrequest,                          --                                                     .waitrequest
			req_fifo_out_csr_address                                   => mm_interconnect_0_req_fifo_out_csr_address,                          --                                     req_fifo_out_csr.address
			req_fifo_out_csr_write                                     => mm_interconnect_0_req_fifo_out_csr_write,                            --                                                     .write
			req_fifo_out_csr_read                                      => mm_interconnect_0_req_fifo_out_csr_read,                             --                                                     .read
			req_fifo_out_csr_readdata                                  => mm_interconnect_0_req_fifo_out_csr_readdata,                         --                                                     .readdata
			req_fifo_out_csr_writedata                                 => mm_interconnect_0_req_fifo_out_csr_writedata,                        --                                                     .writedata
			sdram_0_sdout_address                                      => mm_interconnect_0_sdram_0_sdout_address,                             --                                        sdram_0_sdout.address
			sdram_0_sdout_write                                        => mm_interconnect_0_sdram_0_sdout_write,                               --                                                     .write
			sdram_0_sdout_read                                         => mm_interconnect_0_sdram_0_sdout_read,                                --                                                     .read
			sdram_0_sdout_readdata                                     => mm_interconnect_0_sdram_0_sdout_readdata,                            --                                                     .readdata
			sdram_0_sdout_writedata                                    => mm_interconnect_0_sdram_0_sdout_writedata,                           --                                                     .writedata
			sdram_0_sdout_burstcount                                   => mm_interconnect_0_sdram_0_sdout_burstcount,                          --                                                     .burstcount
			sdram_0_sdout_byteenable                                   => mm_interconnect_0_sdram_0_sdout_byteenable,                          --                                                     .byteenable
			sdram_0_sdout_readdatavalid                                => mm_interconnect_0_sdram_0_sdout_readdatavalid,                       --                                                     .readdatavalid
			sdram_0_sdout_waitrequest                                  => mm_interconnect_0_sdram_0_sdout_waitrequest,                         --                                                     .waitrequest
			sdram_0_sdout_debugaccess                                  => mm_interconnect_0_sdram_0_sdout_debugaccess,                         --                                                     .debugaccess
			shared_ocm_s1_address                                      => mm_interconnect_0_shared_ocm_s1_address,                             --                                        shared_ocm_s1.address
			shared_ocm_s1_write                                        => mm_interconnect_0_shared_ocm_s1_write,                               --                                                     .write
			shared_ocm_s1_readdata                                     => mm_interconnect_0_shared_ocm_s1_readdata,                            --                                                     .readdata
			shared_ocm_s1_writedata                                    => mm_interconnect_0_shared_ocm_s1_writedata,                           --                                                     .writedata
			shared_ocm_s1_byteenable                                   => mm_interconnect_0_shared_ocm_s1_byteenable,                          --                                                     .byteenable
			shared_ocm_s1_chipselect                                   => mm_interconnect_0_shared_ocm_s1_chipselect,                          --                                                     .chipselect
			shared_ocm_s1_clken                                        => mm_interconnect_0_shared_ocm_s1_clken,                               --                                                     .clken
			shared_ocm_s2_address                                      => mm_interconnect_0_shared_ocm_s2_address,                             --                                        shared_ocm_s2.address
			shared_ocm_s2_write                                        => mm_interconnect_0_shared_ocm_s2_write,                               --                                                     .write
			shared_ocm_s2_readdata                                     => mm_interconnect_0_shared_ocm_s2_readdata,                            --                                                     .readdata
			shared_ocm_s2_writedata                                    => mm_interconnect_0_shared_ocm_s2_writedata,                           --                                                     .writedata
			shared_ocm_s2_byteenable                                   => mm_interconnect_0_shared_ocm_s2_byteenable,                          --                                                     .byteenable
			shared_ocm_s2_chipselect                                   => mm_interconnect_0_shared_ocm_s2_chipselect,                          --                                                     .chipselect
			shared_ocm_s2_clken                                        => mm_interconnect_0_shared_ocm_s2_clken                                --                                                     .clken
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => altpll_0_c0_clk,                    --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			sender_irq    => manager_irq_irq                     --    sender.irq
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => manager_debug_reset_request_reset,  -- reset_in1.reset
			clk            => altpll_0_c0_clk,                    --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => altpll_0_c0_clk,                        --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => manager_debug_reset_request_reset,  -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_004 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => manager_debug_reset_request_reset,  -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_005 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => manager_debug_reset_request_reset,  -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_006 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => manager_debug_reset_request_reset,  -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_006_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

	rst_controller_005_reset_out_reset_ports_inv <= not rst_controller_005_reset_out_reset;

	rst_controller_006_reset_out_reset_ports_inv <= not rst_controller_006_reset_out_reset;

end architecture rtl; -- of system
