// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
yjhF9tmiusg2zYcWlDXazovC/zc+++9SVRMQ2hJmFwts1PbPYIBoar+eS1r6cYxjsBxm3shLJvTE
NqFAkLzt+RAIBDROYdGH/dzlCtfXPC8n8sJZc6W1Ayfq0uW1PsPwtq3+yuyjB9W97TRfyTPperrc
ybTH8Bi/NfyGT4PNV4Ei6IEE8q/EbUxubSYSXCGp05qLSr0wIB6YBY9DdJJytCyLji4ramaCFBQD
bmZ+pK9Gtw/GGAU3iksPHmHloY7U961XcTJtVBtrGZoP6dHeQg4fvUpLJluPyaAvghXbz2PG0UUM
YocyntStT4QRbOwsoUWabTWQ626R6sAMXRtxhQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 93456)
CvGjzs81nPj6YlLPXMpwfHLuIiYxrp/oH+AjpbkrGxc1BWhIg3l8f/ZRcjCzwCkzhoTm5KaFlorl
SPkgtx3+acBBgu24oO5Na1i2iWs57dCjMw3rF/xcnhzIEkWapVXpZxKOAnRpgE3sw1CJnLVfLElp
fXSzBYqTyW/CY3KDBaH/O2LPSLawq7MFlQcD9XDfAg2AOBuwZbI/DttXrTawUblKg41ksAotdvPm
TyAIH57ZidINbaUZI0z7o75UdJ4o3bT6wCrkJEnHgC3L9kJAzuthin8I2JTiQelUl7Ovu9VLkCmD
1x0PaKN7AFFIEg2OsRZGlhcx8E/ZOt8IYPQ1J1p+r+3dWoe3/nLQnW5TQU3oYfBHaMS8HJv9iXa2
Ta2CdsqDYp9/crkn8Cr6Mdz7nompZXgicOcWdO81eErWfDgj6ySMksqJ2aRghXOiGt/dHk2QjUH4
94yOoJhLDGj3xJUjyRqtXUBbkHdEps5sZKfSepkXlKKig2fotoRRkNCI4ErLXt4jet10efh894k+
WNs0Ipjv7SL6mW42LhqEGS48L3Tsq78ba3rPdY5dP00bOPuL+aKbeeOFVRt4e7lYeTRzShsX28xQ
hIqmLNGUB1ddv2fKookXxEexD/pJIIZ4R1LvhOp6IrVHUO86+rMVx6SH7VDslK8+f/zECixCej+q
0KBsK6LZedQ1uuMvJUfz2l6lw5sfT+SuwO/7IvV89ae34cCV23md9TNnVzhn3N/6AykWRKFq4FVA
eo6ISB0ra4h8OgbLOe3j+xVa7TU56qrjf5USqHjpbaqQnENt7kZWzDBxR1hDQGsLqafN9XrupTJn
gfdyZfruJ6n/ggbcx/idnILumWuY52tT50f+MbJYV8tRPI1S3nQeepqyRAxtQs5YXwwjoAmYX+x/
RPqwOA50hk1MoJLN3wYeGty4aoP0rVRic0U3V3ynaTNY2+LbblNg550RY2wGSe0VDipSpZFTAuyP
PX5nCL64NQXEYTjxgCkzuXDMWHqS31FX8+jxmE2K7YeuudMCb6O4qbd5T7UO5z16ogynd7gqGA0A
1igve/38M3F76U0m4CTSEcnk/Am47lMY9kfuaOruyEA+KupAA8wkYfgsBKUVZc13oCbUWtaVCqO8
J3XfJ7ISNO/JKhRUw8uANv8CCjTPYp2bRhbc8MIWSspJnv54E2u8Av76J8ziekE7V2qd0WKoyo+D
47hNVgnl2hVN27P4KvQtA/KMbT0VgZCoV5EhEQIkgUpSlQq+3XAADEUgUKW9hgx4/u5itqHEqRBi
5JV8V9BBzEPt/8Czo9uPNNEmllH9IENvv9EWtyulKZIWo2iF6+W2xmZeSnNCT6Mc2fYcoRtvmd3W
ZpSpHNIiQy43YUe6D16bbuHqAovKZJJNUfmfvExpUV01wPb7wIAP+gcPBwoEKAXc+JoZK12JkvZF
j4WYm0N4i4SnsVVS/Ouh5dgndrLglZNisFD/FvKaHHJOZ0fdV2jAMZi/KxYH2kYq18I859Jr9ZUe
y8c2SMGhT5dYOxWOEK7wmU7ZWhSy+S10tRrPeQQOhuLTPSAyWEPs5t/9vBQx4Oq4dyZCCsZlxnUA
5HNgJQ9IZCH56xFjROIF6ldCnOYTvZtWHagGBtq3PzYlsMg7oyZYTblbQBPgMlExncMMJDWYusoS
08GavCxsIU/lij1Xlena1dMcbNOT5N6zhy1CFDCglJ+jh2gblQAh0GXDJIFdqbpH2gZ95GUy+koH
G5BEBf1sdOof7A24Txcg09/kzAlBQfTbEeYE0iI9exqH3s2j96IoeiAMh9WRW3PH1BkG/Z5ycnA6
b5J5uikOOc2wUbY8lAhDz0UMEDcILLZCW7y9+i9Dpl7nDTnP81zGln2eqzhpIC/RrXJU8ND7VUWu
5gWc4IQF7JDYahCWdeZDzwNMgu1LO46Z8oo833L0ZTRUnNyVXB3sLH+5NeW2Vnq22n9Jr/duNKaL
PMuzNedkQTveYqunjkTSicTLMvZ0sRwl67TgF0pUFx2NJ6X6UECnAUS2PE8q7RMh7vSrl99KDi0t
EB3e4btancn8DD7QOMD9imaHJM3uAOiuD0kjrZ7lXUJXanSAh2GSdWoFjcRoU4kDId4ymgVX2XE4
fE4L2bkDHrQbzV3VfnYrOyYx0Z4jeyiDm8gA5uvyfhSetTIkpwFjxjDc/0SZB4eMtqNkdlKoVZdS
tyxx81ve6jKo18nOUSdVvwJuxgGGd1NqeHsePiSGDdkKttMfYjCIADS/x0sBlDNVZ4n2E0l5Lhwb
soXjISrZcKx3S6dcQQeCKpolWaGwAu4xxRLIIeLTYEt+aIep9b3TsZLaZeDZTMu2xA9911KpSioT
wsONEXuTwDm0iQJJX3BgJCPbzohwCflRRnUPPoUZpCqb5qcRMKEnnErFAsNGPMo+l9fn7OWEMFOe
zXATMlmA1tNytlv1EACPBqkt/PHw8wF/sprEM+LxVyNDW5FYo/Vjkq5bOnkHx+vHj37liNV7YpEL
kTe9/KsX0Hvq9jZvbj9IzOBO6i60Gwcf8eHml4fuaoYTZX0fTU9pPNSwp11pDXD3me8fzjFI+Frb
jk0ctwqDamhAFRHIfqH0NMPPOgVXvI7fgU4LJgmNghGiHFTQPMlMqitSCAitc9pUFJ2WhkKAppZT
E/Et2rlyRpx3DCHl6r09qVA1rZ6edr7/qJcUCtFjVSSWLtbOQt4kBLZ/ue18qFujA4XilZlHh+2o
SmdfRJzZH36d5qYMKvkxeZh1RpUcSRyWVc7AkjijRcBK0DQEL6jwL4E23PLlGwE4LSDnuKTIRf0C
IeKeaiR8hd1337DCvwG7ikLDJhHyBceifkR1oW4vk1TJm6GgGEBR91OLFKoJZx6Ufwh40GKzB51M
YXJo9+Jag8JuBjyqDkIdIRyhukgkrAsHOTFhDkzXbIdZ3dtwLRL1OwlLeHsyVcN6TnYzr+iOg+vN
dydK6DJD89iNYA02Vi1DLRqIJsZsA6/004ewgOWVXzG39y1i/cSncSd/IiHjss9thtVHTshrfumI
U9C3UwjVTHACDYtW8O4YJQpt2sVQVH+h1b30hRhEIXsyuMXmR/RH0OM+SmGtrFDpkPiBfwVxEyqF
pwM6Jjv8xRAED4fD3yjY8AMbDtz0h2pFjGb2JvT4NM7xudgYzEHaeWA47Yk/37NV/a2Uo9VqMyo8
VpzGsr6bL8zloEuJO8uMydp0D4NGY4VfUv0jMuWTVXMcROgIpmiv8wQQErPiPMdOG5Fm7ZRV0ejE
iQUJXCHZ+14IODwBDtYYULZliypUzjcys7EAkrKqX4S/bmsqG4jxFwWCLhaGX+iHH0B8J8gIjqW7
+NqIWykxHz/B54i79IQZZlGCrBeLAQ+vSOdRp52Q7wPCahMrG1M8j1cpVi+beuvAOQj02mrsTCUv
vGrX0ZAvW83KjcbyudULeBvHKBWIVFL5XsVrSWcyfWTPTxLrbEkBbHAkpp7AWW8FBQCr8+MbR3iS
jAiq5cgM1nk7GOtZQ4OKPC0N/SGq8nNncfBuzi9fH2BjaBOcusFKvsSvB8YzYzgNrEkoe7FFtz+E
EUkKKRqdXq+DNv7ATK/nJcmq2c9HQ3DGuv0YG9pkib4WyaE/AB0RmudixJq9zI7HleXo4jCYbA0R
lKe7XtIYwDloQ5yY0z+0KGZsO2hgCAIa5rUxSmw2Q1gfRL6fPNwnOlzylTUBtIJRuv5osNGZmUvc
sv/exk0ukVbSYn+cuhGtvpo1clx+sYCxaTYToPV+qZguDUxf4u/dcJ/56m7J7Ph1cClRqGQY9mrL
OXBmAitXAnXDOsu7U9RG41/mXlRy1+E1QJHtFgjvkk5jBUUJ9K0U51Isu5jf2bmL540XZHshbYHQ
a3O+i3qkxVqWNQw1Xh715QB7Zge882cPoIEO5noti3NeYl/aW3I+q1kH4MprEDIuzfUAR/i+smPq
r9d5AG8cQ6t5lHhug0htla7rBzgWBApf2iBOaST77vu1uamyM4I6t231HqfpMhqCKlgpEmA5im2u
TjaFh9d2bzVziGL9j1WT54u63sY30SgZIN8aRK/21/1HzQFUuImca8e9Li6TbVcbmuKAmIJxTxK9
T9xZhJUCdfaBQLrInzprRLniV6S8AIAY/vQRKHvpiT1SVygVP9YKjJjjrp95689oiyI+DhyURtiu
rKxHG2PHZUrZB2+oQ29hJlDC1BV54aki9iK3+QJkRPvQPUcyG6gD16dBklUrjWh9Sf4P3ec7LVZZ
gw0kJDyWqDjeFrL4RcqRHFAW7qS/dcTS/lcRv1JsbdR4GsWuQH7sNxD4H+NzKdEWo47hWjLihQ/5
3F7UP8oEiFW0W4ovUHrW5QhSlZ3EdzdghmPkvlfEJEKdC/IwBiYGcAZXrp2wBskUQRzU4k9fCLqD
BtCQQj/vO4UID7C6daKKpuu1BwCU9cJdPPMBfLPOqftkWV4Q1RAH5mmpiTu16c6KjweCAvU8EFn2
gXsJHho6717ZAgJppdmjB+FKtU5tbdh89CneAOryN0/m8CRvJPvw1A08OL78GF1dHhO9UweinPTQ
r+RJXggmFrQasMuQTymzLpYm9L7GiS/WyenJLSgZiXt9mtLah/slUqgtOgnyUY/L5Rv4cqVuaatD
190mruygWSIUevqSyjKp7ltXM+pip7TkeE263BSKfTrdt6UBkZH2qT+VnZnvmQC0AUzOKI9SObsi
Qr8P6utvLo9ucMHO9/DgYh3oMoYlcvMgMvMd7gMQRkAkeOin6aWPQbmQ4ozqw5A6pgBznJercALE
EVTmIeUF91mZJ6Zqc1KtTPDE664SYO9LufrRgYASJjPp/i31H822Q5LbXjLSZDu5KjK4zDDDp6NW
69IX1ORDxrhmViV83IdbUUZ6z+ium16MpsMK10JcyB2DfIYztbhad1X1JWIe8boWk4LTbwbaEOqe
+shH2BmHlhaRcEvKwv0TEDUJ66aVtXtFzouSzwOz/X9PTVOXcxEZC/hh1Sp4xAyCrUWc9JZT+hph
/rkZ0CPUb2x6y1gvMTmIFGpf1fQqgmnQPW1X7S29U2ViK4QhYz9/J8YGIH8wWvFwNtUhA60IheWP
6CZ97om+N2Mf8tBT73LZAa6LMcTav5zK2nOIPy+L2ET254CSWu+yxu3K6tyjEE/B1yF35WU/d8gz
jfkij2Cqls47PMzz42GRsnD/IPGD6JoBeMCWXevN45rBKwJ194pvgv5/VNPr25hBrjRQyvbeayiL
ztPEip/6CMruXeg3wfTrVo5bpvfAeIpA6JrL37A6JwGzRo/5z2LZ+sQcYUNdBlBhBcAAV5pJQTIu
yXDjASK6+zZxu40Cm35Nx068n08Z/x68NoAyd0pxoZin9MfY8gNXF9gh8guIij39Qctxbr/Ryags
gO+Ji+pY6yI7CVLVyR0YE/HyZne1ki/d1roa/DPJdPhf4oZqedJZqEYeWbcXrhzt8TvMrIC+tGwC
3ksVMLpnyM+o2OkitcI8eOJsTcK6mKBecT12PC3TDYyerICXANyTjdHAOQ97a7OMxnn7GCFQd3Au
uf0soWDEpTTZdfPy8BXUaeMiAdEwDtwbuMdq6yd/1Tn+pUjlavwr8tZZDyaHV5HCA/0UOZYA2Aku
U6n5zZbXoYGUkPgs7qEZ6er5h1c/6cFJCXmW4B8yKIiRPpEx8pO4vBoMhC/5amurQEB3Jd1qITV7
om6YVZCVMyBkgAU8qibUtrTXlfWBkNEl61g3PXCWDEpBHgXW7kE6FdXrC0yVa7LM24rOwKiuzpvw
oZ0Rw7/azBar0ueF2QF7/KCYrC6//O74fHVLRbWDMUhAS9uofmwQFJ0MraQ4myY8n/+c0xCur58f
yJmeeqEPCpH+hIpF3bi48Low3VfYpYS+81mc8RwU1M1RvzH+dOvOvFi/lXcYZtwBj0tgc+hw3gZK
TUURpL6x3n0pb8IP1wbeyys1vBFDSaoEd8/Y9aF5RDio6JFl/0ItHmOLptSXALcoG6d1ebUcokTy
3nDVbSdmOv8BjW1HWH5pcEdB9R1yxl8DH/hJZ9sm2Wq70L3RMNvUNKVN02ibCbUTwOgFehjimWGB
P2FDXcHpFTRGoILCj+Z5RoZhhUB+OsVYtnRjrNtT/Fc9cxGTPyroTNCb9ORoLnI9X6K5EbFve8lF
NaxQgayOXJTZnx38AOUM3ipciIYehtzrubDDUrW0JCQCRgkKBBEJFQ9kIq0RJCvVV0gkgsswXrfu
8zskHMluZrtxokhxxBWVqqZy0fnxzIyv6KE61pw3+158dXySV6XetrDBq8F1Im3MbosIyUF9ub/F
vcRziqegY+2zUAdwv+Z4gIu05hqWPMZgtIajp04pyVq+4dx2h7K+K0w5QrHABeMWKch2xzCU5+8v
bupV3D97w/EXsD5KjmsUD/0gIy683jqewi17HQLikeMrIlIUu4Tb76akq8dzauDOuBqmXnKFCSvm
LZxPi0XUku/KIsaXcw7O8bL8ALnN8lO1y3+pUT3f5zOIFedtngyiUPM27A4SXcqZOSH6FUdJgOI5
GENVQC+lcCl6jNiCVxh1pfbTLmHI7qcJ66qnIPIARzU3Mdtg9u1I+I9UhCGgGfMwM7Yw6vV0iCJ6
9+giMxbOxaOydpsKyzmGkGpaFXQPNxOjrqgo0irJIQg/87esg37iXShWnb1az4lTbmKMhtkhA0m6
m/+gZfAwNUnfqkPT9kBAjY7Ueqh3lXtavQQLl19nyXLRTyG/WnaNGbfcAxkyb7FvsF7OHsTeRm1r
h+jcQe9qC9ka2hOCGes4Cxkl9Q5YjcPeTYKbKC/RAGJP7qXTNwROOGFmbzfRav7WQQGlF2eAU+dv
Nd0W0szHCfCdzXdXop1MEjQPdqWNWyfF3TYZacXiwpvg05WB1L09o+E8IE4YcMC1dyJXrN2kMSkJ
UoDK+8JbARwpZLR6+kBG1LygEn8xe2vkk06+GPhFzoGrJLFp/USrTaByx6cewXyrW9Eq+YUJyk4j
9XMcZV8CIxKRN1w+m3oGJNQ3l6mBvtXhkR4EDllEHfRQSBE1ioLSyhw8kRcX2dZ/ylNsAXaxAERf
kH2zZMK2/NpBgogCkYOQted31R75Vlepqa/iGQXtBVOYO24Anh4YQ+ZuI7RQ9JYPKWTcnHtBTKhv
f/HxXKknKslnwukZTpQC/VGQ3OTFtseBaMs60l+tMKXh22agJ+QbJmMAEC0uH/3LMFcqZX37mXuc
fzXcTzQjUZuNG48a2usZOxEIsW8IA2k9xssD7oQS9QSiYhqU7CV920OpXubczfa8m4f5OSk5y47E
VPNtYNXW8kO7ULH0CnzLvv/7s3HTcnKtzbqsqY/4unpNWfyMBaIvLY16EK2iI0XsGN44SS/JSREr
x+qhc6jgBUsDRwM9CZLtLuVmcuOatZ9lfzeO0BZPi9zmt3DoKgBvspJUf21lIzsa7h+GhiJFJ6yN
SFzPD2rCEswLG9ezR+QIX2BqqqTmTPifL6U0SPbH6cm78ig6CF/T/C1KKGkM757ho+46eaHzJvT2
DHYtmXdW8ffHDVoLLHEb3jOVgNnxLhcmebZJCkUk+utZZ9Qkwf9MKunhYuHEuVZZLduW1XwbkSum
jb5V+1LFI3cMj7tuQXaApFBXNAaIjAMdTwQISKOjxSgGG7dD6aguLr/KBeBppFOhTbhL9r+1fgbP
iSXdb4FKfpo2bS5C/wFI7i/IdMbLxQBcRNTmMz6o2CQBE/IUDNpInAPNyRD2LrKJ4AIuh2fesx1T
j1n4vzf0U8IsEu7ssRLnyeWgp5JHmHlpl51zkkMPDPAc9ai3YgpYYS2lF6tIJA0kXgH47qsbmr5V
3CNx7groBBk58BqN0AAHNEhDkg2Da0wWcilkvUPZiW/Kkxc+iY8+mfYw7kM13PWZNJmlNb07hz4h
crpZ7+d2gNKvasZuLMtRXy/h7qbScd7oov8B96fwbfgBwJzbYC866galslrapdwzopXPnX8gP2M/
4AJvnMafSLmpVkpAA77uXIHQ71sALi0Om3mM3OQor6y0HwPoTyDHIxjO+cjSa13dvHz4lHROlMOj
C5tAJPtcYG7l9opxN3oHZrR0Neh+8BJ63Hcll47xe3AkF4dGm20yK5gd/T1ycoSE3Hnfs+ysy8Pp
YctcVrmqRXagPj79S/7txRLLQxKxdX8GWHxwS81ks5LBVLOeLlSttJlAVWnblJuV8CbiKja9MZTw
8Ia7ypX/ROHbtGBmWJHzGSd5dadNU+NGdXlNL5RwpliAKmxxeB36S53zJBdeFGDgIwOJuzY+8wyn
uVuL6EyhzKkLMrAH/dSWYjoJOtraqC+T64hSXNJbmCG69vB+LO+ewO2zaWLh8YO/w7HRoZooO8kk
kq3kV41nCc83XfmohnG0ecZCHaWY6udGBsZN9jiSsvsfT3+7JFlzwwHvlCjZGVuWtYsF6R3GQCH7
OywyIOlQR66PGDHQfiX6PhFOqLF7tm8WMvhEdbK5Ge0rVDYstukGuub5h58WD6E2DX2vDuBdCUyj
lBkp7srY8Rx0bWlM2YoRdsR9UT6KFjLYOTniEB47WxyVGD94t5vGkb68iGbfOs6u1dUb+RdC22DT
mqQ516DEMQKWtbwC0AL2AZrx0i4YbT74Ds3e6k6MrD4Y9bmLrUFWbK/U4EuxtdP3tpF0rlFhnTH9
9M6s8F2y9h+YflpyHELL//C2IpPH7KAe8SnMEVgdR7WoT8Hx8ewWX5YhMel08Xo0LzBuxpPepHqR
JpGy69BACx2GFP0VDCwvN/WhBFkq4MHN4Gw/9Uknaap4JSxiZMwDHzQ2H9vvbJp1ACNUTD+vQK9Q
jpRCEzDTZBhEZdITWFnvHD0ImdhUbIz8avMEQ/O3/plJVmr4iSDBHHlkPryp4mVfXCRQUymbDINI
TT7qZB1QvEyO5FJRw4Qp9ls8cKwK6b+36zzuCr002huYUUIn6sUCB1qVRcP/Y/AiIIXyHD/F9Svd
HHHdqoi+b8UDL7HMXncoqEVh2u47MMycVvGxqA+vObWjLiOR/DhzygGVmu0YfVnoppV2kETZXmfI
uY+BN5ZQq554MZ8W/Faa5GZdsUg/bcrXLjEV4bxhpHkJvZSOke6oxwOw+02/qtXBwkE7zVcV1Mj0
CRhmV3zcQknLJ66Ad5WsWS3shYsj4d1HUHcXCVlE06iqn3XQgzlfIqiVqd5tOd1zBZa21SK9uYag
dwCcYnBCGS+VgUOADE0KhwvLf3roTXNNy7AVanWr2SvaZZwXU8dE+/FDNwt66ROCuCbB/XjfVz/p
EMkyirwyZCXLKC2PG8SYaM8Gqt5R1Jw1Z9o/DL8TcTvvl/Lv04xtGdKnxvgrlbE40oot8wyakEU8
dAXBr6oXmxXjs1QRWahRjx2y67m42ICJDYd//Aao2wpL1B8oxDALWBDvXTb4BcFqxnCTck6fbuvW
OroXssefctBUKvYRYJYlh0/GTGJQcGphOLTAwNcBRE+bK108f2miTV2dIPiVWPpfsuLDf/MDmUQN
CDyTlzIDVyzYi79jLqsoWEpSKRrOkZb+VMIz39QX4+O8tNTyC5dC1l72hjqNsOKt8+Puyf/pEyaN
tPT7lIr6TGZPnLE1fxWpeGCj2sHqzpiPSin9Glz+pn7KBiYunRbI2UEgo+9hKPdOKazR4KjMUFsi
8aKXWg3lXKiozaaXNzjofLGL24IPFLHVess/LJiahCRjDI5332TedRLvEHrMVGcZ89ZBtEY8OrWI
/hKPZPgY7hoKdy6bsNBJrz5Eqr+r1XFqsYkFRM/YI5mO+H6uu4Jw/H0vARKlHkohfkQepFE9JWDK
OGszMnxB2o3yt+3LChlgLfJ01423A6FDS7cClrqh+9XvlqbieAVprflZ4eerJ1H+pVC7OZSq+Tgy
rk8C+NMGpNNj0Pbf2SYTQWF7lsWHOJUpU2Kf9Vt7kQ+BMiwGuifr62k2nNIGJwbjeJRAEbDV89J0
6U3n9gC5IdlxTScSSWqKddKgX/IQHt27U7PyutbndQH/2Vzm0Csddgt7gfzDScyZ2HAOMyVsbfeB
M3ZXEl1chpOlb7O3uDwGPqFs5iiuTUV1RKqRjF35ayTSSecskXXN/hggoumgDBZ2j0z1DTe/l2Lo
ewzQmKc/Ow0KfuFDUhGBJoRr8n6j9DnQWvkI1WxlKGjYXNZ4Fri6TpGMHgfzXPE2uuyFMfN8No0T
OrELSc3VTP/oEXeg2R/SGc9fzR7F6eeYokKjb3s2EUbNAql5tPobE+cdPBQmWMH+xLEDIf8jQkq8
8ANhKdg7cQx0pVVyL84o0FQUnRxh7jlbTFk1F6vfEU2jc3uoR7oWaHi7ED2Jwcy6Peu5z0RzwfV1
Ns8+bHh08mutlfqMW5aMRzzGZLc4J6zltIQkGNghWgtOdZWnieJdd5r9SOgpVqFtCF5wrjXzeFI/
kCFv/sdz8HSLamdoHidjmIwyWiYSySRFwWAH6EICY1Zu+JHk+qYhay2a5HB8kN/yYKe46vIkwRsR
H4CiRPqOwS5laeyWyu/Kmqna2hYKOzBIwKS4RBdzoTfBBC2AHdpmM7NrZFvjvfFn+H2yPNoqtFyh
NxM4YjyZJuqv1bmilfEKkKlgb29mc9yHiMkLVaxtdmG63o1sxAf9HQAutCtuAL0UWowUD0KvpQBL
2g3jaQ89AvbL6j10W4J1+5nm2rO4O++ygHlBJr7lXUWbV1B1Y1+L4ms9lPDnzHDR3raQ8usPBAql
isj4Ct8s2L6TrvjRjmzNFJ/Arn29g0JJVADDGeVMfddnMpsaoHHokghsmqwNQcaX2loWfPLh18Y8
0ud5PVYvcVrIRkzhSu47E+5oeTbhvHyWn6zShMSSpO1Nvj5pLxMsfniUI65Uz3AQsZOFECvKZ8O9
ygKHW9TN1Hb+6TdFwtIk4lzBUEslo0Ao4cCuCf82XKTeLT4DunKrR4XDjbqmsw1wPXPaDEftDyJ6
1apclZVTvjKIzEHJGLdZ3LqH34gGAiGccmUb0BEikl9+K0qJDo5bjj9b+GIGHT1oO/Bj2kInJS72
VTH9wPJDUb3/MLmzxtoLZa1GrE2G6kSYuaJwZEuGYRJRuNK3M3U78Nkv5zkvfNyovtH4ZjPu/xl9
o994vehSJrZ1f0OAgfXbrJFjvehqBLxla4WfAP6AznT3x8j6H7hMub82lnrOwUn7PsCCOJ04Jhwy
5IpUngPc3KnwjexJE/ZD1HNeMZLhWTCUC5PUEMjCV/AZu0KfUndNikEZ98QFhFtOnZ7uvd1uHLG5
bGY8MtE9QnASIoh06RBaF9rpP1jsBfNr4PoGT3CsPCyOY3h6wjar5Z658kOix/tRWqkdVV3ph17C
DOScIcqrn3brUvoc1OWvjKnVMmoforkk1/60AyHXV0j4BYMgsLfgSYFug4hMhHjNzE4wEFh8phI2
cIpQMLA28kqmoGwHFqB5vEuUJRp8kuWXHDlAaEYS36/w94F6zvfE5jLcsVFTD6RnBgSpU3771fEP
j50l72+5VgmU6d7lLxtALxeXnnUF+tv+65ZhpOF7H6z7PfYq8o8WYQaXEfy+gPaJXxa3quoG7hP/
5ZJT7Dw5VGWk97DDzT+28cYXv3tseYuE05b/1ehQS4FjmJ8u4wafOsdfQcgfmacN85jbfLPPeWIf
9m4U2bnslJe9S9wFogoannDYIMpHwlQTpILCcwx5Nf+cP5+8YCD1P4moxrsVWzpIXpjbY4FpD4ED
PgLTK0r+j9bFk53Qua5x2OzvUvHa0Y7+cpuqu2Ktq7m7Bq2vOVmaoYbxCkLb2SZBlMzkHj+TZRmB
5HVreYfP9bDMNLarJtn57iJlJJV7rLFCATxS3gqa5AltEDZwwp4Jh3ja2nBpdrq6iBaK6CO5igXf
KPNbSQ9vVuw8zx/9j3XaBDr+tje47usiGUSuRsBHw5gDb22vhqbx4m1EFK4O/x+anzPGd43UYzxD
o7Mb7SDADZUaAblbNZBPrT0qYrk4V2marqHzZ+KGnirwCMsVXATKJQ51rhhcVfbiSNc7ThtJi0Ct
JJwEnP8J/KbsL13hgO5at8qPejW8GxmmezYH2yjNrA+/PLMf6XfzVREP7kh/RHB/A2IdixHtHZ33
JVTU0NE8Qs1BUYC0WgQuMx8b+xVWGGaz9sDylbfmcDZ9AKxdS5fxcjUH+dFWtnyoZKibDh4/jvrb
3awF7zWhpka1ebsH/5JwQljKm2tyCEIsxHf6tFOoDYCTTsLJRry1eByV1dqBDp/8/1Ol9E5JcNHj
iwkofm41++e5JooQZJouIt43XBL+lqZR1plGUflAwiqrbHM5lNJIMU1u4Csb6QZzlxiu+YxinVc0
+RGPT8fpTLqQmEFver5xW4Onu+BPJSmtn6Gj9EAGcr6iWhRgWHnr7G+uCLMD1LotUyPJFCpKg6e5
6Gz6su1hZEK6TK5+r4KAR2Drxafp5TXge9I5qXRyM8lSvrdHj1px5jpP76nLUUVjrC69DXjxGRSE
uVHHS+sCHzV94ry/jprZlmdf3GK5WF6dHk4SjPXidnf/VnnDG1nbVuiJEI/BWqMmqATvoEgN5xxS
zG6FemLcyR2Doe9wfgWmale3xqt8afQb1VMNkJJqJNqa9grCGlbS89/qL45IT30VnfasSXVgXPkT
NExqMM3Ss6iXB7MXERlnHOQCxpdL8gK60hl2Ep7JpeoX0TA/7QGZeD3SdQNyTyaQelYIQPTWeyRD
f3qT8OCmQ5pF0xlwsjvgRsdKOu27ggxO7LBsDcKarHm7noDEohXS5dxgALjmfKfmVIM8XpWerHK3
Ryr/PU7jWD+ufOQR/E7qFop2by2t8OtOqNZEJtn9WYcEfnb2E1xmEz0+7SGgnNv6IeZvYHjTg5II
f7RpSJYWJKReT9EAo2Qzf/8GXM5f4Gf0CA7HzxdMQ1C4zcL0h57sH8tAjd8YMks5mmxwI10EZSy7
o0mrHaIweZhP+oEneaCQ+b7wUC5CBSftEEGyjf7FqbZisVuz5zKd1q+/UQhRPnf3/QkIsFO222Cl
UxAaS+DgIL1BjHfUw5iniO2nHrUq3tV4UWqv7ZH6pyI3Nr8RWop9j9LgGp8fZ24E5PLqpNBJwuHx
Vo+570QcJjjNYEfYjSuNiMvDTjQW+UkStiuu55mCiLulJUsisoaHo1uvjHq0avjkNW1dwUUrYK6G
Ry5m9Mig4fibbil6+S60yIIe0zUTQFpUNHyS9b1ty//NN1+uV+TheqzjZcbvRihwgP6uBSifRSYN
RaTnSW9hCk739dGs3DWiOmSI932bqJajOOB6gABHVXn3QPA/wxUqNHX7q0zV+rqYZfm8wv9p7cK5
l9KgZUsO10Hf0ASF9DznVfcsA1x/sBmorbUQ8ACmNoNDcHZcmYxSuaSI4yZn+YQN1nzT2V543Q33
NMiFr3DLgQ54oik9Lae5ILPs3LxN17yzaXflsIVBqLu506siW3jYU+UAn7cs6s9xQDQJXQpq3IBX
Oop+apVDwnxknfcmWn6r7oQjfShincWkRZvytqHIgyjF0AOjL5aluhKPMxq0iItVyLF/pZod558P
zY+dyEaHcKVsFQFxPSGMuPhwT5yc2es9QAbHy8/E1sh898NzmJehTJxZNgr9ExSetvdjRFwFbadU
J4ffQsndoFOu7KZVn6oZEbpOe0W562gwvBJYbOi08Bgv9hjTsEFwPIG9IBZHmsDWw+2glM7WjeIb
yfIxE9whOu6/uEv7oRNpXvGcIuaeMwEItMI6IDwClFjs5G+fUcUwTIIhAnzCxdHyvSG6QjKpujdO
kYAPncg7xNPfz4YjNO9xMxf7cQsXg2Yalt7iKRVv2roNEk89104n0May4dWesneup2fI/8g3BhO7
eeZTtq6aqL498pW0qzrxWe83oWNCJ6In2MK7OmK+fxXEka5iIyTilkW7yFJ93pyG1EKAZl9c//My
rRwEGsiRPqX6rObkTIFBoWVC1eOtBdCjPUa1ew+7jCZhbDNwxaUYXTOZCEpZOrQZrjJwXNsqvBv3
LY3qn56AzdXCBD4J4UdYNo0/hd4Ogi3jfKRj0XlqmGwb0y3sP9TPof6vhlqUXLpYMeR00KrbVGzF
OQeTGbxP/zf8DR3S0ADtkWuedbGS1CuLDJlGqXmeXy76iort7bNcFs6QJvr46ltK5qUdyN1SvN24
h3b1PDULslcgc7CAx+mxRcRSgYUPysBw10mzcf0u1uJAfYIaBmVjA2NatMdOYP2cmFL5QIL8BlmD
QS5lqe0s6vFiEhpjzK5GFpSMse9+hOMjysuszCgSTQs0bqUdqMT4l9U+7cdJIp1YqVmnKjTVVC2N
auVHLhEb9dzms0+vIiSsRlWfeK9i51TjLnEEAYc30zGA1koIfKPKTAN2Ocs/A7BpwCXwVeoF7l3n
LYrdv+O7r4YPGiuLrxI5VmBipb8ak9vrzt1CLuAPUeszLSNju9lffA2sL8qmrZZXHBjIU7EmCoQx
GgBuQYXrNwP98uFwgqSCp0cEuHXBGH4+DXdyL+u3Sbg4xYrM5mzDtzfq6El9eYPNRDYdA8m9gZAt
gb0FV6HWYJVDzzajG6AXeKKuwyhPZSTgFyf1nUO49cLUuVEn8ktWecmaypjSHbX5hhdifP65ihRO
Qqe2HS8bGTwE/6fJSzf1GQBcOrLzaH/kF9uxFbCukVtzVGEGEipN7gOr1NV10ftMAVcnX7t5KQPJ
YVqS1b4z4yJmIkLAg6Haz9GdLiGm2u6gYG5IAtLwRxw+UpYcXTCNqRDtJ4O4mEGZQDnIgAocCICb
nj2o8XDiJeEJDzu3s5qWrI/MjhEYSTrOBZJicRvh25LaxT0N/cUyFkuek/e78mmwQSxYS9R9i62+
L+lf0yDZE6XHdOWdEVAubgsplwd4hTQnsSQo6ZHWrdCw9z/C1vn2Ur9xXpMltslSfe0BqmGtzn1R
NwE2PqRdXdofiXSJkYmrEvjHZC1yrj3qWXezqQ7y9M+csnZRyGu/S41x2P0gmM3yhmMuIRa41W7H
G6ed5Ivh+ah9CKMmH6DWnvqwwLvmEl2Uv/6qdsgsq+2qDJj6YVvhawJ21iajJO74Mwf5Be48EdG9
BYYmEgZW0fiH9aUoZJtMVkg+wFdt18UnYjE6AfwbyCcWPcE6UebXlEixINA0T95lUdPKyErMuVyj
3gmNZZzTZHA0K4N7DfeI4taxARMO2eDw+frYPWmV44ItN3AP7SCHJVpvL+219HWr42DQGrCqlvuT
p1vjVa1PYQfuRELMrOKnIWB46WbjuX+lqT/fd9FfBC+0xRoaXN0J00kvZdLcb1revvmBveA+2AhN
7Mft5NhJNcspN6jrQ6ESFm3Y11Rz/NVbHNISgqrkE+F6NKlAtALqTc4TjMIHJ+Je70AGBFpBrbHF
WWo0ElP552eoDyyO64nlPA1K+Sc8amdmI+NUoaz9gAv9EsZT1PmfztF1gnOIJW/JWTtEWRXrSbhD
5SZ8hbyCqRucdzWHMC8sFkRm7vBIgWP24zqqj1iLkRqIdTD6z3Y1f+iYqqAAnpM8I0rxTpuSQ8at
lNjHEtVJx/Jubrm8dVLJZ51KtCSngEGoiI/YAKi0Sg8RrJ2Ngbc2bxBUMbDoJe6JewVX+nwNy/B8
M45AENtQ9Gp1ak6xSzrd8cLyq9gyL4kGyngE3ExcrHVVq71sakCPzMBNNTqslxtFwxXtPYrTK6AJ
Tcud37r7beUIf978LgAO0nk9ENo+U5FkeK+S0drKDm95lkEKtJ4GmGOeoHexfq05KAj4Xwu2ZyUj
X6HUEehikaahOETcDGe13gy5gThRr+VSMTI6+QYLvY0cTeWM6N36+qtHw9qKuaJzC7MJ5n0sDPA1
0Om+yckeWpPF0HMl76XScHmwOKOroSDrvbvaKmmWVgVdzYS/7j2ZyEX8ic5lV009w+lajfZew4hq
yUwq5jCQuDTZy8MwKyz7OG6zYrWPm4TGCXkR4KxNg/oWxaJ4drJWcUoBr8byisxY/E4aNV8g2w5q
TnMRjb46guvIG6Md5f/YPmyWyqJT/O7fL51jBVDKTMDWfvp/Nvc5jILC8VCOfG5/kjSpEnl0pOql
xAnpJW9+kW9otIGEpoXS14k6IedXE6h+OYT2YvS2tkUgEcI14EL6sNhg51nxizLFdoUc4/cAGkWI
+pWtEWW5NpeuYf6ByOQmAP85rNBPhy/WLXTyZ6yiS9Az+6sn6CJARElsp/2Xr+UCtNMkZvAs28c3
lX2fLrW913Y2LrRDG6UL8u/XVmE25wM6NA0hbTnp8kKYTR9GswZ85I/o7LuwVWEHvhTI5q59HFHE
cVvn6eE+IbMpjm6d/4BGJ1LhfZdAzj1230BD5J75OkZjiiZerE/JLU4+F//pHuXyPoXe3ANjq5Hn
H11KPOgdZ8wRCxDaEo5uwxWEsv/DnT7jnX/ZxewilsdScLLQpued3T8jLrA+rTuKCrX4KhG/fbnk
Yps+k2eNTkHwBj23eYfNJHBaR7Tp942QxPHEb/xT1iKwyA8SSMSTP/3G9N0s0fV6GGJwDZ3GYdfy
a37HaEM8LNecUFGkKbqOdlLwyCxmM3fCxxI1FixKhWJsx1simXaJDSHQDP2J5h3/lZCzB8UaiWjS
1W3uMIGBRos56u7oM7v8gvbcl7JJCyemaRiIdJLqylNmw/WWxJD2XKqSu2j3bgdmbtiq++7TsK1y
L+AkOLQN+JxJ2DkKTnh7L+w0x3e3WRv69p9KJc7WS2hDf9Lt5CPqnm16K/fC6FNxC1Zxhb9zupAp
M7xvILCqhiC4TeonCb7kSvg8lpPQQrTK+9+EG6cTya7R8SUgG750jqvxc2zWO//aSOtbzHNmRjQe
AVuMBA0vTO1QsICwgNrpXjoAwAorrBaarPziRxWQqCyg2GxzwgvpcMi/RL3cM0V9YU6Jcg1VgWYM
xXzVhqCCMjjG//2y07EEFRCRjVspfBIEr/+FxAgLJjwgwRTPgTsYAbgnH2WlSOObFeN/rHDToJ/S
S/MQzijE09s6a4HiCzszcRxNKjVO04M5JnQktHoSEd7ZJjPJlUC81nYy5VoQ8NAMP7w8C3Z+izKP
wAh4EdEszFEDZ/H1SrVbcIC/X4fRzALNclAaGJ8Hjv7GQace/gcIztdapsg5Ckhz7IGuCwdOKs+l
7vG9R/jzp+2jQ2u7lUrhhPWqI05EYmwfCFZUcIY2VVJ6AplBM3NpCHDiagDsGaMIH8dFRQz5t0Sv
eHet28gwAS7q6NduEGtm+wp+v01lK6OjdBheELv2ZNrdSJTXgB+RUCvaRcXRfnG/38buS4nTtOuc
k89xSm3yY8hzuNMFe+xeRyDadCCQWR0/P+irkto1tFDkAkaEB33gMg0M6jxSSdaX8SRtYgkRXnSL
t4dwge4vzs8ZuFu8f3VoX30080iyCVPkBduC8W45oRko56Xk9YbhforSV6Vh5oJlZ7S/8V2R2TzU
P2KQDTHarkFRlu1/Aifulu7aybO6w8aKKEEahNpsSFJqIVLymMfTNf0NbCoNvaLqWl+3Pr8WY2Ww
BLAT/MefwX8NTYKHEeBNKCO/r+AlSSz2EksNvLUKicbMcjFSi01WgQNJUNvPj7wSYY4fs0TQqxgX
gfRicSWFwlAuGZs7eLgiQ7PePgdrRWkBZVssaK9lQ3syCAFa/gY/zex3lljMh6GIOuEzp+pwf/k0
GWIzE2Y1SG3rO6E45zRmvf+4H8ni24ixugtpbE32vs6cyY6njzjM7HVTVuLCmh9/L0LSk9xcO3KF
BYNfbVtxvhYZ/fH5fKSa/sDB4+wqsOaFouYIihNpuw5FZzkTjwok9zB2TQ0pp3GbY+RDulfNXamh
jM+E5gX6d0up+idencdKvx+52qoN+jCkltCmmoGjWfoe7H/yh+eGLCzN2asBG2Ku6iADGYaBoxaG
j46E7F9teTrRgZJk9vnZY4S6wLE7Jec1NeM/vvTKKXb1m0tqUGY0HomkX9K6BRduuuDzFkO+tT6Z
Jh4f9aDO4REim4RzH+wJFB8qkNnHh1fx3wyE6UTS0Uy16+nc93gh1Z1LpMlfHs0f/rqAHjf5k0rr
FDut+9U+fRgGR4hUldqETw4ORhIFnnJudD5KjQpSFRiYHrelqY1cwNIeoCHPaB1OYWLigjKpYr0g
QCEjWejisPo5KFjnHx7FE9Ufr5RZJ0C4WRiin1hMcA1lEZ1+HLR4pz86JXZifrP0CjfzZHHiMa5P
aXhmBXWEZX66NjmSwCV7zLu7sz9r+S6zFs/MbcIKVt1PApsue8sb8yydvs0dqOokOLsr2oaNRWJU
Zg8f8krAGx0He38iqAea2ZAtKjNsOmgypJeweJgt09ydWsSCdc2v5ECA1mH1FxZm/Hx0duZYQBiB
7r2z8Oj4Fuk9zKSbZMXjzHnG5xrldoE6u+rQlSJ9is2aLY2zSgtMvCR4hEiO3mFkXgvYhzaB27aY
bwopkbLSdCWofNZaLaywyMu7xFoYmnlf3w6We7m5Fg9Ya92kacgjf1cE79HVI1tMMIKoL5fhf2h1
fMRmisSAohQslwMIOp7lsYnzlGZ3/eGYoovbfd3kch5EJROPsg3b7MEu35DaG6UJFwpRV+VcPpOS
4VWISMPeiAaUvCP1aaMIRw58DoeUjD4itE7l9z45C4fmDR5Ud92+HZwtUuNQNQ6dSwPYnTuQi9Rr
o864nlahDb7CvT2jSZ7TGzjqZSxGNQ7otHpzr3oo89mIiVt39zTg2TyNm7kop4oeRZ4/30AQdsxd
xTPo06pHvmIxdOZQDGz08/WKjGaB2CxTQJwQthhMBxQPrM3oQUqtuRcDBUETWn+gmR/dZljppoPH
UZ6TWvrAaxABi0vWjy8R5p5CbcZPh8vnvdC0nyrizxftZPf74RRFY1dnNC6igDUZk9ggfhEvy0VS
m3d1Iyc/+NGwsQSzGXbvYEaGexRbXs7zEDljABBs1u6J3i1mi9qxIkISKMP+uEGLYDtatoadQV0O
Fc7PQPnpHpMb+V7mr7hdrZpH3LozjbmZixeC8TLGuhdnN+EC+a4pqxfeMdz0YT4RWKQ04ZyenH6g
2WcZ8rAdc3WvRw7SELrHTKXFM1Jp1KNclmW08f6ZpHHGnTC34uQryXltf0kvaQmX/+pQYH0eTrgo
KFSfX/EKqvQeyQMLHLrT+qDz2N0Pk9X1S9ZQfpazG8NC1VNleaKvzT5g28cgCQCC1BSrjuKF5fOL
VNb86W2ayoRZZ/Bt4aMyv4Pf5/rejb/EC/uVv7lM7ncSxvsKmaIF5NsZgSr7O2rqCYW/Rm+AAr4P
n2RXxlEWNrIKWzv/Kli8JAbnWEY1TvENeVbfs6d9zIrSuO9xSVJDUg9uz+EYObpVUw4S6Vr7h2kQ
9YqzZSFjaPTaYqg6Zlz5vF7pgB2Ldw3L8eL0jP6LIkV/Gt+B0XQo0mpO4dj8uPRlxkEHinAUpPYT
4W0AvyN7eSXkmm2QgzDognPS+hHAFUgcmLvzzNgHIqpHthDp+jxDatoKNJgWpq5Et3psJKCgKDxv
lVVPgVQ9brUa3fd88GNHqjUh0jaCYlqYF/LGJixDT3NRplwFgL2JZpIQNB7bVQBi+kCWGBapOhCq
PpPdVOYXvs9ZK4yyqifwf2gzy3dyGKqADdKlY4L2fGYMAQo+T4au1ls+KDPUrrNtwIYBZA4DTAtE
dkidEi3pCu02ovTxp0dAcjchQozh35Va3fw0lmeH9juUEWcZOWirbB3HXY1SzjYWcislPkQrqDMh
9dyUcovV3zvgP1d5+Tdz1LSAdgezHT5s7ys9Yjgmbx2ISdaJdDfVk1ayb2xJrE+JIHnAcDdHp5We
RhYitelP8mj+qpv1qCfbNv+nrjIpIi8/ShdWWDrHVzLqU1K6/3V+zlP/lHChUOlpQ+t9IOf2ACil
I/Rkf8i6q02AbEV855ZSmS7qqdDQFgo2gCyZrIfnYeXxHRfL8PJzZFzbVUCcl5uE2XFjXs4rklpk
vJ36mxzWDS0Jjr37rTVWLN7Oa3t21X6tEnBwOOys+iMQCtck/FpqAYmJl7nDmm9BeeP2666sMg3c
jZ8yC0/KOmz0FUa1mAX9Yaj0DcIkoOr/+A2LPyyAv7jWLILMtKNL9A8lp6/hBbBMM5HcmlWM0XeE
W1R3evVfViGHjGwvZObEW3mlfWIq0yIiPu2Ak5daT4qiR1Akl7tEiRXs9K+SmiO1wSNA909lPZTL
RZYFBYVMblwiNQLqp43gigDL9R2TA8uFMwZdTuVACi2RVgl2MXz7EXT1Y37eNAW4l67QFCPhiYLD
IrA3SQnkW9ohI8+7okbAosUNroTbs3x6MvpcKRgtbGISBY26t4LJwDTZZIpzxqxrB8TNsJkWEVRH
V2oaxRyyGAo8y0u+jN4qKGTR82wtRnIQ94Exuxqel7EUdFqk8/L0TK5J1a51PUimfzgv4Bca3fr2
Q3qDzN4QzzRDb2g5cY6Un0KRQ5ni1CjGGjIojvMfC2f0Gx9GaP0ySxk3pUY/0VgfE5tGpcafRaau
vcupGgU9+daz93kpI40GoxlX35bS/NbmzFzMYZL0CHY07M2MMSDbaPFFD0hKDLmPr76Xt4GdwREG
O2uHih3BOTIFV9JGH+GLwVRp0t+k5wA22NfXhg6TC/yu6zwtI+UzP8PbwqXQzKUWbK7y8JiyiaZB
jnVi62v/RiIG2G11ix+maakSIl3Pdbv94n4qjeuda5LSHhLkondmxetCFVe7werwoufsWYtDRIfc
K3cTFI98BUN+jLd4FXDN0jWitrZkOkxWTcRiVzxiG1/tHDF1CmQX3ACDaodbl+yJ3KjS4jPS1UlO
A3pYEVXAo987VqFzRzVMjiWRC+GGm6cvNhySoFcdQ9huZV7JRP7IKWzl2M4QSUch62ack/gIWMfN
hJ4smwGkXBSUPWHvw7rmJ9xocH/X1YVDXWARhhE5MprrrW5EASWRlAGX0D6SKjfV2eurk/qSZeQc
gCOs8ziL1SWUvaVvKwdtSqgugNnoG1l2gijNXjyDjzPMmr0jee+aDpzfHAlA+ieNWHRTjJkDBRjK
Dby8HwJIowPCEjbqZQ18OfowDpUt/05EwQ1WIN24Pgw1/Ou9ngGclpSVV2TTXXqdgKv+yGcz2FY1
TIY677sgPAOF3opIla/9vfxgIjw7/ua0K4SJSgRto/4jBNNogbJvoMnRJfbyjDSTjQ9uO/rqiwUb
yhUClxdpe1vUvlxtdSKZVZ8Ur1VK5FTkqEMEbcEpWnF3Q1ega4YTSA/MGVAZw1ApkPR/L4T9u2fP
L2J7SCRd6GdLM9Hrz4Cy25F3q2aiEiPjCQOLQLDQGlyN+CF6b81LDBnexAR73AFvMVtEhCDRU5bA
5YQKIHHU1eXRXF6SncJeAhrEosftTCpPUtCjQXauNtm38c3Tuh/fkUG5BgeeGwRzU3vJCekut58R
R9bXPyHlZX9H6K1BAVDjRa6mqni/ubWYFqkG/d7VWj5q9mqtke5p9jX2P4s1ODSdQhIjpY8iBqGZ
VqLRdCJgZXeGcrS+Z4wxW9Ws7TMyL0U95/1N+/kpccSf5VHvVumfpcj81xP5tiWPozGdj6rjGjK5
V/hQOF6jXv6PWPcSSW14xT/2+k0lEe5zCKga0jHnRCwwu/MaBGCUECf/TC8zg51/2yApGfN9a5i+
pba+sKZ31fhMC2DtU8Q7J8F0ELYKIxb6cS3jy2ILW3SHAQ8LmMs6xjapU4ulXmBjlK+pdogaY/9P
f5+AEzL+eO5ePLIB2ynT5uiBMWStPI4QfQ01gbYVvMK82B9C+AEAGtQAqIw852hGtmP9aHKc6Ord
lsfLIJ5IGtU5ZzsZAzCQNtiVbI3SuTVgBZlkSaf2kTlBRnnppMpxCXZUZZqUT/B16PR/jvPb+R3g
GznvxUDEwy7XfeGbOPmJXCGP1pfgnYowQzmDdJO4S6F+ZKOo1TghtHRhmJDxz0FrHo0lX353OA5t
1m/U20zYeBVvnfGpB1u7LxHr8gnz/DAmv1dSJYR4UleB8mtQXlTu42oY3nQW0HI3hoaUika9PtLU
ejyW2KJ4J7RXBbqAMDyB3XTVFVszRPI58vnT0PV5S7uYNA2IOUybH/JhsB07HlhA5jPz0arydYnD
CKrIS3z+oxje5IOZFs8j6c5T53Le+4IX6OJI88uqE/qI3dk94hXfBOz2+ijoSaCfLknoaGz0DfIM
YgWAx5wLkOmWsJAZpUgAFNaiDDsGlI9XUNYfeZKc5mhAtBF1yFLQg3pKKWyQVVGwbdTbFeEq/Tmw
3Dl+Dn+GzpVj3o3OUyjvwlbee9k6DrFeekDB/XgqdsS/Sl+7H98XVVD71+7ym8wwPz02VE+HuUR8
JYYIjzbFTBToW1sP/AxghQjFE7+GLGDi/vSw38I1rq8E3/aF2jE2a8oTSyICPF1l5E/vYlk3futf
3dIzwW7xQdvvgWALU92Qpz2CPn4Tb5uVAEMTipyFuo0ad2kRPjoWixBU6tPrkp8bx/2IyJ/qjvOg
6LyFDH57ISHWJpobSocTrZohrhGnLX/7mFEOEINacqU4oE9d7ShYyH/x47A9ufMcYmOLy5SEvrJC
tlLgPz6Km+xYM5c/fvcl/MODrIDO8HL0/2STkBzhZTNOh+eEkr2bOQ4NiPzIUpDUd2lRDGcw6vwv
IujefRNfNEuLRym1tf1TyQdlR/WBtIUS11Sjj7Dsp4x/I4ayqY5aqUkBZMCcSSPTlZXVmtv3rJJF
2zrbbKqa8l+c6/MUiyjZDLVDgPdjHV91mpuvebX+XBuM2ubXT1hhr498gmWF/anjT5Imecx5EUer
i+0xrfIli5Damk/rLLHK7jfvrDa4YtSP3ZR+gSA8oDBkmrIP4/fFsecVrvTVT1yexGoLGZjugrKi
OFNfNgxQOdxx0CoP/mXBMtNjtFFqkLTxebR3Dl6WnpJue4X/idXeWBiPPThFwyGV+6jtlmYR69vb
D/Yy7Ie8pYH7Ib1VOeWnUOX0grSFYO/SIpNBA4+/+qiGSp5zD4B5FYIqgTopkQsrjqqT7isVxsxh
3r7we1O4FxUsloYcYadeaLLI21tx1M1oJTyZBzyMGONmkJ+jM1mSc36KL430+b8jJw+nQU4k6MVP
DwRMPFnpWyX3aFT+IlUvEDMcHPB0Fy7MwvZy0KOdW3VKiEJc5DM0RErSlbaa0EKdY93Lhw9D4wcn
/styj9i2EgyWM2qpL7Kcbpupu5NpSLNzP1Y7h/ZXTfVcZXql5izQs8CJ0FoiE0uTu81YY596NC2c
f8OiWidsYP0XbX4HglxFISKj6AzBt31mx2DvDXkeCPP6HlIVtFVoOMP5YjKiUo6+MW8oZbuiG+kG
IgIufzWdTWZ2SPvKJTVGe0m8PHEizp2zL2eCIc+Cr36/jxzJk28AzPTHcXp3nMBv2u73UIgcR0tu
KmsUiDS3am5BthJkkUeqeimzfRw3zPbZI+7IlVBanzTf8djBcHRlK5yMH3JgBNTuMZkCSVaLRsdV
Y/rlli1Bh3FQplY0W8wNkquHqaSwoDpT2gQOXNC+uLVbTQSOBTOr2dhfbZKxDQ4RpryBOpkibQmS
YDUPF7WOZyUa6xDDPeeUzazglSRpiW30D5AqtkI5rDxBIFWR+eYVDOuU1FXDMapDUw5zZfSLMyLR
paKs09P/EJ+tEHcFcSTXaT1Q7rxWxEkeU8Fs4bF7rsEcL1fTNOWTHb4lIxcYnmPsz1MWmPg0c3f9
OdMIPj2ZlnFK7vp59GjvzFceahwpsB3N3qAEaWUQAkwl255QIRh9WS8T1d6A/U1E454ras7Hi1ZC
rR9tcDwsX0qnv7U3AVYYeJTEiMQ8pEmmmol/8intVIUShhS6YIPUH66dmSqa/wshf8kgQXF+lYho
U9Qqyonckk+YiG5RFm2rUV9Ty0f6ZSPnLf2gtfYX6DezNUFYytWubq8N/Fu2pvSbUMdWX+cmQGnw
LA6izrbRBZOc5rFSxgOOVLeEwH+D0gASOYkPZd7N1j4XJYVeLPYXUJCyU1+YsPTeFMc3BsL/1nhE
qlXGI2g75k7me/hKMw/Fq17wjH7VxDRPJ4/t1wnN8DFL17/tnHPgPaGuTWl8o/JPV971RaXag9fc
7fn8Uuf71HYtit6HREd7saLwG1zR1dKvQE0J6lVsAEbNdc1lobw0F/7c13U4dkBHaYBe+3e+28Oh
N6pxx7OEx3tAj45bkasRo0HbpYUJAhMsmMhSFyylTfs5Oz5X5eJ8ey14g+2u3dtbd0zkiDJrPs7P
cNULbURHovL1BiW21SM1E1+alD86iargb/XMwAIAPiLFkChSUEQ5eswf7S8jh3SOM2wtFtEGFFnh
cJ1AT2HD+D2DhxSl5gZXtKIdLLD3rZgafHfTmKIjZZbo0lhhP+K+rNcCIH8p4oXOHISWrKFrUxO2
em2rX7I2Uk5nt2iqp29+QZG31JATjeQbBusOq2m0jzn2BxjgIMnh9Yrsz5qHVSIMeEDmOn10bMtk
h+Fvk/aen8kUjxurQH5e0BBN1EC8V1v1oJOHCWav7WfyTaf3R0TNL3r96voTQd4km+yob4ShpUkB
54yJhnp725zz7FsDkjzn4rchpHOx7H8ocp/az3mjikpk8j06TwwpsPchKCcFAJMcScikd05qohaD
wubhKTk1JTn9S5mehhhJvd/Ajnu0s6qs+xF7A19Wz9w2WPxHIY4INDBic9kDP8omYPUW0TWgJk69
ntJ04edscT387RGxeipEW3qSRjNweop0xkPfjciNzMTbc56F/i3FpL2+v4pTexCWK1Qssk+iKeD7
rgYRCEgsxf3HOgKhU0s6XerQ46M7rSIhrPjyFiMZkVixGOI69FPyxwNW/AC+aDi3FQqSaziLw5X3
EYe80Snf5giAXKD3gmi9x8Z0VjCqJLVqkAN2riEz+wIXRAhAU/gyWO+C/Z7d13DCx7rDQlKa5fJO
Xzni3+q4CvSJnlWdEbwyciowzkeBkZMrjuKx5LhX4b7UmtAZNfvkpviNMzv0kqKYV6OORlgOpAWG
TWd2zmw4sPlznEyXaRTRhqdER/1aBLzPFIVxun1yWPq2P6HA3kZKw8iJgoTlq4tuaVYAzDT55GKj
QXFTlBEdBhTtahyJ2MHiqrnaddSrk7i8vqds6ygqq56sZGZnhDUaCGI06mFumZJC0GjK6cuP2pVO
1V9pvKwZTtpSFv59kEy30F+1FFT2o0v8tNDoQLc4GxUW875CH8/IUrOw3jwJYHqfV81zjQVBrTza
Wq0fwDKImUxmzeY7zWUupFPYLMXXzbkUAYiHjsqRhPTjJL+irXLmYCq7E5ZiUA1nH2Z/ovj2Npso
5oTjf7mpPbalP3F8cAY6Q0UJna970JyPgndhkebK02Bi9H7r2px/qfh9pjNkrIVx8qcezBlFQf0t
tTpiq//5Dhmui+2BCv0XVAM3UTls4Qv8Np8tYvrmVk8favKO6BcGJUApjoywMLOeClfeuckU2yKU
R/1i91XHBzUIlb/y9UAqV5SIV5xTwt2Oqo+jNzdHlk7HoBmZMl3jg3+R66V9X6xOidqYlhXCvwhV
O7Nc3IRGlnZjirRygw3x9a9TTLgVdLpJ/7FYPVeh+uPPafmNeShJNOpleJ0jyq8s1CCG65ZjeJaZ
Pu3MYBOsV9687Ipq9MA8tq1WQuCqaV8gJBPVy2pB6FSFAOVyvfog5xhqcI+EsompGMbCLiJfkHs7
scUk2B0k4G0uJ/krXVG3Ue4lQOwfDh2/XakaGso+r++Cy0LPL0eaEqKvGI7oiJfFEX34SeAiAPBU
IFfgAiMNL/iJsmNyE+Gf2qGyw5Ljcj4S6iNQ0hu2VFce5fVTLQwSdes/jDVaAFMS9N4f01OWUnDd
qjYG2ryzW7ha4f5MA0AeQmnD83kzDcJltCEPHfERokeJAM0uhZUNsWTOjdUob5EG0ojJu9rCEGur
02q0qxeIXQiqGzCuXhXDS9GF5Oth8YAaZQq3qwQ0DeIQmiHpixU4DMEkw1qoMqwaAIcVGdKevl8F
2t9CWaB7ijyvTDVQseVoTQtcNc9LI7Daf54hNPSJw3maOCkNGLwf9CCPTsK7JDnqrWcjS1rgLpBl
+fj46hc8S2jTPXeKUY+EErwDELj3IkvKtgmFzJZ8RDlx0leqqTsXNG/O8v2O3bOyPT/aEdJDkPWW
zueNq1m28IU9Gk34Sry/Qlg48nWDpOOjMgd2hb3xhq0FxRCdV37au/oBAAmXbcMwivFz1aAXE4gJ
kg2Jbq6m8aMQb0YE2WPD39xjxvZNFp2AHFtkQwiJCAC9VdtJvgOYEGoe0vS04tc7tXRWtxy/P8Nc
kAAbA4Os7PhiB3XbkbpHl+UqeQINHP+rd/FRX986pW3azgTTzrqKWWnw3ea6C2trGIu/Jg3dZ3B7
PIY4g5sPfZ8x4APM6LiBufDWeSUMFfL7UC0rE9O64MBNbU9hNZ8OGRiFaMCAS0KBF+7/dkYVBy00
ulSlG7tJMYXjs2TSTOiNbOvjPwj1t5636wzhV/psaykYDsmuX6DM4e7WEX1iDe9XOHmJwngUQ1Fl
KuKU0XJe6YgBDo1/Ixd8VehP8ukbas/I5ZezMN3mZCToe2S9Fgb/t7JhriEnLD0UGjNqMvz62Ndd
gxCv/DaLWVcKn2QAXJ0dXe44CzqTiIz1ppaeMKn+51vHPJDGx4yBMcqT+mHdBGTs0Ww7YDcmwBpa
LVYrRgIH340Fabjm5+yZkdcSX9tPf9QFdnJ3hhK8ntGGaV4hQcRuxb7Iu3DOI7VUwSXxpZTAthCM
ih0CZyA+1k9UlIIwknKV5t/3HNLpiJJWn+d9Lq67DChPt+6JHynWpHImexkIsrOq2/98Z8NSws6Z
G+o2BhOsD+XEMkBggPaMZXxC+KttH7vtQZBBdj8CZLvSthHsiiD5k97autsvXWVqCJgbOqwjwdMt
jEtDhhjO9KZOoYDByWfW6GP1ZfuL8gflT0kffF0h5s2+RAvwZpni0AQ5Hq2C+YsO5F9YdtT6xHyY
6A0P8EbSI5filDjGUkhUxEbx3xfACVegwFRiLpIoluXGUlz23Z6iXC+eX1cBC6midROH6ldO4+H4
tMbQYW/TMMUGEU6bIezG/AsOFeSnC9HChljmb6VSuc2yQm0ShaB6CjWQ8s74tee3SXhAM7GWgwjV
Lu4X9/M7qoAUnfaTwdEk6zIhy0IDrdQnE/gYXxtMj3XHpQMX39lXkeCF36748ilicC0HSLsSTYwz
DpbpRalzWY5D3W5Rwq876Gpv7cgEnffumMuC1RGb7zo6mjJv+yH/kwV4gLWLluSuhZOIQ1Trnbqk
NiOL4KcHOF9Us0o6vJyvlXfgHL0D3lstFjLr7x6V4BKZzER9ZilOmdPPwAqufrNAoCDn25LF9Osv
H2eSia0cI300aLd3Nkcj5eAZQvAA3Z37DZc7kT8o0sBOvFhjGnbYIQNXUm/qNnElb3x9ZOaCFjzO
wuVPR4Hx1zjC7Cbn7BpMfoseL4ExRSAg/wRCfCRunzjAsxYo25tbAAM9+RoQjVghPZTamdQfHHPI
3irNkfwCIblUr9reub9at23q7k4wFG6X4ij1B5csyQBHJEvxgCUJtsPXZNjfK+tSNOTKdoIZwK9s
CPxviEvRSEETwVbqIqpiEVvh7vgYjrwWNrKwgudCy5e6+O2FEAZfcO2yIMyoOR1Ed7BFwgvylAMs
GaWs1AsNaPvyr2rUMkOf7OpfWvsEIS4+ambDMYs1j4yBUJM021Be61IohBQev63BfN6Gd09dZNj1
hFxm2UISL2Rq2qdKYMRHM18zmrTmJURzYd7dblF/vxJ0m9NVORwvgYZjuGJylX40HBu1FCB1FcRd
pikgwNeVVsW0Y5QVuiFj4/PrcQLCOTXED9I2O7VgTdGzKCAFFnVY6rSilu9aORFvHmKPEcdhXbMk
UJfmUW1zRk5zoydpJzX2+NDBsoN2sWHgjw9YvkQJ7+2p0la8IvyoBrfbhy+AUZpN1aTWXIGwOpqJ
UwrmE0z6Qzx9kVbr9UUZn0/zudtPHKdPFNxEuxotDufPMrELjNUvkyVXlTyfFUpwbGv6KBmPnK9I
1zcK+BsciLuuq5zTGgAcfdqPLs5c83Y933n9UoF3HPujaSaTt2N1SQF2R4cRN7khx7C61qO6yIOD
/WrasL7sVYGQ8dt38UT9XvlxYLoOOc8zLfIgfKJgzUviVFmnm7SWZ/qJBwmo5WOL6hULcOEkIhyf
tGiHAVYHyjybreIJfc8m66/iqpTmg+FSSKMq7R9mtAFpTfOwLqgO4IrD+30knF3aJjQny1Zsi/Mn
QRYWDPE6Re7NAJVp2xhIqPQrrAKUaXCciOv5GncEd4zl6suzXBUsdnwS7HMVDClyjfXU/I97k5qK
8iO8agOjEAUP6rfZvg7q4Ltk/W6AYRgKm3FUwj4hpHISOTMmTOx+UGeHJMmNMjYNY2rkSy2gvEuz
s5PIpPJfr+XR/YYFpevctXLEmbcoTj2IBvTbfjuhC9tQXON0qGsstyRisUYb8eOI++gBWdzLjtEo
xaOND9A5Q+mwyILvUbiVEiuIMp5s7cG2N+crx7a6vmYDkgZss7dFoYHuVXyduJ+UOfWOc1bkC5eM
EkxJURDr0dmlSh4GCRCwIaCEvF1/mioNFCi/3g7yi7zv52tVVuS0oTImeQYslxA15nDv2srAr6SK
O/jEBWTTlZbT3rM0Eg/4zBFsrmtLbSH/0oo1pRsLFISznnGqbB25eEt/CJIgTZHv9qpU+bPjNi+l
0dttQj1B11uSaC80hpmxz9RXc9zi0mgzFqarZYrpWZYW9GY+8zSzZE9FF9Ha1o0hL6NrXeTluCcF
D6JB0qH6sQRnZ/RnrQuOEsl08sGg84Wfp54lQxK5uXBIyaMLMimlDAI1+flP3BBCbyo/GNTPZ7Kt
4K4y+NNIOQBfAhm0VSiqZE6u2QD9Cqn1072AQipVFQUgx9c8fpvRkJv0fmUS4+itZRdzSkLmOYVo
zEZSUUTcqPq99y1WeXAz8O8JpJlI9yiAOrC9UkrSZfXm5RCOK1A2PLs9d5DjMeRdBlq7IPr2/Izk
BJcKw4/HMy1ExY+sZljre4ImloL2Q+SE9BJ29sElD723ceR052WQUKDtNR4CKQb8l5MNnAzt8Wnk
VZpFC4Pz447NmAFNIkfBkVMLgLexTvZQ79l2WZCikjJc84AjTKLUQ1SAsXYiLAoOXc0tYOjT4eIT
PAuvhJ7Kmpd6XlJbxwbBnGSlI7tZdVPPfspmAfqAFJRRCPt3OgNOHhsyHcdm3BcThJBtR3N/r2VW
QYv1j/h7miFUa7RqLIig2yiWZwTKyhYOkHp6gNbw5BLfylJVmT7a/FgyPgyYoIKh/gEzOLhSY3M/
BWVw+u450T8dnkKzYryBoHnDCHgHW0JQBrlevjKxMGRimnN6D+LG0mqkMNNuPn1Onq2BAVRWWPTG
jZV029mwVewv/mzooZj/MVu6uwRAVdCme+M6i7qUdKlyTLnplzPNFtxjpHec9GZS6svLZdeMSaf0
fUR10zZdsHuOKQTY5AnAqXOZbW7hqscBF5Nc0CLAWj8v1yGNuC47GAFWIDFLMCI5gCPzXyRHntR6
FKxHi7HfprZhRq2+6TSd0bhRRzrrDnKza82f7OmtkEtTyVwe3J+nsGRlWQ0iw6pp4CkQ4+mrYoNW
EHIr53DrWV66aoaabKivagSoxS2JHNjpscBA4UVQ9qxLi96ZujIfVSI4z0hL60GGO4vG+Ah2oKMZ
UKKkB/DQwZVFk3RkGLPNjMEYw6fBCKg8b6uNanzBL5k3AhUSRt20xLTd8SCOCKmbpuXkBAE/gUGS
fCqz4IEbhOKEtPGDjTP8tKBqzLKgLYacQDZBpP8HVVK5GBC8bhTHRtV6UcibN6FMLpwT0ahLjh8C
bIW9zp0TCvEOnoOp4XEBatqqVK22yBc8GjfEKGUf2u7ZUazrwI+xE+cNSF2Y8OjDH6ktBck15t/f
wdfvc28tR+Tf+ceUu/pDQk/UU5pGB4S5vu5Q76S1XSguKcSYdva4Oq80rfVoAVdnLNBDvoBNf+Nq
LzDnOQ3KO9X0MOkQ+6ORB1ChvVQ6N6nYD/GR1ukO68Qr6ph2dKmZCDJZlLfzLCtVSdjRtFOJ/4ud
DR7Cgl+DQNBPrcN0KbDy0AdA4z8loR1F8y9hMxc0qx30EAfpW/DTgc7qDEJE4+gniObDhZ4aVnpN
pKKShBkL9LTEWoBDjkcL+GUrOJJ6CICFnyJYsqhWqnOOzJstGUDtg77YCKX7sry27S09x5b2pRYP
ssdoSrhDswYxIudMdrTT1OfYe4OeypqiU9d3Kk5QZZGQEB205jDzIwXTDVSTGlEsDPfakfeH9Oq1
jILtcsYg2sM8k5iXpfGdHnWjQGiQqcGtKoX2TVuTN9SXDLEyLbZEwSmpy+jlIABSynneAnTng7CQ
8oITf6jmbuHp53ivo3SH56AyagZiKMirTsy9QxDHMh40NjvPptB+bmgN/K/9jXKslKfYSq8EpmCZ
cqMGpfmCwTV9tWihggs2Rc18shZNOjjpnWEae05DhkoSuIU1g0Eaz8g2B1cafRCobsrvqSbyzE4q
cw8o52/iA4as7kri/uEWBU8Se1yRV9BtapESnq7LljP52gbDF2XWI467wug6ee7RrOS+QpVtYaq4
3EZEfpDZ5fgHoEEGBilSVrVNk5gm5t+FPoyAls7eeuIsV9n3Fu8tPmWj9rLXCCJmVytSAR6btnfv
BetgkL0zzf15LogAM6lecl58ZY8T1LlWmFvpO0E7rgyB0o/nF+kjeQSG28CbvXDYeqYFd8KUs20M
Ey/do9r6819aPDjskjmOozLUkz6cOuBuzbnbkdNCRHd/MredseDEAbZu5qLtN3CIR/lBUc+E/Dwc
BU+ZRrwIE8MtZxgu1P04QONrQoe+iYSD/oFccirhetxZSVQZHakAhNl/SKe26DvgE9DPJNyeCeWj
vh9zH9GwILodLffcIShmNEekn/ysXhk4t/Ke5cPvaUpg+Zi68+0CGYQOstTBeceztW43cqRAAdlQ
Oy6OvIap1sycIxGfvOF8VXLPxkrPPEMLbT/TTeqA8LkEcCZoBc07PqiVo+dfnLfIrWlvvaWXpeIk
ePKnvAgPr+uriq46Y9LuftCWCjNPSTyED428N4Fp5s8sQlruAJoVZHggmnnONOv5BS/brKaQzz7U
7MUr++2HSH65SPZT4pDmuEXXiIb1WjgJitW/q6TifCF4mKJ5rneZDFNgfUS0+0uiuh6Phn3TVo1b
DO2TFS1wHVZJezXe+TpV9NOCpUye8YDVrIDph5QbkddtNGUo/6jqNWJEatUuKTPhdVQHKcSMT4nC
FfIME2aRtCo6B3+OUxzzJBiQLlwDUdp+Tdoo/46m7OIu7umdtj3lxC62jA1YxpZJG1EjHNYlkQN+
pVLh37E74MFiqJ+UJxf7fg96tZUUdVTIclszwkYvZwP1Vt/r+5SjKFQh8jYDsolAUUlS9PIlg73h
JsY27S8iUnBmTlUmnsmUpzjlL3WmilELqMtbKDssbVtSVVJR8q/61GIAyR9kaIJr309qUYcDSYdj
oWv7hrQ7BEz1i2XXqjfXWDpY/XkrxKhLNaqFb7n6m0gpKFRNzQlU/K2BSccXQ2J0eC1gsTKWpQ8Q
43j9pAjn77l0AI8xp4Wfx00rLtO9nLAnRJWakDtWk31Qm0DzaC2gf4r3ScbR50rBe7/PFexF7OqL
75zkCYQhqw8UhPFqUBscwhg2k9wV6HVN+hLp1wW0N4Mg3kyJYB6awOd+ljrZtUZO756+cZGDKKGX
zc58m+irqM/MksO72sGwQpmv3uVcucd1Fs1rgEXWlxNAZ7HCLFv87GwJJvRNjMXu85AXU+9BICNA
SUZ1aGFrY9gN6i21QXdhY87MFM83J8qQ/DWhqHkd54Hp4tvtfTxZEOWAXtczoVdejeLxnx9/Ds8+
9K5+y4pOAk67E9C3aBj8IaOIWtXzUI62U/5UdeFvP/1kSPiQewdk2i3gukEHWP+EodQtcPZMLSgY
T51llW2dPOr/AzhsktHELMTzbHtNMEC6XMgU/40veNqlaBu3XckrF4wZIfIGJ2uQmzv9184p+9JK
7gQvDPorKRaCnO1GNALeMD1yeS6GXhcvOYMGvbWUPYP2H9+YuyVHeL2z6Kv4b8S2kqROv/3WwHAl
pCkB2aGRcXJkh9Gwkv5P1EjCEykMYokG0MCWDi6agN2WnI35maMucuITMC4IdrN6CC2/XFEGepPd
3g6BF39DlS1e83g+WqSFjIoFXdmUOLkvx1zav7KEdxm/65sX/0gO/tPcIRzv+27+dUmRjCuXOQS/
V0Ungij8yA+wNPLSyX8QFc9BElBfMUGBQcU/5LGiJhKQl8ebqqJ+1KGhEdTgzR3AG+7sRbpCws0U
lB/u1bwht1+SVwUWOdGHNB9EbW3iHm4AVZoP1hXjuvpjhikQ8Lfwbel2D0hQ+RudqjtGl0e+hcHf
QQgfd7LQzp5I11lrZLFlbEnspCx6uBwLpG15UluF4eqMjs0LIvJKFyh+3u0YuXJZklxxqHMz0jpv
wqp3GiduOvoeWTGrc09pbLCFIImlwoJFnNltxMwxgs//aKwsjS03lLOAiWWSEcoAZgc4hoPrtoFq
xEnjJImxSYYz2daYAOwYmquEVPm3HeWP+chLhVHJ8+Ip7uxM2OqJHKMKufRYkSU6w+odGRO+CwAY
bs9sFYwmDvbBJN4ybeo+63n5MEKFdN1QVNcHSiasOmH4LPFyV45R5jp6pe3GZFdNPL9xfAZ7vS3S
IpQKjJsZAiSWAu346E9y5RRfuiuISVrIj/3Qn6OVuRzoOLgDDN2yPoJqTZjfH+Dod5rNiTvAl0vt
thd/hGCrWCS9h6LvW5C9C9o7fK4Z4F4SGo8mvnmInkhTfmRaQT0ZItx7jaMizeJMufe+GYfgW7+D
PYTorelbOLiosrHAOFmalhzrhc3PkIylP0C87s8X+r0gmD1h92wOMXBm2vRitNxz+ejsEjLxQ5Af
RqjIZF2BBXzpvTmccOprnrEmimeOjZ7ZNMjxnM+WGhEAEljd8oJjooA+r7kUbTN2GsC6Oc0+WNGp
Fvaq9qmJJuLpv1ctYT91eLNauLRVNR9zppAASh4+MHjTrkh7OoO3N05SNRtTJsZtw+Za0RUF/T0O
C0EmhK39UUTC5Y456KEh7N00vBk04RYfuvRabVQpmuobH7mLQhY2sGCPbNDZkMnTlA7BnJOUTvA3
/x6HH1gtGoSktwayW5KyQUGOrFuzctByByIDStoOPQFcMrfJwR+JX/dGpVjIAZtxn414SuyfAUjj
AkUHEY90hc9scHFdAF8f05vMH6DmYJir4eW1AlzGyKs/BT1C+8YelSNxwU0dS+wg8XLWbo0G4r/Y
8BjPPvyElf+8OLQ/h8aW/mBEkp+LSBBJ8MAOUP8jcis/CukN/S1ZwvtqAtzI/YDgsx0Cy4zQzAHa
RKB3pXRHuF2Q9vTrHERWLX3F0tZrPqmgd14SKXoLYBzKi+hxjyPzZYh6PZZW7d3UhoNjZ6KrWg6W
mJWueFZ7+C8Bp5peUUN18iVb4FRvqP1DxQgKcUjVwzSp849kOqWUYVjJ+X1hfNkNDTZ2ZW20Hfej
UuKrmFeLe/CwBfj6ScmPh1xjKn9WkGm30LUyXm09ZP5Mg7MMuQ0YPzpqd5hqXi5Qn/S1cRhHbzAW
rg0sjXHzgnDm1SuRe5RT9FViKxMUf9kr2q8U0MTOgCNCjH0uDVrCdGqRki/fI5KM8Qarjs96xC8V
qjUDK63Wge1hup70mO/OIz8hkre/rtadHgXGCxaAROvB0DlMI6bDkpR7IOci8VergBI0g6x7eGo4
5FpjfMiynfACyXDlwia9nXwd8X/6eUxcIqLbIsLeE2mRVdhwrdOe8IqM1rUjlqVhqdJYwdCeGWdB
8N7gydORjkOik9v+kMam22WiHzERk5ak8gCNnK16n7Bhc0Uhbnp/GiWnIX800u6CsLS21vqvigMI
pecF7PCV3v2XtWmRHJ1Yo0ueEf9lRaxqYcW4NIoHc/wMz8bI2jTJaj+q/ebspRQITTtS7LtgogoQ
MWIa+NTeUwg4bH/FDiOPubVWPRDOKbXfmIKnOPoj5MC++OLFhCtgiQbgo6V//niv5KrLJdUSL5Pp
kPN1tjMfJau7AN1934rUmBKZta8j1Fwm486BLoZ8AX/xch13BslQL1u5P8LPtFnCb1Kiv0P0B1hf
B5Ip9LC5gpyKHADQhbfyOuHqvVdoyMGpY5rwSny72k+4GvkprrDcyyE9r+XuoEQgGDlTpRM2t/K/
330+65wbEd9WbOfKvxB8/zpPgS9jWG4F3d7X3SWQzdZkdIEpg+f8X1WBoODkk0+lDD3F4BQmQqgY
gyg11bMKVGtOdtkvoF6XTrXGPSuj+c0+rD1mJuqtMnJU7S+4lHCYFo7BaQWcvyOC1aQZ5Evo/l6e
D4NxHNwAhSyXi1pEC75VN5Pfp0QRBjbvZLDgQJpJY41fhzJ7VcaSOBuAVKqHyX/EAEwygNHOy+HN
umI1mbCmHeojWo7S7zinLDxbsYG8Cq5KYrndJkHxc0RrirThQhfnMd31MF24brrbeD3T++QOTi/P
hFS/5BDQ33Zgjw+6hMlTKHxfSOfYFZ8eZ+Q7TjGKnQR6AbAqmni359LrXErbyLOeTBmaU9xoXIJj
8w9uAAV5scOFRT61223GhBrcqSTovX8fFT9k9M13uwTmjG635axnneijWTdaWNG8OHPwfRTSg9Cl
PK7ZAFzmdALrgLA13PYvJPKasIwpzwc5yMTEVvMDZK7mvvzrKI/++jmfThHWW10k6bJ/Bt7ju7ZQ
XHVHE+8XDFkRr330td+LrdwjsSn7NWn69jNGBkbGPbXhIcIoyrkNrGtJyXNqxuMLTAddYnHKXjNc
d0W3Awc93U1EkF8ACIvU/7nuSnt6aORQmsUEFDQn7yke7fskZJld70NjnFkicn1/yA5C8DpF4nr4
27OWyIpsaIQ400MhdGTPefwFve/acGb91WirWCZOYTXsPC+AVpAwztx78UgbEMc33Gv40NGzKQIT
hsowX1LXSioTXYgg2QUYIZsITyg+FmHsV6+Dbjs9OJPqKOBY9BAVpiAvQ0VfVPBJ0icSNZvsfJQl
6bNmOA4GN4qhnAq8hfIArTBYx0DUgjYz5WbHEOfazHciVS2Oqdvfw4naGPLZNw4sIwuIaKQ/tzci
T+xLE81VL1WGh1e1bR1DcfXfnD1IucqRz2vrDw4qpy5UeKUk1srSwWlgpnkd4ie44mJc0735fC9F
odcKn30Kxcu/1Mr/2onLd2Chd8FyF9OVuWAdA1ZZX1C0Z+NAVfmd7x6GRDyhSr3vvBH2YOpCfg8+
E8gjRqNVMPdxvdDna8XPv+xNq43anBbex8GyuIA6QPXNUHpN9CbLcsJu2BCmU/hSti+BwL/TU94A
WUS6K+4r1/Ap+JD+kaC2OX42UP+Ui7S+Co1qVpzxR9/wkghIjRSDKoXW9FZ+J16LzovxiT1KBXGB
J+1HN69sfxp/z/RxmRIlkt1xyPQnYmMyHIVesX93W7bA71oyLrR91q8/XRqsZEBmfhNX6ChiSzpJ
qjbkZHlH7h21Q8DpIW2UvYA1r1zDa/9bbGmt/vsZKmiZ1unRxieuwiOASk0WuvbvOGP47BCg64P3
jQBrfSd/MmD0ODHqqZHd9+bukjTvlDG7+IMKg3Gel+Nymf4E1kINCzRW7ehDyUMVztK4nzygcDAl
59MA90HY8FMhraOu+FB2t+kuqgRgeBPKO7I7VEWjEzBasnijAdT1OS70z5+6jweBKyyYj4FzDIkj
wllXMfvzEgiMn/Ppg7tiBuFC8TOEjGzn046QFvlzJ+slGplLC43JqetITicgFhR/0g4Boi12aJH7
dE2m2wQpbEM71BnwMVT2sl/Gt2jx0J5MDclkOAw78np3dFZI5rdv7A1q375SbtUrzG3wm1MJ0eyt
qLdLl8nBcwIo8kg1SzUOK7GkylhJ63kjjn2Pgizc9GyyKsqUV8aJiE7g0VNd2Y81paBgZWHzmxN1
vX8AX2MqsAS0AR4BL9YWLOzu3iqDFETAenLsm6/be9IJoIpg73ED2c2Hi6HjN9UfsDuTII1Xjfdx
9MBej1L47I42t7mcl5HxO1Lp/Wk5xSaIuDhsCzuQPUkjnI5erhFIIlR2O0yY1HPsn6NOmH0xrmnV
9r79iv/QyOFKqm3wKF0+bJb8v+k/RBfarD3RTl/kCJSpDZDcpl1ojNHONYHka9xzBLv4ekEB1NLW
mFmZXUQRSO1b1mt4So2fYj7gnHK2bA0LyZ9vZbdu7vKrH2c7XPSNFEoQPFuO2jD425jOof09KOPb
DRbcv/VGkGomxTyTFUJ/KrHTVeVwUNRibkv4ceeT4Z+QbEWRni/3PG2yn+kG1p4BvRw8/XoA5erl
a6SOBMjWPp8w7g3QMGbTeOd8p42WeMsyYTHSom750K2nKHDl5cc3rKCzC/BLTCKrgApwDNhxhrHf
LROvJ3cCu34OWsA2EkmP4UEpP9TFF+zxVmd6OwFeK/75N1H2NYagb4M1dP6YcfmfDIsdUVFh4sc6
zuJkPhfT52D+WhiQkyd+2dbH5DmZrbRx9esWbxUNbAYum0b/+TEcHbP6BTrlEyV35JWsDBJmkNOU
jdYyngcLMqI+Zrj1jFpuHNKP7l1SEBe5+tpB3fifrfPgEUk4jCHJZofeMDNG7Mt2UCmJYMR4vBKb
EjvTNXZGZ7NdSJvrm4TmHL9pBd0rqAgJlY7y0Zz9sZd48DFSNrZtaMT1ObpJZG5IrnUfbKsK6G02
27VPucxEaLZJsXBuyWvr6gJRYt/MFCfyg8eWhwIk3C06yrfSVIDgyvRBlEd4bl6d8nxv2K5LNICR
OFJTvf3RvN0vxcE2ejc+cbOC7HgG63p1PqrI9iTgLQ209s8RY8SvnC4XSS8j/97yX1HHLxvLytXM
F0fkOmSYx37LZ0ItufxuU4SxS7OxkJq8Mf0iKThqRkSPHD07QVxz5tR7Q2YsWo4zr4eOKVLdMAst
CWMn8dOSzG+qM+nGVAtH4Qhgdcy6bDG4dsPWLXiYgTn78Dhn3P/w1MgUcivOILzlBkIf+czeuxbi
xDH4cCh5FZB8vAm1ZkyZ/dO7x4SFVJSIW6R5rRTUlmQvAWthedxBB0/6lZ/Eq6dP0Gpyf3nLos6r
DQa0+geLwRgsueRrvmTm/uZuk5/qlCVqZfKHgBNQuDqsD2zMC1HzrWxXWXjJlQrA0hNxp1o4HINE
zyMqdtjE0/mjdnbKv0CCtbWHRaaT49Wgh64Zjt190PdRK7RmCrcT0xsQrhTS+1nfvcvz99WfC64e
yUAObqZXjUYutUkE+jt2t2pQt3qG0PH9Ynk8Rx2JiBbP+lpkyjbk2TM57V3YmJXqIzM4UnD3AXsZ
fgdPh/iy4gYRmRoZfFI6Y7vf0mj3gBsgvihWqC2pNHsVtoFliZ3/8vfGBSXdCsG3801GrVUDjaFt
5FAmuS+f1sYzWLOuRwjwo7SIlv/ML71kXrpd/+1zxSFL3+iArjxr2+K9FTVSajNOYWtfxFvXxXvo
fVFtqfHg4KtBaFV6Hpa54Y5LEx1nwKVX2dQpqLTVBBu829ogvu+NhOtbeFo0wbPagn2HPyFv1eh1
zli5CN0O21hy+KVKjLL6TUAqPwqUymmD0UwgpQb8h1XnNNetdXyyLsOo5EQvtNdTB6aNJYrZgnTV
SH2Q9B6b2AkzRV5lR/qzza42CBUSn7GfDX+My2oeoP9pm+sVfaIZFvAANOpziO4PPCTd8SUOF7CN
3OdE5GyVZ+vnslMxkrwArtjGsTR/Yf68bYDUdMRroM1HQHme9AAJcpgv9/eHwCyJ9apgYCVK5dJv
SwZ8ny55oNwX5pbIY4i8X0F7M8FpGUicxJ8vQEfAy2OVdjad9n2ckYOfZb7qt/ZwoAYzqpnv/6Sh
afU6ulNlZLX0UZBR79jMXYOjdBx93EQKk+he3nTMmAcoy285fIvrpx82HmweWjpexUuCZv7TxKnJ
xwenghr6p8grb9iCqvup6ekxorfJK7Dtb38YZJlR5SYI3p3xiae7Ajv5kg540AgADY7NzHp12ygl
PKKMDSXD5SEdulowK6H6aI/kKbZpyK2h5O1fCLVX75H5K6L8JHoNeRSzgOTbft4d3Aad6aHstmDk
j5Goa3fmdA3HimJV4QAIUxB4n/kRFS/XPRd6TY34BBB2NWQ49F3WFH8POt+Y5DldXKEUfI7mBG34
CJ2Az2ikwCPNEbsRv1GXo13MY8WhypjbCcioqVwElWBv5yk8NwgzRkkJDF0GHRsvTpr78xyiHs/4
pR1UXmCHkLo8YH5erSfnnUWX5Gcx9pRTVxSmeG0VtWGwgvjtP3Pt6uALX+xKpre2eDYmoFtHP7N7
lKpN4y61vN3l2fkRidt/goN3/J0b2HTcMzO2q0X4+9UAcgiouh3W799c65B1mQJIzwhACCRzOu/h
ayak7KGn+51amNfVZbaKEr1lfyU7YeV0qIaKHCaLncLrxupxSCfp9eJPbFz+e6ZnCJpwaRTk3bLd
EyaTswXkGU84ojIhGxsO4SdR4pYWhi53rmnEzEHarAUFBvo9OYbQ3/0UIZ0lBzje4Hq2aRitrsQ5
PkYM0Wfy5+nYc9oM4B8SKYMg/JoDQxfisiiC3u0bz//mdxP3e2pXVqCJinq330Q5p3t9/42APrgX
11ogCChCK7um8DAFESdOrArRzveSepZmweTCeOD7AEYMpehZJLDLwM3pXipJgrTlyJfNEiLKcWce
Xqh1Lk1QGWaWLQu1B5aALueCDM1OXreFysP1ZBKV63PXKT77gnz4q1R3UKdqA3HQ1dNKOOAoG9pg
67kL37xCW/ftVl4k8GIOT5p2H7Wu4yPAXw6m1Dl4ZKX5mT6hSO+3f5u0MwBhb1pjz4yYZm0l1E07
MnK8/r5xSPJfvUdeaH7u44ckozb2gWyZjZTcEkuIYw1DSlv3tDeKLSbOjtbbD/I3FCOV2OrqziDY
A82am0r1bis5j8XwEJcY4wtzdVj1EghhLTOevMsu+Tj7yl4J9AujqzWhZKyu4VHpTo4IbwR9HR20
A+HXkzFAKIisd8irYfxo+q6811MIYfOkhPXf7lJ/pwLHG0aFLcjq9DPLQQE78Cc3gpFftECJeyi0
W4Zv8qxuIDzKVz9BYcpDCvxpl2EibvGwVoSvf38r9LYnKS3i5bi7ECvMrSLGlX/CBbi7E0mxN/Vr
IUjtOEloYMjvGR4LneAqIfj1DAO3LMUXoYyIFoArFzCDx5nYXQGc8KjcFYKbos3KhTeLFpHiRpRh
+u5N+OlZTlNXF4mGaMWUdafVLONh4LtFKmbe14NsbDq22TUPmluC1WDsxzE57gfmKDIOTgcaZsgT
6pKagtrZmbw1hQVOJa9WryAxGaQjjyHt2E617/KFQkjZY4vH9Dek0wVxNJC1PD2cXzmx/oDVDxUP
GU2GH0NY9jI0jPjieSppUCAjIbhTWk/yN/lVH6RmDZqa0j7ba65iWOqHMszGWVKRoJaPOn90Krih
1xWRatEJh6aqfTKh4IfPk84q2LGOTyVm2yX7QOb90fMTrLWq3KOK1UkLnHed0vqKxVqsiCKYerLW
z+rPTj+m6JBUPDc0ujY0e8bXyxdi1MkFmIT1znYeJVXh3NWxLVgFgkq0cdSemBD0buL9H8JDkXyx
wZGvumkGz7TgeMeY2Uc1IVxy9U0rzldx0i6V6i4AkYA/EzYLoiAVZdp+0DctvHhBRcaI/5lg2Jax
pI1xm2Bq7PlMj29HGehLUz/+B2ecnGJ0zI6boYbFLZLO1h6kuQuUb2Z8mRxj8VWZJdW01Afz3NO8
YTJvMP/gvELnj0Vd1CBad9DfvU2oZUT/LKLe4iMK5GFUxw8Hx9E4as2w6quq8272mReM0VMZ/gD6
ALFK5WBaHDEt7lEiLmgtjGTRE8ObcLfOGYexoMmGB8G4xjHeNDgnhAKF5WaVBP+uXxuaE0lUYHVN
zsiOOs31dOKYPWa0LV7pCQAw9+VSeRu7ftOrKHeh/41VQWExkY0xgTN9p0Kpo7XcRZzny6t3/43j
vdMhgdoCNu9mH8+QkHMbi9TyF60+BD3GRmxK5KHAbWxRxpQoTz1eBVJsxMhfoLYZp46XdSYKr/aO
pciluHFencoQfJFecpReMdpnXs6mFJHVz9d3gmRLld9dca5SPRxAXHpz0fi3xmyUS5EicLiyHsvH
wCWeduSnO4C+OUQiMckBfL32N8Yk1KXem52CXKcnU1e1ZDcygE0cOfam36opOl59c40sW44teQqL
DZwvU0R0tNupzA+q+ncoY9Aee7Ya4iFnsl+Nu/OSdrufBUjzLWLkTevp7BQlWe2HPAUbw4rSfYB8
uhbgCpIJ75YFKv93HxCSjdre1yVAeMXKdDEIlYdrFfIzvo4Z4pYPNxqUA1V0KdMTCCvyIh5OB/bK
xw87wXWW7cs9+Qlj2Xa2B4y3rIbQRr/a16L9R1/xjV40v/d4N55FDVv2Lzj7C9CliKzLYDvtyfR0
1TiMyVWL26tAqlX90u7UC8pDiNh7PIPlmLD0L+UFkXoCEiYYj7DOgVPeIC6IP9sfbodR7xUz+e5j
T2DFzxF/lk7WewVnNVbWn2LqRDXsQKcQMrCBiETtVB+sSVb3ugFct1WZ12L8r0sZkI6tV0c/b+NX
TfQlf7Ui9XrCkNBqC8acXvkeuM6H74Qe7GnXe8IeKnuOTHXsCfHaTsZRb7uD1o8syNAtn3BMVZUe
7dCTkzsozzHCvXe4yCPqvBCdf5ImwEKcnkQ4LQPCRTr5g2kwmR2R9g4QDIXT09AEXpCLX0eXo66h
96LH2fbWvhbLZI/Y2CkFDYKyB6f9v7If/IcBrPMxis4uG9xFernW6EmA6uJPTFb0E4nfRKUEC31b
fp9+23lwivS8mRGFeubHIpGrsl7z3+PE4v/xj3iNSukPepSgWJjhhrbJwvjy2Us4Xqppi0PmJjVc
7P7zJUfkuPyNP/bijtQLN9gQ+el1yRM1gPZ6M+3Khx64E7IM8xYz25Q45rjRTHc64jauybsvme0g
UQC6Mytp01ioTZcCYZyQxkV3Ta1z7UNY+JHZdmAzMdbXB0004WE/CoAaUfc+giK+ErqCuZkPUnd6
wIFc/01+1v3DQAB5BkvMex1xzDcWjfuCz0OCGB8lbHiUTvcy6Ejfojrqa+0h8svDmXxf9CyIjony
BYWgk3pKqrXIuIf0jkvUwCPdMb9O5fn13c5ihdspNmZ4GYDBsiOYycZNcAHgEBPM+ZTpmqRa8zqJ
96FvfEE+1zaWe3ESxN7Kvx3ZO+L67b2BNPDSr80yzkDQKYs0dsuub4IyLJOzmrYBuUaJ+K6P50Vy
2rv1SlqSkAEGGSbttmJsdNgfAqGp3JGey6pqP9ZqCKGRjPUdiCo3hmkMK2caKZuVdKfLKxTko/Lg
CV4dFvFBUpZwt1q9UGDpyVEHHQHMRD63kGAp6fgO6PdYtH7ezSHTJRI58jguyC9Zg9f+Smve7PO1
exLsLT8K1MbSUoztXJ4ai4azzEvmFxBfmTovFW2hwTMq+pah/RNqUiTnIh+juzLHUekVrr+liZoS
liy/9ZYJIsESOUUZ1972V5qcp/lXYpjPx8KAKVUPyMsoNzsN2YgrreSf3BMmczzf2d4oES63KN2T
v2BQEAmNoDRhYB35Etzz5W5RTYxKmu+rYMtgEHMHZiKuL3ehxaHDzF+I7yFrSJ1VEeZFJ0ExMwYx
u5TIrvPajHVTllGX05GCby3sFsy2bR5O0poR7D/zrTA6AnAjIHW8cY1La89wmJbCO4Dk+rxApsqU
9mzOQ+3PYTp6bRIrmCZ7+C8hWmoBN9+FI8+pIDAevGjGbJqu8NGeGxiglaJaFemT5ZN+eqyO522G
Wkf49gWgHfM7jqMYmUbfBshOSdx03PjtwhmYW4oghFnlYyTznMmIOSuXcMMidv3jpFG8idSIcEdx
kUu9zQ6ibmOKYIsBNcFN3qtG1e7k69knDpX8LM7ngxSpLArXh5GSBtsvWLSdShkmuO6iSkMUpgog
imkJ3OtP+EoqetrEsA1cyNGNDmDZ5wBEDLrSkGaHsuvacHeuvBmhIDcbDTAUojfrB+mX5G66zxjC
yK8DdF+cPUh1d0ggIIjTMBb+WCW6EZ6v9MehnJUfa7uK0jyxxlZqz/rrSUa6I0UsGoeySW/0ryX7
7cHzsjAfK5pAYivUruYjwA9rOdp0wSOXlggiX4BhueW8Rhc7IhHW+ClYUl5dpN6+RMGiyJl2+QmI
CmRlJd/VydYPCttYAWtSvKIFo/OPCJYw52L9vHvVNv13QzX87etli4vo+nP/q//lyCZt9vcv9YPB
FvTftMNqOQoeK8jyiD6yqUEkBEuPJl44r7R757RrxIVXhaXwsrs0rJdzr97VbM0R+PtLCioypPIU
wuPZxSMQz+DFmkfKyOMVT0XAUyqDNnFb/WJqOU73wPp7AKWkof+IJdaPhpj7yGJRbvM/+UmvRKMt
yyETfk6h73W0Lkougm5MPGjMT7eMNRsoJoQirugTAz8NqN8PfqzHxe/9rS9rFH3+AkBwmvXdk+m0
bGvzJUTPnWXKkcToJQl8LBNAMqubYQeVDBJrSsrWBUqp4i1KapiXop+Vwawg0rQOHxIHPg4IKMNb
bDOHHZYslZQyIvGOm0Yueop9A62dzExNOAlBXbpBu1v74av5ObDo3RxDgXLRPNRYJJIypd33HY4g
/0TkODRCxLn86l+VXQgdLAXA855s9HkYYk8e+e69YNaJSwqNuonaJMvfCYs1SLaHH2FepivbLL0g
FCJfwzN+9DRT1F/LlBnfW3kLDb8EXK9NZdt2dgfTjGVxRMmW+ZPwjNESrIChq4MifZnK5NTi8pyG
X1QbONEWamkt/XePzLrhhArfMn0AuCdUb9ry4+6kmp/qpLnIxUY6Cn+jPUCezv9Bq9jTUFo2ZlQT
qlN67e3jOLSzLxwW8v29SfuQg8jdJfQqYCgV/fkDKSwiRAF91K8iHn7PMICbKmpqaJdaJP2x25Fr
Dz+nl2krD9PsT9EaSupqfI2HhItmC3scJpwPO5H993rYHnSmjye++Ut4GXb+QdEG42W+w+E5bVL8
2yJG4PqhCsJJNkbCdPbQv/6a4tducFgNqtR6Hio1ApnkxPmUrseSzC9pcCb2MOX8h6MR+rwtPWDa
9OJmQILQXwXWNti309ESvdNFZeDYzLq/7diIX4TU7sNrN8h0jcnSzZPqqRQPIFu1pfeRHCdbbhIb
fSpupL6PagLJElz+spCRZHL3ymBFXtzk+Z32WalT2Hv16F8x/XgxIXlsHwA6XtbpxjU3gRGXVto0
6gJgzpYxQiNBrV6Srrv8tpFoIb275piC06T464/ueG5RUgjsCAEA2WoJFtI+KcNfgc/SLa/A2K8P
THs1h4bJFK8qKcp3tWrngXj480PCg392I4CZIf8uunRHWcpmZkX1SChfpaXkYreMDKfWqp7V49xv
Q61wNl0xNa9EOsb3G+9g0uZWc2mjg5+8ykU38HdSCVR+4wGv2R1z58G7cFdJPdOq5WTTGfwFe/5u
XPe7r8rjVJUUazGsCiOqyaMb/Nxaz2CG1ulhEqKoLBAbHStSz6xvd/Q7BkwMvZzJ0tDS3Tq26V2Y
KjNxIq9klpy0Notj33O21EtKE7AJykOYsqw8HxnKqs2mIm7ZRMoWfvIKaXdDDNTZmrRcukxSinwe
YCV2WmC46Dkc9956wuxDJaIelnSF/Ki3xZCRCI0p0HU9a0PBZ/oD0+MHz37YeHdDdFuZ5NPWyn5V
uqd/B19NUlkPqbkAsoe+YOMO2B0pYNphhddAcovrnnAc0ueWdxvQ88u9fQoBieBMKqsmN9Zwg6PO
bg5x4XrCwpggaDNEEWa1T8wyvZlK//Z6+KkET1F9YwCgVuCVMiab2ELNnZFuyWk7c1QwUpcyiPpl
KkpfaXAjA491KHcx5JVP5xjGjxL988oYkMzEfspfjOzPj2TlYamWKhnYPSWPDHgCVnO4aduzNqZ4
TDTIkZVeMCHmoHHhm1oDlhdWdSaa+fKliAXEgT43jECrompOpJcC/bKNxZyxQWCb3g58OEQn5XZh
/ckrkpszWxr7pADzdveJcmz1GPbY1YGPmjKxkdqhTLIhBKKOG7+4klCpUc5lC1iuGGsq9XufY1tc
H7LiyQTJJkm4rwu5dMuK3NM3PcO79B7Cn1vd4TfnVMI1A7kyTH5TsclpTK5zLyLOxe/JrtpZx1A4
dDlaN0bZU0537Av3eHzR70k4rEYHYsgRLsA/63QPHQ+ENVqCopaiu//nVPMOwsQ0L9kntmBqWVxA
iWun0cWD2I8Db4+mjiiMXXQnH/RQmhGkBluzBSwBAgo1F9/t/vu58VjOVspULhItyaxzjMLL/jCX
LXCDUY0CFSiKFF8jtHGJfgsLqE2zyeCN4e3+MWJCbZgqvNSaB4JGLTiyG4impXKoxKvCHe1y4G3i
0HVBiSiF4sOqX3KJNf1YLe/NvxeNLEw06PxjGUsFBk0v9RZNrudhCpvMXxZrB+LmIngRvtPKfeCU
d3I1t/MyzoX7hBes0uZwl3rpnz7Lfh6bbsclt6/I+LOxkWmcMqr3ukdBZMW4jpQ2dTuhQouzFia3
110DIanKeNRBAhlHl9wcsWHWafXatAO275+t5dmuFIkvcF9cjjAHroVBHn2wpDZvVvw5oMAHFHqq
8vBb9Xl4w8SwMoY6RKPFXSdMHbuZ17O5h7Xdc44tBYamfF8cmY0CxHEygAtqhyydgOUJczl/TQ8L
rQS3qGoKAKNNfWuC3Umxp06+Gb+7KsXlA93e5pRyaqTZQ8bOHVopUCXx7mdMU/RpTSCHESE3qE9M
JQhgpImZcczb+4XyetqiuyUroBO6yezx3eRfgwYEXdkZj4/lsrKNl+FCpTr5Rt6WvVWrSnmrmgHB
ALFVBKptX7tWw028aS93rKIyU3Eqcd8i+D2pzkGzwPYi8BX6fo9tO30Llr4vNzPh8ZkESeDBtaB/
KF6IFOUDoUW0LjeO7YvAWxUwDVSJc6QmWWWv/Vox8/m6SoC2apEatMfoPmDSxLEc//WuN5pPpKMZ
cTmbWoab1pib26B4H/VMoY9bVfaynQZt1xfAqNz34YkhY19AWtPQgKHXvzdBvPMp4ksa2q+JayF+
1Dc81b8b+nCwAQ7faihwZyFZBRMqLbgp8NC5/HNOQkvL1ZuJDbo+y7orZrpnqgNhShZ/ChS+d3ck
ARNwrViyr92sgVUN6iPGwYu5R1a/Ztbpm+KPXZzKdXsT7QNoaFkFt8dafBbASX1VOw0eQsO5GgD6
mV0YTbY9B8Osa6dqKrYhoGWqXxALLRWzSGKZguuaAbbPYWZRG1Z72l4+hTFGHpvotF6MYEHkpP3F
ftALkXUa8fVbfy5jrFvavcpRcLISsuDV14jCrcKpkFzcCyZbC1LBSvt4p36Zg8X77Mfle7MYd+hJ
9h3jM3KBiXre4BI40R5XS4skcsQk0g/Q1rCpGB3UFgHY3uNqBJYrM/Qbp4H9R73nZoaU6rABZQUj
QEasPZbMVV84ToaP/hDruwb5dCHC7VmSzYDwc0/AlrXvNyqgWT/pOVn+WFjcfFWWzgqIfbyXgOnc
0XnJrmImdDlNXt9IGzlbDV3FBONYUdfnQa8EkgkcD7PqkJ54jaI31Ld30QQ3LYpgqvqjddNm4tUM
LajTh/5DOVE7ozoBMECUXhm9v4rdWV0KxEewn5u6QOWt1b9ssVwiJicOesYK4cMBMci8Iu1iKfdn
6eJEeIVOhHWZwQNYpNa9GlnPHg/onuKXjO2/Rm5OvGG1jRXOI/MC2AfLiW1iMx1rrSVsdvQzEc56
jCc3kZxvIfaaGEYEymPdMjhyiau1RPPqe5shG8qXYByE3j5x/uozTiLpCuO65ktIe3SoSGe5FrUN
2x6BTxrEOxSl+n6hrelHeO1vRpS2sWob36o++Rnd1brpTyNgOMmlCI3XTJuQ1bt2c4nJxdCT1237
EzpvDD3iL1DnV9rleA1wVrlxuUDKV2piuxSFW/QJE2gJALEe1jKq/5FkFCeYq43vm1A5BoxkVsR3
EDlQ1xJ7Kl1qOkpCxSknf6w4p9xAOa574C3VZe/pjgqd4ZTSG2xvAkP3vBjWuJyUZbDWEDJgnTbk
uo1g7cGG/WYze08dIgiqoo73Lkg7pB0saeiH5KPRJRqmHWYChjDFLFmM+sSOmx73jBfogRhV91n/
XQuV4tQxv6bB5buphFIXi/61D6kTJ1aAMN+UyGW3d35AR1bJe+SqDg2PrFjYAIZJV4IcyZkcCQXV
WL5yV066pR70bX5y1dsgWdfaOR/GT8rjVKPl6/XTjlWdFM1YH+iMxsGtZZpufpQminK/jMXoGC1A
NlCT4hrSYcjYKuqqR8EfVAEBgun+vBUkZB0aWq4Jd3BvnUG4Cu96vcoYY2vxxzXqBrlmXf+fv6nk
jWjZXy4y5qDdGSJSaSXRF5NyHgjbrpoo7PhpoZWs2wowlGffOJw+SCY3CrAb1qfRfpH+BBfBU+Xx
iPx6aW1mLjBrNBFa7wHy/nR39HsBDGEi1u3xvDIlqopkFN1tgM8pZPKjcqb1KtclxIfj7IYbVt1A
+znJ9V/dHxeDlAoHOFuY0ZurZUfwZ6gntHMbrLievHbS8HrthvURTn5dpzyuNp7XHnHWtHmqluxp
GZ6o/cx1bCy4EoRqI+7WRwA3gchkHUE/TR/f0eN5lfQ/yC1I3sz/sIIm8ylz+JFOOP4kNxW0Diq0
es/g09+zxdOOrkocLDg8JyrAath2J5lyj+q4XSCuaQb74PeoU5RO2C+ZF5y62oz05H7Vtfla68J8
szuq6d5nGvud62U6t2fnSNeAh3zRdxgZi1KJt05VP01mtC8FgTf22dYsBCSTaJaB8J736lPYzpnS
YCLi8HtKybbjROSOOdSX3bpYIhtrutBSSi55IixEx/aCo0r0/B0Ywrbv+c3+R+6T2tnyw5w0XRS7
KNRrMGfxsCiQ2DWjNG7qlhv6V0ksz6WNqaCQ8Tj2HQd4ii8XnCCqezRG0Bk8FlLARWggxKD5nbTZ
4IjELkoOP9s9HIBqg2BLlu5QgIQnfc/t7mqWO11ZISs4+gJjDxwIPD3AjkfnduOS79Bvj9YF6b2y
2xu7OZM8mGFlujDysXk6zBUpZtXpWEZo3+rvjEySaVXzB/xjiZT8povoR6xKwihiw55Benb6CnkW
wVsYzQtZj3tVnhNqZWx8VXrMeaouqjnfA1oUftGQ6W39q7Y4FLrBjtx1dQIpt9X1oTwGtHGNMjw9
LxmSjP7JwXNqf3AdUD/Y/gfk8/SsRDr/3o9MnniIlzRopc4NaFO+O+Mo7IMw+ofshyoPs8nI9sep
BJOWbSAe3vNsSIjJMb2cBtYqoUC4dG1K/+F2U+53A9GdW9i1cBdNCufSnbBrulWMI/AhZQiQTAS6
2wLqAzRBA63mYtZw6c630CmsZLJc1ntmZ40Z0k6GnmS+vlOE+SWudAz2haBCSeGWs3BtnMDis0K9
bxiiKnSni3ZxL5Gc5Fi9ca9RqmTbXnZeypJGMof3gCVlv3CK1Wer3OMarV0dxdUzqGTfmYv8cFuU
AVTcmarJ1OOjTTBk/D858mf8qFESB6nEI7vCYzILPBPAnhiVxd29yf9C5PxU2GxIuAvMIv+iF4Z3
y9F4KDTlhSiIctc2JYelI7AMBtCRZ9Dx7pc7N9WQdO6VjuRoFtYDQIowUZZCSoVi80J3iXLuX2rr
gh8b0KUQbsenAmx01y8DzHmgLje/MrRX77JqRmtvFxcspQ/QeFXLBjpIc6gMzp0IIcXlJCyFWeAo
h3HKnx0R6iJs76bN3fDzc8ZVFNepI3c6O54ExRGrquT16eKte2i+ksOugjdd4/O4ZDMs84T++MQe
9013z8JkqaxsM0M+dXfnwPVonwFsK+zgEjCbgcFfBL3Nnk71owJaYsjst78SX+Mt34Awds3Subnh
Q8C5fBkn7wYXnvNXre4vB0iir2/idaHz0Rtvw539dLVmcDw4jt/yjYLknDLiDZCBosTUC5wq5n3U
MqLstAYEe+2Z9DPIcwy1xSZpGqwUSFBGx+U2KwYVGPY6aiNPYoYXh3/rtW9jtHcs4a5F1t4PCTZc
Qst4MB6OiuAEmyf4lH5QdVJrelpNLOSeHKi+/CObbtwONCQ8cfaTT4wY2Y23U7Bx+dZQeXzv7lj3
xF2gywYhiuHyxDxZuL6lEzahhmF57UloBVvOYahDfuMfsS6igMo8FZcOHVG7WJU0dQV9IFsjrUIc
1SDLb2tezEB7MjYwN8jQ86pGG0NPyo+nDoxYaFw0Yo6FGEc30iuEInNmb2gYodLQEduWDTHkYFBj
aN19ef/r5fCdfrSe6256NOv6Z6g9rKsd9mdr7jplhljCfjJqtXu8YWkwVcsbDQOKZp2g2fC7a5ys
NPURb9SShJsXrRNrU82DKBi0v4sY+vapHF5rGQh/0Q1W03cQhNTHDVRLP9ZnIx/xXXhNWLhP+303
u3ALSxcxqFZcNxGhTOI+v7qxtUXtjlYdHj/gxu3/YMdopENG3CCsqwO30A/chAErdF9DQE4pOuvz
NG9gLKLqd9WbmjF6fTvaN3fGgBY7j9iRRhONOONQ2FhUbZZFtia0GRxOC3ZXSoXFJslaD5p2V+oh
PQGOuA/GsqnJsE4iVmEjpxAQPecwWDE8vMayj87lqflGd1QsdmADzj52g1Q+RsXz/0IbydSZ16mq
qyFRA7eWuzjloRQwD1capOUAOVsF3FhXAukDRKTvywieHIQ2hlDX8zdpwHMDqZx0lCX3PinlkyMc
zQx9s8x/3VvCfWZnnoq532zQ/c101DqnQLGd6Nxz73oKmGoJtxhWx6x6U3VmSdBYsBdFLHkDeuVT
2bPEw8Dj1d4h9c++/Tk5YnFIcpKvr4PVvXn3VwmUI2845S/fGWfZZ0EdlfI+ddh23v63bW9DW34N
Hx9Au/iziJFbG4f9nYOHS1eCRNKHYUlvSOguiv8fSZB4RIuJzwvrsJV98GOlRFiYEjDX2WP9GA/H
DDD13FcnnXauKO7gKXYr1QEXtW+yyOzKZVeuwgAiiq2O0Aa3Yb8GI1wREeRFl326Jg/nmQzjseeu
m6ltCkULDGeBNfwjVUaV3QxPS1V4NWuWb6CncGdq5gfAU2leHYh3adM5z/4yjhEdb3sD0ShwDo8V
BAgPlO4I3yCuPq1xjT0XaF95TXSrBKmFEhcBNxoeCUzrRHaAPe32C9M0JVzX6nImFlds3PVxzgxj
eN7BQDxVi5WK5ZEieMDaFyxi5uLfm7y5iJwMdnWdcClQOdr3nbQZkySYVpjrhIHfD9T44EfvHXJ+
WzJZYjJ8bXF+j0X0cnjFyzZ1CzLCGBVv74plGKIEwJ+F9yQDCJGqePzARQ1ey2qeMrG7LDCkxosU
gwbUxzF2A5LJeSFS56k+BJJhTq2ZcFDfJHxgNaWUaViD0UkktyC4TBLPRPwWgc9NpjNMwty3gkvK
ZqXY70q97m+9l3cpre+wde0yyMkDuHBCHwVb2GxuMQ5v0MJZMRykTk5ocgvdBpr2YaOmYwP8F3lK
bd1jo0VI9zrfMg99xre/C0aNskhBRPmE5sD+GE9i6B6DGpnmnwYXEYmaSQE6yu4rB6otF4Ba3xZj
q8b0CKhZxjF/TI8hK6Sh1DTl92kNWz7x9SviFk6+rxhGOw50N6+OLrPGXofjYX6YkquKvizJhtV9
J+bC0OhRQBQ9S3ccazxWCrXqssN2We4vSw5Uv7tWUj/lU09Xp9+vBq+d5/crcTU+0D/l5gwYVR+T
x2Yoal/8IbkvNiAvcWX4Q3NYi26OShSIN+Do0c/lMPm+3s98Bf5CFfZzcOqoB/Ebcu5Jn777/z/7
RVf+QF9v45hHkwWBIaNRIMkvDHJHHYjtzroNIJLUZmp85ov4RZXFwJTn7jU/w30jM6nwg5Ol+A9V
xuqpkziRMtrEjnnz7KTQiY3OrCuAyUrtQgpWTURVPBdJCtwDRSvoOCE7/Yr39njB2ef2bKAEhP1b
ve/8jklMY/3M4HF5rMJpx/2l3yeRMswOn5OU0FFpKQXOQ0uh5mI7cwS2pjlNGYxiJp2NLISThx7Z
kRPyyRlMRReG29RprSdujz28lc7Rbn/+RMfEo5LCj6LxKuJFyfy56meomZQfXPI916U7umDqqx8x
Ig3WioYzdc+bE4b+vJp/yFqs6NdGd4D2xX0jMv//aEUiOryZeTPgf6Q+Q9tLm+hY4zatTGvxUj+6
WUHLMDCAqXuMvzVhzL70QFUBxDqeq9CMs3FQb5uKCdAv5Aluzy3OTAbjpfpaK3HKzoia65B6AXpr
3E7a/2LuwRikknOgCH5Ho6Eked6YQRrDKZLwMZz9vIXJicFYE8k7FMXhr4BHJqWmyvrOoFT7IfWJ
GjGfudBPEOGcMqGe6GJBmJxMtDikhCIn0wvh6ui58HA4/uLJWtp2Gj3N/6ifpnoeYDIqdHhDDlSa
bwdS3mg0MqwMs4LCfteoZjGOSi4BtAxGIgOCrzA4HfS9D/3k6nNyPsfN6by5+XfxbQrWUK8ErCWy
OfTnmecB8o/910dZPx6jfH7vkJeslo/RjZO1XH1UooPp0tRlou+axdySjtmLYCFhaXP9cCedEkoL
u7KIFZLvGAmM4IsagRlqaivAgAvZwkzxxhVkmKWlgvZ5LHgLiZo2sNZ3iDd9OAgv+5Jm9BdH8kUV
10/0jLt5MLR0CHvgQ544OlVHB75hnzfw7eVzEGN4ENrxKw3t9B0F55jpEvcfDzk58t3R8tX/XD4f
LjZkwEdwrsqgrCwXz6HP2WZY3ht0JQj8/omd4YW36xbNeYtFWKnmHzzRvLuz1A9za1vpcdKDzgCh
Td6fdG2mpMdMKk/LO96meoTiGcIcwmOKEXSf87QNZMMz+t2XL2s9k8Ksx8tQOTvzyHm0VIDAYIa9
Oh11tXoaie6y/hbqel9QeLhsf+IqeWgH6697eqdvA1APoghe0521DjXc9AinA1lp88ytUrY+6I5j
F3aHJniaCvLfJYokY3e52wIuBWm/qLd43609ufdHEaOWXVicWVVQygK5TqsABAVYtgBmf/HwuqhT
59WmQSMvncwSEqFvMJkyu+WkFqQDoO0ur3IW3tYM38fYToXSNJ1IU2JgZh0nL2ABJS+1uiwQqwMv
1zGq8FRpIbmIzhz7WrSxt752q4ulxFTih5/e33ucACInqIwzhJQTugZiUlHbtvzqtqvywUODvzbo
U2ZBSOg5JgCimIZhIQSeGXOH75IQTvw11izyJbUHAJSTncoJ+AiD1CrmiKb537mF3/gCzMrDZ5BX
w6NhsEsNv295qIutqY5GXuYgf/fIGqSLz4iXmcIcfRebKD89EkAPT3hD9dzh+bf9Me48Xt155UXM
DbYjQdogLU9QOCwfBUmaYacUwVaYl5NxSwJpdzczwUXFAdFPAvkJkr0gu9iLRBvnA4rHYhQpPTuO
/xhv+IXFhN+MHDeR1DtGtE8G5qQHSDMxwNyBoEqLfq7n7+sdSfehxNYbk29eFEUObHaNP4zR6s8D
/uN5EI7GP/DU9o86WL0FC/Wy+GWuMFI4nKeAzkj8SFqWq+Us8AWO7md3RHO256pV293Hw8sFdRmx
ro73CDVIv2zXDB6t+lpXYUXlLMVyI6yRHwNBT+u40sIlALy/mU6tITGTCNvuhMCfsZ1st+WGlzP9
MGAI989UljRabIj7Y11+VqoIYWaDzAG3LBKE5wsITjqNIGtPCcyWTOWBi/scw8LhWKt+v0C9XnyC
uT6nCXdN8tAp6tStnRsFW3o3DREDY4++Tr9VQJKVytjyAHvBVtuvZo80fDC7quowrpJLplKFcCX7
IRKT/AyTT2XN0zrSONZT8FCCc0wJgX05gkHohgQNQQzygUcwJfEYgR/nLjo5H0e5PQke5Dhq7esU
uuDgtjrKpN/YAfuEE7dCc3AyCU/Q0sa2IDYSr9BxQMgbmg5wC0NejF0tFSudxNUIFiCywJLx6i/s
/Y++OiL6M0vPDO0gtXdqrE6lDhrV0Ts6Wd5E+Q7QMhOk2RKBZWNlzNVvaoGFlwaMW3KHzWGp4ANx
TJ+WWg7EviWmICks0WGn+sfW1ZeWGEV1mv+tyv2yBmnxVV2qXGGa4ODJAceBd2FIHgCO29oEUCzQ
aA6DyJAlGs0c9VrJATL2UulPOkwPDMuj5KhxylzWabwTYmoxMwv166R5ozIffVA/XZ6OUyUYNhJ6
mLx0EDPfdglrVGZUQWKFkSekBasak+z9Cm6eV3O6APrJl/ZMcQEMp5R/s+bt/ukeAp3ddoro0pcp
dGMso/T+xq4P1dKrpfKWQXyIU8m8Bo5aQeubRhggP0dAvW+Zhhk0kc8EnaYCuaVwZ+7U1S8+2/ON
tPW0oDg1qSDk1ToPSkh96koyuGw6JGTL6CP5tqeBKddQDvpEmAXCBMVRDEqkztZPVOO0SOoLXdVT
R4Ob/ZUN9yMXuWp85n7Yfz6PDAmANGIjTNKe6bd4CyG7iPJ6DTsOK+g1NzETfg85n0XSTdgR6kqv
wrwiLkbdaHDiBsSX9xhh6eCbNJ3S0sLCnpy+glMu26/zzUMg/5Q+14gvTcSF18WJPr1PqPqaAx25
TT811n+Ak5cxSAi7+0uiWWfNKzMjKsc13qGVwIRgQVgozzMHnIkKDbzPHIrLlDxWPLDkdrTXLaqh
nakAD1DZRf52zj0JzuIkJVvqproNmxWiYtL0S3DYHdJh4gwy7Fv2GTwgZmywx64BXqSYh3fbj6+T
qBLwPaWu6A4BSEdLHSPrNWLXjsVJiPC4fV48wnkC8unbxJ1sQMG9W2gn0VI+31MO2J94CFzSsS1i
cnAC78MSJ7qXxixMNtN7T1d+x/ZAk9H8VqHx2yavFT05IuKWUHGL09Idu6YZPe2usEWf1ZKAdbvi
H7R1qKLDkhtgtoZs6hr+Cj2wVgZyIQlm6WEgLYG9Es11Howbzoy2ojgGe5+d8J0qp2b7/Lpu+ynh
0Cs6BWMtH0bq5EckLVDKr5UyhOTe1NVHDtefL+vCSea14PI+2OSRV9KYnuL+a+2A622Y7H3893Cg
rCKu6Ql6vp9Y654zdw2l2+7/2Ltpe+7TA/pJFroo6j23lVE9/O4PpPSIXJcIhgGTHPTbX1kng85v
s3R/mNlBs2c6FMI9UpVvQdePazTvwHPvrMk86WEHLFGxyNJJbCBH01777TP86168sTV5ptyRkqSk
at4J7Mkx21K6gS932bxPQpUeQeI7YCEU8Ks3KPBrs02IvAx15b9AQ4b/G3t+GRfvG6c7P26+ZcZn
gSs+tffZxMQws8IrTUgKFBVcjTPe67ixW6hPu4SNrYFVXMQeTYu8Z0l6LX9pBf4nJjvg1J6Wsm9m
dkCRwpjGiq484YuHw+JZJVfnWkJjZc6t6L8p2pE3hqftVp8Is6eKPv65h9qnPEJhiu/9uwiCR1NW
9/hIPyO1MbP4S5hXizQWBlPQq5ke5AZp++L71n/QtQ9hRC/fAb3jsECDbgKb0wtSEnKldt72+Pcz
JRDqHaY+429tq3uIKTNlSUpmCzbRNkorR16xWnTvBaG/HuavxF50mTR01q4cE2ig3ODxaZPWXeph
EZOEy3MIGr/WwFdbeEb0TZDvCEbt8/k/RSwXffXZAWTSx2z+zFAGFL1+Hsnkds0yItZqAEx6nXMN
4AjORSeK1frvpFGpf/RIpNBt+KmzYNpnlDBWSjhgdyMzd29o1ClEa3BlOgdvnBMM/p7qqbhxouDY
N89oV+JN34d2rZTZ+5o0I44uRFXjUeMCieedOX0nNkyiFyeeWTEmmw/Us0jtnp5AOsggKZ86Qfx/
JHHQjYQ4BiR900/Iz0DdoHS79Rh6rEn9f5rjkkN31URF4KqMiA1UxGvIz6CexZPaiJDCJUWmj3xT
6m9GhC6LJYNMmgJYFtTAFYcGeYCZOgKpANiqiPd7LULeh2CpggHiKk5lY3lVGWds84s3PpCNsu+d
ZWArMyek4mQGuP8Q6TOQu7knwoHyg+RYk7KA0LSe1lhD5kMDb5/chRIrMbvdh3M5+rH/En6OhM1a
yzczL5zudDqkUXtmbGXcUkRjIs/7qGa9ISXK+K2LEHyZ3jKEVJfWypuJtXuQVvJCOCL2CwZ5KcRj
90atLrT8Kfs2j4MOjUKibzkAprF+FvFIcNaUyzdUrgXE9uOqrHcqQumnBu1AW8K+wtx2xuvXmIAM
SXASqNnZKB0Z0zhmpEJTn7UIUSg87U67z95pWBCErFz7ovgxe5wCd9onxR7un3T9TJcRoxRH9Rl5
cBYPrlZSbGYwiarNRNGI8Lmt1Zpmda51eU8lduIjbCaL3d92lugIqD6tXbVALc/LC6AeRrn/5SUI
MB3KM4yB4/TiEhwxYOVYwUfNNOSh0vjCYPQPhZfkesa/LnBLr+lu/UbRc313j53rH7ErgZyQdrp5
N/nlwv822GbPS2cmjEVlOJEm1ETnebMTJA2MNvRttohnhaL8HdHsIEJyDWV/Cub55yJFcLzNapMq
9O97ucgh73XZxd1QoR7qketWU3g+HYaKkrjDaNzlY/Zv/F5DtwXcsjIsMsfmCl0SfQC2qAfOn6tH
PC0tf9kdx2ztf5Zj7dsO+EXRb96hJDQKC21s0dTISi+SdC5O5YjfTMayNvI3vh1PGJftbFqnpa1E
BwoNhivX8SRgEmKa4w2mk92wfGLzTV96v7GKnf9BPgDgbDDR60jsYr0fI+Ut1AjCiFjJYjGgyBZd
bBw74g8D1h4vqQ6/TPd+5YzULUJ8Pljtbz90F82d2b1WbkLmL+nE+fEAzfx7immTRFYMVEiAyUww
d2yQkXh5chrnVUMoQ2o9B982wk0ju8qFJUUzsZ360DHKbalg1+eiOelnSUKIae6slec2vlcmjD60
jp7ztInO28zqJUYeJixJHeWFdmvSG0pv4u3Ia6+fE9qOLacn+LHyWN9e8Ax01BKD1Q8tcR9M71tB
1gn/SxSjEQhEZ4UbM2eO40PTXeHO+pEZeR6VxYGJMJrb/kSl4LouF+LvMryhCDypktXq0QDyBsON
+tjkvrToKCR0pcQv7nPCyEL17i021pHvcwz2OxZKKrH1/EATt+1l/P1hXsmbyTZS+g1I4SeKLCZF
n/ETyy0Mngt7c5EYdrarObtj3iyWKR2ismW8zHeNh6W39SE848hQqi6wWam+QgQhII1C6aPiqKPS
byXbTueFY3A4DCO6FXV4ucWJ4X/Pe6jJCdZLwhwBqTRE6RLhLBy3J9mgCxxmH58YXLebQIbXByeS
hb9ncZ6gromjaNUfaiuG4yp6qothK292p4KQTGtcUlHrNUT66Upqs+WKoel+6pRjfncFwtt6+Hes
yc7GJtZBIY0TrjGJJcrxXq2l9VodQzdMppA6rv7BeSdFrBnXOS2BeSaIdWE5h04nyQ89kHlCYPPE
Jct8UcRNQ4okB4k+xyXWQoVU1ixLOMa7sG3xvL+W+7d7ceZRkCktj+jUjMHOB4kl/WZi49xifazD
8cTfyi4jsZLmtNOa0Mx0C7MEh2gy9PAMsKLA72nrVdQ3PVy87iCoZ1genIwZxCL4ITrQeqiGmHkx
ymDB9fsNecg00A5QxikKs7Z4C1kl4JHQGja0xERWbc5AJ7XrdWRBqe0H3zQ4EIF49a03pO/QUfCH
JeFdm30aB22ZaSai0Tc/qWu4r0QHxPZsBDzlxr1OPgoDrD1Om6mhmCX6JgY+SmaVa/OV4W3iz4wP
YDlpjwPM9uGBnpYIppnYnn9QIBMCgdjJCYzh104t3FKCXB4qs/aUU3ne2Lkuq2aVAuOsWxQ/gDdY
NCheGnmUX104jK81gm01ceLy0MQz5JuS10+BlZtOZdrxRLv6GYNkX4FgLe28ukjZiSwH6QIyaQjX
neYTzsKO3rvQafdTEhhStwfyKkaTQlHJ4GEvDa3seTqD4PXCdpULJ+sQ4SiJirB0tj8juT3e5tEp
b8l+wpuizA/s+KfGvZOFe5xOZrFXmBxO0/hP9kWvaYIqaV2V3rr+QAPzKPOt8rUEWpZ4LvQ1yv3H
MQ2Q4TTVQam17HtrQpvJEeMBa0ZsWhofcKRyv/L5y9FyYU2YZ438h1ICGy7rfg0lOjfyB+LuU5Rw
p6XaXz8JJewC1wxEP7Q0MAMKo5VwGeXiyC2yuFpp3XvoUfdApnjx1dUuAdqqGXhVD8NTfDaErciZ
jcf/033dQ5B5A4M7KcGtwWDLqfpjsGGwuBxUR1tqVnaIHbGfk3ZYFv8mfuYIo1J+q3vDYZ3zegm7
sfDDVnlXPyEl1pGfds4JlfhX33lSHq1khNigMOJUTsyWgkIhlDo+NgiQ/H16iIhy9f38QBe7UqQ7
IDde/Bth87MIQfJ3hoMX/DcihqbPqlf3nTSh+Q3czjDonSEUrLrGwJ1e3rdLAIyF4Of9iDhhxumr
WxuVitHLPeH7XZjasjW/wVN+ksFUdtfwrPpShrd+Ix9f4cH5u1uj717TmAZEy6VZRxnrgtuQtojk
F17B3z7jR6RGXlzySPlXnp3oZ31mOlOiqmMQ6Nn/F+h6D8DiudGJnvlukpmshc7FB/xZRWAJlmBU
W6JhCWgHr0x2s44dzfB/QZaL+SuSRKdAe9lcv82FMDOo9YtYBrrxeOVDjpmmxyjKt4La/lwKHVPo
Wg9xW31BhqExtqf3ZOPyzruEyDJLSkHGJpKGHsDzXBgSR8Pkm37tJ5pDA31jQOxZzr2RHFVeLfQR
nnF6gUNNOrUv9U75Oi/QnmgMX1iaRzwOybz6mou0baQ7XEKdG85giR9iID+HdvcmEtfqyofYEzTG
vnZmnzytZ8bl1kgYp6PV2Oh476i/NH76Q9iLGdOsDba4D4HARZukMNrblPDtv3rKPl6jgAuBl48g
4xvps9ydvyRnJ1VAHG8TgZScbAMN4K1ENWGGT6Ds2mjV7ZFQdRCbatQb10l/vvDPUaqiYf6GUZKe
L9hSkfIA8yo8npS247+dRc5O6n5jh0LenzLrVS/Az6K1wUCOuvuvprSjsggz95O9PAfHfPHviDGd
DmFJjPF3ONywnA9Kk7Et9iOr6M+Zs76/Jbgv21eUhc5rc/PBriB2kPg6s+hhVZLd1h5paxFt8fav
gJZkB9w/840tkEdCzL2h1unbLvNIvgypjPo3RY8K842QBfunn7CvjtTloMyeW90PLi8zrk/5JqX+
MJBoif2AxMVxBYkL5s6D/CYVAdaqF2fdfVftmN0XZC3m7SJY2mV0P4My7IoTDx95aT/0jgLw4ipd
gRpuWxh0AcbsqKTHp37WUWARbW1C3/7teQ5KBYAD7SjMkMjQ0KB7DA7875eHkCRUsXPGKSXk15Uz
TOwW0m7yY9rM321jPXM1YOr8a76/EVGFq/O4nwdQBskFCZS0quE3Pa5dm7YhrPF9c3dowVWWOv0+
8wSjiBPDEaQkMuEvaI35LeZRddR16o4HWWO2F/qs/h1yoasiy6EPh3CeGuSTnmqqdiWdNe5YV268
yX2Bm8GIu74Gb/fM5VanZ1BkzJ62dzCdO6MXiK17rDbdWtgQ+kIiLX87VtAhyFqLosR0RaEfgIUk
pD4ToqoCKVMlFvJJMpftjeAaZC0OPL0oDaqSVV06BDu70aPfWwYRm5CJFsxfGaMmm39RABrlQAWi
r36x4jScQXHw2aWqSY6nyGabq7KrMK6VA45WxAuTXk5ljqtgUqHv4RbnKDtUDHoO+q3qCCmwwZVa
tRmjUuzBchi0Z0u174SuKDYadeyM7wg7ZsJiM1UmLEkQjDf4/8NB+VZGKE190TV4c2BXZI4g0Ti9
u/4QrIQQzJU5lwVtmQPg+7wfDUSr/XVLxG5mQQkAjUpp0W9oBged928SIr/y7S0DrR8NjXNL5MlP
0RnL7yrody/Zl3UkKbX5XvvlzvlqrUOxCkpdnW1Qd0p44YHqPZkoqUa8O2ixmR7nEEQqxdvT8g4b
VFJ5lPZMo9Rlfksa/jSPnghoamnfKNZ27QTW7K1vuKbMIyYrEGBIQc5EFFl/pZ9kd6VOZctOuSKc
a4tNqC3lIv8TzJ13lgjdLY08y464muR6AMPU16r8ErN3aV45Dbz0s95nXjcJM+6QTZB3ir4yj40m
ex113nVLcDcwYCS++aP/KugeB86F7eSXzCPMNDznzcW2ZhJP5RhwAXrJU2w1sul3DrFyE0nxrX0W
CMJ4QoxfHC6qVUBGpPeLG922pFQtXPn9xsnucIvSXx/NFCjB11l7ejF0Zab+ZMGbeAt3n+TM09tE
HYp1A+pGVSENvfI3bcwSMxTuXBE2DcU7XXOPWbxhQ2X1tnT53R/Nm15F/Dv9dEADVbRxk+TkPx8T
awxfM3TnEVM7tBXLoFGos9bh/YtCCCeAYecflWKmVfBxgf6+yN2hIpwYDo+Ap2HETWDXuPjbdGP2
md9oK1u2MCVGMx8ddEl6LPPtNKGF4IkMVJ5G/Yi4KZTZ4lf3BnPajGQjo7wuKH/0luFkW9BhGMKE
P51VenKuJJZ/7W6eGLotr4HtHssCeKpikbL/EBteeAauHw5ptuiks4FXgRX5r6WIfInbXZnmPVwk
ersQRnMVPZKPEhu95kDAipKUST14c0ev4QnY15/jaQcxJgPKjnK4j9/LqT5fCU4xgbJVaa837CLE
gx4zaMeVkgbgkgydmitn0FZDF1r5Y4F1w+hwd2aw4QRraO/8eIbU5y38TG1alLhURXZ0mut5Rvhf
kXBVmUWmSNE083dimMS+K5/VdghKGoRHqRqdEGFeBTnQSKshJoIj7FeuLq7NwOn+YE/XmI+fnk0T
0fu22dh5hLyvFktL0vPD0TYWT3veZKqIGxKn2nmtR10fBbx8kzaXwXCVjXZQ3y2uoukaD7y9KRds
AIwSor4fgR5BSffTZEMwSGl709bcS2H7yoyCtbhGzzu3vrgBTNlqryOEejGvI/D0OafhjTyBc/N4
0qKPIUFhDFyxqp6jvwxRtQylasUtNL2HTv28JELBr9Arr7k7oCwKCNhMVycGIJ2gTSxf89rBG1AW
Zzcg3D/4t75GdNo7fQA4albIK7SVDalOeUKPeyyJxdHLIekOF/yppPu1QqqGxXP15XzBS8kC92mr
LlrrImjr4sOH0m1h5OlLTUb+Rag3CbK/TxwTK+dIHN7uI2rVgLqwAQzdJgr2vjxe6y/RdVcdpG29
8OYihRys7eEpNgGVv1CdGiSCls3DY4cH7ZDzqDiABUlGNFDkIssPuKt1sXV4biwwzU0VDZKb0Isc
l31hTFn3DPFHyLFyP+UQkjMONchJICQM9MuKVAfHssv9XCOk1r0b4AaWfPmeHCDD8f3LOE8Dw5pI
5ZJNnYfoZ8xDx4ez6O3A8IS9TaCrKYzu3JY3FYYbePjget4QY3AleiDebdc/1/sN4ZMG3MaNG08O
Lm/H2uGXqb8FLTCP8Dk6wCivda29XwD4Wq/HIlM/y/mhx5cLqiJhXzf14orM63J+EgyAFTpvLtMg
XcDnSRXZ/I5q7dHnFaT8BcLvT/DqzN7IZhcLK/qIzELTJ16aYZnh3/MKyNSZdZDqsKgmWno/dbcG
sIEIBQB4rSXcbb1Mfdwe4x6ZT+3zLtgafktFq4GEFr0ni8zqn3Kr2dOM3m4Up7+yLeshlIB4NpUc
dbFFRMYrA0Bg6zt3zWMDg+RlReiTzDKS1/IHAFkP1n6N6oIUIaSDPTBvN33FNyqPRpNpF0uqn0Fa
EU3M+svawpX47BuzgGY0Nh03GqSBUQR+wLYwsfo9fhcHZjqMwAJ2jHweu9xXphls2IIVuGAO7A0g
hnNV5Fp2cuKsziD4OpBOQ7wKUdwLMSxdXQHas85gEbbRoF7n790udS92i5HCB8mUCnq6y1SoxORG
vQX8i8sCVKw5scCwdFeTShaQflKcPX8UQ99yf83G8zkpmQstmu8rVkgDzDnFhSBHU7pghz3bik8S
mu1lY5Gtfm87LQr3oLGJrt4ZhjhKJGkFZcs64H5HNo+fbUQfFXmeC5VrfdmBOZO0Hc+w8CeoaEvl
2vil3wsiRmB3BveL6eqMrk1XT2PHYFHrvFb+/lJ/7nmmvSpWWI8Nwbdk3pRpeZfuILCSfd2CvReU
4knwLpkjJDspVYQmsJFCMeB3Y9E/yy3i72Z8ZNUlhfNvn12xAa3Zd917ncJGCXXFIGo3zjreqhXU
Yl7YtIE+o7GpNv9K9c16BY7wmHqyYO3GIqdmmWJj5wX/x1nxXTyDMBX3Gv7YhUlLYRQUUUMDVuXq
QGZBoDuket4nlj67y72G1Wa0T3uJq9VaZAAvk6qesxjA+s/qW1GLb+Yuf2u2FNdQBvkhxLHd3pbb
Mny4YREu6CeB6TYxO/+T8PTPJ9vhqCXdiO6RlxGPzqqovSUxdcDsv+enyP4SlLc55lRSvl8Dmf2s
ENEnALazyGxFWd64zkG3aR1+5lU1HS+m324hG6U+RjVG34kWhlHQXxqXWD99u7dig3oVHOTVHflz
p3CbE/VJQcdMVehdk/oEBYKziqJ50S0EKcYyRK0i3CH0cTjvxNk+X1muARAMT6b5Q9azQIPaCK/U
r2pJgEKxECAc9ye/4ILcWO1tU9bMj8MLLBXDRJm9tpDqP1F236OJtRSzR/xH8bTYUO0KvB2VqN7D
3fcQ2ldeUTF/rkxIthsGxQI6GGYV30fu7m1HwkYvXHCFF7WQMDReEcuQIK4aiKilLM6jINGb96fi
RjfJjqhAtPx/FAzKnEf3ifYPx0fEHfqa1d8A2lJmL3AYDXGbPMUy/cCVu0Lj+X0hlw7Uvo15ZBoZ
nV5Ueu/KEKk3+VgEIdVUhNhM1G2rC27Gs9jgsPmSRKXw3UrcHD5ND/x+DZ4dxDRkx8CEc5w+N4QC
Ri8XTszmR0b/SRNMr4N8o3z0GQ8oxcniw4IGd2RVYZxckWCUKPtauBmU/2exDKcoHAMKyCRJhiuy
hc6a1Zi2XO6wa12s2rh8w8p07jg9SEVW6hYk/c7zpGrMzk/q3AiB7Ln8HV7PXOFsMyUNg4c4uzBr
uDdQpWDlVh8FwnZaqpAnZ2QijliePnPPvo8G6GPAZLVeIpWEwO6fXWcueZJpaKX1nvizM/Nhvq9J
6tQRRkR0XfI3h2/TCEBahDVOd92yqOn6UlOVKTblMXQI5y0PBS/SqId6GhMIrQSDNXYvt3f07VSP
Cs89MHqMVe5jm1BqyPcUhnicUimu7AHKnBfIKadZYKa0EsoCFlbjvlFUsDJjF/EIP89c8M10wFBr
RGhRIZJPXW5S0QVWRlZgRMHvLJ+hQ1ykP7nCbbx9kcutp8IuapwoVwzcLkQTuVoqAeMCnHDlLvna
NufNgYivTDklf4delZwoLQPyMEFc0aXngUtDPkv95IYLeQsccN78QeqWcCMjIfWVyn8eliGHwe9v
BWU9eNvQh90n7E+fli7ZwS1BNXXKKd9yEKCKbhgx+F1SyrrrDNiLrWPEQivkiMrGMWU5O7MkXZRy
xRA+B9kAjYjyseFw9Jaua2oV/Y7ltvvKmdnX1piec7Xt28axqZHgsCyxLzwRddatY2HMk7NusUiY
5x3RhDUCSNnBDNRDpnMrubyDmUCnIbGvm+mLpy+6xFOXyjl7nAoiAz/7TXSp2uuCdpmjw2u5V60u
EpGp1f0B0PTftUCfjo7gZV5m3kMgfBVMG6T1eei0i9JblRrVPMtj3CFi8fihDNDLg1W5vpJQ9O3P
HDYPJuUYuM+3zgVmAENcRKa09Z/ZqfN+SddmCnEfVel6AOX78LHrqE2PiAOy6vEEvL0b+xPWp8kn
eJYAPXt2vQrGmxjdiQ+nYHGztWzTpA0nJeocs5MzuWHKaJ4aDh1XNsC1NhhVefKF9hozP5BOE2YK
Xhbp1njPlFp4PysXCMTa6zBAZkz4azwQvM4Z9vMY6kAYZd+REFf2GsoAtgBFXUHY3QX+O4Dc8lzR
Z7XWbfXjU+wmgGgVWS7h3Oh3Xb9n6cP6rYs2K2Q3pNJnZH/my7k2MEWLdRCwn+TFg9AY2+I4+qeM
2b6WVxntc7TqfO2kpyorMC4Il5TkUl5QbDmQBSr091ElgryVx97IXFglwNZlDfICgZLl6FYTovsD
aNxlNQMM8gtZPQh1R9Xj5KJIcGKYuSXvXnRbx8ZVrrlxdwACGGNTHKqmDXm4CDCqM2gZ8tZcYIu0
QhN0YpfJKqNnnyIzTiTKTBPpu7P9ijYz5DdrrQ8D2sB4fwum0/imIRjWJe9XKHbkgFIJ9BzTBfP2
pVZMtmQtWqf25rIhWxVpKbtZQAoWVlds2UrOIdAOxNksVQ4lXu+UEPhKIKFeymemVFaKniS//ILk
vyTiREEfqHQjIvOOu89P92iW/bB6FroK7s9Jr7r34JpGlAfh+/I5HgkNq97a0QbV54AefG849Si8
zpYR12t3KyDLGtwdiRzQiJOjpFWRUyGUIya3up7410Z7v7+GKtUEDQVCeB6NPU0gJuzoAAQ286Ar
/khfVwJZ3UDqDAejkrGjlFVDQdWB2+qbsJsTAA1yQVbaqxmFvQqmqbCDLRkNUtXfJwdcUEVVFopU
8d0esz2pLvj6BoaBcUXHTtF3QPWkAjgDmxZl5dA7qL2HMk6TsSbJIh6J7RIj4ggi32pKIV0OqFOV
i4Sq+Tt19HnzKpk2UeNev1ZX/gWykMk9091i2pVGG+hcBxMYuCzCQTZgNPCuVrlXy2pnBgaZ2N+m
r4r0t8ZeGOhyi34q4wHgdmeyIk0zU5mpdbLCaKF0A6hpOFsXrbmSx5YkPqBunWwsNGYhJ41VXGGL
7AhvSR9usgcCvWXRkBHRhBPXvtVwR6B0xIWmjoTFZeFzAyyYcaO7BpPqGjReX0oVD7kxFvmB+Qp/
JAxDZBRtxPC7AY0erXC/wqsHVcqjvJCo+mnQ6ji8k8XtYzqrGw9EsjEFyjtkPwkzC8m9a1pirUAb
VBbqEkqaT9fYvcl3I1pv/4SoHuMQC9EXA9rODw1sFOp9FfQDn15ItX5Ig3Bq9HUcL5hM6ev94OeK
L96o+bGV8EGSxJ2lIwnfOSFf7Am0c0+OgLPKTriyjFymmhihPtrFiaKq8wYSskziMJruxgrdCvlC
thblw0x7NfJmZ5/lJs+ZQW/QCT1sF3ZzJnj5QdRvUPFGIWYzFQnW4lEtiX627m7OUHaMDRUDYLRH
2TCkSAz5TDyiSeZPtZOrbHiVTnQNF/ebuubQqhT0/5W0UVyatQ4jkfCWstTB6p0qDM+qJssUbGZW
MZuSi55sH3pJLugSkEp9W+gjIhw3XutUqqDGq+raqhfYp/iZyqfktO4h/aY+mfgKKQ2uPfpr/ZDv
e2yATxY3fzLcW3gim10huYF8BiE0sWbuMdDVpTWAD0Ko83dNCaz7Jcgr8TZ113AXbGYV/md6Cluq
38ThP9uCgItkT54BDQU0AhPbI+JaMDVeWZ9UJzYfWuVMuPUaJei7kg7XgYgEIsBdAnZ7xOj76F59
EZrKPA94s13WzXw4ACVG7Zp3G3vsB6lum+mpJ9zbLJDLev0q9BqHlF0zjk1oqLB4EyRqMgOAatUR
YIo3OxKcl22GHw9IYuvUBG6DJxaCEhrhjlA0xUmdhou3bYYyqv4tNtFEjR1WDUPmIdqNmHiqSTDw
43XjK/3A6mTEtvEC5DkyPtdPbuI9oxkpnI/JJYAMefRnuqA9Tez/8AHr26v2u00rgClag0ZpgqK5
YHmvbO1OEd9bk4iugrV7iBvESNjh85WE7B4iNba5sQ1a9TVH+1nUPFtPJx6kDIZ7myckUrfs+5U5
6E1aVUhAdqG1ymVBcmRzNvujbNAtodutRsZdyrzsVwZZ3ARu6nh6Owymx2d696PjxPzovhf3/Ub8
ud8r6LO5eWXAka3cPAJUAvFxCbE8HMIUnG6U3wpB4NxTvDqfTSofiTSbaXDMON4nO36p6q7VnLWW
jiUteglbfZXtGVCC9kz1QrjuhsEqcOTu9Rkpbn0j66ux4YPfGRMRnPeulYT97z7biJpRYNhenbOH
Bn5GGDGIG1rfIVa6ESVIen2Xst8YI2vHZixDvE1J5H+b46/ZmvNnkNRniFDoPwIo/K36WVCquN4U
rGqHZxddLYgzt0zdwaKvsooNzVeC5p3HR2MFbuygPUTU1y0Slxy8Ifq4BtPgfevTJXJBT6dtZzm+
WxDVfYkfmBmZ0S+Rjfn7NX06x+xMGqeXDS8gyfQIg3+bAAWiFabmCL/PWAXtZH4dKx3eyOPCL0XA
1WxVqCozWBvTAhPhFPUKHV99useXvcZovtvw5kUQAm+SnjyqzYjTDeeoOEXJ3BuGx0XnYwAFCd64
fINDs4EuEv7R5/ShD5MYcE/Rw98TqQyEzR6d499bR5rKCDlQs/k7pRnQtQn/RtFrMEdLY9i5nvDd
KZH+//Vtoljy45AfdfwzAvSFpAWDreDjdH13fsOwMzOIrN64pxa9gD1kpFXuwPWyxU8ud9iAvzO4
g6rXSlMrz9Wk4uACAFa96p2VGJMaeFE/BYBrbinDAy9xFEQleGquqSQ2ScuaSJRJeVViqfdo+05B
OYtitf88ZNWx5RURegLXD13ZuAb/IaZnKzJteirXn2dPmWEivEJymPHacoWvaRnhhc3y8FGPe2A9
dISb0Sb8ZCLivAckH4KnWNJU/H3DxyNVcf5BrZQ7Tpn3OTVf/cQOS4DSsEoL2p4Q2tA8m6SeDTz7
YuQO2Lv5MpKXKih5VoCJMqFhCNnhvH3EGHiQtA10422jiUya5HGSjdT4vUriM79S9f/mhG/eZqG4
ErOnmmeRS/KoAaJzlRuzvq1zU0CdYOAFMvY8AEdM39O6V4IeH/OSgI4rA/b4gb0yHEBbqmiiJ0bm
wxEQ4JVPeVO2agqTbgQ+MYxx8MdbF77X0VUaxqa3gfXJqTRMu8hl3eg/Vvc9CIYouKn4s5oWsNCI
mqGx1t/FR5t71gWdwFxdpwzMoRsVWo3mkVvuSoAMJ+gGFa5GSEHNqOuktkD4b8hYg6z8kx/1Qo1J
wSJjW9yvKYRrHt8p+TQfNRIwUI5NCRw8LltIF73stnL8kJ3+LmDf3dJG5Z1rVU2voKrLTwtaQpGy
pUcbYa44AIRZF9sae02ch0I00iZezbKgsPwginFKnDxOhvWTNsM5eqPDh9lhJRjkqwLMjYOPfHDi
mGsj1IN6R9rb8IBGy5PY4cRjlIqMM4fhtiW3b1ujHYG+1EiLH+nASwKMKFvww1MUsrdWzwicwOXO
yzsaRUszNgpni0CdX3pnZccQgOcQCRalfhZZ24uHyT/tGOulX/+gOxcERhmH/FksEd1hk1alOwoR
wqgxPa9uD1wd4tiCPrpzsJCXIeOBMhIy1DDYqU8dvfJuAW9Fts/Vwi/XSmdfNcdNjLAfycLEbk6k
yD8J7q+O8uCOBQyl4orK8cZCFqSz6og3gVkRChcSCNv9gxigWaGwpegRNcAuml9mYoHZ5A7XSslV
O8v+liZGDUoSkkmptG75lfkSt7spg8PyHNReSi3SVINZSxi5xxqjhZuMhcTZXPMGimry+W/L1pVH
/BwAQ+8wMN8stL/lhavdUtOBA63cMpx2Andx+dxTBkfjAVXIt30DzlJ3zk1P8/6SZXMYAmbWo1Za
Lk1f9Nir2dQ4PIT/kwTUAnsk4x/cvxk8qbapjr/EHnUEJ2e7UVDK/9YFYyGMsPgnyamqsp7nCRuN
bCN3tu5hVv7fh4gDcETmuxbwIQDnwoN2I5Z9/0dfbZ9WvRpBKgU4cmHJKQ5QCW9nKUDzzI7QMrkW
vhrksrovKymjDjA7FKMQ/FRvy8aO1xB7AdgqoKqRdN0ju8ho8g6YUSCzU1iCpT8VVdsRBH1pUAEk
fzhM5gih36PrbrjPd5+ffMUajZZrdl7Kt6YFxou9MF4Kqc0gi7p5fpDjTz+halRemJ4PkCKC1aXy
TkTYUha7sKwL38b2iQXG+7OhIG7Abuw0wj7/GBKR0N1tYhK5ax7Lk2ITBVTAP3CyZI+IIbNBX5qc
PeIZVy3ef7WkQGRC16B3dUD0v1iP2kLmO+agwZELZ4s4w7SehNcQao3A/IdrhDykh0hE2mtvXq6T
JmliC3bdFTFYy5G2o9LDbcSAhaNygjf1HmfeWtjhUuI/w0vWq2QnwV0RXBmopq72yHX0InNoNoca
0n19y0cb81Lb4M2X63s18+uCl6KbTh+Vr0YvVvlcNNhcS1abMF/02EsBeKMT07ZfdUWC+dBheJEl
iw58rzWN4m3uV/a72diWYCatfYsymrpUgi30zkKaZIXALx/do419OW6z/kEZ4vDIivIi1FImsTe8
apiWo7D7TwHmxYG+k0vmoEpHSGC/xWq4mpsRd0Q/gMP1Ca0FTPYUOk9niDbmeDdMDcGZ2EsY3HSr
87Br6/dfe53tC6E0RaduDMr7CJBdJTf3SD/n12nmixgFA15yZQikQye+KPxj0sUQ5bmWR7GfBrc+
d85gd1kFQ6ktTzlN9NVQ8Iwu3ivlMguIu2Bdto2kc5+2SuQnLrDBleQ1oVLzuV6Myjfhj8bdEsQl
uJ1vQZt4ZQC+KGBlijCU2vW45j8BXLqNkve+4yErgLkjM5Q8Qdre46FSpVUEaNWmIOkrfKW4qZfF
XjpLiDvvx555FNbLVvnT+YP8ere2yW32JUJtWKL1itErUlkzrFGLORs1pVTGEGWu8DsT0VXqXEqu
SKcQUYknAa+soz/ODyDTTBZjnvuMVWbBm/Eqmd+6DZfENmD0Eknz9oGV4Ph1W5BH/toKr3pZn4p8
bJd6sKCJ50oybQ6bCoUiW8xHJlPmtLb3UN9mo9SDjyEfRx08LpIqeRKgz6XFFjXJzqcdAC7CZVpv
3cfowiPKnf4DyQazFZWKS3k/9xLUBQxBj6+zj+pPrZlWg97K0k4USAeeEZkkP7h4MecnfLM6ZAJC
mKO1awI+J1+Odb3sy0q4QPIYdrGnKIZoX4XSGs7Fe5NmWxM/I5snc6iM39AnrQFx+syh350sHErx
wwS9TM1CR7XOsecUrr5gZMwKv6iVEFGW12uYV3IwCoQPUnrZZ2neJoL4aL3U50DLneLFMMoRQvSZ
p4rR1ZC38p0wGzrbtuaSW0U/iW3tuk2DxLc60JwF5upAfSKPZgoK0bm2sdU134CovmwPkceKQfCJ
Ck3b2qXluoWiCKe2fijHOKdJKlmnZzJMgsYTpMIyfsdzq2QvCKg8mu2kmMW5dutK6YNdR1uJj59o
7XPQPpfmn6KqDJCQddcrvVF1G60WR1OVt/6zhNwj6lsyp2BCeJwM2irgBi9V9sWrjAqXGK8sxA7X
04We3Ud1AN/cVlABpIxqE+rG2kwiiHTKZW4vkrKMtm3AuVaaPw6azAzkwn66mh0QwI1HC2mGuQ6F
noZImMKUNg+nJ9osNcdwzdDczxqvyQ2uBzD6d54HLDvmMgLN6YVA5uMzH8uLfJeYSfSce2VWUCRb
E7hc7t8njCw/FhAXK6M2A2trDQRmpbISfCiIWcpBK9Jr4ow1qX2HZgrkgkCUWn/tcLFSR1/N8HAs
BoBPNoUTubIlNod6tefSnaY3zvgQyOm7dqiKuDglPSy9UNNW9W0KydZa7AlDIad3v2GithHuJiQE
YsfzVE4AG6ZogNGPnFEHQClUv+TkKWEDuZTqsTRRFH0jJLd2VVD1yr0Dqke7HdeiBIRAnnLlFLny
V2yeX/luWPATFBb990y7HbeIyEOKrhrypUOInF3ww+Ij3h9wOnLanrMQIzK5tnJqmBEcrATpSHry
QcEnoEa26GLrq8TrFMHSu2FZqhPGXQ1noZFdNGk7s9/eD3cTSwkQNl97uUfYnTLlJIabYkFYxoFN
jj+Yt7r7D/nrPTAZCSex6Ax9xYkR1CJqFjtNEPlQPXZzCO6Io799uN1/o6+4GoaVezm2O3X09cvX
lCMqll2IjVrXTNE8ezTn57xkzMDjPT099NwoCKb70eFYHgpwnGecnALHuRhF2A/QNZeLzg/az5yB
5+UouJ+QeilrzCeO/8oMYWqV96oQGUo6dAWxwcm5aZ6IFi/JULw2xDkcLlKGX3pjX4W0gf6aRgKG
MizsFMDTrifzeXra6SC7z6NoAjC9cE/Oawz6BP1+orAzD0Z3J8QB2wN85xxpIv75JuqXao76r5WU
PcDDzbSRWPrPGYPcCVwnOY/01ge5kpOAT3Om+8IJqfHcVVog5dwJt7SVOH5PiKQkHWPifI6DoyBV
5cw5qvg8b3amzTFaYeS9SEo8uGOyKh7U7bWbORuBejE6bGVkKiYMWq49tHsyN/u4OVa24uC+FTwi
HQccWLllXYqe4wUA3guYCJC+wQQyZhEnhus4krJN1s6UgstgR6HmahTiJuoRISNMGm/ohZgQThzv
+/hwcxyVloI+REwooVuPH1ykm7ook2u7NVOKW2p6oLgFuICjjBnN7Q2FOldvfmLmxSJGJljkEXcb
gc35B6w3uzgKCt7BeNFpy88+Bdt83fH9G6z+Ny4ygTweXa/dtT5j4xUREtdiH7c7fwsNUCmkAkWq
/KkTWiR6sYoAZ7GDSLSn47iPqwQ+XmDgv0vpMN5NTCqK4XROm6n85j9pGDqnZVNSnhqRfgK6qTwL
VxOIW6ULse/BAh/SQ/Vf2+I3RXIg8h3LyPsRvy4AcMrJDpuMQwNj1J51iIG7gjHsTsWX1o3D2PS7
zMwnyqKy03kVyKrsGXW3t3zvT6ZhwMRhvi13vmHhmkHg1zDi6GZl/ao0MMazJMEJqvCijKfDewz8
NqIgsS3Y7gSJwePJOb+6SpoTXNVCAzgu6KICcLIZ3Yt6L2SevauzicyZynNn+/f4NG7NEznnarGc
Qqmk3EkAwrXmzJNvClRnffeaRyhZLWBvkoar/ZyoZ/lHDB8/Gy6I6xgCUCNVVi+Mac68DIW2XZZa
RHYK8CS20zvVx/UNicHLonVI5V7smTKqBiE3u2e+rAtNq6dOpjEnqtg0qO436jPQh9KKtixchNiz
KFCJPHOkOK4MHli38SlELQF9EmRGE5VR1LE27qzAjcD2HMmgpFCq9P/DGasMM3vJaXgoUXmV1nlX
fEv1MATw2xxGNw8sAH0DJJ55Ebq4CJEA+RA44QcZmkQiTBikIohlbqfPViOWaUTw+Gmz6GQv/60c
9pwKbCaYyiw32Ht2BjSxN2Aj9KhCtyxg0gqdOlK5/n8xOnN7/fsti5d0HBxjj7RM39d5pT/cbjQE
Gll4l2yyQ10z069FMdIZ3j7IAoVhMWjU4g+qrHp8lJoTY4KQfFAexPa711cT4zLpajWa2XEYNejR
er9MptqsrTvs5tzfeQQNAH8brwTH0fYMpDnCMJGkdm3nruUA2axUuzaK7u3+RZTCc5sGlRsn5+Tb
I5uGsIMkqDmiewWjtvMnmkOycBm1ROpdqq9Vyu5yB1XqW+QmwivxjxjwiZthgfxI+xC+MmTiIxU8
NNZka89w9Df/sigcxR0oRVaPcflPBtRXU6uKu8smgQobFNmIGfrqmQER2iUEvT9BbrnY7C2cGxEK
XK/zjPaPg1imr45uXKBLW5eSULD7U1KPVyhQHxeZJ8j+DPLBV2HvjwebSTduFO2GMF/sUfWdWi7r
WrCqFUzyU/fcsL1Ds4rpfrUW1i3+Zan6702STR5cWpbDW0A5rEZaNfstJMUH+DzTLZGr0iGiu7nY
9K4TBAxLPrUd2AFomkeGvBR/uh13mK3dr6NP5Ojv3AP5PtNnfgct7bOYuVQXlaGYsmoyP/sA2Hc5
Gg2GY+11/7ZjVT7MSvBTVo1PifIrbMMSt+5jrniUOu4J/RwGdabchea98qaEGlEze7hzdMPoe9P5
u5s4+BlyqynbRaT98eEK8mEwi8fT+EP8LOYAKXLZt8inDBlY9au4rTNq8ov6re7wWhI5Oc8I2n9C
bt5LeSUyRg9GDyznB2vCWsGbUUUbF6BEY7YPhtJWhshTAaimECHINHN6eiMaCNNbJge2rdle4ztB
jteZlfJlNub6lbrZbizto+ecQcamblNmfH3Df578xLnMSztVcLRTY90H8DjrIiafVZnJj2rEzbjv
9oE52BiGaS/EKCYe/fXHg1SC9RtlLOW8QBBDcDA+ruStJZFd30nBo9/0HjJa3oSeFZl0mYcTp4Tu
RDUskFgMmkXu89YpNFpGTQZkhCxX/jw0gEfn+Kt73vGeJlb06F252W0VWCzhMH8FnE/9TQD3hB1K
fmOR5n1GqMADWS3Yvb9bjc1w1iQB/Ah+VOBmQlU0U8csjF1t4QzWUqljp/4yZPpUx5C3o0LTQYk+
mGxPW1f2JZ9L0djzGtuHM0ANt83IXlzWKumHpNKdm8i8ZN1dNauO+7QsUuaxB/hI1npwo/B/NE+F
x3DkOAVzybUbVamgv/DjHVyH6OB0J8RGttIUGNS5wTCrdbeklE2nGNihFfDamEkx6m1xQrF4jl0M
m17ilYKvazOoe/rVaazycR0Yl88p65VRxgvdluGoHkoaV4VEntBnLWaQe40NuhEoLpF4ppIMSwjr
0gSLcHnIol9MqoXuBbZInbTmqboWoqJf8PwQyk/M4dGPqxtrs7YJYuV9EKImj1wwdfrrSGN0sxie
zBXBkSPpHITQX2igj/skdf3OlNfF3QnO7vD8+5JrIRuvzwc2awIT7U2jMK6L9usECqucBDyrOTNh
rpjKKS56y1VPi/mhB6d/ZIV/kQYGCEQCu8XcP82La49Ex2iQ8+xsQ1euMrtRdC4uPFAFUFbQGFId
evwnhvrjnPo1r3JrUg83ApmcM4xsxzul5CX+foOQKf4/YKHUIckQUxvGE5DeRiQObk0Q+6CpSvkN
oW57JvWwv2sQv7WoaHpcGQEqFhiy/vXZZ2KXocDRPoiD/FjltUJDYV0vMMnKUaKNpZtCT+9A3UKp
urr+/CTLjUauhOZmNaR90vby+tLD4qAKgnkuu1/3VekecBXNGbTFmv1N5O0TSm8yk2oY20Iibdsm
RHYDhpasojWKH66xodHVBxUiYYScvOg/ATDHDiqEZd0mfSpdai5j5pNYxE/AtUA/5x+KMFz/4+oy
AtNxQrwXGvwUdGxH2VFtKTt1Q8ihEo02Ur9HB+37A08tpQODguhzzdpijrp1CcgtVw7nos+EOzLu
SqipV0+Y35iAsFZ03UgBYHaOqq+ADvLZIftlDHD4cFOKjBkleVMb7/K7kScN1OYYs/2d61obZAnX
cX6Cv3Unu7BtyWcYBJMK3526C4g6F0GsPct8RKfAjp0XxUJlCPyqoi/qI03ELY/uEOGVZtAj1VCl
RztnmPIjavLp2PRTnLvXeGRvB3kTXH8qZDEEWCttlg9AvWJxSQgg3s8wTxT8l38X2CM2yuXm5HkA
cWJYN5cemnqzVaC7jcI6ad8HCeMEYHwnS8dM4Gib6RdSYSYpMMKPtDV7SeGRD9Z5pCd75suAtpEe
ABKP+pGRvN7Je0WxuphenXX1D06GcIVyjhNaErg5zMguWmXjj/Cj4g0uz7uhRFyyw+b3nkFbOo9F
JGGHPLoXjLJ/saMoI50vnXy4mGYYboeJvNZWTnJziusuS3Tjys5wj5Sdm/aiktAD9cz1PV7L8Tj2
7XXL2sbuno8WiupK392GY0WEnQ+NFV1T7sUaDvazLLjDgdLm19B0ZnPHJj06dKrub/K4qK1q/6q6
mAfi5ns0DQIVwFXzeXVVViETRrMJsk7f+OcdGJrBqRl6+rL+a0jbXZwCf/7/kwBlM4I0W9au2gJo
LjC4XlRU+4IuOvmHFk3AuSegW3inCmOLSiQX9JNDEJWH2/JFbXpJ75/aPNwkc2ubs3d8Z2aw/8If
oH5k7hTDXvvtuviGaMnNB2Brqv27Q2OE7QvmdMnrFfYVLLu0EjIlzAWtPiwtoxIpuvCEHumxqHQO
nNjC51MAKTo227PwmCPxDzJsX9VElWBNbAtZAQrR7qAjuvtOjr9S5CD5VNyQGkH5nqI4mQM48CoK
5+Rp6LmY+G8Cscz8UVITEv2butGxeHZC3OWGMJAssPxgYt+KJV2nDhtLX85SWrgwmiJ/SC8g2yDu
94vNi/YDzwF38Eytg1uNBlv0ojd83/M6SUCOePa4kGqbW6EXNZC5s/13jkSH3eSxSLmjMz4wZElz
ogiXuDFsmWde32N+u9LaMHGzFCMsBj7rNex4gYmFbIqE5k3YEX/Q5XbItZP3hm6Q/iUY/C5Cp1nv
h0OEz8hiUVmqKR3vpY0lamtlCmZ3BlGQVUz/oyaUZFwC37nx/hOjEW8LGhM9QHZqVjQ3U/ADTfee
szIfalKdmbC2r0XnPRRXs2XtKEoHpmJ16UXMTd3XIYJ47LIn6vIBX1K3y/H2PIA7wXCQXEHpZn5P
Kc1ZIXSlRBd9oLrcvJS9nZN6v0Y3U71IBJQk0p7igZj3jdmczNPKh4czB0FRAOVKm4aPO+p66DJ+
M/LMyVd4EmMHp+Ci1Gze1vnrG3r/dlqTGEmOySaxdGid7Nvp5wzcQwXtvGq6/uJ74ji3s/s3eXhH
wzXE/sxVKbNYIludTLysF1mO1l8bQ5qJCczbmlL7LrcpG62MTKSuPVzvqvNa1mRYLP9V0MXoHVL4
7a9RXYiCetpPWI4NugY3b0mH5XLvmf94k7hXDJleyPzeX9XSMVZzpxwvll5rOmfi/iOEpGTjTtgy
X+tGzHH7f76AqVpYHakaC4Fc7irUnIBfABm8ZdO96WsZ/QprKh9CZt0xkj8mYnwDIfj5gw/GcRZx
re8w9xP5iEAdrIQaypyDMpTTWMllR7IDAnjIsOMPIVDx1JlwCrO+Re1bdNnrIZFw8zTE/rNJhnfE
pDSRAJezpiUkpZZY+y3R+2j7qwwy6apT/2llIbqUeHwIoo6GA4WV/MdvxHL3CJf7lgZMV+bUZZ+l
wc4tEsRddY4YOnYx9tQw20EktYfE7u56zCx4hehPVS0ulpO16oXKZloY30kJttN2SSyrTyinI8gh
1aS6Zbif/7NmR4NG6olPx7h71/rFxBfb9FrTq7+uneoDdZuSE7z99zo8+cHemWlzN7dmry6ZyfqJ
e8jq8YI20vG3hQlJR5Bf7Fc3zrbQeQV4xDDQxn4jn/aByKHKxA+n5LuZWcB1LhULdomMV6lziSn4
lc6odlPRcoHuNH3DmjxVqr0FJXciLVLl5Hra1TJUkGRDOW+/tZqZQMTRN6jNVvnRSODq+0Yi/ArG
yWQE0f34DG59JPISOb5ZLBqSox8JyRu8lH4844UuBH/pi9B036KYHznDhF7Fj7KduiWbEdvqpmMB
fRVJ4KvU5rif14BqZA3HvVSvYANckLIX6kPG6fVRY94j6mIPzQp+fdZ1MnB9bxYlDhBH95tcKRBN
FSjsupoIK8pfOUWqADvZpCOPz0FrKZWZnMWjlkgTb9warEvCFt7t1jEz1L5A4AReKmbwCHzYGPjZ
fofW3Utq+7Wj8J1Y7wEkjL4Vq6K3bDkHBJX4lF/18sqgRIuC4RO3S1dFWHqRP9A+VAwl9m+bdlFW
RjHsa1erEGPvYKkZrmpk0MHgZIzY+5es2lq42Pb3AXcQGKzEFdO4cirSNcHXr8kE0bT9Gx6BDUqG
qMdkqVmeXO8jAjLcAId/9OxS8ND/lT5gZ1ViFBBKKg4BMjh6ol9MGtZuoo7VfCPWs3APdJXpL+A4
MLK6sPzS/OL1YGGjuOLFpGNFWgEExvbRNydze8dCloxxkGVDvIYRm3LeYSjg3xwNE1q2m0n0ud5l
ijMkohtJyOpEkIuTc0engrPf9UdFkiHzP0Zq8yl3AG6LQZjnAzfyWA2YjaqWx3HrQG9Hc1nQR3Tc
DAJ2UPlC/Q1CmJ+VVsCyyX+kWBZG7UFqjJ6a5ZfyR46WwN9wpEtD/pab4nYXdmtN9iWZl7i/TwuH
/TpjB7BKODgpWW8NiNfc2T4Y5B3f7ZJqLjaYBX4H0K18igtzqsdHoLnp8Ndpb5PruYw0ohW7tD0P
ohubQzp6gdOhQ3UWUqLsPTVoQeIJ8Tia4U3W1c4dua25bw5CHdlP3ZndbAB6N58oRdCZfdwNb582
A3Tq2amXkUGZiHqP2sy4kMC86SXRO0gsVniAw8XsRmWLQwra+Q6Tiagkj6NCRzjyCWlvuDjmNJPc
uzI6U08V3LC+Ouvg0Jk7yZrKaL5vecM3kqcKGu+yXuKPLOxYWKfPRZi0pCLw7gSbzec8SENIvutN
nEBYTKw+p0SAdXewfT0W3DW5+uxbZ0ObZviGOHXsVcn1hAsXvI6HFfGZR5Hs7SXy+OC3WAQ0Ku0D
JY9h2F0tXRK2WZ8f7ZmKINbohvDaF2b1fodGiQnl0xOhgUfv6kDjDXrVzOEBUs4K+6iWYQViQHGr
IYd1hzL13HCq7Eq54O1OQHVlijUdGTXD5l89fOJ1WcASxjCceXRNEjfecML9hBAr4LiW+8xdI8BY
ff/XwZpfihMkwviFG3bk5ss/pnsGLHeevzVoC8JSL3a5fwxdzjZtK3veDLNku1Ka0c2wtSzcS759
h0sms3GW+dFglrb9TfJaGLJ+AxEGdAUM9ck7LYcyzONKIpEUQHKzNa7FaR6IVPTHbwnxL/klLr9n
4SZPo/+M+lopxbx3WpBzbJ6uuGL2F4eDkgMOD+La68y9VhaAlGC2/hYQmTW+M18E12365jMB3gqF
uKSJhg4l9y9NvGrfoI+FREKfVqUdxoA/vywhYaYPntNYOTKPvrfGL9njf3pQXL+hIZg6G2cPvanZ
z2XCyhwZsydojUHvsGTOOcf8V6pQtqXccS8PAQAxXrpEGW+2Rh+ljtXApV4VuIy0NR+KhEd2Kd3b
HioMeB6DW5nH7pJYUDP8y9833df2tE1R59HuhmhhG8BarOAfwRJ8zPdV9FwNf8I0/rtyxmxSNhER
EhuBNCjoUHbjmhdFp94jTaLmvhj9pgNHP1P51eteDRgHUvOX0HEg+Lraqy0PdV42cv5w6oZr5GMF
sB4kYvQQnKpMXTu2ELjxsB/5As1hWvvs3q4zQBTgGGBfg+CvOWxr1a4/sIC+k7eg/Z3duVFzBFeW
HyOeZotW/vKmrEHu34O0AwncSS+gIWJ+ITTcJ5V2YkD7iGzkUEZSRm4bbtQM4YEGX9zrA4C9BU8c
YHdhT/dQJBVbyJhUnR2ZvPs8sMnVBWxJBS+UkIKTPS1g9tMEhPyBob1IRqxO8923GmD/v3E6G1Rq
IDyyzUS52uzBJSeRguBC+g1dmxumJ8YYGgYZ3Ng4v7FEbFhGCnfM15V4Q5zJx+KEHUrJM9Mlm61S
9/TFx6abRjHP6c+FHCssXb8A+6jgoGyQi6IEo/ZTGR2cM9Gl4WZZvWGLQwUC/U+cyadhfjggWYs3
VSzhuP9bykbtnnVtghHGaNiOausf/x0PB1mkfQ8xbkUkocGOOY0kNUJUzuGrG1ryiYQeAgzdv5T0
sRQE6/54NqHEYKJe06/f3MqTq/VG+3ZoCxiB3l6h/b0HSaiebEHYmGAXJBY+FFFeCsKnF7AhTihv
x11E7XifoppO60D3nOzFeGijpazx4lrL2TszqKXi4n9EqEZLGLLHIX8WdrPFn/PQiRJggA1sZ/Y4
EHca+wgI98INUCWLeXu33UwfmzIllASrXnYmpM1V/gLMmA96ziOjYS1JFBBm9EzAesbA4Aa/VKXg
k3ZYprEuG94UQVnMamSIc35tTKFzo7H+VBPZJefQFbN/8qF/UxMt6UiftpMNR7kTvG9l1V4jvWi5
iriD4iGBmOPzt0/4Gkzh2w6pVOhxgHHZSNMEx+lyzGjDCbqc/j/UV2hOEsAoo/q3hkTaZ8nydUPo
8r3vFqfUJZ3l3MCi6ai9uR5M/1RYXg+ycEbgvH/qdRRfaxyhLn6aOfc+3MUmOT+0MmnOkFvmfSHz
rMAbdXs0n05KkDv49udnmTFfiYDTNslHl2E6innJf3iyUgG2WJYELzknDgJQr4lQs524mvrLEOvz
eUmOoVaVOqoclPiVlvsKM8vflaPD732WctUubedqwv6qPEnzjl+YLzJLlrVpCXMtowP+I2STl50N
qGy3/n/DMckibSaevvjxqR+bT63LbhkhLDd4mV8B1fOoi/+4PqNTr0C1p2FDshH/75TQZ8E2GYW6
qYuC5v12DHmUy1DxKnFojUynxPXk83RLkh2012gruYpQqFAczQdQ26KpaPT5IQt+t6bIyX2UPo3T
AdeF7UjQPSpMz6ClSnLio5NVlncqK1oJZ7Gh2D56kn07LtcWx1ff+Xq1jYufnGw3s89MRL5kr4MC
DLIj0unaghgRaeepKNaTdFQXVkp0k3APsnyL3NJfTlr1m9RriQG3/PIFipTfWRgntxNwmyAF+Oz3
EI7Fdd2T1DVnVylbQrVNgHb0XeypRsWc085RTVHPCVVNB26lnwD0kgNW2vg+c47Q67bOnuZHdLac
LVGrFuP7JW77b9lBKNB/TnPuB4SeZrrcEVzcCeq3kJd52KvoC7pYoTbZjdnqP3FU4qvNMQCAecP8
F+cWxownFiGUQ3qOyVsQQdDAuCSnlKwp5ve+kAdfMvKTYysLnyxf/LcAbExd1gm6tvwOa49DMlVt
ieLTWxx/fwe15ZU1CQcE1MmBlP3pTel7QxISpOw2NyLJwS20iSLL7AShRl8+dVe1mL1Jw6Q/sF9N
0esDy9Dhy2vgevL3t7PchV8vRuBB67KN3FyUaEwPZHZRQtxAcbSnZCHCusLR5oZbzLRnSesO0siJ
ypwLn3pL60+CwLNgrZiSkPJ7QH4CLCDKE+oi1DEQfU2w8AcD9uLHh9ERQRNJY+O9I4cuU19X2NSG
ly92dQZQ0t5WoHd5D9yCqMOV139gyb5vaupWpBrCbnvbupfPLiiju748E91MkiAHSvpXnWDK/cE7
kEpCZU6H/Qu3oKCC0Ie9mctsQSLBxYctDZ3k9bt13HaALyPiuFpZQFykjWfMKh9z3euIz1mYZ9Fv
V7ePr0HCJ5eOFbMXwg1C7O9k1YwtPNmLip0fG6LGxsyqzL3o7dqtJcbKM/HJyALj1dAxcKEASkzW
GKAOaxdmS8TmY/nkkpPH+gin2oCscJjqu8GJdhWtj1XYUoxYFh85Lvv7UWw/zdvB7ooNH8fmF9/s
lyq0RWH9yjJnxEnwmqLLt3ScOlFgeVTg/eKSxaUqOFvPQcdUIJvwn1wSX3wRiavwrVXuRYAP91mo
nscwdVIg9l0HAfuSIcilG9RqLYfIOIYD4ShxbL+7oveLwKVu4uNF15ZljUII7KJm4BVVouTAEmL1
6uCBeB6GmFALYM21XRxCO0QZNT0KNPpCL98Q2MKDxd48Mz5qf6gszIhopVWZVp3hmPLXUR53p1pK
m/MG8IdMk60lLJEPLJla4TnPnOWempf702U9FXDzk4UsLkThqrl/PVl0cWPZoPuaiajOsRvY+nEf
xaH/El+rudbY02MrrC+f0LUbWaezlWdkAizoypo0Yezv42j2e4ND327bRs5uwY08y1gWTT1yH4LE
GN8MDJmhoI5jDvzZxurgOGpdr7mVbU5Zkn8QVJr2lliQ7Vfbh4cPzQm6uxp42OCJy38uSiasF+J5
jRjV9MhlDUxj7Uv1CgpciidTDQ4xa+ocU/XDkqDW2eiHTXkbWVe2RQ48Sh7GMLmbXWJRWNdiMoac
lg4K2AIQ7QsMaCTXBIPKhVFpI4hLXWhjkXc9OQZPaPffTJjLjowj4koN+DyXRnXuFd3+FEW1Hju0
ZBp2yfoyeNz4ef6kgvvLnngE89JapMyfm69CGgCCqOESjvTb2eG4BaZnN5mwVfsTruUaBVp0E5u9
c+1v6oXg1BPx88YE2WIkTDLoWoSSxutYv87rhRczfptYmhW6h8yVc/+2AClLGdMwcPgttPrHec/v
SSCl5xU3QufsNUmV6Ny9/pJAVk0I0WJFVLbeqy0XHakC7pQXQ4vKoX4BoZETNhRz6VrQqGKlmFGS
NXfc1WbV13d10mjdhIzuhEBXWmo2OYZVQylYLBBE09LhkbsvjihDx6p+7IaBMpq7Ug0+vDuvPSGi
mlxzw94tJhxBmobFGAvmGtbI51zaD9Z/SzZQlx6LdaYmNiiyUTcfoqP4J/fZ7MuOHLZ5vjBQNrME
/32A61FAdvObJ6CnDGhGYo643eM8mz1/j8T2/+fHe593ZdQWxSnujQ1ev9hHCw7NaXuAwYauQnK4
McJ2RG8gfVujqjLcZ9tV2T7mQvn1izMQU12l0JQU1lWv0gtnUQELGWnNAwfqoKJdxGdFIZfiTdNX
xTGSeRmN4LTu4QOFPh4WjGQwjIWHjv8Z+3ekuuGwWEw9TYtkSpiK4MzDQDF1MnQL5iMca0EriUU3
5yAa0A3y1MXKewEgkjzde7XXWVJI+0j8Yk8q1bnXtdrqhzOzfpcX2zV2hnxW6MIPE7131WxVbOrd
5bWdrXBvkyBr30pHwuV2F8nZzUouIz66rgBosI+DIz9XFWDD4H09fbpT+1AR6l/zbJh5svEUIhZO
Bd93mJJEeINWdEJkmezZaDv3Zf5p+dP1BYEy3s0ejkKvyDMzaWvlUsWDcgKSR2cBvAkAFwqf5P5a
PSieJifrDTzIbTgaIdhGQZJs7Tf7Ye+W02OviqWd1XyTOuHqGHCe1Htas2ragp519A5lYtoZ+YV/
qNAWlLaEDNkcD3rb5zQHFxqbvI751hvH4TIIkdPhDWJkFQAkcOHztXGaIT4RQWBCZc+viyOcY16T
AsuvWTU7+ycNY3PoQz+omfXHWRtkI2ZV5SXKvg2K/3LXzQhCNbAqT/YTZAxJvzH3gookSGGgR4hO
gDf/dYUzKi8EF5Q22TVGwnM+EvtTrz/IUzIpBhoLmzEq8th0xTHVRhkniqwkXfgILyuSwbqE/XnY
DUwKoRKzfsH21bVks5S9aI0Hi8wbG1MGMtw6qxF/DgErI5Bi3HYjGCETrn+KL7Plz9h8zYpWwj7i
PDy6ZTuTg7jlu/wzd891DqCztyJA36XghRWa90z8ForRwIAmkhxRP7zPN1NN8CV/lp9r7afs76A2
KzBORrXYNzfB0sLs6/5+oaOknIH5fjRoW1FMFEtOE5RqPBj+xZkiCJn9S/aaOK1X5f0Re1iC3KMK
8ULynMtMgWKy+i/gK8n8hxnC7tXBNqZ+Mnw80f+UaWh4xi+1XpUyT9weCSvxs4v5JHIlf3vpxG09
iDpA1BCnxUVlPERTxHCMy/M6BVfizOmP1eSgw+I216rxM83S4Ic9lGNl2obcx1k6NjeruHnIZBT6
BBzJoxEg2Gh/JMbGBVO23SSTuiO0sS9EEcXcolJXiyQ2EI1JUDv++i02aVzZdwQk9JiQYIEUQw7w
P/CPfakn/MH/wCqGQFFQAyO+m0vznZ8+sGVtk3MBxFE8CeiobbeG7QDpd/Xb4k0yTDyMpIIg/PA0
FXAk4y/oQSb+UppnwSXRGJH39aWkLqh9yZTDeiDmLoTBZwYnSJ5NmTTWUHM0ueAIeRBYUUmvAiLQ
MSx3BT8H7opem/hsAyBCLufG6M5n84cttZaYu1ePS+4wcwAFgd8r3OnqvenOFT25VkEsDag8cQUx
kt6jhjxQfTy4khey9YVTrhWe5Vw2AS4mUaGA04W+99O0UxJCMRpaQrplVkdutgGP3/kjd7C3G29/
HBWQDsc3vfItnN5+72h3ln66/w3PbRlKGu/cya1L4dOLNbO2pc2LQXgFDPC0EznFYkvoKGxrbFBO
QEUegNeEiW9jOfCgjlCJG63RsTrP6LLBdr1whW7Ao09lGWX2iEjWShEARoXJ7soiz4+Std9DjsDD
/rfp9mQwoYvrdkN8g5c5qtLvYiR/6LH9HV8GtCMdjdYrKqhX3IpcwadQslKYMWeeL0MIdz/3HmZr
f2BUySOdqgOknz5ar+N0Ng34zEPeNnSA4TWKEmlaeWJxQUuCCaiP+pVsQCy0S+ZFuTZoWmGlAgbg
7IGkvtjqasc8koJPLsoSguaIeth/8ru5Oq3jrILrQx9EpijUgSR0l0al1YKaMDFW0xtjo3nMetXo
J3gQtcX2lDrAjKRk2ZwfV0uwozTtxWRbKNpl+9Z93HFFEjkgGwuwRpJwdJAQzi/DUz0361E0X3uI
rFFdrgeb01b02Mo2ymnm+PAIwH2oieSjZYwTkAvfQntv9mW3VPv/xlLI5Chv2AtJbBofhA3uQ6CX
zaXTrskpmqhUaAGZ1s/duhom4FY21HM6GNFrGmg4mWFyUk80LrSlf9WSk8JQfwUPGjWhtOmY/9+P
W2wqz1U9VK/+cBRXaxddUfLTipXxb8XMCo9aQtwP6j+oo0bxqnfUm9Y33jIaQ0nbe6+hic2xtbg8
6k2RNPZz7nLTHrwb246CcN11W9o8QJenCH6Xou+flQHzgBpCNgtjsBUNh0LL4wbcug33xjSOlcHg
GvQHrB6royDeY0mxQpNBoXtRuEuScuAQTcjs1wkn56S7OtyhCm8LrbD1OqEOIEiIkUNJipylSZoK
5z3qCxBRWWE1p3n1snZUCeXoXxV9X0pxNsyFlW/SYAXY50ElZlBS5w92mGc/ekf3CcSEtZSxBj7a
Jg9pcIgRMaLnDG3+w/6vTySmijXih2BU22yEYOKIH8nawzrDTdjYxJk8dnUsbr2u5yi+V1mElweW
oxcwqjrLXjQmTaNELw0pTDz3d08ZXmWVQ3KsHUf6gk8f67Hvqs2ndfs0zuVZeJZHIxGyK70e/8xu
eAMemAI7Kyf9nmGkjjD1cN81ft1H9XTyEA8qI+jkUeUuCyzH0RjECKhP5CXt8ezPfemreIey3xcR
y7h+tJwewh01Hj+wa44rfU0eBFhIHaU9j+LFFSfCKTNj+pW4kU7HN0Qgt8d9cVAM17VGIySsPzpU
Z4MHAJpl6YwKHYECCDgWCf/PfuqxuFI9LRWdEtgsrv44Vg1qYWdu+LMnBJHbMCOXyGBEEwNP92O+
BBIENRzhoqRwkURRu9kDXHFZWHL1yXNPjzDmOf1deJualn/tnX1Uh8GMkwAEbTAW5TX796CUWPnZ
fEsPJG4Ai48e8xZsbKjSFW56YMJu7RZ0NYm6IMj4jHP9U4PYWgUD9bIc+0LbXWGs0uA4BsvxyhNt
zkowWVjT3iZ79SpKj1ye7tWMIgGsjzHj2b8AZYGkgYFBqjrISZkjS0ePbPgDPg/mKTnoZNYduRen
oF2kMcB0OVPkb+3O4NurUFeyMrqYIniuee7oHrYfqZRfVWZZaN4jud3u8U9aBqdfcNC5wTeVvlOb
V3bruw3iDwipamtyOflQ9ojnysAQDiUF79IoZxwpgqPQuAK6tlwt2/+5Tn5ee69rbH470TWWHLPt
kG+TYVGX5azjbbSGJBZcjIfJlEXKAniclY+8IKN+4c73UQpDu8f7WwDTaJ/J+U8+J85DPlOHbC45
ZlVEcgUF/5mxuTOju4DyUe/YAYkrUtbNgMnSfeBMMuRYn/KzoinpEzEVy6jX4UcZNw/eSWSldMt+
FeO827HBQOne03+Pi45aKJS5DhVfN0d4IwGWjav1BPcCr64vTHsicPGYzYIneZ0Ti1e061CIeRPl
oKb+F5S7nRQCvsAq9brBhI3K6w3UF64pWE1PnNRNbJ40tTni//JSI3ntUIINlVnQljF75APKXsiG
+iW1UhCiy2FcImDRrUXjuwPhHgDjNbdZrb9+NPkImx+3OWIMiXPK5bFzlNKmxObVBqiSM5vdI7A4
0sMrqs37X6I+VmJuSjubeqgh5vu18WQ8er2nuHbykP0Aw4qG1GefYRskbMvXpIhmbmYUHI5YMQF5
cB9PvwpWSfo0pdRstadyUkRf10bUSJ/PPU45q8sjFulEDsf8WRRH6Ac/V+hctP0CjintOIJi0E4B
hvhUI6LvhOxfsDw7ZcKc9dwFyatK6rdyKtqpM+SGHUde04QuTTuuD7ktzy8Y4FSDyyIsDS+Q6Mpc
e3bCtDKzcjhvD6pQl6vk5+GObbXeEubLAW97NfzGC9u7xyq5tm+iWJe0Bw7uyNGpWVh95z7eFy2/
mty+TliDXg3hNTX4aZsAxJSBZsEA/uRDm+JqF8hgELP2DAl68O+NqW4E5Hd4m7/qpIGlXQakCLZL
GuBSr0rNL8js8lHIKDfgebHhCxPOaaLZrMTb1iwGzq7URrUDE6QpfeGdHVYQ99vTt9+ahsWcbuuG
aduhfnMjVMMid2C8chLulaVkSBjI2BRXCcvhdtZqKD1k1KU9rufeLoDmhmcPOGghMOIlbx6uHlCG
ibLajJ/zsaXcsoOchADe1XSE+E9DIuj1JzpfgVIowRalKn4KGQbQMDmsgKNaKRcpHf8NlzM7HeUg
M0mVnP/D9r06VVOUt2er0c9rYHuklxxXJkgFsRVRipg88Nd8tQjZ1cO95bhmEPdFy3tfSYgApVUt
Gva7buDHazkONXjGrSrS6pDdJdmb2c0ZtdQWhUpokFtvJL7zKHQ4hzNOLJ/htLFi+lSVdn2ciRxv
pSjMQ6bEKZPxHQ/Lo9ktpwU9C+z9C+zRFpic0OVf9ZXAqd/NY678ynGYASEIc0gHQmViYfs07XRe
tULhgoGs1r2RClqeJfTKzOVqqYw5DUUweOJwVPLMYntLoq3/DXajgxhTJnBH3M/KsFFGaO6QbZOa
uiqZqcylhVen7go4J4ApxHgR4us97SUI4KTG5euVmlDc5bvK5YDTamuSAk+R/R/cYAcRiKGKugch
GkYDKTLbnkSIUk3jj+6zUmDb6KgoB3SfkuuiaSi32fEDyoD+iRHRzWBjpcep9MKuGFb0Ez2CYw23
kr7spZQ3Dh4WAK6A0xMn3FAC5dp67GGUw0Y04XOOjvgx/G//aHX4i+9/knAa94hRW1miRY5Pff8p
kDMJi4lC4PT2RBF52GZfarabi4tn4GyyhfSpOm/3xUwIUgRdxCcX5fn3CaFzximIcsSuy361boij
vCgHoYMpRW26PhRAAoJIM7EZVVp+yhIlyLVABXn1Q9n7hQR91DfY4oz6m8xA0D/XXVtAcwVsZFZk
pgD1yc0XQGC/J/f2vNqpLdC8TfIenovRLJOaKCaFYcgwPCttQegp27GRWtkPxVjlJ4F5mSGVgFvC
5LgfFBrPSMGMuG886znNKdzeKc2EAInJUZM7N/JQIIYSxAiNLiH2AlUAlt85l3tIU9H3F4io5t6S
4Y2+7g9w1fFC4wctk1GbCW5Ey9PdYbFqapAfrglRxTxOZzk7N0AlVgVnGdKnXVhGZ2kU4j6Qr9rS
MA+Vd/ThZF7btNQ0mUVpGzPr2o6gyms0YgJvGmFR9458A61pHMCSuQmKhP9XHw+lPQ6q8hfm7c9m
eVgv8hQKm1Z6G8j0VfUQo7q3TfW7ibAkVdjw5K0Mx3AEH34P+078mF3fNGQorTRNbb/Q/6MCa8ix
ZkTELzR/vv/vd5RUQXmCjiScF04R3chcBR9QJnWlwdSAOjQcEjxABzdFo/bqihOcxeKGjvz3MCCV
ZmRigGb3f2j2chZ3pHoSfmjPUsCRasPM5RrWio3xFDFrXvE4GMSfEp95jmIIF8o2iW1abNYY9LFn
JKDoUO8Y0/ovbdk2s77tVOCPic5CwccOqBeVjoaafAnmFbSD9sEuaAQg35MdBmjcaXVUjk9isFAm
hn6G8fhE4FB32iKVXztBWZ04kdG2hNldmPQtAxMItfakMHYUSmhSt1lBfEOAz9EPkj2KrFWPyXo9
it3WhuRD5ErwlRRJ06fDBYzOopktV9X/V1xtOLnyyyly8tdb+adQ0k5qWSjDEKsQj4Clw+e0pR15
DDhbvY4956Ui6gFMR+3asYgu9GQzSMF3LCawrLQerWmBk7LKX3JUKgeM73O+0F4abYYhoH8rJ360
IPLX8yQQbdAaIgOmXZggswYFijHBPJCK0ShAIccJBjAjWlvX7NEhPiwM5Zr7YcJmPpeZ11mZNyks
Fd3eA4WSQp9EvSfwqwak2exype2gcbtJnQRTN+cEvGioV+OjEaXnoQMfCRyXZ5INrlNTZqBBiHR6
LqjWvY6+mJtH0ISnz5ebl94Py4ZadClz/Plgl5wu70/IjXARQdZhoYyhZnVQImi+npdUPpS3ewbC
ZD9e5CCi6xnUeHnQSm+CVObTxjW84hzyeKY+uBOtIvYY0jZ0dyP+mxgVMxQf3U8e3kLOJNgW0+za
8XE0ZoMlGvS+sJWIwbBi1/GCACR12nKIG1z83pHHzJXHH/NNrwG09H/iP1s4L4uqMJAUHAFEy6MP
bB8tFKrsQ6sDcYwLOCcpFs/AYpA65quWeHeHDZIzQ5N4xclJ09IpRetLBE825KW4WsdMUNZnmvZ4
jFiTJgLtXowMorsSrShxZKNyqqlLe8Y/I7I6G7DCSYQZUZYMdSWegQvmMttM8mlyc8NbkloxBifw
ivmf//iArt8hV9segoKx82+B0TwpdsZl2f5R1VATK41hTMa4BYwjCHKaYDB89eQ0cKiIZyziKalC
SNYYlly4lEk+7nqOitIzm/YcY8/dI3D3DDw0flQnQSJduP18IlJOCjDaQSx+Cb8yhIRjRRxYZlU5
JC/80BJc3nZDWGaaqw3K8O4pll/PWEXucwp7jelJVubHvofaSQN9lzuL3dI6ICxJGnmQwX1UoSBp
ipueimWsyfMtKk+TSbolUmlMOEIT3yYX8xw4/BCUaY3ZjLbFZgm3Aeo51T7aGsc+nlmj1K9gWQGr
E+6MiNzWVedJcOk+yaSvE8GRO9EUCzy0ALX8oEgOctXZcUjknPJRhkd5kltuiWexc+LQOlirOxt8
tbPW5ydU2jCFZmR/Q59Bo8o/aWfnbKkwW4cDayAB/43dYYWShcpywl8MnOSnq5Qvc4I2e1YTQsDX
YKd65cXxJN1Nu0NPPxhbPwY9++Ax3/fkqx36/lFRcNFTNguDegVzgRsvPFULHHRCW3sEHWGMBVMC
FFNKHS5lkuG0sDFre2MzrXmyTXhMSsn6g5MfwZ9qKkSMXjMuEir3FrLgcD7fjF3WbHdB/UpH97Xc
sJOQceM+GTIrvnr9Vcfr63pSvZAbrIJd8ahxcTiXYo8reNl+yBteKat5/GCic/ynjDJj2B0pOqCU
9RYzn31yMT42jzTr+PG2lzJyKsc1FL8f11dMYKmQ/ULKrS48WI9Iczw9PNEzaYvY6c2/NiA4HZ4E
8pbe7mCDkJf89yHzTTs2nnwD1t7pDvDPGYyT6+g+ZVhXyBSamxC6yilBtumFkJ9jQr02wuPT3W7q
j0CDkUC8lDVjvmD5gXOzLSyK+KkZtVshLNo2K8dXapyOS0nBMix3JlL+u5pzx99NZJ97HaHjYqNt
UUENDpVeZJYXQXnaC3lQ+yS9Ob4hqCBG+qaOWR7xxY6CNxWTFv0fN+CQngRGD56UQMLVMIE+jkBQ
OMXxwbISYNvKfGitsb9BlBf0ypFG1/j8TgPF64oPR3nVpMl53giiR6Bx1qbXon1nQfHGUzLFP4ux
DrblJSc5HWofejAGj/7eEtdCFb9//VJffew22DtSWTGD4XsqCyyE4eVQ4bgDXgqqmCjMv7yf1ooQ
045ZrIf0nbtinIyJocvtIN4qbdSA4tEYXLloXeP7e0YCsuV4ncrj69HuzqPtHocMpRZmpY7Gb9Gx
2TnJi5N0LHTFj2FINROfgz13IL8/BAWAdC4ZxjnTBsyfiKyPdQLF+BdcYVIZWNuNekLYvbqxm2Iu
aOrfi72DHCIcfqN0eScEKSDMIT68dZZvUSrAkIHt0Y0grxVBVtrglIXGM048rWtxYCNPFGwOVX42
ScIAxHKi+LORleO8dTGcRpB8q40bcVEA6+Q4Ws6BTtTrLcHltQISP/+W6QhgOFeWoUENeaJIpoYN
m6AA915a9mdF/kgpk25vapbFR6TB8+hcIIgt+CjnFMSyIQ7yJ9K3oyTGgnBl8P5ZsGe1gSYD/PVn
0zr65yzNAiqXYKrkSHJLDim6m2skhdvLjG6ijuSMNrhuAZe62KVQp0IfWm1TDSWVfm92zjo1jLaZ
IxWcWiB3nIoc6UX9uYTn7Ywgj33nm7blouSjRgpL6+MXSVshfd6uen3YxcycAVnwC6qQ8iwt390L
4rdrCmIDbbPIy6G/vnOnVyeY3GBuwlf42pfk4+qnTy0PgWcG47I+nvN8MIIt1wgpEzbZmCct60uR
dvpk43vJJuqEZYeopdX/99mxBbIQ0UA7dXa5nNG2Dx+KCwvQ1CQ8NaCcSyKeGk2/3h4FRSbkkpok
2YLPJkvM4JpY+gABoMFUkOoLNwSJw5wkINzGcaaEGAYDApoxFyqLnvGv7squYT4BNw2RbYxOVLcF
EiF7tGGKj63heD1BFHRbBkujxDZbtcy/KZjRoX1dJFWvwpf2DGXR6RY2KBh5xyJOFqcGCEmeUc+v
nFuEOWlkKxLhn0ppulHPfgOpoDhhnWZ5F1fMlt+BKegS1Xjjbhm6ScP4p+8VFuEtLXc8ZmBlV+7V
A4Vc8wjTPYxvFQaUIAr1BoUXe4aBLJcCLbCc3UCpd3q8ME3HqnEXd3jxvTOd18oPNW4tL8f9eSds
zd+23/Za6PB+oDz5DlnCnR28VTgGJvIh/Ydht+v85ZqbwZM1lfXidFJFhb3NU7wFKQajlLsxLwS1
1lBBhfsFLqkfRzMBxhp7H87bx3Q+nLraIupA1uUb/sgUN9CbRLE+XpMKn6OHVOvmejieG88nUVlv
0Ig+8J05CkSuTEM6R3eMPQYCxsNkW85CsiYRTtME06PB80hTPNueLJ0/lwF4avLqcnsDRgQKgX34
EFrGhHx4Q+zumxbfxatWTufWNxYfR5Mt3J/2wx3Wm/871RDpGGaTNm1reuB7TEEDCccibb2B7vtJ
aoJVKbK34/JrzmnQoKVp9+HnXOBlXjM5sJRa3SBeKSMxGIM33FujXKH935g/R6CrwZt631t/aoPW
+pbbw14fVHyhiynp9z77K09xt/tfGms1pDqOtfbuFL/U35PoqDdY+9ouxsv1GfH8yokSG64i0+uM
ozaMwQSsBaYIc+ALKT1SmJ/Nw0sWQGAm/ST9JYlieiF1we8jsleRS3acEDc6zLvOyzMQB+9zrFV/
3UdXBdrJ+sXkv1Ejr4wuf9RGQVHciGPEGzbDb4YR7ST3zS6atHLiHKD6tyq/9/jSbqWQc3HZy/al
d7AhARKSWp+PT1a8qatBHuGLZ1dtKPdxbBFyr1i7IaR6jlZCRQOGR0Q4eXW/fbUbQsLpMQPCgonk
3HJYceoYUyuIaA+BAOnEW7XIdHSTKWiTQR83sMCTBEVDrE4mA0nMQbemmIogtGjd4O9LgsnI9vmJ
Zrh8KobW3NGNGygCuEwShyNVGxdEt+c2kxPuWyItIN/KNezobJNK4U6KeK5NXhnLzjiueongTXaw
aKW55NFdOI/or/MsruS4/wcMEDhp5hu3XQETsA4ZryFAwK1RQ6c+CDjwLyFTXlVAk/56QWeuQXnd
LjSs4Nbx3W7ogSviqIF7Y1VFB+Z1RvMZi/zC94GHODuIdyphBncvZYJc7Q51aycCdI7/kn++wjIb
3jg23vOWedqm4RgbNWkRWwz3d927jxa+FSynBFAr+BoC++E3ksUc2gcyl9lGvUf5Ye2TKq0FJCM5
kDkMEk5Qs59Nfg2I9eNRAl5u3bJ4CVWg9OahGl7Zv67iwvPQANmlalHW4r8Oe9qYof9oXNv4uqWK
BcX9RTaWbk/3dWqhBsVVNb2xx1/qFf6jnJAH/1BKT06q0TfLTwVFlpjVDAT7/IOLsdrOLO+vB6bv
ydBs2K1KDmdDdDTNIPuUCVB1fGSwP+m7YivqX7E9O3VKxeepHZK9ejFvnFA+Fxjq228XBYe5Mfuo
XIuR1M1TOe/g4T3c4LB1fYqIRHLcA2R+TB80W20oviNCSrx3METfUU4m+0kDrbdrLOs29zoy+KbR
FyuQjECVsIVywll5hCQI4ePTwzRh64O3nSDSCxRT9EHeEij3YiSAtLlZeprLfuIA4dpYceb5pBj4
apyOLXkqUHrtkGMuwLB/YK20SA2lKCOdfPVGboZ486zEVTMiHd1Iive51fPdwkpIIFHtcF6HG2mm
gBUaTqT/rEtSjAg5g8eG7sp4krqEaQsbh6QeJHpzJTOOBI0wxw89DRChtixeSrRkKVwfyBEB8Iso
7S4jvtlBQfKWunVo86vJjCF93jQkf+sLz2UEWk1gHn5XVvJ7IDfrySgAQrLJIwuKPSUN7YYMnd6t
nHND0s2w8MUoacIbb+t8YTNDUEKvBiJDdJwYGnq57+O08z6llfK529LNK7AOfdFenIdClBTv7BbR
/JAiYbtWHBobmWddR+7FRaWtWxbtLhu4gXmyI4UMXNyDsGOzeFameOUtGzHW19WylqryWhpQZJiT
JMuRVhlDO6zFlptZGQVGluvHexjdJmFK2kw2lUeD+vxSWMqH49ydiIaWW1kCj3khfUxEzpprF57R
emRVD8npSzt4kfEVya3d4TOEuYcgpuct8vRCqZNGxZ7F9Wqa6a49ySrrywbsa1wzUnGsoZ1bExfG
sGKS5yK9qzY8l8D670KcQi9c/50VpX4xApOmp49Uv7ePjNwWeDpGloy2SnpBe+maQqifFBTEU/rE
/fORHE/Mxys8j4gCHNDoFfBca2JtNfhhr9JNIm4Fhltm+mdxLIwaKyZCdUj3R5jClm8fQkTzrDjO
CpFRGF54Vx8Y2tXVXeyGsE78A4u2x197eG4s/herze70lEVr5w7WTwlOkC1+5c9IW3zTBzwRthwB
jlULlCEr7CiPn7QINYXXshmrt4KZFlbAkT1nwpmg+RXEEQMjPRqGea6RyQKnbGSorDliurazcs4b
HIOUeKHSsZROsF55qDOIDldvgqez2jnMheVsQEHdZd3Myo6cKrPkzGdeyQ8zlWxLAfPpI84Fn2cB
CKU0O6j++iiWNzSuaf35UMGJEc645Im/kFZ/iLrOA27MFUmZkRUp2fR4e7bHx6cyipWTPw+2FUrG
UXp1wZccYfZv5cC2VI+Cg5AgQOXtwEA0yfq6+khjnyld9/vH8JMbDJWZD0Q4kGPhA6tgsh3+7+df
biOXc9pGAyGTbrh42H03xTfsiLBcjKxBbyI/AyYKgqxjOgDY3trYFTIKPR2czDu4ers5yc+dhm0X
7G+g3miSpkMD5UiaNE9TbNyxtQ/f+ixRK+sUDXfSY3RLfUkzV5iSY+xzORqTYEuGgucwlY93Xx6T
FRtEvz3mGkcaKG8Os93Fs4QWnhRDCGIiNXrO9d4Db8pbwOnwU17J2/5wqzEsMxQbME8SWX+1QJUs
/kT7bp3hQkud6FdAJBfNtGgiJ07oUAHMjMvO+mnxH6EAbzwkQGoFNnd9rHFFQv8wIx1MUUkSkswP
uq5cwxS7sl09/h6WhCqxQ+PAYMntzkR5B8z1nZ3uRDoqKwH5VI6Jytrja2nE2gTCZpzAdiywapvF
Uuvq1ZsZ6Tgh2MnpYOTXSZg/mS0Pd3HcsLNIM4BeAKCaI9gu33zNqY7KrFTXx3Vmcweyp0a0emRF
MUmkWKifRB86XJRQgTuEJvmbrO53iaKxYJ9z8AIlMoXcLowXY3RxGOHx5iawcUJTWoLTnFQLDH1y
ylfyEF7Tu30Y0EEuyfvdHSUz76WtiBJBZiklC9RmetFAG0l5Bx5LaYtMQOSEK8aYoIXOFTzxsKP1
9Nr6KIlce0SkBnW0Y1JfXp1fGpIOS0KwD7nD4OwBXkuwLElKoe/830JqyScTGx776+FZJp+G5oUG
c174hhVSFNPUa+1vhgV4oBCVl8JyPnS/9CiTpfe9qp0xwSnc0mvImezND86WDmV7cl4amDzx7sZK
QCeMVkD1ktcV69NonhvP3R0uQ77WGgnLKfLu1xwD5aDvgBrHKILs2j5JbWxyeR3CY0PYl/JVfvPF
Xklc9cGHjt4nsy3nBfyzxJq6Ra4fW6ink/78EJp3AwStFLsHqw+hrdsLXYsfHfScqmYCRG8LAB67
Ilmv8F/5IihrLYM7BsBPyBjS76TFsgR9E3G6GH1s60htLZRPPPtnxVaDNNNnPYDmtgf0n/9f1Tp2
4TfFmjvHaooTYUiv4PhS8OZeH/PnjlphZYZ167D64nbum1Gmb+KA2p/iqvzpzjxaUnxHHKUp3p7Q
/iOajiFQ4/kYPusy/DylNymHcsoaJp1M5Cnp/D26vyqIdXatsaeg2BnBFupnNVG4PeWHl1G3EuCU
yNP1iZjvtMKGbPe9KFWbnnFmPmtJR+iuMHmmw4n/0mxQfy0rGGEEqUUPrIrjgqck9IzbQyOnAeaN
LnSUUnT8zv4mAcoIQZlKD8u8+X37YsBC9SLbVC+N/M99ezV0oCxFdAJECTqI0TvU8ykqf3CxPTlQ
Ytn7JPHAA1zn902B5CDNeOy13aeCAC+ysIwN8nLxvgndwmLPtPpFG2iNx6uLhTWqIdWBlLbwIlrp
5Abz2cOBHzqJNft7l1eUIaM5s9qU8Y3GYioBRaYTZ+B8pVUVvcv7LMWLtwocxRceJ7HJhSX3Jc0+
2a8gsvMcvXWjTPuiQ1R7WMhJ5dJYocneY7CCC/ojLHxHv+Z/njBVtS/QwGvSuYIVdRu+rPMtOotF
NnPmpgSqr2zbf+K7UUxs2++ucQRgH8Z62lhCzCb22Xl7H7SB/Z8gNJv5pQrN3c0QNSzgV1h4ZiqF
bZUrASAFkNQthWumT257phDU/b5cYDHknmLt8Nm8NAQIuY9v4ny4Dg/zt8dGsikPIdbPqmPlSZVg
UxGcPRkomHkqv4/yQY9Nuak1ETJIvbniptl6o/Ufgj/nM1Bi99A2DDsMEIPYwqSgzQPfGrTifOm6
wqndrArwiHbp21ry4L/Bu3eElt2qTFPQFGxLowkm32kRNPV2EDejsobGQg9IzX/CvD01lt78oXWE
ID5RnTxV9DV0n4IzG947TSD3wCNVHcchTdCPRlfDihCi4QwqVMVZ4970G8+9UbrGsrFxc/3ka4vI
Bk0lSX/l0gCCFsA62S8xo3CHI+jW/zeJsU+dZwqd9GHhi/ZYRQPRvBmnV74KSVZUcoRLw6EbupsZ
b0RZwJdueDUIp28+xUdVwnekRXKZAmSCk5ZlhzkmEq7Ft5zZ3KG+12k/j5Q9ntMnfkJnCmgfGg/B
EqC1ObH6Xi22tjo9LrkewSNim2G4sncfoA8No9zxG+mfOHw5n5hSDudDJKqBMmJpttdoBtauh0QF
GBWVbfvLEBnx1xDDCukJxxiaCxncFid8oUmGkwGxYavvbcmt3DxeG7F2Gnm26Sl+LmYbONUGrzOx
qWkKrSC9bY62Rz6SQMQ6hEvxYjU+UdGXY2cH69FvtlMkVNvKUW/pdlf9U8SDcP64z7hPptPnndwJ
ymEYBRN8wqoB60p5/mPGehpwwwwNZ4BarG5aOh5AowPn/51B0VPVj3Vvfrc4Aw8A0EMD7Zeeh0A2
PRvBrdFBE0tHrS9H93DGjB+eLHxgS9JMQxeO8q93gpt9A44Ncsw0Me3yk75U0cEOPNWlKVqxL0OE
xwhZ3GkemZkTyndUQiGMYeiy0z+A0lw/mVH62wSXdfAfFiwc7HhmE+2lqNPGqrgEljODHZDIb0Vq
iiXCRwRfyhHHH9f2pPeffaCtuYSp8v62NJWER920UY0l9LhAR3xIFle/iEWJR7UcuNHdWJyI2UgM
MLqSkSUr8SMiHYwP4Q820s37RHUSfGOqzED9EoeRTUQdYQNyUKa95yutwz1Ow+gI3sTQr5Hs6cX+
s3NLyDRmFJ9SYAhiqJd2CmufSWqZeHAaTB07WTVtaoN/sm/xDxoErCtwoVU8LppDGuLggdX3CpI/
a8k4HyUDNHLf6PUzfl7tPG9HR3+EA82whRT+WTBuiRcokiDiGxL3wMQLG7q0QIXmwH/6iDRqzX7H
6j9W5oeJjTtNK47k8a3Nb0VVoWXiPf0zC/VP4PGs0q1Or/dgwlkxBWqFfvvF70Ekjy9NRMNkNLcb
4IhqKMB0WCdcGuUPxXfG04YoLo4zO77MPicgp8asCa1O9n8Ybvp60htioa9I1MzJxzALX+FGMD3w
tutq0n5JeAiUXpQpcWayNzrE4k4DMiE+W/Uo72uSNUF/u5rX1oxMNAoEFqOLp/lhjUblR1C5uN2n
OJjUGXgut146EXDDEWVIBdXjkmNln3ygsOhQ+VJMe5DZ1rcE5ZBmpN8D23ufeGo7EM2Lu2slnt70
76aEu7TYw69HksOwDo/FdSrh4OnIi+jp94+M2/1LePFhcto7Age1wP51NhrYT081ulG4GYFeynm8
fT2lOutHTkfkzt5/4MxWMPB5rzJrhbaZdN8EKZw7juh1uDCjBEK5+p9S19bkjseUxK3l7WghfzbY
pfJr0vNPApclR076m52/vpq48zRQakDaPP8rDUAs28M3y73SEPibVRk41wpDjJjeq3ZT40ZxaOPa
TKIXGU4riFIaRq502HdKiU56AXY4zyn+8ivz08CLExemLMlzlZWjLYtQGi9U/2dqaxKwHuWUdw3d
wvOlURi1ThXkS2yCa+S8BZF9EcqVAoMFYoGBXpKi0uzitdCBOaltGP2IDpFx7m1U+QDUEvrYl1Ra
57XZunTPdqGqCVnyROUc4k9wPaU6XRITjXUz38l2rNdY0xZrdd9vwXzGPaUDczo8vGlC+Ne9vKa3
a9KPXlhzUbX+fdFm/s+F9hiHZaXGNM/RvzeRJlx1DHesZJs4PWly6+hpKJyTFwe6RBckUY4SK4cJ
/EsyFj9JWFHGnHT+IrShjz3coXWJpOehjw4sN6F1L8QvdyqCZB+tnmCrtyKC9Ku53NO5kCsTOyxr
sdyuodgK4tYczkhyan49M53oORM9eR4qaDJpMez0DDrPG5FEOcMjMQW65HlJTUtEGZgAqlEyzcYO
s6kYkRFqdUxvwwsjAHfnym/poGpbUmlhztDuXsLKiaiEcHJ9NSUn2z0B/c+CcL9HiX8t1CNHculu
QKSocbvw2H0s5ESwKgJEZ9fQTzNHuu02GiS6RpsJ9F1T3xxAMhU7SrIovV0IbKYi6XOVvN3FZUJr
T+aCJqGvDhP+YC2oHVKlZFjTOyU/k4hgXeRm0rurDv5t/yW2XHKsoDjrgH7uz6ZTTWFkBDYyPl4v
yDwy6/n2WzUe+dMi2XDndwtcuklGjNfX+mD4bgAX6VbItpE+A+K38MJIeNKJ3eTyDnrMWHg6n6Lg
oBLBRnzcd6r7pN/Q0LBCSQp9vSeztGd4CL55x5mrFQCL4TpLTv02btO3GE0yP6G1Kc01+3jxhcGD
hdW1ebF2omlNPILwf6HzWKLJCDfPZO/P+fObUk6tSiDWTQmc2h8d+TFyjtBpxmo5sJ3AzWi3vGsf
xFw1zZCGxwN9fxRh+lCKuyCd4gOiXYaxe5Z02A1ZIdLBypQ3pReC698bOI25bp9qBBhB1QfM7DMm
QBSCbyn2mna6tIvx1aUq17Muqkz/evf6jmujZxOjmVXvZ/EXSKaBg2XFVBWibKp7oPXI/x+DdkBi
cP1TobqHx0DfjsLPb1qmieLOlbEyzShtu5aehCID4Ig7QZi6494qeZ6tsyHhpwMaa7Yf24FK+wyd
/ISniINrvc8sbA1Ae7RsUFXyQpEbnK/gLvGiUimQfYbGkN84rS6MmTAjdnXck6aBOaC4YHeam+T/
jIzvniJxPB0w4Tr6FPAkuXtFs2nz87LDW+P4qZ+d9zZC+vubDgC5FNPTMgUzJW0pH+MM2E4il9qn
WvjJ89k7UELutL3DwjTsXZ3dnhF0od8Hr4xn/wkhMYod6IAamv1MHEkY705eQF2ig2+7XjSMsHfb
op5hiYk+gckdpHD5bTD9krE0prdGjqtvc/E6GYMOalAL/lIkO4xrh5jL44O/IjLuEZ1jIZtcAGJP
pJ2o9+hZn4Z8Mo9WL+x7XyCMO42PxTi46e/9u34Ow2C5bmlnGB6GboNt2Rg/gPjR6hZDZIabblgv
9iFxavenNBCbkFqvAR+Ikqy0eoJwEjbMsGdwZ3iNcHxn1lYpKUNwwYCMdnTMywLCKeYRdGegnk64
8hYQ+iW1SYrNImsjeX8yTTqI4u3yDBf0rnmrJYn5IR2yzpW99Vy1RsRnnrX9ek9hG59Ueo+jnjcX
FYQEmH5D/ONrOi3v6v/4/+LFe03EXkPo21VQdJS0msT9vRl3WQdfH81wpeGYLDgK0Xt5+wf8YWGF
Q4p5s5+jPQqmWi2mQ4w8sTTGKdCes9tkgWNFEzsFH53mf435JiGrhVkrZfLiDLDDO/7ZfTwuF++T
hh4JfPc9oq2b/92WtMXhyPx+HpyIoeYPlKjdItrzCrdNwBett59Apu/kVvzaL7Oyvkk0EQlKcGGB
dgkCPtjoUdFpHO0eY8WZ6/GO8ua+MTgOJWWwkiLMheA7YHyofJjd1V7jYxxPifDFTklBBEjpqxdt
MWDoSU4gm7qlExeJdsBpU98f6Dmhp+yUFRFbcT1T57wUcwwmm3gk+I90RXAcifLQKZhda89ve0wE
rKUrM6cGs7P6AxJzm7Wst5jKM7WsupUls/50u+M5yTG1Vd9c7bplHTf47zZx+iaNULxuPaXPSMXN
BI3ZxpsXP128kAeCRVCjZq8BNAqnNU+c8eMhdy4O4sPkpKjm07F4uP4pl59LwuIgE9uKnKPzl4AZ
u8BYN/lRJANxwz51XjfeHp8kkjyDEM+uRepflxpZV4OQqEpltXcHlEWNjOcuWIlNNzRshSX54WsL
SU3j2tJbjkULnPdSyezQmn3FafeDH/o+97lwNKF6f0QIWDGPY0T2mFX6D1N78lUZhS5GKQlHTJzV
jo9AJDR38iNuiOQlGAR89UnhLdOPnNefdzsNzYXMQfPGEzyRNCBZUI11gxQE9YU1NwXBPCrm4vvl
8ijzAM2fNtn+FJ82pJlIWfIfPVkfiORtoQVyRCOXx0PGn0IKvY3oPi9Oe9gdKvTOszcH57HHa2Eg
p1sTDHnxbtOgYXB6YBAr8DvTZlFpbxW0JGOdbzSa1JL/5KTTIMaCF2Zyp/sWnfzHb1TPMv5hNvCv
aIdcYrR8caweR5z/vRy6KDwJCtvg+zAvTq0+oz37L1++bVKRaSb4ffhNyMyIUe+H+k3i985ei7Fe
nkcauad+NNs2Wu3JwviIb6gAc7fas9fHks5/To1xm0WTpmSFDVSywezNkBgWgcrGk9aIaU2UFT+a
CTGHAPSvcWM7tE1/rFUFroTD2GGU1inru10niJLcK5wGK4wFVvLZD4zbEZpWbkwrdEuw/aHP9lRZ
fsN3OP//AI/i/FuudtWlAE6hUmkdRpJnkKRqmK6sRujiRkAGpql4SLcLZeI6kGdX5MgtYBp9SVPP
CS9uKBJxtiwzVUF+zCrk5wvKZmjhmNZsj6uNPYGqJ9/e8S4oGJL+G8NPJT02nXFAXdiVj0ksqUo5
b63GAjRxGGf/BYDAC0j3oZX1X3tiwQcVic/KebJcwaC9eC2GaJOBLGNqhvMFYVWlITT/QHzFOgdB
mRyvBi1r0DGS5Og13M/RfbmyvD7I6ePo15vPyb702qhNCPqL4KVsvgA9H6YXpH2i0VMrmSQiWfdu
TW9cDr4+dtY2SRRl5ws2q6abVyKU1tKoMYrXc6RRw1ixCElzKePtO/GH1Oh/0Ab8nKeKYYNp+zuh
A3TGhr/XDTM3h5JwRqKtOpTqdmEQuU+9MPbJo68/BBmTShIKm5qsdxN5794QvmBjEjyAvW0emzr+
u95W6/U6vb/nfw4gvY+iLWLh3fs6OXRpwchhsZyAUmTp++ChiO9wNceVYS8zDA/XxZuGolHSzRs8
3R3r6YXj/qCDUOM6mEUbQ6P5hdasIA1G5IX5QlLmpzlzNJytAaG5zO7pn8Q1Rht9MHlXxQoanZrq
F0qRFyR5nKzG0gp4ZGTtvUsDMQR91TYatwk15FqcEWtK88pzzjJSNSugmozoXdiPUo3d4Cm6RpwY
bmiUjzzMcAQgEGAIUmPsUBMXp+VK03QqV0UUxomY+W/i7Ny+gX2TQiv9cxM65nX0wFA+A/eudXnE
w1pcN7Qn4X0+WDogjGASJRtyNYH7ha+wLvQ15l7/C+M83b7lOMO0bTcxOnZriUb7ufwH1yqTyPAG
EgRwEOfbUB7KqcL6/pOd7S6/d/4WsSmCQXkgNf0XltsRWRUu1Ha5mcTaRl24JU+X8693OGxy9dfD
5ajOZRFz1sUUjtUZEVfrXc7dXdJF97qNuS+xFM9ICb1jQQ2uP0UswkO4FlolVbyZpd4Ppnxbec/n
jmXyrKKv7US00EiEHvoiRLaY4hjXFznfwXw4rSwxz6njU+kba3lo08pTsXt9KGZenLaP0WbPlgGn
lC2dIuoFTEv56VKUviDrILd46g7z50QBiduiRvsjntRamikl74DpureRMVkEkB8c9THKQp2BFEdJ
0+feweSuQsk7NmGnfV5TKSEGOYq2NpLGbf4x9ENiEPdBdalmrBMWuz5wU73Bi+EV/CgVXUQmPqFb
3+1w8vN9LoyAGeV42j1fE0rQ7Tq66F0C+YrEswEi9MGCP0LYZLN9Bz7RRbMyaAW/pbCcFxAXHKXR
0jOJSpdqMAIGg4PZZQpoGGjV54gJqvjmn4dS4ZDkjDJtG+TbVwRpaLgNwqqxY29D5nwHtcNVFPku
2Y4Kql5BxJV8GXw0Wb9Zz4eDdwnwYszQTF2EC78E9cr37/khcrwhzoHVLy6ep9jK2kSA09oAQ1Ky
9RpD+v0Z3odcQh6O7ET2Ukh7UYvfHDPPSa9zd8jrngxX3WVTJ3qKs4Nbtj9bhadZAY0ImrLjDVpx
B4e0fvFZoHoIA0Ri0OwWe9cSPaxh657LNI8Ekvjthe6ZuQmEnj5+fxEM88OoMETSLlfj0hhyJnRH
VK/BslFFv17mKnM8jCJirppCMGR8KHaBdpANiWGrFUi6dbty8BQjt9ClixwYiSTSjGy3UqWyVJRm
R6NN1iKIg7IqDBS3zKR/Z2++e7O/1JvE2sXIdLCDuWrcr7LjEagHwtI+sNCSiGvmRTAgEAwikpfp
jLXNde91V8PkQmWdTB2Oexc++VUxhHKUhNexItZLTSlWHVdYyyNst4FhRgnie+vphU2kywJ9liNG
UmAgwhdHwIIeDTNSzE3Cpx+lqmII/EW3GdCeRsgJ7XgDpDTzdEpqndHc533LaYvh5Rtv+X2eWooh
CD/fFTbbtH2H++qnBrmbCdde4MWTI4BJKBG8J1tGSuGf3w73/SlAKDqK1WbWXvB3QSIKpEfr/Szb
lSaNfNsRsESXYTO56VqjuoPAqcbFkqGzPL6ziqBYlwoRk1J0h0XHx5icCSBEwH3UIVttt/4qxUNs
uwITBnurMC+a52t3aYrratHWFKYep/q3lcyVBKuJUE/HDaRKguankAVLi/Wp58duMnYfBUamwtdi
JtGWukBIZ/NEpLNDEFCq/BQvlgP3eWAo0c2esQbwiI4ofn0Ow1jcGntVMq2/S8pxg4VGK9VrCcub
/yzw7EdSgD04mw8J4rmNYUAE8EHxyfa+Eu1R6zPxX9/CCtxBxAvxiiY4Xh3Eef02XCo5oqlJvhvL
AESW42UplsoLTI0LaFTZB2TZQep572O165KI5dnxKNSUhg8ZUMvCwZ0Vw+Jbj73aK+Y0taiU2Lxa
q1hG/zYoQA19GzaNBZIaDT6OgvmdAVKUwD3QdQXhgzZlsNPgN5es9LpGWqSCB9SNINLskQ+vu72z
eVwNA2OQJish8yqMZ3Zdz2Y5wOqUJGgHlbMuRwZXyBamXF7da5XzSQVPA6Xg6jLaggaC9727x3K0
D2QKFCM5jMKYTMF5Ye+mD3TF3TheWqFrpPZeOLFB3hsdsKra7MAtnBvueTqfsZ8yrvC6nBvmHVXC
hl32sArxCkdn3VlfTBFDnJGhy+XVKavZGbvdwFRH47HTMR8z0t6mpWASKZf5kDy8Y60JmeMR+r2K
u0+olxyAsyT2Ji6trYc1BOp3JriYBM89pFBIZyGD9WuXYOY13Pc36cEQl+CwLXkfOAY1ik5kiZ/J
URUgLrL9cKk3ajqPzfXHf5hifVVd/iJ1dACoSOoaa4ovoHsj+5CDfO7wnSIlm47cogWkk/wy2915
ro8UcJ0gg6/IWTVM7GKFLoodUzncNfcOoV6wag8YVZXwJ3bt53LbRFI3tFfHDlvQTi5f36FCjWIg
rgVAwJyMWv29tSQ5ktGLOwumiOAfYHDVgKGFN3HOejIuHU28DoZTYamt1uJ1rMSw5+7A9bs1OaX6
OSgm5P9YwNeUrZV2nb9Qqd4mKlA/8ShfJhQRgD81sbFg1HtSKjpuOBnmXF54R3Jnrc7V0yeinBnH
embPFPlxRxAg8rM9LhnoKwJil1ZuHBk6smOTP3GtPXIWve4iTvmBrvNOx+/qgFwVtMIWr6/gS0pg
iLFM36HAvNb6csaHzn+SuARVUBDBAZwgl1jUnMnDhoKT7D81m/CQg6q3vd46i0/tdgGA0iGV4Gfr
5B5hG0wP/Bglb/r5f0nSgq9aCnFPgzNDkOtb/CWRlgg6Zs2Sz2AJWj+Vkmhe+drFDtHSJ520W0OF
+DCSiXqTKBDvh+V3LARZ/3diYILSyBTtzmfLUNSycu5zJ1DSvhiehwThz1VLCKOjV4qsoXSX9WV+
ZW12r72JVNY3QLgQn3wOs3oKVeWYe0VZ7Y0UUZezgdimdCBTDXcn4K8C3lCrOt7/c/at9mVFNsrl
OirTTbG88kgI2n4GFqPzIGL5VJ7+n6NpAFL1b+ic7Nwz97ni8NV+y/Ozy/sxj+5cwsKZGuXJ1paQ
R6vp6ZBJC6QRlCV0BLqXmhLzZDYwGSK0CEMXhlgPSaJeWDVn2g4WIlxbBRISGi6QvM/71xYiIg5N
Qj0uJxfMEkQ5N2VcoDQYgGABzKK3kb8jmUJdT7cSpqtZh8t+guWM6v1enKtcZHREe6bfVgZn6daD
pw9rH5K6KIRU15BlLGHNMf2IZwFtcMq0ZQrulhOiKm+PDehaSIx5cPS7ja54skYmp10zr/u9zW/i
ASxOzbRZBmrYsXZ4vk+gB2B6rnkIhyB++ngn25/yKFoBVnpmjU+YFpssCwvorAQgpmX/l2cf+0TX
Kmn8t6NEHbqkFNJXUgUAsTCtA/e7g/wKWK8q2SurPKdBl4FoSico4wvWC9RnHhkoRRyQNQgU4g0u
6YoUtFv410CfJFIl6TxQDEl9gBLDB+irtKlK+kJsloNJpMPWx8x3jgG45y3EavMxtwJQ/qpVe/8e
f3IrQ8ZHoqXQ/3e3MQuyxalR4NQwchxte/1acoos6L+/Vxd49a+xBV50ilD0TxQ0SkWI7CpjkrTC
PN54cqWmf/1CdkBv48SIoubeXaNjKOG28uPXqwIcKqNXUi3y4g+GR1BVzqkSrSsI0EqAjQOOb3fn
J3o80Sm7lUNDe1z9qB146dk4nj0CuU7uKMY/isw2acAblJPPgXdJHOLKmoyvRe/w3CVt57rHB9kM
q6Wo/+VrrtvdeeLUATLhQ3C9lKot2/vkqL9LO2cvDwrp3S0kSGDIoS9ogZ/FWE6lIUr+8y2nyP52
GfCPjOknomI/Y9gKtVLBbA4VPmJWvhfsxSXBHuXSflKOv1jQ5QMITZ3jOo9BLuQ3GC9u1pd1YocR
D7zdJqZJxjU4fgl2lx6xHc+3kzZMsPy0dRGnFEMmy4518Y5Xeeh0ctc3poRVNFEUJIbn3lnjPIdw
ZkmD9zz1tWMlAShG/FqkRspbhoABcJNjVitgM2C61CKXAfY2KhuFPauPhiG73/09umnhUy733EhA
wU5MGXuwG4SE9bbOnTDORq0tUHi2p/l/vVKe4A2QbLza8ojJT3nD0DU/GHSkCHDX0+TyaiFAUR1Q
cAvGRTfejq7tyQCDPowr6/k+qwt+C834WIe58mMFqTHjggo4TdmT04jscnjRtNwfIe7CoI+I6uyz
rSpQG4ywPVoOuJJI8NaGhyStBTkLiSL7+j0zQv5kEFEmvOb2MOE6+K1lpSR6xPhuRAu4aTal7RX/
AcOOT0ubXH9GTnZ8rkmJHhvQXVH29ZneZF0+34fEnXy+kga/46rmeVnEIYP32Ju12pFtIUNwUMV9
QdWMpTXVT3FikAD08ZdyCGJLKigEnHwNCGkD2l7SU4/l6+oifYG5lSXPeJTKU2MG5+YudlmEr1Da
Lm2wi/DWIVV30Rc7TVNqdV5DWdt31OPGNrmFALAl16ilmirtULdf/OtILgfUH2/tS+VbCwC/A805
kwRN/c5CmoVWcvZl5CboToYD2Dea/iiRD2DHiPdJUYyRiH+jSE+IhYfx54SlEApYCwNEdd8jWThe
9NppYyD4VKjZGeexyFYQPh4ilFNbnHWhbJWmUjTzyGoZdWOCFGNISBZJlwVGv1/ipc47qLjsbGC8
Vz19fZbDX0a5FpPRZvhkG7aCe7QJd/5PhbifWmRXOUDLuKGh4ZYpA8DmEJt7a+0Eg2xXcPYvmUR4
/mTZaye0H8Gz+i+zSH5PPIOWuuNXrpFvG77ljWSkKQGdK2cKU1KdmoMRTLgW0U4Kod3TXjq0K4Tl
Dr7haMkggJxnpqbjzXtMsd+lS0jqPDtBj1s9obxPSw3SIDp0A7RVuqXoWHsHgoyFYRnnBjQA0/1F
NMX7Wn/dBGPr5WID2DFwqtR95HGX+7j4ytNIXnhHY0ieNkVvUIyY/mbDIrfxIBww7O+lQOhKb3O0
TeKWYlN7PuTZWNnXsSeLPuGPrOM6xl0e5YnQQM8dcftUI3L3iPFb3kSEQnzMW8rgXG28fft2hEgm
tY4KMy7RIPU4peQcQqi922edT4aTcLAAWLEIIbG7PGZUiMtJ7pBrfvnX/iitLr+kUr/N41ePAwom
nw50zV2QRanMWkXx63khgOsWD1VCA5lvMHzowCJUuEd5jHymzTT4j35Qx1dZXRTuUR4LeO2uh/rk
bBLGWMtOIKDNDzp4FMJ6TVQYJKyaICrPV/P0ElXB5L1JghqUb8j0X4eWp7rrWQ5d6ai1DUhqrhcv
BzfHYtTxHexre0AFeJwXuxU863sDlUX+EUHRkN9LLGoOYjnpAL5cvuQdqpXNr1aPS7zKNKR2c7V8
RD5TagrQ7DKgCdXM0paGStbuGUJZ5IfPxQiozTyBSJvrDpQwARsa8ywsWf7Ddredzuyvqoo6GBcq
meC/mKyi8EBgdBCk+JYByx7fcSAXB9eVQgW5ElHwDbIA+JQQsbt1q2eLE7AD+zof3V/62LIZp2kb
+b2Pu/r6U9z5HkQvAvfqYPBsu4HPV5hPMNGbA58biP/tftLct6GU3vGnbdIcjKaaEx/nTmzzTgo5
yxYioVQ0UkB5FJX4ctJmiYKxLs3+x3qRAbnl5MRZE4eKvGKsWRKzHoar4k2So/8/x52g5Tq2cjmq
gaYPoqdLIwFQpd0J/ApethjABrhfDNZCNb1rPWZKOQis80szGUK21FUZEuWQWi67JIAWcGuRMDbc
R2cVyNHq5TpGm9tZCgbvHDkmT6SqpfdACWWz+/foqxaltLNLOaJ2h9RvzeapkwfO6ag31gj3J9m/
WGrTFvOBztqN2TdYSZ/RNXoqg4vKdD7XJXXl54iVsSFsGUKlMxLTrgRlUC3x9eEY27gLrAaLxpVV
V5a80KDQrj+KNjHY9xkCbfd2PiHloiyF4bXnExHAUX8wZnHA4gXNNOP85uUq7dWUCXK/uRlAPmhR
VDblcZGwG8IDgT3u5tXCE7zQa8u9RwwSt+U4E2cklPbqF9AIsXgk5u8t2zesIpMXF/kVKkpGZ+lc
LXQr/UyFXQBX06uI1PQzcerO3t/GqTpABHJh8jtY7tvJmgUUTz9r34hkJNvD2UfAYSx1Ms4u8SDb
dxzyIK6EGRLFsbBGvFstKXK2qYg+vhV9ldF/McAUfwBEM5OwVnankyIWRs2LvFDP4koqsbd/hW5x
nXA90lqfnqPANb5C+F9yuJcB58CFrSl/j0NOdf0d558aryrSoY4rcnqB0DMV1eQj+32FFs9i8mH1
CGjfNWdEfm66zK/wd+yypzRm8zq0pcHj0xU3n06lC6rdHbdK2mAc3RZ9xS2HJBumCjvXg7eqS2qO
12CYvPcHFNrD3xMqdpLJvlSa+zPZGZ6MmXA2/TCO0o9qil26xwu6qNqsdjOStftpNwwTrab9bP88
BCvB59HiTkhYz9xe8cfNPEpL64XnPLQwyKOdzVJSSRjrszbWDwYn5QUPSkk30rjttUmLSzJxLBmG
KiGq/BbEGm27/ORKcxZMR1w3hGfJ2I0jMc8qIqW0TdbFvdp3y/6rF9N5tJVw2MOV5mlStYGgAPGv
h5DnrqV7+wvuLA1ZF4EkGGxP9GpHwbuyFgQhO6IJ5zaAnGIYXbvmAAp45mUbwa55S86mcUtjJ+CU
oAqPkmcJZORXWP/EAp7aXP5t0rq067qKhglkodJpG7q3Py4gCqJwWsLfsfi+RJ8rnx3bdrrV1FK+
PmQiLQBJWqtdZo6CU3lKVBmhUDV9Gu6F30JlbCTs0iDhkuBRKbuXgYBjihDe4ftw28JjOtGCaS+D
QB4S0PqdEETqoMmWMVyRXOH2beMKhzh6vWXT9o/pc0psuQmR1shy66kVxI7kNP43zsnIot3o/f84
BuJqaHDbFpH07fW4M17maExv+3LpNUz4XIcqx4vtEBswez+AywuO6jIG6k4K/YDXCi9hqD8J4/hR
noIauInOV5wpB1DZR7V4jShNlolkKasJxOPcWlcqQ7U9Nu6igutTNHtA0GoGolbtW7wdPg28MubZ
YA+dmvy1UJdhWpM72rVZkcuKPMQyimUDjnUXOYEnrM5ApjE9IUMfitZsBdoOFv4Gymql+hB9Ebc3
czQjOg8aC1s6JuzBCYEEOEPhSS68RNVdk19nuFKHZbeOvoXDNELqM2Ac2pjOYuxT/3f2l3BX5Gtj
5+/K/yCjulIuMPuGrHS0+q5/jLX7GKQcdpSBOXqUI4QCB4rsq7San9x4IrI7vzyKpm0XeAiifBtS
ytH56cNDeu3lqU4KNL7yUdlfiP36GtgzFQai+9G3OjZ8CTmLxLlC31OkCbWlDNF7BTa41okAfK2e
o5mDHLqGpwKyBnODnWSelHeLxbT1hdOjm9r41CrffCJDXb4jHA1n/IULOeFdCWriAspVsuA57XUu
ZcA+DhcCYIz6L965IrJIA1GEg6Yd6dTBlH+WWicCtKtTbVkXL25R6ewN7/F1zowgMcmxOLzik6WO
fegUy6qLMAo3lQ78CMH1zPsu3/UegSk+GhxTVellq8kEaHUmgCaqFbBD1l8zSp7MuIMOamJdCM0J
w4VKl2cqzgVt8wYXi5c2EGBVprgQ6xUTVw0zaFPgAJHOe5l3z08Jr/10Nad+qhwmzwQLK4Uk+J9u
BciO3a+Stscrql5m9ZJzuttY3atO9jFlK8p22tsVdViY0oIe2DwQDx3j6Aq4vDi7mwjo4jzj7Alf
GWth5y7ivmkC8PsBH4oK4HWclyAX0hPzvM509tAVraKVpWZugBFl5XPeB5u2iR1iZR5KL7c5sIX5
91tiyLznAmpFgkO5Pg+zYOcpcPfcgEZ/i3aajsg4ZkFxGUzYT1qcqjDtD8n0KCUC7Dtdb7YODFG/
tKcJzt2L379s8Co8psLm/FTEiR3LVLUr3/4IxZJcS35y4Rx+8iA22BhkBsji2VeABzsPnKQ9/VRn
7V4Yz9/DJRS+vBjIok7HuZltSbwSCnekVaHsA9T7hXWgrpLaKE6gCXuMMr4pVc2bB9tRJY45S6ne
cC19BwAUGXFTAYxn/mPpqdhn4IrzYUctzjH59ARcCy94dZoavPElOhGfzkN2BCwEJM/gnhlYP9cW
jK2kfjcdK2whGHdwobnRkClw7T3fJQGdz2yRLQtqfpzha5qmiY7HhASRR2aHsLX4cKUoNRx1HnXO
KKGhQ1vPWVxAcA6M91ntDNAidIWhPdXOjUJ4c2VmgVkstbZrn8t2P0nzpkOsB0SwCbYu71YWLNqS
rUFy6VLcpVT1gnJ1JuuI1UcXuQf8+VF3MxGebRQVh/JsZYdo+j4mPVHnJCX0EnNB367+PtFDW1qK
khiqmIBUsAXMuTgoRm7d7wZQ/vOhqqibK7DaS72ugIvbxIe64tVsamtAaXGP0mYwfJedwAoMq3Hg
ag9ThcyaPBI0VKxsotVpnkVNN2oCXoLyxmczHr/2HDvZtklfqYhuYb/y0i7Tx0xdLOZ1CMl4huqG
0PTm+DiE94VFtQIBwv10Wnfa9rgWaxYk90UKSgcBnd4oPGBGFgmrbtn0hgiZbt5SDZ9RAQ3s0/aq
aQc5CaYkSuorOgbRj3IskR0RKGgLkXAAOYVa7gFMYak9tQHsELupbd2J/TgyV6Xiax2qKJSNA5vd
SlHCq5Mc07LSEJp0UuVXwtCle6wOI+AinsRA4E72jovJpnVhGDQh2SZ2cwSOa9v0eBMgNKHU1lqf
Zj59hWEHnQzEkHD4GjXl/rmkrBCWe2gZns0VmfYqH8ABHhUElxQD9sfkDATKOdxnJ+7RRRa2scE9
jptyAIMsosqOerN4/9Iju39I0ZLhsyO9WFcWlu+KEhcOsVUP1Lf9qqYsgLkmcgTHAO8mSsySKv5J
SzTASM4awBz+otikOUlMR8CRoCD5fPZ0zXSZQuJLD2GGNSAGPx3JrUPC+SypTaGeOLlnt4hWIetF
JeH39ZbQZKQe22+FP3s4+WMiLuwIEuQBLKrcZQ/M0yj6OujpBWansmOUWvBKSVXfkYZWAw/udCDw
LAQYR4H08ygVhP3M8XQYmLsFsOe+eAA1mLmCqqiswt4ssPgZ7iIXK2r9QkGI5gC+DmpyrtdFBQpV
DXNlhNz/uDdwPb5skNUKjMwIKadK/JHBMoa66HoAPkV6hChDynZ9pq1LuOXhhkaHFvl+TNzxba41
phSUqal5TmO8mEL6X64reQnd8MdIavXm1zT/hyDq+V1GzNOOOp3lL0uI+WrW9ExlX6vBs0LWwNTI
s/J5wkZ61sphAL0ZIQQbQ2FqQ8eqFES3W3odyPh9oaYahP3I3swmJFhPcSXsuPWHMlVcVp9Rr14D
4jRFF8peGjK6y1L7+SoTBzpnETxLOJNT2xSIlo7g+Zgsp/oWOz2gOJaXtHZvT7Np/fXMgvHEAcb+
2J7g+fc3wedZmdC8fhG2k6CFG6LoMTda/7AFV4UUtPYAvtBMMeWPESqMUd9llY2Y1VM+XzF9DSuM
PqXkykz5udwacnc1U1oI4CVR7J/eiS9uRgFlaDS0hTl2XtX9fuxJiTk+LizHB7GSSSIOswn3tl3o
vasyEy6GsqzAWF4diyfbbh5ospeUmjWtJGD5LtR9VssJb5LlRZ4oOE31THoF8Is+MsbvsC2mXP6S
EQsI4RkZxkDTjkuzcRZnRqwcdleU3zVzQ3dC+Tfmvakno2v8vxY8uzFmxOLrxFuA/ygCx0r8q0gh
BXCWTPY0gDfJ/VY/WAPFhz71HGTQ+rOrT5/6SHcIiM0xZdmj95qRZmn+arhxO2COMw/d7Sb8sOjd
uD2+Su3/DRMKWZIFemVYozGqKgYvUczeO70w+vmcvpEKSi6UDbUhj9/HwGvAgeaNxP0hCE2KxnY4
tYh1k/5B29Z8edsfw+YpSMI7EVKCiI1zlA/4Z5uhcgZNRaukLu6mwaAm6cDK6p2qt3pLU4KqDuo8
L/ZfQ63ykhnCbiBQvfkCXdoqaS9OFO81lkvdew14SssaO+enl3StEJJPVe6v95fLM1c9SNTuKHrE
h2jQuHHsbn3sVV3IHxdrNfPCCifzqkS4IbZM1Oua0iGdP4+Xr/4Y4sa3ZBw0YfWxmpzp98n9oQEv
tP4IWp51VwNUQR6HDmNWT37UiVUio/Uel0jIVK8LwXQsv92n4uMwacrfu+8PHs4X8yVZAJks3H3g
YOiIkT5ruADyMJ3pC8nOpVGBdgDmdjuzFcytN35vnOARclWWny1Ng+Ao64E4qS5gRgbjjn0mugo9
Re9FrCii0lYSJJXKFr29IybcZJtXKg/A0oyvPPBuBuAMDH9XmyXfTf4POhZ8p7pt6i1HzejHsm2Q
ryKCy4w3ZL3xLqLSiS5xII8ER2RfWs+lnw8QkJjleV1wxq5OYj58sHJFBTLe/Iepu5c5VQcM4bji
bnH8ZcIJZPTBMM8VqjW6oxr0wzyec+HcLnK8f0SMv1o4y+hwrqnvbW1rjNGs/C/eTFHxiMYXRxgS
xiung+aBgJdLRBQWT28w9Kj++STMXvmdfaeiXuRsyphGcTsDsIf3I4O1spQNxDTxG//U3pJM19LU
n9kIaMqSnGC+nKxmNvU7zBhOWHagJ7yLeF7aAAn5sMrHbk8wkDtV+ceYKVkirxyflIb3AihwOqqi
vvhNDeIdLdfIQg6TOOmPfa6QxcOqtPi+TUwV3ffT6znirJ7H0hmjcts6FzRZKSMAjm8yUBC4wNpV
R8tSof8S0hQTRPCvrrtTUYwXLpmMbcCP8BsxsU/Jy2wSNDFDf1Ahtt5kJpKCivvZX3mzF5sF/3Sc
1fJFe7yXC11i829/y7f+cQsnsHQAEejKvQrSAoqwPPoIRj30r8AGkEL91WcWT1xVWChhj3XWLDMX
D60DwigedLHmI/6+bVdTRYAfXSOOLEzpVMn9dfAPKhyhU7X+2vbkL44iTH/GNXb+dXm4UZ5tUXyA
VUlBzcLUjd8ZIOGf7q1j6PKb9m/79isvgbTyllrWoyL3uANyS+2Hcwj6Dds3s2zw7qQu/aGyGAkb
o7Spb0q29YWRJ98Wq+Fxvyx+U3wdRWz+PUPWiTFMkG/ezqDCeMohRMOimR1ZyFnOg2XWXCmYI3k1
KK6QoCCa7jmhWC49VDVbHp2qCMlA3FOnJcLNlaPnZIeBq6TuTaD/eA1EIqOZrey4iIld0JtbS7c6
ByNzL50F8+xN7OVDqWza7FXKU3YRLBnPIWf9FLp8djUeixatiSSO5EjIyRgRg6tjri3uwOrAaU7Q
TpH/nOX4xJUTUAWGsO0JiIQZZywqPdx8ZL8CppCDqliss5/lw9GYBadPBa/pKSAOWYrqX/1LWEaV
JheKTKW/ko8sEqGWlei1sEnAq80fnmjgk4+4XvkG/mXogRWGiNushBMaWotJHjeNQgyFK+jcHTJK
zYrgEg6ZFkVLmxIkvDiTB72PZDowYbXXsLbIuZzsXisEImoFG9TYgqoxTff2X0wK5Ns+F0CO0Ieo
eRdopYdHaEF2hHrpQh1hBFdJ9j+zwf+t/nwHKZ8saixFDYnfAx7Ectrw1DhnaYBV/6R9vOYifHWi
v+CrgSYjguUM9BxaFpBhZGYfzKdg24PEPs3EiwSDlFmZukQ5KgGfu3cuUXWmNjW83/m+GbeBvZ4R
3AC52WF2h2zFsK0Ut9p93wfwQGEJwwqw0YzUobQi/YVIISxkYDySoAyIhJRDmzJ4ODnC/qyobrHb
+/2YMW3hb1Q6HhKpC7o+O+wlveHzY125EKEir50siNXXgA1X6GAhfBvA+wjKMEahFnjQSLO/9u1V
temP50LPQMX6W1aUa82tOgG1Jgu8fKDNRPCFWlegktFGVqzcziNxn15TJ/v6v8yA0eV9Xjoik7JI
krEaynYLsQc0nQp5f2zzGKWtS4gyqCDBrygB6Dak0c2Ahknndg7fhU9I9RBiXtGDNbQ9s70eEDfg
3dUgltd7JlX6BElBMrhfftxIDlwFLKFoAl+Y8OjoxR6XA2YnvlD+IGBcat3UIj5igJYmUYAx4gRp
H8Ls4ZiaIT4lVJm9FTU0z6Sekd10QHOCOdtyZ1A8chDkcxSdr6mtYjvxUUq4fWUKlTxwleF9GpJ4
rPxfNddiKEuvSjsU/x8tHGAcbe4K7mf0HbhAjHtcf07DHdQPe0syQWGyQwhKd+7MN5s9VzCnqzi1
vjv2BzOQYckl+5Tsufv6Lh3B+xKf+InAnqw9iMq4qAQC0TyiI69T2iZKsGCLbBWRqCpWehHiexy1
GDMQwstpgh+PzBaadv0HgEEY+PkGb9MxflX32O63H899ZyswmI7mE89WIV+IyLcnf1wB7SSlnPGn
fnHL+q08la1FqBqGWxoYIcQaO533ERdY5RAh8tlMpM8s9WrIAgUqKZm6YHmwNvAQBqBgF19dpjqi
YjTfpNHBdz1FRBWsKuPu7MWIaEDbgLrQlxS2nFvJiZEUea159ImJqFqj7o5eCbLVrZDUhK1CUKGJ
qwgoEqv610WcCDDvOs7SgKhE732LDMr1dBXV6KV3UELkbJn/ziJ1/17B51OhIVJWe8XXYF+fEVO9
5VPLzjuwr/DJLYoinTCtbBbC6hmu3Mqj64V2rTNPkrwDZQYcnoEOJyNCCrrn0YgyGwqETddYsmjr
TDV0vIFcFF/NjOgJK8FV7kOE+rXuEC/U9kv0ak0mrxaeTgFdf5pkgFoTZXcZb8zmUm1JIokVoDC1
nc8qoxutQWWsNTnigdq059trlQNCiRcgSpD6QX06qQHwnNbUfocp37hHbY7ZO2g3GlCVVA3B0OB1
myRoa+KzrdpUTC/JhntPl6lImk9whwvtwdHZbCgNugaZkT4EovEZ+sAbhq0v9ZrRz3zO+OxElVu/
WEFluC94POiGWdtEhGk++nvzbaAzUx2R1W28hxnb9zVxXpJjjMqm0NE9UKrFobdNy/bmmAT+HoBb
krIDD9t0gNSpA2TzRngxUAcsi9KZh9pMGF00uaDnco1X1C2Wvp4s+RPL4+K6c+zTt9zbiYA5Lg/X
kg5mShozA6CILzhyuNnQxBrQCxebz0XW5PYKBMAhcMWtHRswo0YDGxv9jlxqreuSXbVw0FB4CL+h
e/ChVAKZdF8BIpv2eaG14D18cEKF2dBKIf20KhRFrdcDsG/08UMXl2Y6MOsMtSd17M2ZwkvsXot1
IL2JjaP33JaFa1KguyrOvT2rXaitrpFJMytDQ9smpLm0zLU4IUCY2JYMn0pzrwp74eODS3upQYuB
8UzyPju8CODXuIjcPGMaUy4K3JbsiKDPpI/ab2VUKtpOl5GKaHB61rOEUN9tJaALrZ8wiD52mhKr
eoXrfgyaYfCiod7phfP6QlfXr0jWJ9Nuqxq7eWF564LbCItzTF3LueaubdL3D924ewZJ1RFlb8HZ
yjwPdLbA+fHa4+q0RDoSBamEncL3pAi88nTsQlFjbGqt5G+QCFuqxvOvYU+JvaOh5BErggrLalQN
1DsF9a0uUrY7yPkkAH6k1p3PrijEAm7Y84HiMeCDoQ4Lg7a/d4CNApcX5ci3A/KhFxHmxAYoag59
5jQgPn+ZhyB5QcYOKPgsKYaeSqpqRBGPg7FzpTQplnxtriEEP4u/QQ0KdLSCKTTl3ERL7kU7dk8i
+Kzgpq0mlNLdKx8wN6KZznAvqg3sjlAT+ZvKWCLhHGkjI9k5PfkzfaNqAqaOBl34IBiCCtqGHs6N
Hdix4kHI3WiQsjb8P09L/xvVyHkyijLnTGKz0k0NX5CzR+acPw56lldNdm0qCs1/TB6YD748BR9Z
hY3ca2P6HRU6pz7epOUtFRX9d1lU6hnjwtsnqAXSJX/ccI6wpvhgXIzK7aQFbMaCRCQXOfOOP9M2
MSk5+syX0FAflBrMieBI7ODoUVdx7UajCCtFKpsvAo0e9J/lyFcWeCXK6HhQjixg+vna1OB0Khz+
vpqzQ8WM4l255ubfwrMFlEut02oUPEdGnzkeuUF1WBfhuHz9oC9PaCs9vlGvvBF9+p4UeS3NZBnx
rbo6oxPBAOH4IWsCIaDHRo0I86I7f3ZJwSy67+fEl7Xer7Kin8t9zFt+VCkDdYzfpvHA/7auJSY+
JDCeKHaB+K3aJNOPAskxM1PDtYxl+JEiuU2DYGQS87n1bdOV7aH4EluU8DHl7QP9Dqzmnqh8+bTO
tFpWI92JBnX1lZiYVo5NJou8fvpbxfUZ8zOi1lXjIqRfOG8DhshXMaWYC4CdwixFtq7Byf2QFmDj
IGntdAmIGRehu8eHgjY9jeAd0sBmJBlxG1+fKiAXGNbXLu0adqzewgdquPSh7NVGJ6TKxkJFvdFW
qZg5yPoTdC0GjkE3mw/UcbGkKRmtoxNqM+Qwl9l1ZE2KC6fUzZ5jgEwrRVynjdtsx/w5als0UYsG
fgxt6SPlk2XqHRiJhWquUL/msRAWb+RZGEi7GY/ZD9VEzEv5JNAvfq6GjDu5fq8Tj3FoKAgQNq1E
R/MWNfeU36MlXewFZCFDP8xL4EV/XVjQfZWLXH6j9rhcPhtNhhKqkS3BbmsDLnoZm/hu++Dq/bhh
QUx34M2VVispg1qnmQiMl17785KuAbzYb/MCVO4yA0IF7hM+KIpqrN7EZ070Rq0Fw5plLBePdbFp
oiC9N868V95+gBzt2HU6gxmxGcR63bg0ERcSqWrgOYSq/DFJMWYOelhaMrIuMzIu1PXpeooUx0WT
sgLiVTW+wAoC3oJfULac3Fe0Y2rcRMbjRuuQhRuYTk+AdiVmJlvxee4Hla2vAOAp9HL4ufkeOqFe
0wBZ6GK9zlpT+Z99mzb2UJxDVhWPtXq/KSXaHwoQRJald5pHj+Kc4bjgJEK2ZdnKaC2yz3ez5XDh
Quj33zAT7iSorLmGbNK81U0nH25tPvtdZFXT7gPMqRM1XN6K4J/HQMbsCzIVtbLfRGRVZ6ZYtUPM
3OlmenXkeItqy0OTZaM3KOllvaV+k+azRzrNAI8aOSqmrwCuSSsIC64pujTXDxtqd+dNySOnYqvV
DDmx3gBkPF1jJ4mvnYMga0cw4tRlgEQJeekzoPecatnoSUCy8jE+e8gqHbIj6JMqALUU/r71hTsN
H1FL4IRLpOzQo8BGOfoDf8Vn/yhsZRjHdO99FBhYraX43H3BPAPGSrJ9N+8ST/2ktq+3TtSx00DK
mc8zEd1/4kZmOxRcDSVmNFxjq789JmUtYoXckuzOOKBx36qnmaSeqZiZPA1tqC9LHlupRoI30UtI
GY15sDnHQGnxNS6h/iCdHV1J6yJF2kKdiceGS5FZDoDoYX3vP7RjYrmp/fFWzLuDmZQn8Awt19t1
hqwvFHhEWk3McZcu13lVGrz3b3vNKKrBJ77IKPcVq9IlCvrDCeOaB75sC0V0DKTn1BndWv6fSX3Q
tvv1CCJSpUo+g9qo5RKJgfgvoisH1Zi2Y/Uc1KX9IiyCnJjtylUDDvhr5J2PYZ9f0gC5H3SMHdC5
uPWovJB/cXxYCo8pdyN4ZUBf03yfIF8YkdiWX12Z6uwhu8e2qAFXeEm84kQPVlI2GBQ2djCC/ED9
s4z3FPdDkRVZPX1gpTFXFygFnImJLxPy0wj+TXveG25BXrMwwfzfjBFH05AbId31v1XhKbyaZiLY
LxYwxoCLTYXwGvYt8Dk3pvjY6uzcnC0pyhfTKbKNvuZw3DA9tyincmaXsi21tLsykI/n2Z/sqAFO
b/O4xL1fPMRThH+FFQ4LzdhmkGFoV21fkoHT0R0u12356jyBHUihJKzZZgy/rjaXPHCXYBuk+3A/
IHQkjwH9YcZToEQWzGWeYemwT6z4KEpIoHk+ZQxzHQHni/sPNuKMGlzCtLUW7LQJu5yixMHsMbwA
Pj91s7XXuVLu3C/LBFE4rnRe4jnJv0859gJpk8AX/leQQs2InRoDFPy7O0X4r39tzYZNSMrNAt8h
kHP15/fOqXxqtZM3TzXi7S2zQ7P1z1Zk1ZllGJRQSO3O7l6c9ZIwy51y1kcKDeMok3usT0ZbD8rP
pUAl/LhyEgAkFWy77eGKjtSZa6IycsGdbU2poUY9DO04GjmE4rzleRmg0IVslL/OyNpRmKQngHxu
LbGnwxOUMD/ro5UjES5hmTPqfMeA4J/kwQxPFdZQRj4/w7Ir8FWsJH2VUczA1NyJtbLm9dJ/6hsm
dXusegDVVXoDgjab1hGha34tjl1JX4nY0quXYd9d3Th4sFhw7dge3F0oRqmiL56jSKNdfa9bpqj/
Com+CdN3o+Q+eh1Jpx8ZHc17mH6PQxc0Dq1nbbBLYGX3SR5R/ofsWjojJbF0ap4Q+99BuqBJ/6fR
HsPf5dc2FVz7FbMtBTV7XpGjN9dIaVCuvEsy4Be27gWohW0nQpm8hRcg2Uj29S5I14fl3Q1f0TxC
fe64BUMZVYpbn6cdOJF0m+8XHBNUu57gSEch1T2Xz3i/u8aogXHPmWQzJckzTqq0iFMOJJ4dmR6A
Y8JEzNq6/4crwTAK5hD9gfllM9K+qIT8XNmJv3jwj8sHXHqsYC0EbEcN9S8QUiRP+IqDyJVTfLhf
TqnZXq603Aj/HwdB2YQWS6neXj1K21fBNoNs7InW8273astog5g+ZjRARoycrbp5HXqdM/Ko84v9
2aBgGm22u+uUUGGzylpGMDxr4gLMkb+Gbl2y5IA7BG1iZys6ZqF11j1ZMXGphjNQXCj3gdnHBOko
N1e8VmBTq3VkQlwtRstyH/aoEKLWV7hhjF9eGo/1teVH/5eKUOUdrRVDSHaoGoWw3YWwtwQ5xJ2d
8jZUX+AUpKE4DHi2gW+joC6VZAk0nwo/vCukcZQtZcSO4lR3lJvCPGjUESQhEJxnv+o3KgUs9IDM
fcb4QlVn7W82P0fhRvwFqQQH/t7V5ZBEhmKTlOeH6zITpE3IGfmOpxK1A1EH0LRFwO0jURJHYvST
QL55Ua7rQt7b0fwzuL0Sgkp3xnxnArWgY4Ll9c76eloIG/QCl4G27pJ8p8w23lzX81eEaDtu8/Hn
OvlAj526DBndb28O5s94gwJeiUObSSf2lkndTosb9jBDBQascOV+lp3PoH/J43dcKeZH0EyowoNP
a+TVZKyR8MWqKo7TFa84CuDqYMMxwgmnFm1mKzmuDAXQWvxEW+/eAGpV/2eqA8Iqg2BJcQkhx73J
6gNuZlMIK/bkHd3unptYA6pCDBg/iz7GgYOt6eQeKfAs6c82oG6AoRozr2Z2OFGupukW0SNilac/
59zckkauGJ94Lu9ACUrj0S1ywmCbO5FipL8+pZChwMcfWeZPdEWVjoyiip28e5B5BfXOt8pMwIuF
aVKIs8n0Msr40so3y3Vw5eKeh3W1JIbvYZ1P2gT90kNa8Am4jjtMeJJ1FDEDQrpXSVjJ9WBKbirl
f3HBXdntlH2hgNcAKRclEZ9qnyOFSePVNic1nwBnqJ5WP1soydFQTXDsuYIQTbsnboT5bj+uog0l
SHRO/J0jvoxwV3nNzyUbuaFBtuNRDe74XEoamKSFNg7eZ3ggEufqf4Y3L06lOD6TuSqUncWXGYMm
yR6lr0z6hf7E5VtliYkOP0DLm5O6SoiqrlodIgVdJgYoMjWql17WBmghAMXhPrB5fMO7pugk8CEE
fYuMUCa+kOKCnwckOo44ueno9EXPK5cJtA4TqUEynOzYv40ZXjrCijgJocOm/HSWz6WyHYGfC+8x
oJZ2SQubmqVxt1ykOamu3qvq6UNYjz9ia6BD3kAfNgIdChRO6uKVKpnSr+4/YmstMujpiM9NpKjw
QqgxqFW41KKvas5GJ4nBFMCqOAkdhWj8GNNdn2O5QBJPI6UUM+JPh4pc3nzmGqFymefyhbpn3r8H
4+2fPBmjkkIZK+3eZz3W2uTbLuESMwb9fYjhgKPvo0AQTadII8OygmwcDPdC+dhznsLcANT00nMa
iyzv5HxWmxeSMBeDr8hkYEcVFofMEuHaZ/bvNQCudBIpHxJQ/e22TR3iJTvvMWbyIZVcaHu9mHld
bs4EjWse7Tl+RwPA1+71UN0cvC5lqTzu5UVDoMGgw4M9EDiujDuJxG/PJSKQiQHtMCBCAmMT1qIG
CFCqzQ5RGTkXgmHzWWzi980d+uNeyn5BaDCOmuvi2tREzYOo4pYG1eWe8WSbo5JGZoJE8oRiWJur
pCN7Bb5h/MSA+aiqSLb04qQhY/RCkQlMBp/V7XLtPitWfXKcvn2dh9TGGjPYlw4b0q+4u1VmOaUO
+gMnEn55l0OyI+i6RRaCcczN8gczPga/nP3grcQqXTasdcW0fW7KJ93v6yXUwnqUdOiQBrhoa828
0DRB+bIwLECrdD9tG/6qa7GdDYnFZXEQBmf5rtCUyThEZwhqO2zwtouE+enhxt9STxovz7pkPioR
PjWqpWNzMofCCPFcfm2asgT3WQAEcRA5ES2VlP5PP7s8qgXUuKx50H7cvzIzDVdZ/hEyYNeHB55l
7UzOupgVT/pjrVnIWjR5c7zrxePLWw0iWtiZjn4pKNF91O6gn1QhRF+07tmPLj5rJ2uQL5mFBdqP
XElyL5smFv4msb1f0FKLj9X81NUuxvCzSX9IysxyfEr15JZj428r2be/0KTRAcKMLYk8SYdR5lcD
y138NxmSvyBXai8FM9W1sQU+TXIvw+5rmcZszleHF/KN2xpjOF/Ums3tr8iAlH3XtWUUXG24RZ46
tF6ryzDE2uJxZr+q/aCQNqTWjZtFW89GtxIz4zmreJr/weeS5Vn30quAQIKB6mQdtPvO9Cb3JDXV
k6AWcMF7VwKxjIKjFutINlF1eUSfewoOvq4Sw0WVFsT/xYM9lPJERD89PXp1S/8IWobzRj5AxYRR
8O0p/ePBlU0OuMRuZjT0tPtdmuw0yWadzGDTqC5Xb3RVw8/UFwfXqHlIg7kXlMR2gXkA5mh/PgQK
OqMbIrH2wy/KoLdUIA6hqTpazQSjR/iCF6snZAkXEAD4w6Kcb/yt7bdXAhU3fvlyY3Xg2GP6wYdi
iJ7flmqKg0TZ9C5J7BKMPgrAI/2SV2n1c5vsistRhrwGNBpkYVaTtCqd04iGitvRQP/EFtOCO0zM
1g508K2EN4qFfidNW9VtpAs2dxhzTPJQKX+DeM+J8Z0vDZtqMg3V1BkrtsdyDPsNUwWA31J20k2q
agHgu0ogfNMiiin18BE/o8l7bnrFIO1rPEw0CaJ5jFiSOdGcquHKd3ifGstoIYnDpUQdekAe8klO
kTEdOIgf9CvIKYGooQKu6gp8saH0dvC3Rr7+6gOeBwDlFp8w6Ih/PDpbPSMEke3D+tPcNmQzucqc
dPCBaOXNBcQ6iJA+cTid+JDOjr6Y5JXs5692fq1KdPk1/1vo6Jd1zBhA9E7lLkYTLbysg4GSlgXo
ZCcVxpaIzD3L2osppIIcbYdpMdUuMfL6PYL7ihdFZ8NNTrC+Y+w6j9WTkbem3ajANRUphefGsrTe
nx6yIV73fZLMp8O7r7oppCCq8qa+TEaYAkiq4FJWESps7ho776++avuILicf1601oUYp94ADEInn
dkypOehkdB8G+07+kyEtAMRkHT+M1UAVbIBFhrvMZbFOpPfBVt5nskC+dJ/a313d5N061T5jQHwR
ht3CVNQNsfkVW4UeFmdQ+PvTqduaYUpcCp45LERydhYGBnC8slGzGmTQ5x5FzStpPwIr5wNOcR1l
6USvsIAv3q4nOJ9Cua8eG/xKN/mWRr3VRWEqsXkQ/YfVnEOqho3xDjtibch3b4fX8ywJhP1URAuO
d4qeb+av7vQtjh2YKaaKBi/WiToYDWiLNV6Wv8IJRO5p4UAnPjXXUicUn/gQHFwf/sCedmSPy9Wg
6yYRm6JQlYW9+sFnNatoh+6b+zpTUkwRLD5eKzdEhfnRaPP9D3D3M2tHWeBdmYGHxBG3JvQA21PN
DyzMwe+qtWRDFdjptxnbLu7NvWRcv+woW0fZnE4f8z9dlG4OXqGDRIjPCxWLiMVQxscL7GYI7D3B
yqJQgIbiYb5xynJpzxeyoTNpaPm+7EyBmUpIeSw93ErxWwf+atDyhbtA7QlKc4OJUyL2c9J6qPb7
DfeR+WKRPDlJjDIJxi/GGUe/8dW8vnC03s2LjDDbH5Q1Q0Q+abrdDQksWgBhHMn3UcXf1WXT62Mk
gRDB8xzSwxzQIggQ97YOWxmmWedCev+HnsHgDhOnwqDaylTK5lyLc/OubZvBoaArI+lWCaHSPo4B
SfRChAgDyuqGnsE0LuqJas31McS5qPvlyW7gB80EeZ5fuI1OBXb8od3BcNyTRtFP/OIIP5KxLkhS
oftBxIYlx+eP2Pb/0JqYr4JYcSAFVjqe3fPEI19QMR4Cg0pPs6eqfz278QzxRZkcqFpDwJKbDra3
X1wV7nx52G6aSJ651ajGfPRVdSyH6Y+FmKg/i+BiH9eAOe2UlqUC54q8fRdCHeGk6hZt/Rl1gp6u
1watAWPghuA6y/AnjD85dMQ0fmyRiTxA1kcW1hWPQEm2VtL3uW6d2yhCsW48GBllipIYBV6nLeLA
SJSYuhM14/0bxO8KCclVuYiore/o31RYfBm6XWGgMwNh9VDK6eWr3r9WxDen1T0lWgT+GvH1w37O
8IkzQKxWuO5Jy/RIDy20myixtcnUBozhhoKQ1csN6IXwkmI1xiy/eU0nFc+lt3NXJP5M0ujCjqpP
mDvRGR+MLgLIp69EiDPvKRE9vTQE3MdwDD8T2v4//evzQfOzrYekFFdlgcb5m9z1M9vnnGtNsLts
ayuMreDzc9Lme8CTPbfGclZBQviHcihNd83NnKNH75MuZXpVfg2BFuWSSTPqNrPRZCwrj9C6RrJM
psbSgTPngNABA2OrMGJuHK3rg0SF4xKfCs3LgJe66gMF8MQ5BzkISKW6yY8Q5hovD+rgmNmTbptC
h3OhJKKoIEflvOLzdnuFdNHlWMWRJfKxz5TvPO+TuSD48f07xKWPCUeDOuvOiWLZTggycNdh85UO
4v1pEbL/BD+JV8/VmKVsV61ErZZSIxOau6n9e37KKrNZ45zOmGSFsyuQeJgRoDI0oSOOnz7bHycp
BdrGOy458BWyTdXkkfANbWZQ/uQlTlJbn64BVHYS9RAJ/WoqHkl5VV1v7aVfZ7KJLZB4ON6Pg5K6
GRdUVv/uQDurGVSa1jI1HiErSlfB0obd+LJJADBoHeby003+P70bEofbgvCINo1K07DF5OjeZ1wV
Txb6LTFmzs+G09YAH3xdSXizvHMiBhsShusujCdg1mWz9+wiHhyQF6FRpncX3Iz10c1C5mlkeyaH
6feinRwNn6SLx8yQmktfDusMuGLBfecpa+BK7TzbmtmzYhoKAhs9hR1OV5lfePDTGWVfiPIrv8Vc
l9jogdbLFL75Y/BmfUEml+UB7VmBrAgtN3bJX1nWxeidFRRQ8+xZQbULBjZBjCqxKu9b8qPMSA41
nJmWdWfm/v8SFZC3b8r8w8crP78o0cg/fl+YSmunqXCtROk6F72fsZJk07mNYTmcsb06IoBJo7MS
t1gnjsYPt8FFBbFi6j2deyjZvbc/563gU3AsM2iiEW6UWMVq7JNpnTsl/3t1BiIxhEIQJb9y+tyl
HTi+XeiUNC3ODeMFQ75B7AU26CZEeopnSFtxhBA5vDhUxgOw1nXG2GZCwZNQ7mFg37p6JdRWqhwE
6KxEPA8ABZkw0MDvb1CHZuSDFDxnw6+oORmfJ62mNdFn2MzYCDDqq8VMl75hrkcIjeVlR19qmBIL
tKcc0K3pRuV2Mh4f+WBMoC4pypoueh03qf+g1PWDlJo9nSJjOjxgoJMGAbOsqAaTKbi9v//DfdnX
HqXQJoLWPOrX9ajN5RQONXyGtBcTCugKOst/ERijmMhJ+JBRURaPexx1GFhGxJqCAaN2ynpqNVlF
NmQq8lG83C1o+k8DTrBrHXO+3z0okEQc9JvZhfayV0NefZHe0Sy4SOUhvy8GBw3GkT3+YcRL9YEz
Tc+F/FrJH9ElrlubS73BaWrhGEHZkHmIdxUsYEgs0WIM7y6F38xk6f57++byaaDnGDe6WYwpfogi
xxWnqPCqQ0FIKbyMkJ80vSM5+wI9NqOoLrCEhbFLofIngzKK7Wj+3Znrt6VgoqNPgtaCBIYDM7bD
P6nWOLrlHtft8UBEvhHo0wEm3xzO6V58TgFdoRlkMKb/OAK/NTa6zxEQMqTlwUoen6p23lwhyaHN
7R5zePHUOlDAme/G9T8y1oxVqrTvWkqm1nj2YcLjtAPQBEHGjT3Bj+CLo/E/K9mP3L9SeGmo7BAS
0garLkwZ45SxxTaCSf9O/GYWGxGoJFVz0erY+UlyCcPr44qJ7w0ILO3XFIQM/ejQ9j9TFeTMbRmJ
f9WwqAMXR7JkTk4y/AfdNwx9MijFW34ANIAxCztZBwIkj/XijeMQ5p8CRFyTCCe8i+esvDXmx7eC
I6d7S+CwARmw3Oe5AygjACEbbuU8HTrmHYnjv2GCMb+8ZSrvjrmNedl7hXiQOcwlmsB3CfJ0KKmr
EtFfcnl+tLlkPHp2e25HY+gzMak3FqMjqhZgzGgL8JFvJ1rml/TotrQLClnm9A4rtfcstVGCj9XS
/xOTYbHGRWtuVG8rQ8KjcfGse2lY44zqSwWlOJF5RfYxJXXK3pEuLc674IyQ6uQ/wwWzSCEF6HaA
HzOAWEfKys91vhmNGD9HoWOVoviWNlK8dH4EmHAgiL0R1aH78vBOMT8d2YqirRqgRKn0qOovXYgF
5y+G1k8BDgwpyh4lnuIUT/1iZ9wgbzsHbV8RhiEnZlGy00fdFGtfLtfSOsP9jgdAcIqsNsmjtJYU
JFQwCnsiUht/Ha4PfdIpiDspw2TRh/k3r5ycXItciUZ0gch95pj7zlGWPGnx/+/uk3ROkQXaINZk
1v/ygbV9VbGYksW3yYYRQJToXYvxfryKWDBbr3AnqrNVyJoOMTHXBd/zKFyvhgqQb9oJE5aOrmif
FGVC5uUg+V3chw8zmflLgr9IcFWJ7eaCYInnreisjK5tijwGu2w6FUI+2Q+6dGzbUvT2+q+9e+5P
TyPN8o/u82CX4IgRADetWELnOO/If1SUBrXvHIvuEIJvJh+gsCfFPQ89LkuJceYuUc0E+kSaZ0UQ
3udbpYDgqZ4sJuO8Yb7K6iqBvlpy30kq1SvG31JJjbfE7gzS8i/+kq4KSDBE10ZNoFBQf5mG1vEy
Jj1r3xd/bHvN3kXV28PsgcOB+eh0GKk4Xb4qY7RLQBiXUg2kW+OvR+8mu+Mi5L2iE12gTo6AfHG7
vnQjvOF6Kd1YsjMbe3ns5NyFpDbay4ZVfGjuUbQdWX2kv5OdB92vvaryfnuF2DSHIu7To4K1TDdt
SOykiuggPkGelz3KNfHXpjaRBVsFKlVUHHR0mZRxurDcwOUMygdhd0mdKR3OrMATC8Gc0Ba3M3mc
kZaqovyKJbkyE3cc2+zacQs9/+FOeOjSKzEk0TTFPs2nNRgnVOshfY9TJMym41AnA7o2vdr6Btlo
6gr5QTjhI7x4FVrEEM2cUNM+hrhDUr3M6TRdRiP5ivG2hpxNJS9enOcYTsxXL0THEJ4VBB/NSIKB
OVCDBoQq8gCtiJobs5vdWmxAOukNwJfNFgHsLjyawM2CNPTS5W6xEBz+aftg9azDz35LCaCcmQHU
ouW7L9vzrPIGHNtjSNaeIxqSpJXxfIYKyzh2a56NOjtnZ2WFiOIQQ9AxRZ5Zadk9N3ot8T7bXrWj
0RHVYs+MQ5A5IebSY3jXJ13ESHXBeXQExsjOPmYiHDvxiM1zWWfY7pT88jKXTVQQRXASzrit2Yxn
0EtZz/sd07qGPwZr8gA9hADjauexSD01zjTIIjOik7JTOzBh2kY9jrZtE8DPt8gq3NOSrizz0OpQ
un5Qsl3sIsxYIwf6w0aUtVdZUlOg2kG0BRCXZIAyLAz1ZQVWGcc0E5Ztv/su6N5gjC0DQdMCj302
1nXxGxND6I3O/h9SIRr0gPV31iimcLmlf6RElnc4Z/nNFIv6aBt/3l9Qsiy10HHK/YOL3KkCSXpJ
fAzMqaCCFq+KOPEa1ZS+2Xyi2ErMamZr2JILDlf0vOoamfUduiiAE2Wc+6ukdSjF2YxMdVulfz88
E4kyJ83SzhZROJ1QC3XKf03LLbtI7ElXKfAwi3m9KJinXM3lgsH6au8gvF3aoCl7a+aQkAwn4P1E
5zqzhYKcI4h1+Za+/MZz1sTxJwZ4EXI2rreQYiBVzgCrYm/cubm4hB6QVvofJNreA6ZfeVxEZkvf
HlSkps+mNnh7TBwg/TCsXP7D5ss5uXnjBJTQXT16DljrrbAnuhpErDfiix7Nk4rplpG0yQk1c3CH
Aj7OYT8M4ibEyfYnUfF9Ufb0rAaMPo+Yz3vdK5a5m22SHJ6/RofIGUO+jcir6zxZbm7DvtzhsJ/G
FXgKrxnYC3U6VmYwE+lJGhQCWS+VO/lwbehUYKFHYVnZq6FPKqujuID4bHWZuWIzXlzdF/rK6WwL
rcPyEVEdY4N3qXOBLTV/5uYgIYCmwYkSMcdxCL9eR7ZkYx/VoJWkrFk2tL22ikfWBHpQq64I5Rpm
leDuL2nVc+/e8oslbseRHaqIO/jvLvtabF/czWtndLo1ozUUW3Rjz3aTpe84c2FudW7bYYTuCi82
phi0hJFmgp6f2IoYGijQoyAJPpCiajOZIsDNXQW63u5j11ODwdNMIJlgPUMAav9mjOO0zQLg5uxj
is/PHWzC2kCBqSaKqGTAy8JpxCZeC3mcGVuoJNo5sOCU8t4xivUfuaiCxq1hu2PlMcRbBurOVfCu
SXW5Q02swDjd+jX9vq4iVo5Q2xX0YImZNy5DXKiyS8vh8n+BEWe8WPuTgrKP5dJBDbUnru3Gdfbq
ugSHh8dPVdPxdipI22t4vdWNqR7v2FRAGncGD2Vcf57hfw8ySIy+zisBRN3jZOE8lb+8oXQcevmo
SRDKfrE2lWzbkDdsYPuRR/scTnIv0gxPOmMwxK0pezAq2K2hw0xBITFv2mTHhtA5xJuF8bNszcfb
X5lOLvTM1PwNMOXso0GLHt8WLI027HebB1yxx9kgJuZzLj9swXOx5dwNW/U/ieqiJYjlBIRDNE2H
+eASNjLnPiuLH+sPBpvM0emXNo51T5XDZhWAo2TkVZnW2MjNGC4M34E20MI8LFbwgutXPYTw3Bog
YD+qdCGvr0Lc/wScyU/nBDLFseCs5WHnnSLOGv+s7nEOp7hEj9K81UqJqal0Hr0ttpq1tBZjFJNc
ZblMVtfcvN7TZQahR1lFBFEDCYB0asJk0A7GpoxaZcSdHZsZZzD+O6BGS9vITcgMW0Dym+8s6oki
EoavWiC9vDKrAthrMu2P4VifOm5Lhfot+XoM4vJpqwh+1JW/B/EjinLiYtCLJqdmEoyhEBz3F0MU
A7toeLXgBGAfhZZmA1RdwpyeBBdp9VXQQf49YlmyQr9SqDg+EpyNf3/G3dcGEtS5W31Y8IA2BViT
foLx7hT5PvLt+wwopag7NcSYePFqFsKkrk93nONK/d8u4we1dRQt5Ig+598OBEePVCz0uv6xbiQP
8+VFThNnpAvTevD4JMynPvV3qsHXRsaOmb5BgSwc7iQqn2UuN81sPtA2GcN5LtlBF2GqTz7ft9QX
ESjzkyQYH5v8E8rSvzGmqhcoRA0rENHXrsLXYzgyPFIw5T5/BCJqnWByhJ2w7944Cyf/xKE8YhUI
PYHuyctUwxPQ3O9JTe5n1OKLpUKkPo3ubIJUc+c3tZv/ips/X4baankfXk4hLtlkGGUA6ElNyaoz
xGwFnUawWwENh/wyLcqb8s2Fzm1NCjZ+n83SRywLUCA02ox76tYc2xf2T5LwPTUHdmvGEVqNoZvr
SgUV5QXuWL3kQ5jS88QzAr3r+9cHCxH4R+h8iLbNNhJDGiLaMDhwp/LE0Y9kPJ9T8wOZQGTSlklg
p9QVk4pSnLlYzqalWOhgRLRH4mn0tiZSMVZuY8A82gZBT6oIagGN8UsA8qUbkAY++38+sv0n1DIz
Z6EuQ8vG4lpJtnfod2o/cEKXnHZ8rcig8m7+dEBh6AYcMvxUqMQJuC6w1n8be8VxKYX4ku6z0nw1
XDeIsTBr6Wguv+7wQqSklucxRKkT5ivOkltvFia3NQcSPEU2Ct0Nj4fxg/Tx1mMbIrQCh+JXntFp
IA8PhXRYHE4NdP7DOsfCC1mh3epDXd64HhbEvKelI+bLsM++X9mcy/R8Y3DKHEKyZ9pHoGbREJ03
dJH5Ml0JBfBQYfbgkCxZSDtd22LyQcikGjxrOvzm1EjT/GznwORN4MMWVVgxX5A0O1biCPqyiXJw
iL3XAttdD7L49l2ADvXpQgzZMEFsShgi2k7ql/EV+IVsw7nHH+snN0A73sWN/WV/eMVN4rxwkvOD
0p5vFWLjsGllEd+0wxuWEyAgOtCeRvwL/zXuFTDDRehgMsHOVtdMJ+fOrZ42SLKM+9D/o7sbAe37
HSXvg1LG86CjJ54YUfC31EhXCXH+3RWXdgBQcPNmQC5MzKjBIg9X1zObBC3mjRtz8HYIMscB1C50
qbwSq6JNYtXg6EBfj3t0THp0xZXFeEAJtS7aGYge3GhZzqrg2Nq0rAITMUGHExGfILctJuqPfpHY
z3Awl/LuJzpu4Wvwr3eOsiNViv3dxuhxjiGwzMeKBrAsQRfBxf9Cqm1cJzvT+J/gFQkImRyw0EjM
jIiK3eQceG2tZIeq84B+DMF6FVjfIdsN5FgMq3fevT8/5ueQD4RFAFBMPwB4X7znbL6PLCymphYa
viflqRbNNUjCjhTHhwyEJOP+qcMWJHPRTUzikPyZ2posLhv++cGiMIuLm7vscFi04YfZjeCyT8kF
A4kvP06Ufq9Sbm9z/x5mTahhoxskFan4MTfuaaRW6IIND7WttMW8JHnhyZUbxC0xbZ1DvjFiyzel
/yJKLhvS0ot4WrXrVptRsskRPOn85+fmhEfnb67qclRUbqypE5tN/SfNiHsf0KOh7h1Tp/F6Tcpp
r249l/4RXetRll7vE3uUAhEjhiNXmiG/qYHXduWX+BOKdH6ixZNFYORolR+XNPR6kuQGyPDnVeJ8
kYyaaprKzU8swEaK+zBHJYTjo1djoENhLWGOOHydUtliJn/Kxyrb6Tu/dXeAqI9ziYJIQ/xWiAKw
vVUIy0WWjtVDBswORqFeVAqBAQMAjwt12zADCoBfRTjxU1ypkkjFwjP1jM2+SOfVQCsmufwqUb67
OBCRFiA8rrZM4zs4NaOJtT4qURfb1XuZEIcZ2QgUUekk83SygujaT/IJqY9CV6TNwfiut8LFOiTZ
jqXVmO3sVTXnWko7RCH2ABC2l5fE9HDUvoPG+hfuNp+FPjrmA08Xmh4GPD6iPAKZTIpyCTrH+RmV
mhxUzZA/q1nSznfILFZbPjlpgURu8Ws2ODaGL8cKJfZEycP89WAatASq0Mu4nYF9Tz1oNsqrapG6
fZ9Oyb9onXG6gtZjAKkybnrbGlYTu/raOk8UIbXLA1k5v2mS+R3lDrAzw9umdwddM5ZGVh75urnA
g1U46cMCCYpfiYy/KdoeJadlJkf8BX9DC2+Krj2gTcg40EL5bHrHpdSoo032mkS379K3IL26KYZW
LDpY4FYFWq65cRaxKVpxOCrMyZhZ5cPNAU1KqljIOAr0EjSFqwe2oSZ2izwTKtXKGCeLm0YSHqOL
0Co0VrTxrCGV9mljyRSYN46WFDm1r/FRR+i2Vwn40kcws1OyRvhYjg5kMRO7aKO3MP8DjG3kqdSG
q3poMnFxfsdrHZuKMgrV+BeWXQ0KE6zb2qd408iWzGNOJppCUeU48KJ1q+HW3GpvFchH0ERX5cZ9
Dp4gMaX14Zbot5XMYc/vpEysdoTorzpGCRmLAcVKZBVbNc/qJJsVb26FR2fcrWF624qM35OQM8Ru
/718vPyGD/iEjIegyzj+av5T1GErLlTZd7I4trDPi0R8bzeY8uYe+Mdqbdm6k+iXYKKG/xOYlYjS
eBqyXavejFE5otR0iiEIw4jOj4fo4/8AULw1bXnMkVSu8ah5+S1/MFhSwih1gVVHRZRoN1TNG0ft
J2Jci32K8MHFKjxZRG1fx6MGUFjGbDF49rjt5kLbG4pOhzmd0xuFPqm72B1W8RCAIBfTn1fK9IKm
FlEFRFoTjlKCERFf0G6MMRtV6AGEC0nuToXdyAqqaJv2BqMeH//rCrefzC0DBNVpkHNl+WrTmJ3p
xKiRL9lpgYa5pqEFr1HU/fmNYoKDwyFlqoEEiTZTDDf6J7lvfOFmbULbb4LEZ2+gypnySsvcnayV
czOaVn1tes8ad+3PYN6zmjqFzGXBt7HFIzB/ONsikbImwpTD+ZklEl0XGU/oES+xkzNGAYEgK5iS
9JHEPzLmrKWvw9ttrtKrSSqrSNrKl8dxCZaqqPF0tP5IaQ7Rec/iMcl5V4p3HrikqXAxYkIHxTdj
vdNJ8CL3ebcFibTRSvjG64o5HDbdMb0WOvGgQvenAae0l9B8VJnuBGc4kpk5aZzHmBHf4UFgIs7+
85rVA79lPQMw8q6jKEoTBImEBa7fDUSwKPyFb7bwyyYckLQMQs5reKDNALSjonCreCiChy2dNrxe
A42CErABv8pu9ddUamwrvmNjsV925wj8gVxKKJ+OkclmYE+HA+OWzeB6We0BJ46qluXb+L5U9O5W
OIow61fwbJs1IfzpyX+K1UtBBuBebrIKyZQy41TaRH72Zcn8XoE03wbzlBi5EtwicYhCU7/X1QEH
tZ2+5cv3O+Qr+9aH5JxbJ2qaCaGXVbZH0MMX4E0XrrmwkKxEEv5WqmEgMRw2DKAhksSbspskQ3aa
8SPEqRbjCrBLLdA3apmJPFu3dDLkvGGi2F6r/aPNuouUQrcmAIIZ3motYqjzwKYNbcDo99GCXt++
/H2CnP35Scvbf0Wb6ZUVgGYn/AAh2miWB4V5iZurktWMPkVovFvgaBm4Z+WF+1aSN3cR/0Fu7iD2
kN6X13rsf7lbu1w7yQcCro+MV5UGeDAauqdLGjfXZSzeHUR2yMxrj03j1ugL3DAeVeOxFb/kRUXk
kPlwfa+gVxXRVg0KultQ7DqtC2qpU7ALySf6ae6kh7E/KBW5Q37iWFovEUbuNftvF47sQL1lULox
4QDgqDLTKPHqXxFtF1lEw7vkmPLrcQcYWO6ln+WxzZo1Dl5WuUx2XfHYOjoaOwwfuRD1xILAiW/v
PPCU1OgAg73gUz2mVCUn+d8vBCk+rlwtzWwDk9jF3EZ8Vmi4FO+18tAjeOk5mFyRu2pSXA4k3d7Y
rXKrDqb10sdltoAH1OT4e0toebNdSbOHjZj4Pc2VlVoObBOmrKzEp3pT2YXvYHqpp9jRMbhjJJIO
q6h0k4dZED+GtDRIwUVFLf3Mlefwbz4oVjPmRH02lcDlY0vfNi6nU/r0eF+phmzfNmGso2WYMf7h
wmeeTcoSMKejBkD3NQH0lQwtTUk2B6bTFuFxS3IiFA6n
`pragma protect end_protected
