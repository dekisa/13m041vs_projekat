// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:40:57 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BpY4hXZK4Y9c0gGeyQ6d8RMcUyjHqgU2Bxktls3p74/Ief08eyBE+CWn9ai7QdKQ
yTB1QloGbJDEXykPkkmgFjKbqTYvY3lq2/Y2cCYbc6CRv/p5MEWajm9LjDtQDPCE
MRqtzuneO4qW3kpUlFydZ9JK4r9Vuftcs3s1s21HYvY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36128)
L0iIOGPS6JgIGGCgoK6czIzO1ili1b1mc9SsaWYqxdsd91ot8zFX6b+xmtRL5rgI
DxIaKqTN/VV8wXJTe9lNQsZoe/XRBppo5Tdul+Ba67s+XBCjtsBNgtsXTDdoPmH/
uY+z850zNNpADFeI1WEEVsMcc08gj1CEAbHgCiJxKBA4/cI9YQ+CFYkmahfhgqcj
qKOk2dglR1E16jLhsFLuMxiKEePcS2jiALoZexBD031W6r74uPAViEGlRVIi3UGI
Hvbotvnjn+1TTBLgEz3RxAA+BPiambN8YifD/EEK1ngmJTcR41cOSJLOz8UqBWPU
2xWUnepe6/f+HKPd34KeZuvYe8eVEPu38HRFEo4GJO5hsAxtrxK0JeGgnjIuZ/rS
6ZOciXS2gjArQ0Mlifk5mOcO0cFby03v/u/AC3ctCkRuUzP/un/oAYaAGVdkaDsh
6xNembBJFPD9y90b/eJ9Hw5RuWRT7zTVwficX/THwj+Gf04PlcbO/JxAyvi8lHzD
CObuVcyES15PxCY/+EkbxKLHgJyz80TgMrjFBHyl4xhWcQslRKu/Oszo6CYULiy1
MUIYnVULqaQ54Egwrk7zRazZgkdY7RGyytjvRTeavDPvzKFI4OQqUXmKca8F5foW
juz+OWOGD/T2JQY0ysZHKIQzEfUBtcAQ28N2Sj3Y04RQDnYLJckZkjBBfUArrW1Q
NLVAnPtxxqEp9GV54bvhlKmvRLnlvLQGFFz1RcWLIFhv98FEyZZt14Gha+n16PGh
d3EYd5te1lZQDAMYf6mqdWGjY26PKFq9ySNtoB6EQ5mqTj5tO4QUgJJmx41vjpHP
Lg5eoH272yZdYvnxSMG0qbYlo1pIf35oAp6spV0yYOIHiFUixcVWFL8TYJwOgx4S
zlEwSv4uIT9AfkGN3HHii9Ww4TLlurDRQ3SCSJaux0OSsjaslpabv1yoEAKOkBn4
eTiKZhkFLo1IBp+PQwaoJiFwNhVhLCnsP+cl3RXDVZZog7Ii28QGqPr0KRZdaqIM
kEvZchc+5nQCRsU/JWK+SLsJZ8p/FSSk3+vRfGV3MtHVRgSkQk3HdlpYdlrUiAyR
2Ejj2LpmssMGJe17tUkKsqujZnpAftdiWuO1nweBu9pjHPl6wqDzxbj1n8s6I/9b
FdLVvhK3osqPCJEpxYE6WRxgDlWysc0CH7PLAyLQKJWQgE62wG+RJb3ZyqsmeBiD
22kq0MRCpR6xXeI8TlsmrceoV+r4TSSzJ3vgQad+U1TVviO0VQjig61ramQf5yrk
4VALBs6h9PM0QBuop7QSdFQKTMwWtZJzAhoQTp3vLZpKPrA3jIkhov+APANjcSvc
JZ63YMn675lwXlSDs+NtuGNeanFFisfHVprpMA2SHQrahGG4SylIkEnqUsRO1TLJ
UF3p0j5ZwsH8utRrSV8GflIswLa3FXYhHbCD0eRksiXZrFKhjaMKiNHrwnGLHTri
aDnGZe3ry+gD/YPgQTgCaD46hTnWxw75Zl5kt1oYA5R3i73t7vJ3KsxRQjAHWa8R
rJ56omgTsHUGW+YU1r+FTQFxfYXBvZ474iRkIOYqHrPfOZmG+nTJQHeae3zHGm46
5UHiAMsRycIFBaXv0VUTVgJEy4CFrKg7UkqfrH/lqqJqRKgFSXDCOez/r4IAxf5Y
ST3OUKTAXwmlkgGhTUP+c2jKLMFkT1/BdZ0CaWDdeJxARlEzOuBriNDIMospju91
Plk4nwZwUL57+OqK6HQvaiVVghax8xZxrvnguEy5MPH8dPz5RXVQBhniEDF7O998
b0qLfuOu65AASGJOqGODFsH7glJeElbPT/YE+UjP/F7fykXDgh0BecznyaQKNUxv
NJpNewsdDJ8Ax8GlS+6LPnEZtzydl7v7cSU05I9zmLU8+EMpEhncG5D/ZLk28eov
3ol7dShih8GvUn2yaC8xhFmHvwLNwRh9fxpwfIqvB/qMFs5VhqLRcl0O03Xcmbsf
8hPVX9DGV3jBR8UY1dlqKVRIayYaz4KGxMGD2uaxEomQ3XtQyv/y5tLh6MWaizGV
qlObkZ4LKYBpCmqgqXEgc5tK0wP9AYyBt5hHSQ+hxW6ByVkv+WbFU/sI2eXnU0oT
KVVLoAh44+bvRDGElFwCvuvji/jhmQkJR7TuafYcLF+/PX1ZXftyjcHVI+o2UyGB
mWyERTmYjuHnLMyxH+ZtNetH/WEVcAc0XFCENhtfjFh7h5X12spClszDlZStbIfU
og0oR3EB5lexGOGqMs6Hp9HSg9hHFhhrbltQJdWgDD+7clRgBumyCLk3sSSGGQeh
/0v3jXmAwE7LHvFWyFA1NKp+H0GbTZhS1LkRzBkGbcdLhN72tcse2AXqDvzcECvb
Iu9MFJTf21ye0eN/urWv4Yf9AVVvaeRcgiG/Zdno/RThM767COrAY/E0Yfo+Myr5
/zPni7ySi6UnYkfEwC+uPgLc2Ay2sj2vn3ZoqVt2CDQloEVJEWop6nXrMTHaitjj
UcknByLQ4eOEgHkDiIaguV10v0Iqy28bt3PyCi3f/3ug1mK6A0Z4a0uVGidgb3e6
PjXBykt0rj1l1PzjYu+cmSbY2POUBpxcR05pgogxb7VzfopulDuW8w46B5Prc9FR
h2yOZPYr1g8AP7TWcXvELuzVQRBLIjpRp45AfRuQyVz8LI8VbN/U/wUb3bsM3SgO
owfIbObjEL/RckcIdjEGZT6OfqYrsLtyV3g66DbUBanQsYgv6kbUYxgMxx75B7jh
Hs5p6iMl0rebsGUS4cdkwtHp+bc8ET3NRs7SJQcQmZBnGu1XouKJkKm9AlYcVfJ/
CqxGv7wDLA0eWSVmD++ee+hwNHSm8aMlodyH9Fcm+IhDcLhfIJwJBg5mDw8XzwbN
bCsoG9w4wHOqnnH0cteeC0Msujwr1H1isvXzbmgn0nnSpjhyEPwidQ0HXeJSQrUj
HBBTuE0ig6L6RckdciDl9Uaam1el68oH9MIM5Iv/WQXvYIbx9nWzuY4Rt1NwvoG6
XHufE7OOkC5a4xnCE7qFaFIEx/+Yol3StNzxtQ+s9YFetBsJtHH3Pd3F3lNKo4bF
YiENQLRbwh+diV3L55bvPyvxkb9QdX9fbV8SKnOL8WU2Fe1T4V+cd1iQXCT/BZja
jKwfH9dZkxLKYnFLMfCvzQAOvPinPoz3QLeK/oTc6D9prWND2esD7D3rt/InqU6O
1LkAIj67oQ7d9TdR+b2ngAhUXTfcfFIlhNkBwsGww9u51GeCfBaLzPMhp7ox8rL6
rBw740gXsk6O/SFjgoVXrH7PNlrgEpl5clJGuO8JaLHMSa2/hXkZR57hIRjTZhTL
1PDvFACdrMt8vklGBGpKVrIMgs4pb+W2yFwIpZIOmjpRLS/iN88RWV1TDpIa2g7M
bVJct4MAKicT/Wu5GDtUYDVr3/2wiFQtTuB50MrHQc7YZnoHsH1uctO13d3Y0bfD
vnnEhMRc9Lx8ZsY7b0OnP3qjb8CHh02kPcwfEB1mmID+vPv6P2hzfPBp5NwL63Vh
yo3IvSFiu91NgC1TuA8Ji8RoFUFUj61pCx/RL+ViLJpIjyvXrIpFLevXc2CcDomB
aTXlbVT8JyhTmhMbZEX4rX4GhqKj9kP27VKH3GhBuEdE3uN78y0Sd7UC1d4tR7Dv
IJDYAJQ5NGabxj7j6c3NLs3rDGsBPQLWOBG/PusyUnEzrmr1msMFDy9k+6DQ7Avy
76PjzIz90pStBrWbwBFlni3zsjaYfTFL1qCaKpqb3z8brv7D1hlKpg7oRFmJ1qFA
1/QLpLF1axKqvHLQQCIAY6TCcI8m37J/2Kl3cqMSvo2LK2vfQP6Lkf/5ZSBOqHqJ
ZnHREF+/UpnHOewRKVs+idlqn4EC0EmJtO3XMsyMzmKVyxM3CkoMzxAdNgqlqszX
Oa06wjIMzaVTOK62Owc+8Kk22N5qYDKcPG+ltswTU+ORCXiUlww9B0MxoB1Mlm5k
GPipTf9tt7ieYmTjoznZ+UyG8RUN2nUky6o+TiQm/AJjh+4QZM1G1fH2iVfcZ0P6
/fq+/iseg9gxLX0FJ3aSAcGeG+7yYwjdkE2W1vfS7EONCxMPoIOBcsxWo4irplsQ
pq1USw6p8pv4yr12ggssluqcEHk3iWfYOOjQ6sZe+/ejFEs9FbFsMglzeDeeAhYH
BfHQ4S5IDuJ8/r/QTsDUVn6XRAGNeEU87ah18q8b8RFzQYXvuZIxntaE4vUu6NgI
a/BCre5lLA6Z+s7CGkBXGuac6d51bfUJ3mqkzyMPIbIq0t0Tr0eZ6NGpKDtdAbZJ
6PluTABNrg9cUrvbuvDubBEbgjIjNGMlNBEMUJOywxdGRY+SWoV4ViojDtEmcXWK
zhK619yefMBCIxtZm3Q4y+c2k+XR9DFY939Y9YUcvdRCirM711hyCLqtiHgHS2f7
ROHiOlGG/lXpFHLSN68+R+fXiVqHer7z84cWlSXW88QgIXpLkY7Pr2j0qdFOlipe
PTVdCNvC9nF1J9jf3tiS7spZRGvb6mOZj9r4dtpaQGKPA4MIX82r42SR7/6UyE/z
sf+c55qDx/fL5M+JqukBCpdg8E/NxFuhjRzQPg8Wb/8LPMitAf8Z+/vTwXnl35YK
W5lK/iurA1RhHlcm6RKiw/1MB5M+WfV44HZKMfuzX/e1yTCH2wPJfqxQkpVP8b2c
jn+w7Kr751e5ojmzdhsYIU0iD053h6siQiVvfiPJYAGyoTuVkRMUI5ZUicSym1ta
CzJrHBnrICw1HygGaj1SOkNxjvRbtkA5cIFFmMvALFJacPzqy52Epgjl7tv/Jos1
GONEc+CfhQ+2JvN7LSpFmfGkM6NCnLLPAVyFFpqO+05O3zZQQINrs7Vri05mA7e9
zvr7hup5KqMr0+UoLcmgWwjjBdJwA/bA2Ok2ahv5Fu4MMwcGDJJZc0vYHtIVbDqd
DvWMD1duVjuaXlq+bskxfGGE5Seb8ssmvv7sF9pdMct8nQSRbb8At9Q7HgZ99e3u
LXeedLX0a+PBxI2tVkn8aASNfM3jVukpkpNVW6zxO6QSN+1KPx0cD28PXYcYYXdz
VOL9ic20bxn/3IcrJG8h7Dm+gWJ0UL283V629w/wuEOyatxvTdS6J3y3naNICv+E
vQM0xdaYo+BdTeWy75dBkI89uu32oXmY5SzV7NWd2tYLNuPa8mTcJOYsz13TApS1
leJcFiJxVJrwXP6Msczg6DyS5G+LxsJgg0UpAtjcyCCN16F7RnsNUJ25NqEBATUn
QgkXPhY1/qZCs4d8S0eaxKJMiorWUyypSLI5eDWTvwWd5R5wmH95BMPJBlKip0Vi
wYuZkBTl6sYyYSOZ/Eb9XTzvNt3LTW6twU9KlfXAQ2N3ICXTe39h0YE7nuckp4SB
P7ADGOF29f1wotHhZrpWyqXzmKrgLUUVTHV8EH/hk9KuykNV36awmycCHQXbH7Yw
hrxqRZ2maWb3NQTTFpMbg7abxJJw2XbWv/ksf8evKgRC1J16sV+z7uiH+kEVHKjN
Dy+RGYfwEUGBS9XtQiIDhglmUwME616VFYrsBojSHVV5BklV0YGqi/cK7mPyk/3v
VRv7aYhngXfk9RJAX9z7LCZ4RXT4XjslnTaAhGyERHS/ZasSw7VPqs1gvTqx/PGN
o4DsqExDSDs9Uxww7n57AFP5XVu+Bu1CYRQeeZ5/bPL7re2nP8lcsc0dkZbvAK1i
AbLJ4YwbW+NsFht/vSwa2xhwu+JvdDfU/u+FEVemz8llmvLqJjBtmwFztFPEBBVI
pDU0L9agsZvMs9p7yBjxPzzOBrHKMJaasLaERvuOIixJgh7EF4uLbFxVmVgLgefg
jSIdudWSH5BqzMAowa4pbF/2xN9Nx6y0yhaD9SRLKDsg42EMrl2Zw0ItDtQKD62c
yJZPW1WGuT4RRH6WOhkgpDw7wWysY2o22IxvoDMzmSfOuTxc4De2VbAxUPQ/dWNf
EZlrPBwz9LK9QTjwNSgXE15boo7CXao3X+AGI9n5PAKAwpKVie+TNMWMiHKPRvKI
uAYxTZi7q4svpTG/ReH1tQ0RGNV7453Jku3kHPXI4+nkAdfynlQySAYzl+SEEKCV
hBCX80OKeLrcj51/9hEh1D78wMx5MpQ+ZCblcCkzj4gwuLX2qprAr8qH9B62FPjg
L1mhwUJcEekMxm7l+kHtHtNcanxw0SFJ8TDN8S/tXwol7VSjhR+X+l4V2BwuG1YC
Nu05lkr9CjrziJEaQLy/0IMoyHIjynFVZ6Dpuav+lcA35qOA2qZb8SmdChfpkidk
w0pugxzoE96cC3dTBuj6nK4btU6AAYO3S5Ke4fybqFsS7N2grH6tHK9z07zMnW7T
CZ0ToXRdxEw6pt/4k/QCHCQk+EkSflIaKYVQfJe1zuipLXDWsT91+a/3gz5PFBBL
UEgSMxRToMg1Av7zPUQF9sAxM+VoGFoWzjwi7NOVJA9Fciju5bD27EC32lJVk4FR
oWvVCUScq6qKS9eSyL5pFMexqAsI9RQKfVI+RQWZIbDGCCi68Wpp8S1KfBSvTKW2
7yx+ThLlFzbiiGqnhzRb4vejzPhZEkA6tN2PCkFVK+KBttXfaylb8wqGtINZ4+w1
e1NMp7x9hhnl8oM8K0VA6SKyfEqOsVecYCnYikzWojQ600mnZCKD3wCmJt/D/+xt
c5TdptKzJ+QuS6VNoKgiu2S8Rz+tUWun8xg7W2ZQ81tc1y6gisJLbSL2YSiuNTzf
/lW33gf0DKzL2N1KbkOdf1ZKtQ0bfWbR1q2WkclmmzriTVas4qZaeDIKs1CPW+MT
SXGHcOnmSMehchsrF30FTmPXayK+Ydz+F7zx6CmZ5igxfLAWJ8wx0T6AyY6o0P58
T7E7LxFyzeLZFcakXy+w3xomZnj+JrUoXmnu7LuRTXgHsiOl1EdCh514encJBIp2
MxjtBitYBpJTlAfXzXKoh2HGHvhTJgAK8WtoKEeFcHwpCvHvfzaqhegDCqgInQm6
D+BVPPncqRJNaxUD5qMNkJH960/IBafyXnnYNWgMft8md8Y7veyrYi7h6tDfj6f7
E0iyTXFUgZzNeAWI4zFDmfD6wiRwJP2qhsd3cHlkl8dMSnLdizUH1XOfTbgWYweB
ZzyLFL8kYRFPqB/1L1kZJZe8XilDpu2e3n6PWRu/QQNrbpS1X9xZiXOrB044qVWz
Pjgoi/cA6meXhxtXxgBaCpxrps5yCxQtoENf0X04TJIfmcna9FqTKJ2MOM8qrqaL
WRU7TZGZ2Ii6GfWr6XErwttrLlZrVSrlWUs7v8ioSIxG6WHSwcHeI88c9Pe26x3N
nPn/Ui968ds1WtTsZSdDESMJDBSImoalkMzIVwd13v8ZTFxddxC31+1svkBxBEWx
vXXb62tgFkfjb0eJKGZLFixzbqV0V8R4LazfyvfTYJOl6hfPLwxFbm8VPvfzhuVI
Gax5DGhRxxTFnrrv5JN/LDHEuc4B9HPJ5V2ksJI8suA3iFA6QiC8CluzqEs0neKR
NlM8SfBXOeyDB1TPOAP2rgfPa53IIQpTFzTIPNk6+bjUbuooY+mnAOYnCKTASxKt
9ceaDuVGbzun2WcCn3MbHylE3dRpc30i/7WtngHNw1nxkOqzirrc7IZCkq/mVDM1
ZcfamWacH48SAsItDH1OcvMfaG3NWLTyldyCE9MrNslsnn4bjr6LkRgLaRAaao5H
h2Kc6jyNNCT9NcGsjub3lR64lYH9B5CnQP8tSc06a3q296895R9ckaCMq9WWVZJJ
cDilXtxNyVtMI/0b/I0VgSm17wx3Pdmhk382iHTKncd0oZCOKjprE0t4QasVYo+7
+wZVOiBnlymVJFTf6hM+AwotcH5/JMNiQS1F61pRqrv/P3MtIbXDq6JcVXoglKaf
ql+td1BDxE0c3nlYWl0wR8mHmeh5qxaedv1AAKoyZOMO+qEnCXZijNHXiq4//uyk
yLvypdL5MNaE0WZjUT9TxkHbfLG1/MqSfgJ4M5vWdJKqXFxclAXsedxDMfC8XqX/
zd+IDl3NSSv7m4nXjw0c2EuiAkNSYxOZBcSo+2UgTSkqOq5RYnINBczBA7/JKrPw
zE1r1im8yG0IfufpKeeuYJ33TfwpfOSEndtc7yT9OJzTUvkn9W8A7yJV//bYiesg
7qGFY1yFz6kf9Vu+n5/UHdU0wDCHPQlBEYRKw2KUosEA0nZpu+a6fHADJZxEPCE6
lr7A6D4/UROW0cZioLoRAxhbtDnVGwrCWqm9dlF66k28/8OBRY2A8HhHzkfbo0BS
xVkTuPK4yXAnkSe3B6ZJ3vAw51VKs1BMogqR18Je6a7R+K503umI5i0IRzMtemL/
LO+d74G4jqiwAGpI2pQmYibaL9GVB6VW4VqChqVD+N/9bM0h+I82mZ/F+Z8hFXMg
MzpijG2GgAYWERyRfNnfEcmtK8H6syqZcAbidsGney6KkXYYqfSi68DDSNIQVV85
DmlF1h7RaEKOWaZsKniIxenditxUSVfyOXAT1nx5tPFeE36+0HpXR72yLKRvKbIx
jGrcC4i+2LlVyGYnU7JJ3q6ZgjKFwJW0vSyqXWbT9hPHLVubn7bs/l46pIJ+LH6q
2yXSMEO8af7zqmY8+s96CpCIbdcFzmBBI+45Te/2VA5nR95Knx1HQ/2WQQQ68QRh
bHkdHBg/yUjA/9Zh1RSK4vo8DyAx5Tvg+102kob1OnPDZxitH0O/Qm2XoDwZJApm
vnuJzllpjNRHZsV9nVUlhXiwc41bBHdXTYRxd2i/U1+/ZfT5UTb/V5sROQuV2up0
gjTRcp/gwab2OoPaOKM8IcfCf7Bi+1McWVtMvHnxXZD4jomESjClgNSsPNsyQviW
iqtUYT/yuw3AV45YJP0STuoxjUhWL5nDI/lBdB0dI8TQ84hkQhhsINXS8dd4tvye
qJ5L0Jlnuxwzy1p+LDmJKNbk4CgPfdJV+kG0ibvwpcA4M+KSns5XSJogYpVgvo0X
Ws7A0YEaLhyloQAqzk9+P/4+vLj90nE6mYckT7CAjyzUBeR8BRnQUdplF7uYt3qZ
rwX+hcXCNvZM9eP/XeRcVpB8c918WVgtVK6iptJWBypYOudV2OCfjEy7Qjs6zuUB
4rawtjFI3zKGwvF6vf0YpyCY+yElJH1KkZaYsmeseVqPRG/kxfRVAw+RTQCWAo3g
p0OdjTxpDM49v40Es58+aY9tN1d9u8z0a1Pza2bEHFDTVl2HCeR+fwvCz8khX36f
vlPFOdym32j+sMFgfz5n1XV1XAEKdXxlT3pzVUo4QGbtSMNcrKLx2aXF+iXsBK0q
Lq7P//UVEtLUbxFpcg8fM6tlqK5RK4+guoTzq4n+7ENvYG0pMMnBuh4PhRgBwcNu
N3qr7yeMHhuSPNZOwl4m420Arqowc0ySzAAQKACo8TkZ7BFrqhSzzbw5O5XTpB7e
svAzuWxMmfDnmdRty5iuA2izQ+EySrtfFUFSXyKTYbGJlPSWt6aDV/I3cudGuu5+
6g9kyU4u62NkMuq5eM+0Z+x/274LxLmVloNum7cf8f6iqgtYSbEUNJ2heoztGC5b
XxkUkk/PEjUrTLZXdpPXPDaQayAz2XpxCxEgX0l7+s0fhEih24xmQ+aWz1F4wXTH
ldba2Hf2x/RjLn/aNmraKRdxtHJg26Hkf68EwPROkG5zsOHjcSaXPQYKGsiT1wOZ
RyliTUf34nPRFvInrSK+0DQuAIfPwV9ItDLcTFV3A8Ykrxw4tO3r6YMJaXk1mK4R
sG5sIR3VpBnncHyBP/IWGnKHWH14jcCgdk2PcShPCjhP4/xkSlTLUx+qYiT3T3tl
JeeYexHHfo+nRCb/5mhDgjfSVT1cOPxWVUqoayVPhaBIRRnb8ZFvgqfL20RiKQ+G
ciW3TtVFsW6dc1JQlclyC/qaiy8oTL+xsVT1p6D+cugxaQV3m46B26U3L3LTUyIa
vg4x4lzE1PL7Kz4aFX12RsoL3qJ8+XXxzaybZkFurW516WOunZvhUCBk27sNtC0r
t5eKEyCoZNK0iz2ppmIhPnFaO7XOfS98LPQZqv4hd50srXlSZ6XFj+qheam3cRGT
qurkQkqt8bSB2XrI0mY8WpwIfefHYLlCM3dPkV00NuUHZa2Buj9ovq1UTEPUINU0
YBUkvUSzzlRVhHiPOOD1WfR7PkQIh96V8XCxTUeA6K4X4gcoLaWFZ4wwBWgPllSu
BXbmefc7/KE077Mq0atkdQE9q14PdfeH2vX7rlm6dAY1Y2h/FtqaJH7JRiZKLYbw
iooJ5V4Cf4oFSFNEu2Z6D2uf6LrzYVyhQSzX1Jmm7+/oqRRhT9vm//0A5+ykm1AR
2h5xR8TeBzu4ENHqwLilOsVfzt90ORKjCYZ/cESgZZDguYmAQQXl4dDmoGZohaiT
N9jLNm++/L0SyCWWAJCkiHtQJBIXXAPllWgqwOTkMTPZgUAZKr0MfCieCPsh8XyE
zQ/RWGk8XTG3x65+J27GHzK7pfQUOAQ5DMX19POsUYgW+EYTYzRhz6SEKd40hack
ODcMdoS36130Wwvg1X1+q21WrGSbh50UD3kEC61mnaeY1MZHX49zK5o4LYMGBy+G
VY8bzHWYSCBSW5GuM7ckh8axFv5UfH4wPHcCUwmde4IslNFlqJbPoFJI3xkJOM/Z
cu0lyDDqtA3/oFL9MC86aOqX2VLgWCNB/UUNYDzUuhpQ0zQkeq2tXaPQ/DKTLlDk
Si6NE1IsHYKI3fJ7i+9jp415tsGI9ago657Ez1WS0FWu4dChEEh/fipmJL6Rmjzx
/B86bOYLZjTtQZ1g/SFY6eoMKH62Ebd53qZ/803GqQw84sc5RRqg73CmAGp0sjcL
+W8rC4UQXj6nfsL9L4X/htCL8uHm+7glyrpipnLWYxsuqzv0QWCiZi9UrneT2fYb
+KenKjycGpQDqukFCSeNIuxBkUiIRaKyEu1xpdGgtdzY+EGM6NIRw+i+6BQb74m0
a4Lfl8YOqYj6RCgFmD/EVXGts+cbKnbHKkm+FBtSFcOOuYh6kklKdkMp6EuuvaXj
MWj+vsg/SX0qAf+0n4HOlxONBakslN6HUq6PvaZ+KLTWY4bt6HLS/d31w0wjgSx1
HXBQsCCaKSu299UoafGS7mV89yqqV0wllnKeGKd5XYcz5iIYP3GwDy1XbrNQe4J/
YGiYIcfAudjXRJ8RchGqnqDcPFpa23uqbv+vbjPeeithfoFKvCAE0E3/CRGISuFj
Uxg8f9tCRKRQye+s0oRDB9oonw7wfMSsAAJKRM1K2MTq+bH2BvHRELjRsuLFcC0s
aElJ+ezzPxU3mTw5QlRr8s37ALifSVUgSME7YFVydGggCOfWuOFRRO/lftryAHs5
XVcl8RpOTO4rWs/Y8V1KDEn6r+VFf84LksPLNXUVNg83r8Y+xFaEwfxuoCOmFTwg
CNL9dxC06uxT83dAg9NoGt8tN+WtObKYm9Ds1xF9fTFPdFjosno3AYVgVMPttf1I
uyjy1fWluCJakWKnagOklXzhZa+TihH3p3Zw6T4gMZUS5p3AhdYcROBpfAKcdPTS
m4yx6gVGrBkGtthF/kRxwNi9wDVhLpWrW9/V/2nxRfAqV8xfBovgrH5vuDrR6csx
HaZo9fqK4ez23V6b6ChepEHzHQhQ6ruIX7+O6zS/5Qs8/KZfe/Xc2B2l6fUaNh8f
jNV106HVRthrm67ARrwG3xOMFqIHgZSGFJ3nHnetZ6mhd4OmSiFoaiw7b0LXR2B5
LSNrOaswe3WnVB2eprFUiLjkw2rIccM2AwTf1fof4re0SxfDSazn8ChUsyV+JyxH
tPj7slOEiIWamBPfLK4DX06JP88sGLu7JcGSqcKQPDhoGjoTE5dtFIsAsbSGSXB5
RTvMvtLwktHS7iR9HsX+T2ckyv5pE2aFJDzonWU60gYby+qnU2IB8F+0MGQ3+/hQ
uGEN9QK7kHO/d9PbYpXejZhtM/HNreHu9NEc/5YF+43CfDTwpCIehMxpAACi0tMY
S/4NdAVN7dE69kmsSoUygG1VdmlsJl6fPMr1QZkHbvgIO2YnwFc0Sgk0LgZ1/UbA
E3fjAdg1OBVn9+qcJN9y/L3GQGenv7LPwhj+Kru1Ac1rfnSywAF6ATwg/52ot+7r
WmGiPzx11/VlPNQyu+hIbsz66efHRuucJ3+O13opPSDMCywQDsC1YsxdY1KNOQmB
y7HxZEQ7Hf2mBNmli1NyhiPCjaamqMHQyFxbvgwxytBPkZ/Kj3mE8r6/ZIpzXuKn
iDcLp9zLiP4zYYe3ze1jehenZrUQoZNcjxjxn8CwFteSlFaW6GXJgWntRK+U3MSJ
jOhwdDu6lTUJbCEoEUN/HwWvcwNIs9JDdr/L7cNO0fgaZrkZLqSOfuwBqSLWFt0u
gnhm3reRvFTVn0POXykZ3SbWoi3veemvYBHh1mSf6Eg7mj6DHDSeonNOdMRjNZMG
2hUtSokQLgB83ZwfVsKGHopMimeXvKJYdc0eXzA0P+S46ynQMeQf3lvuEh86Tzx3
boyMaQTvQeSC6xrGL4VgKL8eJRUPIoBVmV/idvvbdgv7y/9tXNVSJzApBP6wJuhW
1qw/Clwj5RiqNeFdUAWRW3nUNxdxZq9XebRgmyHK/5BWckiEIBwnr+d7PwUSrV1+
zCdS9wO3NKijIkOQf/JmtkQ7vQGB3Bz5zdse5Gm2gbCplidR1X1BQSLz7C6li5k0
CuppGSdHL5hte9qqOrtWrbuAzXr85uF9gRFNRaxbGKA3xeUKf98r3ZHDm9YRhk2A
mi4AFmRocalSN94Iu3h4MlOMXwDXOjbzwx4T3MqVHGVNDCM9Md7PCv7TYXROmju1
qg6hhRWYT5sTXEt7f4aVHZjNk+vJejNJ3FCR5hwzwUgc1WFnhgtvZOesFusc1+qf
Jr3qW3G2YhnL5exsGVG0f3hKz2OvOWHLmMx8ixCYU+8c8f+h5ttuMYQbrzzZ+fRC
7YeLhN8izMgfISvDA7xNNICFVjlwsW5t8XM7/VdjrsDiA4M/DTxGxRynwR78kUqu
OxSK9dgL7YA1sm0npcMlorFFAD3GC1Ow4+3/QkYAPAdS843eIGaaSUfuVJDqqutx
6bKLl8cd49+EhAcj/wz9ppvME8obOdRGIvHArtmrqxGyGuErh4pZnbWUGO5zxqCF
uMmefDGywRbwqWoFlBgwOKCnUd4xeHw82uAWfdlDrDxv5NVRjG0x9tYuFhA5GWpT
n+KgvJIfM1+KV/vGYZVLZnEr6NbZJsPCvWPwJPYIjg37GzdhqhaR4W9wz6AZkcW3
1kq+5ZNqiO4eerNZGgFP7wwbk1SwbhZgGmHXigoMewGrjd+ae1k3QEFAgNtoQko6
PhfdNZemqAzbeC7uzFHmsDeoWFxvPwi952+7LAHBCxrSRnLVX7ivyHBcNVak5DLQ
Q8+/mijp+sIcpQlvi3sdbKjQxKPaHBard/HLjJTo5u8jkN5Nb6CgwusiPCUZqW9V
HOpRwJK73T0lcNK69J5xgHPV/oUHafUOInSXS1NUD1o+LOCXU4fogjEGidXRs4qZ
Ks4NnwEFsmdQ/FxCzGXqnOi+M48cprNP5NkqUnOKFOWZ/AQBuO6+aZnQQ36uomyS
h5mxQdQKZiY36emKFFWuHUxOUWBwxU5qeNZvQhQRxN57HWM8V1b8qb9sdRtQSgjK
FeuVt9QHhUWBiESZxBjycCoIM+vCg2yM9UMEA324cyItKls4MfwRAMXEgwIlHkSG
rSvaTiDax0a1FGBFy0u7Bv7y/QD4eoX4eIvQ/vMOpUeYll34bXA/AOGrCZdo3DMC
LKateGlNOBSqMqv33qMI+3IT0C1L9aR8VsCbls+sU4JWY89e98l9HueHhR7Oemwd
qQCdU5nu4JTkeg04qWqisdp6hqzn3c4AcJ/j1GeqA4die+aTu7shXYGs8n4yHIkw
ABEbEjwlU4Wez0qppj1lrLnB9K0F70WLaIJMpychY3oTrIKhp/bCwNyQdnNlZ+KU
WWJgORoAlVDouUjehSXeehTxN7ZzJMXNlUbkYsiuPm5TQmp21fxsS3CyObC/sg/e
Yaa7v6utLv7BmEwO+eRNJoW0jUhe/knIFVdnImwvWSO+uibuEpZHRzLU4ATnAI6Y
NiA926RlxnJKngJ8EAETsSMO4/bHlLLEC2hZ4u5mWwpMhWl6nNfqfq5u1jQi2bRY
HRuXqpsOyW8F8cNre9mj2GxFaQDfebZmwsV+Tu5bzE+DJv4K4aqdiNZPFQWTCgQr
flkMKh8T192XaCDzRIjW/lf0EEAreoq70vVJtjei9h33wYy64knseSyb0zN84g7O
nsoZKlP2HDPU8k60OErgNLmgt/980AFt7dy69Q1FFAHPoFqNH7gW0B4kP9ET92Jw
8SeQqBOJBi0P6FAILYXel+6CnHfiJxUsdj99CgYcCoNPlra3u+VjIhWBrMl0V7o+
wgMiY6cxOY82ETS55I+b/enRYNhqTkkyX8N5I26PsWN0DA3P1ZYk2nS483gXi/4W
QW2eLGPdswOu3vfcxYA0nRW+ss6lKTEGzsZNloAb9oXJU2fnBRdmLifNWh5cPGZU
Ynro7IfDtEQ6oDQRi4XVLu0PlE5EUEa8XGszrmnjDc4z/09fGlikWwQW86m7JGp1
i2bu/Y1Q217w51pFbiDX+B5AOrlFZ0AuRonyqTbUgqyyADA+/oOBryxF6BT2J0FF
ftmbl0Aj5m4w/JBUxm8TlSpYF+yfXmlwMGHbqFVbVoLfieVBp9CrY4YAQcSGobuD
MgsS5zh9LHB+YH/CKQrPpV9c3Wf6PRolkErlT1taYa7D65BXLe7VcMkTXrb3D/1L
cwih2K+l7CEmpKWOOQMJflJkKj7v55I01qMboTqxtQyua1pnsutJJabcUyRfO45+
+CyT+Wo332FUbDGYTpd5B3yPcmN1GAyfpvoGDMM26jCWk4Bh4MPjhV6ECFnDFA21
SX5A3dMTfe6Zqvod7RH0seMfyh1rVQw9qbgOEP4e1Hz2wPsk3JPkW+WOIWevcPe6
VAJrWHYO+o2dXzIz/0dSK+Oix1VSzDKWoRtwhkvRH94H177P95fhwJehlmByKe3O
zsszbaxNP5+0tfMXOpjkT5oooNgHXFWhIg5jnaVR+YOrG61emNnIypHEv4Ruzrjq
d2NwFaQQp8E6VGgaQk9DfWWt91kK/SeeFqR9Yoc0VFqaayZ2DgBrpz4oGCZTydU8
HuDyakZ6LwLgcZ4XXEOz5EI997bqSQ25ultNIws6B35XUwdROB1/5cGbYDfoyQd4
Qx4HaCYnfdFv9iKumX3hwaac9KPoYUQHqhFTaZa5fRSDWYU9vPpvyBmjpIVfqq0B
AtgYRW4LyDc2VU0pIbYIoyms/EEEpHnRu+1jK1mkv9MmDjz2qC263YGP6NZuK0qc
cfsQJeuLdrAC49msUUVUD7c6Bi42C1jtYwj/hEmSXDg4mZFNqMEnCVDSFm1QKYc7
XwAjoWE8FsrSPx++6B4xeSvutE0vTr3qQPnjgpHLgbKO/7sDsdEXAbVV4RoTE+wo
tOBr3FUNQJ1bjf5JsPz3V63E8+DG/o+1AzrQLCzD1o/WjNshNSBQ1A+xJXWmvB6R
ReTBkwUBU2PQ+K1XZn/RncufGiMGKAUdcbt4kckhXQozEoglE+kwHnEhJ5zFz7+V
tMfUpowXJNuzswqvifOMILuX8zJF/bcDCdmZIGKQcSf8O4wFSjZZOdMa/HwI9HdO
K3jFtvJWkdQaVk2a8x/jSRpnI31GzegeF0z+8XCbJ+Tetk0ujokXbsRD7YrQw4WT
98M9rieqhM4OqYvOwW+8F2UsZXiY9u/PyZtyBYTOe9JAQm0d7dbrVP3XJe7s2kVA
ZWEMw1tH5SVuoxLEijREFOljXBY10sVW4tFa1wWR/PTbs5EsCX8g5ZQhpyp/2v+Q
Mz7+lr2MzLe6mbiXs54aQF5M4SOSdsJuKWs/dxi5LmIXm+5qTfHUYj1pc4XbvwQ3
Ao3GePvYephof3eJMXVvwriObnyz9OVH2G8Be2WBWNUqW6CBLqzA9GJguU9T2IfU
pLWJXUKCfsQ05rdIaWT11LZRggD6E1hav27FkVMMxpI5Z49CPLTyoJYAoQHRlMsA
C/e5l7pKRb4i6uOhHjWAuTxO4yZKIs7cNmdEPfbUWJeg3oyhxZOtYzoc2v8SPW1Y
L1wYQjQg+U1d+mVCZfbPSqrjI1W4RCdswojnlRwzztrQ2+JjHV2a72xV8Egcw1by
ltjq5Nd4roqkZ1lAWfCeKwBEd4c2rpC7BfefWBEcuFgPiuY/r60IWjkkoTJ1ZgYO
97BPyQAiZO3rOjDFRgYewOaUqtfGTP5UBipan9aGAhn87UOIg8Uv88hx3AEEDvZK
prtuM0gQXG4eO5KV1Pj+Zs5NLv2KFvg+e8LBF+7bDA5AbjX0Osa0k7bxfFNY82NX
s5da4nRgM0vUqP6046VnLw8ar7Xu7n6eNnb3KBLYyIN9Q7/qRIISYWqlfN5HQwLG
kJRVTWAvxQvMCtiz+D4VUOgctth1Ocb8Dh1GxKb+Z6zbT2rgKz8jqMfxreuIXNpN
ti+swQEQ8oL5Q3OhYEmpBkR/CZbCWrnUwpqY5P4HM8y5cmgiFJk7dlkgc9UY6Zhp
vOTN9Z07ETph42bNu77/ka1JJHekharNUvPONaD/Jy/2ggemxZSXyc0Q1KlLa75C
WmWSE1UibK0lH79RLszw1JtLVKoW5wWVGkxna/7L06J4glChgNA9JcCh9qkzWmjd
bMkWOuvZ4dLwA7TK0SeezLvWIXyBcTbG9e4EjGqr1EZ1dSUy6bxKUoZtwSpi6FKQ
lQPOTRvlc7bh76y+24puRjCVe6OWnA8PxKzNpv05NYihMD/FSuETNt3q0MX3MYWy
p84VlHi9Z7xxwkYTztsAwDkyn5iqnR2gtR4l7KRZuI5UWwqV1oFt6kkpraH9XjQA
IP0aM/6vw7guYQsXhV4zFXck/f1SeOXscM9LdV5BdUrHKFdyTlLYs48zmeGF0X5H
4La76lmbm/aem4HJ3ZrPrt3SEWVUR50aNOjR/5SXhqBKTnccRK8TquO7/mR/sQ7N
5Xmz1j0XS8w+neJUiNdFefmpEYzizGvPl32PAi9XYhrLXpaVbDl9g5dhn8fWl0hp
FqI668MIhgJgX2U4NsHGIee3DHrV2cSMBHaT8rCK0Zhq5s9DqZrFzR4ph6idL6S7
ZLF0kYe6PBqoagBJdfpEg376p2PIYfkNBy/68KlQER8lp21eVPZk9FXmHj/kkl/R
JhT+rAMRn5nKrc1sTvIwBkPnZknbNGb9U4Da3sIlqH2UOnkUb8grris/Hiv6P51z
yKFIe5yUdtal3ByzDIgwLKZxK9yWd76qbRklBRMfDormxV3DwWRlN66VIHXe1z9x
KyCGi4TKUkH5uEpP6hqz0qLu5Iml9LOQIeLlSKsLqOXzXtu+kjJ9zxr4jKjD0ghK
gLUq6l9OLVy+yWud5y/EimFmLJxRtiykwlG5JnT6p74a6Xs+06E/RULq328mnYHA
nkYUCk2nqw9cAVdp15WqpPHaJOLvp0HlHFHO0Sqjf26FptuP8jYPPRQHJchy0DkI
pfg+R1RHDzLPg9o0z6PprRfHrP/QQ1jyJW/smemrmijq9DaQUk2Gs7RvMkkgv+bX
ceClcSsE+waokV+X5cPkeNvC7BFzE78VX/t4LdcuuyLerhNCc1akkVWjxQzTOpyG
IcyCfjhY9RCFdR3wjsetK3ugS7RJN1fCgfvCVv9/ClUu0jFpRLYCVY1/n/r1ZssR
eCnJidGEDtbOwtHE21WKapCCBFIHth8AxVSXGb3D8EsNgECoNl6YL4wBERcU/k9I
ZpG6M680qggJkUZAp+2MbWuGOng2HZbq9UQVrCVvKKVmfC9HyI8P8rfJrvUDHh1y
6JtyfZfvjEdegBqoB7i5wLfmY/3D9pgLC4wyZKEF8Wk6zGZzDArUh2Hfy0RPJ/Jv
VxbEkwd0TGg+htv+/RQpHxYudlBaU425oFrO4/Q2xIt0Ne+rbu/t8LT30TN6BVbQ
44p2FyS6FisjIULkojP1O9ICxeWVoxczbz7A8YP31+y8M7j16HK5M0biW54xU+VV
xQsgvY3H+9bx7hbtlLpXxComUE7G3aaQiei7J3iCSWW9h9urowX5nBUOXvyuVWgJ
MeYEAM+bJqFO4IK+UrzgHj0kYsF8XlEzllu6MoWseTIEjhJBs8fOEkKjKLQOqLO/
TgvCZUmmhAS1zx467nLSKm+M1RdadRWx4Hnj02ecG/DcIdAFVtdWyUzPCxG5j+SE
7kRzj531nC7fgbTkIZ1Y4rQ+4LOTcM4azBb4eYubLkiM66wIu1tOz/FBjNI6rEHp
B6fpxKpebs6jG+qUJADH7XRgTx0gmuEg7QhuP4OQHL20APnchXjmPBzSLKqHO7dC
FceAM+5l9GSSfoJPJJ8/QxGZ03NUyBFHgAbkiIhgI6pTIVCeLeoE5QUgqDxcUmiQ
xcXrL0IMBtORS1TDEoitam689qJq76PCax7Ah6rQoqaM5tup8cRrmGnIn5M11X1Y
unLg5ewM/L6JG7Jo4g1v+daJ26SuKTCSnfVMBgmvlzkLyYKuKuR6sbjIv/90Atpg
n7XwnYz8hOgna9ysYkYabi9lW4WU4Go7BKWU7vAVU+NZBfsM+ogiqFE8JaZ04MZ9
7n1v2DM/BMJglx65cwQKSzs6zdxdE1+34XyiyhOoO+/45L2vEt5bLNy2CKV9YQft
WqgoFOUH1NaDG+F58N/Q8hoJufAl7Gf1gT3UcuCHRQCdJG6KJqLidrte1CRPypU1
2G9r34sbp0qZa8TO2PDB/A7Dqb5eJQoiCca2/Omd9L84dUI7dkL09rrgm9sUmLJ1
jnJbykhZGLV7NbRXEu1HKgYq0DmMANmGnD4b5umtEvMay663lW7T7ojprvZWz+oJ
5/CiztYvvJVUi7IRCy8/aoY5jGRbjysvtJhPkipgZstvD/DqaPty221zXgYc1HLm
FnurV+4UeeDnPiShN93B2oUrgQWo50FuEkRzyeavTJVHvHuLxRI/k+ZO4qU7HBDw
CL8D7y7cz43HhA4NXD9bvcxXCeOymVLO98vBypU8jKObaOCNHaTN94MaZIHL9ZfQ
OSS0ySOjrFKHgcY/TKZYr/JGIbtdkwnY2t0OZ/acoqEy6DngzxrwI9PwQoBDXg6K
8RF5xuZka9E6vU7xsOcGzFyOI7dI98HIBfpviykCinEGQ3R1vwIF5X1gMgjkeTWx
AT+lh31YYE+ucg5OEzVweqSY+QI5yYX9gFYchQG+Ahtcl3DClpg7iPhyULrY4kFA
wZueGrZVfgm9aJFuSrkKnk2UNkwrXj9E2krSJkD73SpawE3h8YqUOzI1S02f7X5U
VS3DiS+iphpzHI4PP9AqNfofjSyO/O4LsW7aXBzJ3AkRoPzJL4dxI6HlhTqwlCMG
R7laA+VMKfOX9G2Y/0NGhYJobE/4bxZlc2D5jKefhm5RK57WHFKOxY5T78eNUTwB
sEyFkg3wNvPLJn+8W+Df4TbPX2Pl94WBIiwoiEp8eUxuyw6Jmv2fWZY95kU5k1mN
HhtJiuz2AqRKN5bXM4v020zF3fQ4GfDYPzXoQT9n1a/coAaERnFEzdS6EEd+Hyw9
y9JTZEFrB86c8+J8o68aIJ7TwDJcfhsE5DSy1LKd1rIilWHCEaH3v+ewGOwBiHtN
zn4HZ8/Ae67c9vZoS9ccPO6abeI2JwKckTn5++HpPoQclaqAIDSgBIBYfkkTVP8l
dlBA59R9lNfUmQo3hu5YPCIc8GstYa4gJfe7R+cuK2u+4UJLTu6AYVJL130lEE0q
7L+OCC/4HNenat6ZGiwSbOq/tDqMhiUyY2ZTww7wDwMIRC9UOp7CnWTgyGbpevfV
pdfzBgE8vcFfDDVJ679B42LYb8+4m8zBubgfxbo/ioxrEIZC7w51cW3MXVBLi3xW
zOM50q30bcpagM0uunlMevdFf/V75RLKtZNuQtjaZI0Dxrq+B3sJFakZfoQLaiUr
/RgDvPXfaIQNsuKFAsgrSl9j6aiesr26ZaZy/bW6X7uodkxVrjoyzXrTwc+VZEK2
E4SqNK2k/Xhu6iCt6gfkN3RWgOaOfURu0tbW2BITu3zr+QXWSaKiJlt5CeGg9e4o
EQ836Ghhp8EwQ/AhSJxHKiJe/moU3x241dOuM8xxAKNX70EIwcuKnO6iTVVlXE01
37BMwZ45qknTCoEZ1YC7zNjBbEm5Ee2MTa/HWf3UQrKnZO2mxhNrejzfPxTLJyiK
KZ9cltJ8kwuKZQktOOR614o6uUJOCzMt8P7qkR8RXjKuLlMVcc2QFhp+xLR4THQO
HFGrqt/Jf5jMbKZT8NiOMIJxWtuLJdlS6ufYGwoUnIJR9y4kudachFCgiVXfoEv+
FSKRwciMpA1J/k9o/fmOABpE60SCVZybzr0bA6v71qJKiwthqLa0LZupA/DrQ+Uf
CZbdvLvUFCAlsawq6xfjJlG7wW93zbRbdETvMMq+cyhnYmhluLcipf33fEnviH7e
tvB0Qxjxd1qO6O0OTruj+7qmZTKslpWZqHUxUf016GPOu2pxuUOG0DqqwvqOsJkH
ceUNxcqT/26ugrEtM0ov1PciiAbWau2Cs808UQW9HF42CHuNH6gmd8M5daQGlxtZ
hUnzqZRVNzJTtVYgdcO0CfwF9uCKeWp5ELOS1NnPU/AIjXoDtYUIdGWN5tpdGN4p
GwCZdIUV7rl+ZoOF+maZrEIlUaJ/MFsBYvFOD6TXHOHW8PRvfWP8bclJHSK79sW/
0xPR8rjeAFgMCfuyKxwtR3A92NJ/1Q2wAo4GHRg1RviN/OvHACUjL/aSreBKUhVQ
4o80hL7OV64VspiBjietxdlbnIizAkVbjKbd956LNOUegtGcvo4zuIHU9q8m8KTM
uQceRrQuVZ/54Mag6o6AFhD1W9qKDduq0V2MFavZ6h2g8vCfGdtlwVPpffNhZfi4
eCZbpt22BjB507JXpyBXwRGs+yRAA4vDKp4+j5JNM45fMDjwmqSprpsqNG83vdo7
/x4du8agNamMOR1xBC1XRCfCwKXiDmc72988HGV6eiv+RJemaqzjXlcLH67m1oD6
GZOTLJYVNs3wiUXCHZB1kUF9R0p2VY0BGIM9eEuhFvnpBl8yGz4J54Jlah8MderM
nOZDOdJG9kguPiIh/n6p0C25DpjrvFaYWAS0xwS3RZQ5V2JTQ1aybVptb6yoVzSQ
S6Y/9M0xRBkqCZjacAHbCIXzkhTiQt1UZISq7XA3NSTXLOu+DGXbuDWipyBUEK83
a6JxCaHgCJJiP7BbArmmqgRaX0TSZAh0wmnnwCgiOpb9t4Rsc7HfgvYI/BFnw4o+
nPIsICQsqgDI5kVxILwi+d0YiKd8nzMK1Jhr+IQmsdaw17+2o+4EhtCt0FjtCHXr
3TC03IfkKdkK4yoeoPaiPltQBKU6jEImqBvzraUaUg82YtaQaxUZKcaK+okBmo/t
RM5UKzADHWavnMIAaO6VgkvdzAWGWWYUjRnv6tF1EOiH/zBKujGsDU2TPgnkMD5a
JDDKgIhR/RU51vV4b8vrJ9DmCSUg2oU9cimDTmK9yEh/mkTYPRRT3l0ZnotTwbet
/EnhyGn7RZABX2uZfE6ub+5gwiK2ORt1Tg6QS3W2ZBE334CZmUujqlO4Wr/qqjf7
kptjiGJYc04xFcMicJ8oE0LbGj/MCUDR9WY1bVuqgwGnH3VVeyoN8AJN9twgKLP8
yDRYgFZ3I717/PEnztqakqZjM0s4Uh7C8MTVldL7o0aDD4rOESqbVbimrcM2v5qy
w7QfJgZqKE3xJ9KeHMCyRlY25+YYdnq0VrqfZpH7L8ymCgQ0w5Hs4+fa8H8AQY+B
pKD6mN/cjs+G3X+oBBlxPQK+zeNYt/jgnSyL5xQOHMo5orvLECrwkvZ68CfQJxjP
/jTQUECLgVVjbY6EUxoXjdpGa6FxdslotEuZrGTB5XkpIOl94SD/Mv455FHMLoHt
3mEuxs1p3IpLBn9VcdGPYQ7ecpZnnTHCmjaO+3UgeObr8v5qudKHBrYQ0EVl7WAa
ot/A2bLsDPhOgeZ/6f9AYlXfw6fVcq7djrOgcswOw67vMzwItRxX5lpvevrZ1UXe
leRx8XZYbo+bSod6rIa2il2FUuZsMSkzuInndabejPPWHYskBWQHf5gx7KkmYHZf
jLg8KSVWnYdlOpcJujZcGWaexIQa+RQtEh7474u1fLJQS+I5wqFx6CvWs/oEqsjH
ok0+GNT4N4lnO3MeG9Bo0Nn9qbbg2lgwvRjCOlKOflf9x50r+hU6Avf0BkXgtH/k
ucz53luPLKmRlvA8q28yI9L7MRWeOqaRAsAnttF8mCodZ93aXRL0w3N1MY/cr/wp
JORMoJUa348IWAjFu1bNzwEwnyfoLye1iJHe/KTGvMwK4lTGaB2EA37PvGBgLO09
6TsexJPTF0Cbc5aO5NEOr//4qO69vI98bR4Jlt76EtplFT74wSW/+eLIHFjrjxsn
gyjes9HD73sgm9dpYIYxR/6m4Pho3b5erflZfiLkCXbUl0fBSAaBedrzYahEFGZV
ZsCC6B5DTUvAHWJBovF9uem/HApciGI6yEu40OgauT3ISRCc2yloUmoQdpIc5GKr
9IQm9siAkRyceUTkPrTb7AD4vmd0FGIZEsP1Gq3ZgJQCWmTClSkR9xEy9aQuxd5k
7HWx6nd6RQN25w7PaR1doaaliHwgSgn9Jkvjcx0MDJ2vnXlL7nv9m/YRpCvacdMI
oyt6u14aSF8qRXwUG1SAugJKPbojm2W/5ndfa9n3bR9WbQkIKnNMLhnwqVoo+G8s
AT/lNliKxms8xBdqq+Yuuy2osDyCBziwyWiZIvbJH+yk8Wqv6Mtid09BtnAMSxWL
9eBDzdeTNHy5qZmTpReFCI1viLVrtopcc9Yr75Bi7Rjt7WUmx6LmwAnepJlLiEnM
DttxUv0aXHkpjAc4xJ8AlaMaPlIuy/xRJ5C/abVfjYWDTQ3mu9zvKk98nwmGInnB
QKbPOpZPnSjU2Ly/JWYZ9rUogk9FW6udQF6zEkJaNJ1g6U27qVIxhyPPbHFfTrRZ
MGNxISM//ZXOzTQOu5d3/kyeOpWzhrUhE3/YGFob0rWKWW5OkVOxZkINtpN8YnLv
Icb1M/L1zoFIL5aIqeJzlNUAbzgyuOiDcLFwSvcwmSsey6agV0Vc2Z9Shy9tE2vM
iC2k7iMCpQNnTaUktr1Yf5pEuup4j/sbBO0ZKvTaZ39aSdRHLm6IQEgZrX8C/ni2
HyEgdcHANUU3UzS/PhFB6ezykKaUWaI1wtYGR+va+enjHGMK4Emdl/J8c0iwF5KP
et+guZ2ZtO1wnA2jdN5VnhPB0Zuq1ThH5ESvBK/+b5B0cw33D0h4oiZBiyNzjuJA
WU3+i8tbDDAfhgC1woSatcDxWw8zuFpN1LZJkAWTvuOK8POXUXA2CK8xFS5BF11s
+p5580gk98+DtIyYvM/YNYWf6L/Oeo2EtB8KlL89voKq1gahQV20DC95+7uCYLBQ
QwnQ9TVUk0ihJjaf3pF1V5ZMDOAkuBzbkfEaxoLIT9EeOOrbMSpuPmKsW7bW7J4V
HS4QaMBxR/xnCeWKOONKIT+pghoimzTkJrIvb/Me2sCiJAIv1WrC2BgutiM5yYn2
fJSivzzeW6EVI72VJ4+7v/htlsRXQS3RzLAYYLJOaibrfPiY33dFELOb0xOp0kM7
gjN5Jmsts3uzNFQuQjYwTJtW2EqkXjo+wtpM8+fX3qIKtmXZiXyVrYgZQuGQ+kM9
OUA4/3/XX8TCfzkCOsyMbziIntZ84dJP1K+lfsJc7GrJs1vn2/8hK50VUtffqCnN
9vEpjQUXmw8RbuCZK4ywDOQpEScpOwcJl2RBWD/rvKjgKdzuRUfL3qanoMfLTVy/
LuCx/VefoSLNeJ4Nshe/sIb+IZk6oI/KjeC5CUHgsCMJjjw79gdzRFAwMiaDkHRR
lbO2xdc1wMK7SWJADEeA8pWTL0Hibhzh6KvJ9pR04f3mpepMcvH7RpZY4QEAaffd
T4xf2r57CL9ek+L9MD/X8DWJwLFHAKx0WIN1Ci4h0kglj8rl5awyRGBR7McwDQ9u
F5s0TsWMuq2NaCEPTpFYbEd5olOjjVizcIg4iHi+M4TT5udXzZEGm67RZaRs/Ard
GjWEIDH9zOagxhAxHQuLFELoQ+Dj7DOIx6btszhXATkQB9O1krwhkddYFh7jYu6+
2vJJshZQj/ab2ILUtlCM52b3fcbgkpB92Uy//FFpDb+19A8MgBAPet1ES5OeMkVr
sDgOdVIHOOJwpo4u1tuPVXhxhH6qlcXrDBdAInwSdLDyXc1elaKoPH7anauZk8V/
cNQFUD1MukLZgggqVmnfzyhcAvIvZjOTl7+ysMe776VuW+GPSg6mO5SQYAEIRX9F
J9PssFX+xr5etI6HQDP1HLlvWBz6tAhSfnueP0+wq8OEwfFKBse644A1RVM9XBZ2
M13DD5BJvcTIHPPeQ/xEyHaqP3zw0h/q1zmR+y/VFcdwp8TaFLyPX/bCETnpdIyW
7emjj4GaxJoYok0Y8kKsCsmOKWm9t8JKjQCiQ8s9WWhww8D6IK1GqlzdV3MsT3VF
WT5g1FxV/cN1UuHTd2aYrsEwQg+lju0Er0MroymtzQ979Ev1YndNlMUo/XNZ58Hu
a6dNfLAqznKv+zsQiKS+jA9Yld/zn/jxDcnLAtGxmrYwTpgEXDdf8Cp66B7TWvQs
OlfqTVTWGUxaFXCGkrWCPO8q3VGqQvASJO+tZfMv5YCSngyxn6Jnx7Knd5qTEACk
AaTHBnEPeYJt2dB6QgcDAPqUGr8F1bDQpBOOKckwpMEb0ypkd6kTF4vmD9tZ3B6N
oKWNp6K7gNxKi9puNI112k25WQFMeiWnzaTgLBqb6jHespWJM48PaMp9ausqwlCR
gtCvUkdzJ/B96d85Jl7HuuvYwvAv6Va5Z3/Eftr9RmsymorQVJSgMXKlIioGOAUz
QeNUemxqV4Rh7g0XyO+LFUKYyrIqKhImHbILa3hzmSS1G0EbeZYELkniOBEn72P4
EQlytxvmZnqPIUsdTAcdkbnFdZiwVbjh85bO6/j8IOE+xVrZKN1px0DB91qpFhea
AURPw3GlmvQd9P0EQFuDfAWgfiDV/CiFJHrS4MaVyWjYrvI0GMLiymGKMhdZeGU8
qCHBHbWUGkFKcx5//0XSfIMirqfB43daRseaPr1xebwlxZTy4NBddbwAhDqfdZ9u
c+vCQ1ci7nuPhHG4vA0ejI0DAcsNXhOAdDguhvYU5B5RfnT2KxfSLPVaS057BgO1
oXN9i2O64STMjSq+2LoV8WAbXQ0gSXy+cm/pwQmkhlw9CKo4zp/l6T1aikZgkMc5
EoWhKJYMCrqXQqR3DbVQrwV4/3WO6kEwevVC3Nb9lSal3m197FX1iO22i37Y7a1S
GnIPP1wBq6hM06vKbVjGTjpSrBEcscD4CwatPtLs+tlKXTT7hPIAymIQrPNeu0tp
Zkk9jTN8CQLkvqeBGMAf38ckFt1Mdm27WkN8Ysi25rfcGkBRwE0J+Vq3Aglga8tk
GIp7azD3ZneRLOY61Tu1le9aIZF+vm6KVXA+H8RiuoPOjMwTBxtAkRT1IZOAW87L
RGXwL411muAVqEzbTOzlFdHV4RDk7chK7ANQZ//dk7ls1T0RXs9z2E9v5HM+Aroo
EseBRR6fIklY3HKvEP0uM3chNA5IxBQiM7JNj6JnYhhcCjVH6f2SOmBCZsDC/OtX
LgyJIcSDFHhddNKwn9UPB6cSKtuS32DPUBHesIbdkbgh4C+LIb4u4AE6ioiipsDz
8uhBFJHzB1tZwJ47VfHlz5TGgdO7HXt+HHKDjyemYKiXs496shidE3vSVNDI3NQL
pOIE3c/hQXDJyvjWG4DMO2INCIEB1fYIQcdd+ZsVRl/MkDO+wRVz6sWgpRkkqWRm
lTGkmFkbW3Z04KQYPxGZm9MioKpZMY2hlgcnvOaA9c2ruxS8LP/+LAIe+Nfrw8Fj
7z10fHsStdcW4CSj47jmh60k8WWFDjQnZeRgGNm5NWEQlTabV52nzbuWG2O0y06n
rfU7ooPbzd0CB5mvRCPY69PZm1PGNso8e45k9gOzFw14zKkstTNkq3qxuv1NTfKX
4zNQNh/GCjKBP5vmethtMaNgusm90zyEpgC0+xPNtQ+IERmpBdHPIw7e/DhfAULP
FpOsSd1hskqtN29LBbwc1XGv9N+dLn15DbuWDHrexwqRoGlgyRw9x9z1XZHYK8sj
nIhgHnwDcP/tMN/KHqNzXsiJaRoA5ywIpI7kIqsvmTgznJG/23ltwry8tt0U2l1Z
gvIefaEsDWu72cZkTUtBBVXSJiHMIbY+ihmpOZF0vNduxo1JNboBOjtp2BmlnE17
zPdcLSDuPbcPBZrr6OINdG2CSSZsYCBTmrYFZDAWNkogjZnOT23Lv+p1HoBBDphQ
R0Cr67+y/8DBOam9E+32g4ttab1sD0UxVdDjLTlAhrJaYazA7yIFDb7Ty48xplgs
Jih5dshfIqL+7YBbHnUxKU+ZId3PgRznGF4NxFY0sPGXmJiNiL7kR7+MGftLH+cd
Pm6u21OiqNchwWUTgYewbXbS8TPjuzwxW97tvNLIC5+0bmEyU5cbOmhCLzeXg2ZZ
YredPepD2gVxskSfy9UWSo41BKBmkiaclTBE0RbrBFLN7B36E3TOkd0APq8iGezu
p9ez4xaHEDyOEzpvBAoUAAMIbIQ0/DU9tB9ec7MD4EkYPEI3PJlqQBHN+Cnf4sAq
GaFxSWmCPxq/lOLqFoFOqIGCDIw2rXWf1HcsPRMxgg+kEK5XhaSOqYMQAgTzyzGo
k462jhHeGfBEWNdixXvR4J2eKI8aiy5vcsZ8k010eFU0Bg0+FwK37rvV6MVfpch9
myu9XsFbZl5TO3b5TuXO4nFdO5KM2Hg30BlqH20HuZARAEmoLrZUSUnwww4wxcNN
nrCvYecesw43HAVRX3ygoSoEjU0ja1PKZPNpKSMn4k9X04jK+YmDskXj1HgebHIP
ljaSaB8qW8XIh+jMbLr6JN4y7CtPyOxeGV75tSgKXzQcAUlNbSG75padyML+ume6
4WXXQVXIhepPvVDyo8rn6C8FLb97tR14bInhlgDfAYDhyOTjTpx+jZnl2VfpWruY
lJZDLq9EpoN/puufMPQigHtcddYFQNwCkAByGlYLmqbxVODA+qyHqCK3rgEjiesv
dbWHosvb4mbqkz5DJVJlyS5+N8UPZCP8seVI/2bOcdRwtgqTMeqDD95WclFEC1QE
pAwhPM7w4IYDlTQkJjHz2ps+LGOHOVRWu3k6S9lPOA+xu2+Sv2H3f4CROHBrCkCh
JX3V4VN5E0kw0YyvAv6bDkb0jZwlrWmvj93phRFzDxvSQ0jg2w19TGcSbRFJ+uar
e9XUprB0T3YOZTsC6RJu33mbTv91CZYS4llKRLOR1/bdViTjD3YqW4ViW2Xe/Q0y
ZNcuFwqZ0zWzBc1Vrt58/otZQ99XSZfwin5og6VzM8kMjEBRGOs7zjsBtUx9cJQI
cifj5MrwvjEyNR2BQwz3WGv2g99za1WMyJoVwkMsTK13YHJQg6J0R5w/OPXjk5+p
L+1gjJU6/uWhqKvuCYwIad7stXLk175rnSLP0QpKCUveEuqOVFEohNYfnTNM0VgR
XoBjRtku5bOzrLGWaUlsTP97muax183ASK4NGTQk806ZnjVa/Q+1wja7A4/S612G
Yl+TA4nNPe+KKatPTF3vEeHWGCgnOOGB9KQuhJnfSfOk/2xHy5xJb+An1b78AoPV
0i9p2nyPmxKk4V0hD2xwSln6rLJC6eYBFGmDAyvewaDjIglMjQqz7U7eW6BTnnbC
qYmSM8y7D8EC/J6bzprY7bCXAUiQW5C/e7jRp1Du9+5n9td8eDv17MBr9KNVE+ER
oiVcgAtz1qPz//Cb/xtySekhUJ3I++bKirOBU1DztKIrk/mfYi/qb+Vrbp13fe9G
3DIY/bDJ5074gr0Wh4B5q9tVCKTbahdQ7nRnCWeR4WVwsksGybVOPN205WlaI/AJ
8f3FCAjZ2m6ZzkTkBppsvExAiGY1ZsgLlj0OHr5VHCFfSaWf399t8WrRmaKFDCMi
3OIJ+45HPTfuIO0sPNrRcjjIrqmSB7E9WD/ejbKeQ/Vsc9u6Nss1fODZpHBVGDBS
1zMb+gap8PzXJXnI0mc2gdyrlfwxynPSSqj6RppOmHgbGtUkWt8Tx1kWHvu87wu0
iXgcdhwFBSGwcv4P0RO4Mz+yLcJklCkuhQE945bYYWDWBpn+qM3x2arPDs2hz166
sV1gmo0Fpl5yALj7jgYd5PDRP4qTxtymgJf2TxbZxD1dA6t8WzcmJ0qiuqQJjvM+
rMb5RIQTF/WWwV8Lb6MmqWK7K2Qxuri5tQQ497NsW4fYx2/aDB/zzoTYnZoyMZlt
5Uo7RU7Z/zozLoV4ir+Z6S+bIkDsqXL1neQLFq59yPj3s8owtLmPVfdBn6Y19Hba
dgDAD1lZOPXL7nFjJlkhAZUvE/QtiUjMxg3Pot20QFeEpslUjahbnTbBYRzwZIeU
EO0+jlmjorF0aKV2h756QxiiWuGd9ugNQIBBAp/3Hfcsot6tSubqclieNGKP1oPP
FnBAbQMX0z+LKa6w1zvqXITCwgKGIKQP7YXB1RKQmMLYoKYiCdSBE4062e/zpGRF
sOSuguUlherzrkXbEs8TM35uOuAIDYuDgqY+RJ4AwRQS5wqis0F3M9fNWZLiawjK
A487Lab9DVFbriLmMkX+bk4EwptTD8HVcbt1HzTWq29ynGuYOR653A9o7FoQNyy0
Zk8GKsDnNE7zwV78BIXzFdLD/r3IfQVLDmBP+4blWR9Hnl0dDOgTQZJU+ktP2TYQ
29TZstAFkhllV5VMrdqjf13UO0MbOfrWX8Xo6Q3jEmWFTyEoa2AQpoqVfs7HtMSd
J0XDWMqV5uU0t95op5y0DJZHXR8dKpezH65pqAiH51npv55GLCFkzECBQgNwFnHL
R7Bme1LHhgmTSMfYuwBIrphKP9oXXKnCqZoG21hvVH6JNlMYdTrDI3PtFODeJJeZ
b9LP46z3REzdl1+UtWjJiwe8vuOr0vI8OTLsUbD6N4Fwa/QTF/9I4PhHcDVQPDdP
guqJ7rtFEU/LjM79OPE/XvwiMOXXkOX2v7UaVhtXIJhbSEngm529Fo0TrimqPEWk
zJmkcTkQluMHYrzFhdeOGkhjLWFjVVQ9jv4ROYXTmW1AGSm4klLd4mXvNMN308rS
W1uQNXsK8kRTWOtolRV6tCYG4Ln3s724My32hCtJmv8GKE+8LwsUamlY5YeyXEn1
/LrK7CKJ0a/GgUehaVuw1/ufRfuIMnO+WoUycbM+Zmdoc44ju+opeyQjU33ch6CY
0RXbye4bPaSThu6ZyPlJ8tjyuxgTu5srQhENYIE6oLI0XBDFX2mcGXlA44og2YgV
kUmgCD6B3+LF14qiOclPsAfuk+5Tp+nqEY7s3CBq7Pgd7cSjsnoKQSlJVxU+4uJe
0TuXIdqbrKWVgVYW0dOfit+vuG/iaCTXtcE4lSgVYYnAmO+8Nl28Ba1Q0Pk0D5ol
eI936LW4fnQrkQ2kMH0GEUKkSELiPlotR8go2+mbdJb8H592BMjbbPFKphW9sWkX
B6rhBjLRLqV10BMJLYn+V7zJHyv8YjZpWcJBglcIr30wF9IVGjIlkya3jLmZ5D9Y
kiGGXrAI/3BdzznLl7WXK/X6ign45oXff1q3s47RvPdVkJUClvxMPTQX8OoBKCSf
yA0rWzCQMLlTIYPlALhDQDljnVODfvhE6ZpmX+FB8Ql6VeqT2JmQ05SnLU2Mq+Xs
wMufZ6Yh4Zz7x/pdQ1T/u/caDQDu/e44erlJOd+d2qUShCrjax6Odokn2sNiO+hw
EJx/TDGtVGlYSdxTQxRd7j9Vpr1xdkvxVigWizbZV62wx6Ru148ivoxhxiQd6OnD
Oh1T1LztZ5lHxsXsrwwP4rw4NhWu1hzZgDnfMONVPX4ghzXD3eAJnqmigx/ByV0D
mMCY3Tq235oKXD5ykVksALQCzgGYeb8QkGjzOcfo6czK/KWtP0BQ2eJkZa5sm+z8
x//ERxbPJfvp9scvfZuySyFdqoNAk8J9EJZxL78peJqmASwQxRKxNaYbo9ek/Zn7
htWANGrNin+xCMy79jhZliGB4FNwSvqBj5nZhjbSxa4dEs/wZ6WRmjqXGuWzdTTf
ZWHnoxh+cmLRTrSa+eWZq1tzpCHCMCZN10iLQfw4wVoxjCfMc7cqLuQHZyUcARlp
CBSR7+O8By6WKRIPLX75Kug2gf6Eluw8Q5v6F8XUHMSntAEDEdNN8X8a0rANp3Yj
xl1Pi2K+VtAGEohxCVSk3LPfURWnzG7lEUbr/iYGDpjbtY/22/BJl3Q5LS3ebYvo
TbaSxG6q+8gm1WUIdbGYGlMtvi+5jAExa86dlog447EJADCbNfg5Sjz1aJxmy2iE
OCD3/MgzcuJVZO2OEcGuvZyAEK+GqthbE1Xesf+I2Fi7r2kzVKTzknpw093BT05u
3IBlYba8WLIePM9NV9qfVcpc+1JGc+80Bi/5xmu7zZqOP0ExneILDCGQG+vs6O4s
BUwWMurrTTzCBJl772wkOCCyQ+Jn4OsHDIhozI1UppUY8Nz7aUoeGCpsx3Dh9mxI
oaRsIGX68CNZT7RcGk9RSb70/JQXVdjHpiK9nHBI7R4ot6VkRSIp99hcXZS1dCJY
tMaX75uGNKesnrmtopybCGuuT8tb/NLi9AiWOQpyIwm6r26vQ4k9lnLl23citMXC
BOXgleuCivBMQB5Kc/2tZ0mzo6YvN3notrSKupAR9z0IbYeSCrxhF7QIfNn0XtJT
RchbhNkXJ1PG+VQ49eb8eZTV5lrk/zCUMqQhHDy7H6VSoUSwYapVQmKCMTj+Thcq
4kab6kfjJavlmJgp7VQrhSaiMV5x+a+eb6zgWY3koyJDX2UfBt/4wE19MSeL/4cG
gsOp0GuClCSJZu87nSBHxm9OCKBw2uoZG7RstE+/DAXNxBYi1Wz45ke6kjs9NjhZ
oJDQmwvSD3HMhjW2AoBfAGkzYshFARal3rOauWP4N/5HCC1gMSb4xDQgg55kCEUP
s4zRYnryh5Hl8+QaFnDpvMa6fPtgwkTSbwAIqVinlyhPXb5OoqpMhbUaxKrOgp6R
AVGqUyOs5ot2QYGdQ36Roc1C8LkU4jFQUaM2DfyeIfC0DQfe5ZTEn8BHYv8JHvlK
+O26Vl+0ehLMgu3gWP90DQsqFDqBMnxbnJLcdAvm5EPAG0Isi0A0u5/n1sRtqMKc
yx8EWcMQ0NSodIdwhDDo7vzhq4ntoY/XJOD7Bi1ErtlgxCik9y5GmrvH0TNPtMD3
eP50Ug0hJMTTh2UaCGldHaUNHrppidSlekOF5oi/mLyz8baaSTheeWlsY5HAZbxL
W0+PXspM5nyr0dC1yXa7ZLVyOUiq+xdt5ERBhfMoo9xtw6NE8fZFrbYTaXeikG5m
fcao4bfotE2PcwQh7e+oYHu9pSeK/2yLteFxGsMPmFzBWVe9lJiAqztaxpSBkNIo
qe4NzsUqb+v0aX7/Q4CAuG4sxaAgAdH6PTM9rPN8M+D7wXapJe9c4jP5d/pqR6wb
y3igi+CU3KUm+GDC7HRoKIDnDWDqCtx0aHMRdEA4+8rjuD0cpYvQJNlQt3KERZ/e
vtgFF4cbApGtrkEQly5RwliFgbaE5nYsz7+os5QL5/PYiQA1SY3clGUN9ccTGakX
HRHSm2Uew1RSQOr/gzL9oy7Yfjl8j+1nFzWfZav+MGZjmCafsGf2HLtl+YmrcSB0
d5zU1NKyRSO1sRCionXUTPlUWT+NMAY+QhK2L1Unys5lMRQ6084COctl+F9H6VXd
zjycXp0ACDN3EcV9kMIvc1Y5JRmAJQXWJnu0FGdxl2anNnXvC2KBcs41pzXhLjk8
wwYJBW12Nw/RaJFzBBWb4jF/+9rrlyxmc8rXFGeT2Y4MAFOpGTzUVqI7Fv7OePsv
MhJbUHZL4EW/YtaRKrKKr/jrruVbJGuaXb4q3fY3YiDTW0z1qahpcpCvhC0qz/2F
Bl9+Sctyy7ZB5I4ya1sJ8GGn9S89UOF2tceFWmoYVdC4ZpMijQJ2bJgh2DV+FlD7
yGo/Wrisa0fiC5MTEdhd7U8DnCpB3bjatq/ppw9o+bzfKU7PW8G7GTiC2rD5YvRD
UZjl1g7TdEz2YbNut7N96lACxOhpWDtA6T1a764kXwGFZpCloLLb1bpiOhlxvOHL
frXAMASUtSGxTRnfm+dHCPTHxHb6n/JdZPXUijmHrj23yZXRJvjNuGv8jzWyHzCz
Ro/JZ4J761MByZ/NIBqafPS4YAuJ58ipXxwTHryJ4M0mpTamxg1Xj/wGox2xZF9g
f2CDrLVxz+l/qalvN1mNDUiC+OQzrQt/MrnvjMc73CnrFSU6u7IDdL8U5mmRdtrm
9tSul7Ek2wbBVmki1Vy07SHk/FRZ6ROxkyItqQaaoJffpc2EXlRpndXqJUPRs4+8
dxERXNRzEWiVlSzZvf1URaAj1Vtn5Ql4xQAphUu01AyupCpX3wc8bA5K9bKtuuP1
ZKnuRTHm3zOEdf1LMI4mz8mM3ZbRSmV1r9x3uKSbbUYtq3+pV5rEPmdQrBfj2DW2
EwU2FJ47lwMNUm38V8FkUqh9dTuA76C8qLNnsePt+cKohxA8aQUNXxqmw6K4FfxH
aqIot4yPb9Yen1vPlFIzwIUApvKXYQynt9/3UHLpYZI3+pSCfy1SUNitvz66Vio8
BxMhTrypwFaA6nqqWZP6QT/UNdJKB8XoCX4bVPxLwh5rtMgLtL/SSn/+4/cPAd+K
snWwDexkatnrIGViFEao7+6+hRMmuqzbsD7XxoOHyIggBiepQj1AJxzi0EIj/YI+
rSB15hCFneVe1rcVDbfbv5xiCCPzthksxE3ReM9kgc82KcL4vSZxw2TRV/6+rlMe
NXIRb7BqKuXLBkJ2ZRbooGQMV9c+4xdlfTsSFKnEIUsBkRw/BJkGyhrPZFBQ3uQ9
zLS0OBZ6NhFGbyu6jDcWSCwEfKbZW78CurUgoyvm2/9q4JY6bblv6cukZ8rozr5I
KtMJvsZIbJtFAPElRXZY+jzLoZc+NX6TgZ3LRRnq1wcZZJlG/OYB7e0zK+HGfi/m
igaUIWBdRkdpYbq5nfnHoWNK62wNzLD2kPMKIgKF8qwDF2y/WOlzbYflXlS89hkZ
F7N2NNWiYrEwZ7zDhW97+fEhFmwYqRQkjozcvQWdWTOebt8YASHcBYdMgatp5XPk
qen2BX4gLFT6DdVkyZBs0LLqfSAArGNtRtAeMAdlQTr7ZoLemx95AUYJ0t7YaDyn
O2AspNRDjPeI8zKaT5ntAfqyeJawta/hsjbJIQYkYttxC80RZuzYkQVjfsyKnksj
Ia3amvfX2eRamNpJruAu2R1+j8+QgYX6hcQd/4T1OWLp2wiKZFxbdEaH586ffEIi
aiQmtJwMT3PxJVa4DTPA9jeHxz4XuINeVZSsi2+dAAvOtX398AhAyhYT7iAR3mIz
5vwva/qiCqQCVXsKF2BtZikUzDcv0gGOikwBGRi83okt35op6JX543VLZInoa5RO
ZJFibOW0KMpa64skteczX1+j+NuzJwEVTarr4hHiWb3D4gVmGiuAzJ6HgRT54qT3
+KNV9EBwHh+P/ROOLXPf2CXQ7esNFjWVHBdN+HGx9/FQJDVPOCXYNPaGn6B1Xlb5
V8CBKW+w36xz+yf/1wIEdxo5CKB/PFlQ3JYxX3evmabxMz7Q7u+meJKE5jEiU5di
GvJL4Phtj15QTZLMFqOq6rF42tMRJboWbQ128hWRM6yGRl5bow//c+RV21JIgLTp
c7Ea8A+Yb0bul7NeRG0/Xw/bq4Nj3QSA3pFPsT12j79YpGtSQvqfxBp3FEQl5A6e
bariGyo3CaIOT3DDTOwwHs9hyDrJnrWI4XTNiKmMabAsSY+Q3hrx02EQyBC1JAcJ
9VGxfjrilenHYmLAY6U1zfDjfXsq+3GP/dTJInHRGqySV0JuxhXpA0KZpefuaUVP
6dCFaE0KQV/vvGGncjk+19FImf1BMHNcAhmrIWnk+QFOpB/5rO9El5vAeiyQ/wUL
XiOOLpieKPIv/1QBnF5Y7L/gf5I8p8UsYu5clz1C7bNYaJlAqUTAlLpTVvOkzm5Y
6Kc1HvdcNqbeoBNtsolSNcSnL546HqEB3oBBfgC2/s6mXvrJqmrUMo3r2eBtT3Ph
ICIAiqtH54uszhwrrISKjdqKs3DooymZ4wIunig+Dli6dJlC0VNS8ZZ3Y/CcjqmG
9/5QSxiE6kNUQ6vVBD6bR91XePXqAA5Urb425poBzzU4J1Bzohdpi7cuz9iOEMS6
pBMKLHpb6FxwVJHN1rrjTPqRmS3osVltV4Eq+qFXG05Od4ojji5pNUQogk9kGA7+
sMurMNc4Q5DrMntvynkQvlxItPft37JjAo3249X7nlxWAVe142GFmSeLfE8MnpB9
kJeijJBa2VxsVLJFJZTAhEtLClhiC9sInZLJlunf9oAJQMQ16fIsNFSdDHLMeAmT
G2h8JsBOHiMOWMf+1nxipuCHPUnoqUAHUqIwnTJOQ+GlZ1Kgp56ja/qn1bB0xZpj
1Nkpp7laZGfjkp3VPMiYP0ERImjNKTT5tvXPb03kLW6lRO9Bx3gx49nzHTMlIl/c
S51V/tSo+AMDk8GpayfnjNhV3caXw0DCvGtLcmgAam4GHan/44j9GDwzQTmb9Rlk
g3q5R1zmLg7JOxxoHnVsHweAcBbhpUbSTBkgwhCau8DDBifgE9yDHwM2ZMAp2vBZ
NTii+AX4JYYs6TRIVBlMnhrtqR0HO+Rrly/SbmpdLvkm/TsSZScUrM1KNm7/0c0S
BiJNtL5GMSmvOOc5Hl2cRXWHC4tncV4kmfSmJfX5sQqtvbB7Epi567z1OgmGoJcI
HbRbHPW7rln3IPokEINnVk44FS5WP97cUtgp6G8YjTQKXV9TIKh2CZDw7NkCFwGq
zKrxvc2YGRbN51uMHyk125ukGtvcOS/DBBwxur0QkRluq/y0c7WW8vDwPM4DlPsr
SOTikI9aZF93GOOowaAEkCz46EyxGi2NaDo0fQBoa/T4eyM8vFbG+V2CN0QEnz3n
Imk0aDmJhqwntIOqoRzfgy1Q8lLXTFpXTU37QEFqbKjGq5myMHvbT/oDm7mXR+Lx
80gr7swup+X9Iw84ZscNtOTLUkefJ7LfK8vlxDP5uyxG5etmAB9LTyrEy3jQkkCp
7fgU7iWx51b/1Zc7TUmCOv4EaSO4pp3CRcvlLRQm+bukQIHN9ZbX63s1+M8gQ4X0
DB20cmsyezcPNzvJcaG1k5YsFApFT8pf2/d2Hogp/gRUzG708mb3tmdqPTQkTOC1
OMb8SpRN2fjht6RBh5BAzOU3aWdW4g5nJIkSEaEiuIPRxAleGRJeC//MzBfw/lx0
G27tMRLlOeGommu/zJ5waKB85X8i23WOnyG/T9Y5NDdMRFVOm0lItiKya6QesbqY
T6/4fpERbvD0wIglGAYaTZbm6PTbVPGJTecSi/VRuMTMRojFw4FUQOJM2GewSlBY
AtrWvL3gpDykGAa/06ulQ2O6HXOOo4NLDD0O6KSFeqcOaLYdFW5NKssoHSw5BZ7e
3ldeGqKzZIyUA6W8y3Q5mztDk888WJpF51TPtoIB3xtx3sZIP4NuhamKP0u953sV
COF8jScmaG51n/ZvtFjXzOJkwTZqoXDguf7HrGKzXvTwTehUGuHQRLNejNmR3/NJ
bT7jIaWcrmiHhEuwcEvlt0LUcM+y/C27PYfTVuDSx75XcvijXSE3tgyDLXjQpo0a
VYEZYeaU8MzP+wC3UA15JN7+igPx65aLDcL9U6Hz8Nac1vcMsrgxNcgFmI4LjPWH
+yFq82oli48dCL0TIXBqTe4UCcYU2+MYw2mZ3nXNbHATfxdzjTdpgNSqqQC+cysT
/qRLUEuTFGXZ3YCaxPpilzwK+xYWR63ZS2AfQL5ZgM4X0RzZLdcvjIly5w6j1FYT
G8AYiycxgMEPgCDcSUaptYiqXNUvDzJBVP3PYAAVZC3nBmJAUWHm4bW/IlB9HBj7
xCQORgk3XD0w0O/9GDv2qplVUuibvJoH4nOHPs3qUZt6z1Ewqum4cOapJmaZQZj3
xuOFKxHOER4XzXE2NE/umC65JROmIO8SNgkk9oUZE51/MYwVQsQ+iAHmeYlZYTeW
w6GvaMssZvW8Pvwer0tZNMjZ7Wwmppoed2cbcyqEOVjYecpmPUlkLbsmjUXAGjod
f3+oRjEosyGrJzknXCgzj+neIg9RNIKHyynUwlwVs0JACXUiJpaEtOb9ySpIDy0a
iCiqVWLQ6ciU8/djjyYCp7HGJrKqsrrqj/dNbNDeLZUdmDxkH4Jpjqf8WupL5e0L
M/5b2Jsg7LUIi0Mj1sF3P1L69vKONb+b23g2PU7LAVOhz44cCbv7EZQOYW/dOwoO
vC5GlyJMvVL7/xOhZ3adSTSJAKisNsW6hbtcpRJYL0PF1SlwQ32BKAb5PRKq7Tlc
GOG8OIBze4B2duaHUDTFomh52Blo3OiqlEjPf+USceyRKrNN9c85r8qtlqCAkz4T
dRaUowZlO+nUHpQK7JFM2cmVpFvboZNdZ653OWpLo4Ku+8b5fAi10ZkjGUlWADzU
AsL9uXeEUEwtToAKunmz5Z3ksBEeMlK03sjV2ky6H1y6mY4p5T4AtgQgGECglAvx
BiCIsNOiKTTUZMycRbsqFhScTUrwqOXuoaK7Q2+vix+6gm4bL5d3njtx3F4k5+zd
nr1RWgs9P4RDdl5eSVl9Vn7tpRGjHWKHO+yF4eUxqPapDAK8RAqHjKwb38KZE2iV
yfjrJyt//IRfz4S93WOKFm4yYkAWpE+8dmbP5lzJ6swmYW3jqAbK/KJm555LDGSm
kDS3EHwu6YwZqNBEESULOMx+kf2Ehc5R6Yt0ZaXKALk0ynv9o4O8/3cvrgOQaOIr
H3pilz6RNwuQnCpdzlQfGWGNpnGt5terptLEA5KR+JqrGCZXI623k4/0Bo0mHRHL
W7xnvHiGHlQHTng5DCRizE9dv9Ec7TAKYY6lnSdRcEdRR2H5GcBps/5dcJTBR4zX
XDWwHJ/rEoqki6Yhl0U9cfzVlUNrrwEVcAf2Z2WAi/kQvVd6RiMBK4EL2f87rEpZ
3UqcsEXZ6ZLFW74uvBqR+lKh9GFDVy0TeuV76muaQf4OpKl9B1Kn7IbO07tU5hVY
VLH8O8Dt2gPIfNvxP6qNPyZroW7zugVcpcv2WqNafNU761QTAoYpEGdrn9M4RAqL
gTrJycIW6PBK9Cd4rXQzEQxWK6/pOC3tyUODX1Ei27lmHpDRcLjUOD1cdj7w65XH
BdbLbbnbX3sNrDDeddpvqeckcXyMThFdkpnQBF+sl2sbGNr5LwHjB96Xzg8k23xe
xtoElT46fdi0lJxBjp6tNqou8Ft1R2MjrTJLmWaX3kLKFrneKtuDQyyiBjqQJLBY
luzv1Afrk0onaGhxGVwmRJ2pq3M6vjnTDCuLGJx8kXd9kJ1jeeynRP3OkKlNWywf
jZsd4Mw2scimZ/Nt7YO4j9vulxhNCkU4ixO+SaPD3DvDEj8CLmqLV9bT6hoaKRaw
Vkwj4DAzztodrY/DJ1BrPoPKV2vafjNGU/cAFLNsyAdt/hBn7gT+Gsqvbgz/sd4r
I0G29AgDseVzVGTZjcdNHkvnGRsqC9dYDs2b+PuRP25g0H+MiYzeaY4iqJ51yudV
HOYVC0KHqXna0g1bh/xo+XphJixBcCDVxg/HSzJ4LLhH1bNBzb6zywNeaONOmhzG
QHxEQtxb3ubXNmuJjcNGe8UBtNsvSQurny2s/G/Bk8wB2IVa+jabJXPvGcw4lWup
7Yj1wzRn7WBPBHS23VXq8wNsmd/Mfo3ZneZBWTFtci7QNzvw/EX2812jPc0mxyTh
pTIfw2T5Xgeug2aRuoSIPoWzpqCF0PoaqTNWvF5ESuvjewoPW+EROknPOOy1Gj6F
8AS/b0hXlL27ovnP9XYigQLVsqWRgrEz5M5N2kKvIdTdoUVle6Fb/gnLyBzmMQKL
4avE3EtcrU2/tMKDKcXEZVnYoOSrJHwIyZOTITT4a/A99tBprDqzaAe8hUmA9yi5
nV6tOc+gupS4PeoJa2IAgDfGwjeCeAIr5Q3HQ95Wj8lnTmTHvNygHOSEYV9Mm8Fe
0HYJnri2aHho2iWmlarXNfvNFtp+V2bvFIoJwgEe/S3bsgX9yx4+7L4dDd2baaGA
6rlPmIqLGRlzXjJa4pfvRNvMMcOuPdQ+q3YfiPpZCcBAckicQX6ib+tI7+7Xruac
drDZKUMEjaGiAOqD9X2dsHQfBj3jjZsh78Td6mbmGjJn6ykqoe6UXpgbaeoYt7yu
neUQnpOiOQHP8/WP/FIquc5Ocey3mbEXwvBOeoRQnHjy22LqC/LnA1YpzNySjHsX
rkUprb+Hjx42YoWpJXpEU7sDn6KxLYVZCQDFNWrNG2D9Ugv6/9+3OLUM8Ahqbj3N
YK7ZCJciG0KMKeshLZQnYkquNSrkcTyJiV0wyCre5v72qZEXDklwNS/QwUltDydk
8vLRsPxi5rhNQ4XDJzYjUHnqOvW/VGFCH4GZCQJvH0egrFWZLjHBYhKeS+1H7uil
JqhSRw+1ds5Za/nhlJtlzWHUeFYM4t3j/GVm0WvaZ3Le1sg3fGYg5VseS0CvIAqF
fMdLbsfxl8mHUlBsP1Movxt7oZpzAw781fZWVVbqylybR+TRGMXI8gUXDONmjsKA
S8iAXQMm1PApf1Th8iCclF0JnLjvpZDp4vhy37jzPWSb0gPztcZrfniFQPa3idOF
3MoKYrtBB+9E9yW8CyRKnI9oA3PkPLsxAudrpjCdJS0dgBP86S2MKlp/tZvgJtxg
KotsZEPZvuti+OS7hST+u88aMyPQ8rkKW8R+TAosUavn7THGBs5XdEOeS9n9TZF+
N0Xt/FSSOwD5EpcTLhxRf//hWLbg2Cn0dlB++AjCfs9+IFdJK4yfsS3dJaz7HnUF
FU4+X2S4vzB29z+COH31UQUrb05rYNVww7SOnnn3XbZl8mbHgVYuIs2ZqvInDfD/
WqcnZElnyOfM8arZUyipe/p0A2wWkNOMDXBfkDKNx4IrMBh0nmDm6yzibAK6IsAF
o8tMlQfu/aO2Ny4l+2b30WEZShrBUUXiAl+I9R7tqpg4wPcwehLCA1hkx9des5EV
Jed65NgvlC6rmePq2Qz3RyX2eq5AQenpaIYteniTyHV2LYG1MdgPzIFAKzg7rXkZ
23n3JD6QMWRd93882uSH7zxNbX3GEOM4LhUwX9fastHf8IhHg3eJAR00kh5eybFC
vGTP4BaiAzZQv5+edyAaAPAz0HawuYbIojGdjju5lZ7n9wo6lXI0yHLMqUdyZ4uz
0tVP5DmlZh+gqqHsU3JFqWsZWZX9JX033uxQ0sgBppDB/QAOQUzYjZAVNdU8lYUH
1qqzj64zzh5MHciRfLZoqhbQT9pTjlIUSnLFQjs61+KeMN5thygJFojQ/Nf8gQH8
3PnRr9fRz3dSR67WctLvZO//L9vfkBcf5JK/fD3TydRT0qD4ye+PvClcHUIIP6pZ
b+4xpREIHFHt32j7+7tbiFpoFkirnBPoc4RoyfU0GU4sZfUpAaUOuK/BPURHs2Kp
fa2W74++ZNpjzQJB8CdAiY76xI1px+OHDi7/rMcxnzvmH0GmsI92mVdymq1TuPTZ
UQSE4ksAWwuPXJ5Arx9p9EMSSYXRbKdh2FiegLutvHEW6SNlXm1/mpd9ZUMITp7z
04MSsotlDAlzbDw61r2DzJKsoyBMArSIpmjUAhD7C1XesnEdmu74CVB0e0+VZ2Ew
BPHgSZeiftrzwDvE6z9ZDyVf3TKH82E0ctG9/KyLflPrOOiy3nxNFooQtTO5I209
eH/d6fWERa7kwPKcjQGNuciGXvN8I184r+Yyjh488IBSsI3YvLNsQgGSCUbkBOmk
n3zUHmk3ooVa6hpSVu8kXKollwPe6aaKqpvN4OktYHQ1R5pgeGD2q/Q0zH8/DEfX
khgnwiLFgwi0xRrgUjV4L4gStBHAlcoj6eB8Db/c1WW7nxh7OwO9HL/2ozATpZZX
ZgA8dwtdZF5TLOYJFvuvIQzzh43to+CkQQi/bb1UpojV5soHNYteoJV9NGv9duED
2cebRacIXV0KQcdTgoK5xVu7gqakZ4ppOXj/6OfUyVxaOptSr+chCTPq+8Fugu+F
xPGB4V7EalmmPD59132Ksm61Lwuuys85VCgnR3znwtwQI+E+EbuWKy7DnSaDGjMv
zxvchsAcB7XAFyMEvaxPZOxZ24aMbO8I4BNatyFlnwCVf5XXJEnZbBEcql5H1nxA
XfhPOZMqZ/ecmDJ3gwfpwjJYWdmf8uW6EAWYBaxVWUxoVEoDDUXpEPY+X3fBT9Bk
O9W6xId/q9hlSDGLWaPO0mJ3Wz0V+SKIipKsA7k2jhSCvWw1wScmIb4cJ/9nZtMT
qTOsbpnjW+bvS9tQsm4XUhKZF38bS01zttoUbHWbnbhiirUuxcjvza3oE3XV9IOk
oBSU8F/E/qPDV6dV/K7mYqC26KqhLc62lQkATBium9DGO4jIuyF8cZ5oTWLgeCd0
U3ivSDNDCEf1tSudoihw9HmMGAfvWBrZRKclY/1rRAj1tBhZPBHUYFd0znWx6J65
tiG5ORuFuJzkTcNmnjJstRzZCwAB58lSCkk/R/KJX65WZr/4eIpJVsv9FUeIKvdR
tCCNDhLVGftBRehhTp8HBJ+jh+xQujeG2CZyiHzNSMDEXMVuc70tcpmvhRLFVm82
E22HFpo5KTYOqJcpnxi9QCcq77NaHow+Kcl/HVhmoh+0QhhJCSUHdXpjr6p9SxZp
M9Lj0fUPPndbMI7tAWNYJf4FQNK83gdzYghS+BtpWBXRhyNDX8GT9/8ek/g8fMEv
zJ+xvTHOElpN3R6Ic6Y3VG+pf//P0fjuy1xgMj2BS7b9knR0dnPDSyfnjhaW3rt0
tZV+kwS6nHkZDvVP57p3HAc5nt7WP4zrGY01J80hf+ScEj8MF1XBboD9lqnrHRH/
MLW04pGePhrQldxcy7fF6FJOee46oss70TTfwMWQqPQyp3Uv/S60Aeiui4gWzYiD
Uba3O2v93t982hPlPlrVRECKgV6zC0YxxiKZYHSoWV/xrj0cG6R/bLdyW7tcP3Up
GcGqp9rmfGwOQzgxvUrICPS+iq49tr9vWUEemQ4rzmxcyRLFz7VdAWKxOojI0rTO
KNs9PxKHHzIm2WzBYGXOiMUvVENZuO5VkxHRbXRk6x/Wyfyk8L50+pNII26gVMYc
mqJCYbh2DpQndQGaoH/3xEIkjTB7zwFFi3uJQEJFwBT9YLfk06wYmPqeYfNoPGlB
yVx62GO2WAhb/xQG0p+RdFTrnJTnKNFj1M1NFGzlItm+k3aE+OMqOEUaR6ys/0z4
rfNV6mwV2bW6RzKZPGzL137pyvMjr2pReUDihzwKnPPF4mETM5Di4xhz2RspFKsu
LsWOXrKcvop3cjxOsWYLgjsxFGR4Fqh0EHgCPucKNkd1AE+iEzj0ol2ce2ATJC6U
4CwpSYmU77quvf0aoebtSGce/QgVOJbQ3RPFHQUQYDn/HeBeFh3fXYPw3+XbqGXf
hw0y1mo9WE3wDmAXGjWRMrjtwcq9sTphA5sZ+ZosvNuxMnWbk71VM2ohzGWGQtAe
GNuPjbCdARHDO1BWzRvUv6bunoPk8tCbg3gJQB9BWLAGhgBUR+21FMx9xrvec1Wz
8FZDV2tdr65CigHtG8BNJ5YKCGcHQHcNteu47ktekTimdKDlyh8BcbSj9nuKvlHg
+IbWewhgr9bCToGjx8bWrx3zmraE1EQj77TL5SlZmv9RLl2SJfjYcZMysdYpx7Zr
knm21HD9nQNxDG1dsrAhW6oPfk1RG0qEflqxLUDkVnQ6Jzba+QENiVWYEpvUvj09
UlgnHcWqFoaBD/UhwD8xogVeLQEekKtBuwpVxfzWx9HPlWRlBxaAGyn2b8QJGh8y
pluOOKKdPoisCCdi6HEU8b8uk2q0FP2KjRpXRPQoPMTT67iD5s6hKLLUXE8eyG20
mN/Nu5dLfXhd6ZSqJ+1JodUkbTFnhq5DZ33KqaNLm1zLWrYlFmo8fZI1bGEsAJsm
6vyrduoXxu/6tEpFgUc27IeJGcoTep3VmnWYCmECcWDKUw1zpBSv/MWH+CUGEsTb
Dm6FbmucQCnlJAxcvgXizuyHGO/pS8le/6YN5Rk/4gay3EzzXyQs99Ab1dLrK4zz
Q8jOqKFBIWwlzG4rF/r0mNoIR7H/sHbE6JPInzc5d2kHzdSXRQXWFlkbxr7fFFQ0
57ChF/Zc+0n8AhZz6Q32zYmwDyZpaF6PKDtoKTKVgJVP+mbgN04JaMBWA5a4VuhA
natZV7k+CEVb7Kl/DHPQ+bmUW7Dq23XLzHDr+VuyfxGskSSRQj1rpWHZs+SyUQNc
Mbr+CJ4yUrI8km/L8rSSWqPDGrRhJCR7IqzELJLhnxgorm3Lmghe4iH0DuQkxVsp
IRmnkeIy9JXPSH3/wHs6Klgs/iFJ0JXNncWgbRACR7cNAH9RhCfcW/AGmHj1MU2B
/7mVmC5kj/qoBpRdyfSJQ66VEbHkCfjgVKs18tS67k2pc5LkSuRhfN82SwSZFbDv
5rcHsBsVjevBoPs2xaLKbrOyPEmLKNMB2ER69wBJSbU+uo8US0VzpZLWYpGpo0Jk
8JHXzGxcL0wo+s8es/kgn8eX9AE8pi84DAE7oL5T1dqLAIxuWLdh7bW6VCQZeeV9
M2F6U2HMoz4C94kG7NVHGFB0TTovsZebcmAFUyaAadcylK5NKeZlt2MMdj/fO11d
GTItlcC7mXw9hLgVZHc6mxaaCbmaiYbpz0fVcPl95uJaoGIMXbFqLsMnHAUZlURK
GcMOkNu9hMsk2p0SMyOF5Ldk56X2A5Fvdcnf+Dcrgy7DBVNsafW4Np6MwJMbowmp
yyhxJUgG1g7BVxCWtYvZ8kr5raPTfQ/h7+YKdm/xD0d0DE7Ne8d2Rs23fqlZOINs
v0mELneIcshIluQh41hQ5WPRUUA4SmWmT0b5vbXAmG1GJhQgkSHGDs13/WSe0LOf
fAYYJ1g98ipKSNgXYzuu9Dad4hvBt1XJyN2O3fPQt/HleIwu2sIDGpDnRA5EXNLk
7gbsug+x7JY4BfBRu/tS/npJ/FzRb0xtDpvA9MDjSlUtyqtk176mUa/vF5eY7xJK
fYlv2QgujTMlrtDZPD1jkSFDRjFhsz9tLA7u2UD4dMs39qIZKAIrmEMX2hGWygqE
FBkr950CycpvJNH5/gqrhh6BEfdaXf1fXB3ECo70CssXQVleIjuXxohIEo9cYhQu
epTDnwfweQWdPepCEHCuT6vve0uwJV0NYo00axZBrh515G2w5Q81AnzvCS9AWdVn
UMAOWuxQYMrd6GY01A3HjU4TJm5GuLpnIJHJiFOxEMWDRThD32aD0F55oq5aEv3z
ayDEctwU4IexEhvUONaImYH5kx9XMkOmx9FFDCFp9S4hzFgjc5iuK2UaePDWOXjq
6ljWtyqgclbY04EZE9bdPgUSU/WmLi0pab0L3mONbcA43YzKbYdb+ysGi1hrRnBU
oKirQ6+P2u9gDdJymZR7SOtKd2POOQC348tymWnHwY9RcMQM7P02mrFl/6cXy+4O
V8uWFIZatuHhS9+bj/6hltrFAuNsoaKUyO1vLmFi82UaHRJlgBTveoq14IDRvfbk
EiNgYDOi+ydbsieUl3GcnKQlWnEqQUsik+kiweDsLSX3XGNiCZ0Rx21XGaQoqB0U
CIdmCEmeLEpXvPPrx7rg6TtKJ9sZB9dqo54JmqmjPQ/nfvn2Xux079pMgQwhKPng
hKfrQUBGTddHNYcFWZyarMGKpuzKyFQKNTKzve/N0UduXtfDXz4Jl0a0Pg9IfRWE
pkXSg35sonswYcMyNQjhk9gOH3kitTYucTpwZayqmW2gsv/Pclm3BhzXyzCE/Zkr
YTukZzkkjIU89pZIOd9IT3aNNUyioW9h5lrkrzqDOUFLaoo3hX4eP7cfu6wlem9P
USwVg8P0pmx5qfCE8WkCS1neKfcBtGu1gwE+yYCMWcQ5c3a8QOxq9IDk8Nk3YLpO
6iKtep+AvvnaW46bdJDCFlijmdT53z9GYfP9w0qTDcOUgviZOoFgAxI7Sz0bxKt2
J59JBpzt8mmR3/c0KXPmc7hASkLFo83Vwa7olF0AFGKUJDuxWVSqv73UixzjKIB4
OI+6kabhR1lQo1UVHvBZ4d+xuYgnqZUUHUJAGtmslV3rgwfniAJhOzCQ+vVYDlG2
OXzPUFFjRYgxhX9LUNeaRxZJTB24v0PnUCAywDr1UOmctm1Pt4qQsD4XIT3VYdyV
Ljdt2qPvbCtW29d9x0RANI/lKOCBqGhPTrYKId/HMeIBc055C31Ki2LYkuX3aAmz
pa9if/z06q8i5cRORb7f6cBFx+bqSGMMa9jMkmpeShp3yC4Tj/SeMhbbilTC9lPy
kflMI4SUCno75ilkD8IxoEjYc+J65B35q206ErQr2PwCWVrKyYM02iJ4n97J5zhq
fw6VG8Ol/7v+hnSklk4djb207ccysFpAquw2+3yFTNr8n6nc3KTw2Vm2zz0i1dJn
3JlGMkZ1VX9poFEpVjktt4li3R603dmwa2CLPcWtyTpe0NhhwmotPjXiL/oKlIL8
vXr9brQYnH4hKt35etyIsJ2IHThG7xPu/0dKS1OFa7Gecb9pPCxIv4tYJXToUyEC
VoWS5icKn/P5e0fw7YEN89lzZzxqz3yOGmWV4GSifl8nVdC6Fy+Aaht0Seoga2kw
ncy0hpvaVp9KxJnSblG1lhQBxuspFfT8aDWXai1OdQwdV//xo1KMebQm3E2L6yGI
bZHeG15G37R+nCiT6ec5R+2NoKVq65apyRXjxBKj7dr5tuWp3A4UOlQzuFeg29rd
o8dg1lMa20yZFCmZF1Q62+gXgZXQY1quYbx/9L9V+2+OVm5MfzTJC26pk7bfa9Lb
b0j84BLxE2z3YggnONCv96+6+QGQRE+WwC8W0vZerJOqXbvGL/r4FNe+XFKUUA1C
KlJcTIMUsL95FClACR8UggSOBt16mHAnbsh7793R9LPIroVWYbECMkTlTEpElwO6
wza1q/Ed4OzxJ9V0i33J1t3fyNvXtTla6ucTv+wMaEUqf/Z7SEwlJBgzmNVdpfF+
35HhK8ArjXqbFY+OU87yBcKi7ORVLzg7JYZ482MZb51vt+CNxihzxsWFKTaERiWK
GL83v5mVxCuYWtHKD6n1dhy0szxI4AJ8fsYNZ/2JJ1woq11OmhGaZXqy3hgm2pCW
2oxRJvBPwIssKYpkB63gHwTurYIXBFaIkW0gGePFz8I0llEdQNdpS+bwE8bnfpIa
M0IoC3RTnyDiiNlKxe0Qobtkb1QJJP7UK6hyIn0T/V4O6MKRXqu2mu2jfNnZgdTK
vzil4glecSbJoToon+w4+B/rKBwUPX/22aO1u0Nw8FztxDSP+yeeb+aWDGpPOffp
ioTD581Dn86jnneEXKMmLGMT3yHMElD5vo5DX9cCg94D/Cki9X61GpM+Lsf56WvI
StvCGyoUQw5g/fpThtcCn4bqyDWlbMr+f4tkWVCBYPEpw3ODyC7xKZlVn0colrt8
l6pbrRMHbth5DZPMrXVLcNcu97gTYF0LZADX6XIqdXwYQZ21VqDUwxT64e7CV+uJ
/jG7HOOfsdad7AwF5Ihk7nN9APBFr1tyHeVxdfbBibx8KEGZgXMwpmYtf6YcOqd7
SIPitc2cvqd1kURPe/61E5Ho7JGDkB3ZjFUbs+8RC7WwsmXf873knUuD1OaQogGp
sVExoH6NzTMYAUFB/lpldOL22yNxuGJ5lf8x1kcSPb1otCs3xz7O20r1zAwZMSnS
PCNrVtySCI9WTVFu4/eCaDDwBl0Xnxfdt+qOs56NtL9WgWTDtbeFZDraaS7OrUUu
ZTOZAKK56OGL+MSn3P8GlXAjZAtH+xYbo/hHav8fzFLUU/GVzzo9n/PSyBXlWORl
w8G9YCD5G58LKtYIdIdtqfK8DowlDmZ+SwmUwEgvAK2sf32w6TERitLUEQ3xQwzF
xdx63Fazv51Vzjdxq310hbaFWcK4LWQJHOUaJ0YxvLgPAbj6D6myP5GRXvvcg4NF
iwOOcwjUAAkXXhJJy7T3Js1v1R0Tx1Mf9c8XgfFeaK0bSB8W0MFIGxRPOgbmNcBC
UGd3d3Q7UcdnGjUd3d4+wmAEc5E6Fgi/qyayw6+WNOwvdEzAeli6lBkbC6S8C8uz
ae1Jz0M+onUegHtPTd3hvDQq+qj941ZZeQVWvoUAOill65BtY6oO9kEiZ1Si2+n9
BG8keVkJK4LCtuA5bbDoWUCrl8Gh/g4pGeOaZT/N+fQ8PC5mCdjzAlBFuZOC6t7I
UIE1tSP3zKIVJ+6IvNjZAw0p/fr0JBO7+Jj2btVxrHcrboIvuaaUFmzpHVwSeZ6b
+jdOl9/dA+8T00O1EEIS9IBrnkjjYitkgSbpjclT/uHg8fT+MMEwnoZtzffi4KOs
yZdtC1w5hiijygXjQDwVtb2EkBb8qZWIOtZB2KnhHIse69zG1omGh5DCvuN7+LMU
/qbpZm0ZTSSUtW1a8ZicXtYooYppwdW7eZu9Y58SUFSqnlbImrB9tECVVAWVg4U9
z2IFPd+XtmyBYM65WC4bp37zG+kAgy1T1SwBakn4oFABx5kz0tBXBYw6cwEpMqrw
vVXfwpKw3fomLvCo/1xC1kRaBcMd6OXXRdwkepQQfCm4duOaNbm9E/gQ0Rd8rMNM
JjPl/Ep4/JOMSqV+bd+RvEDlyQ+ln6e2y4lSa3iXtisfK/iyskdw0z3er1bH7V4h
av/nXVeQHLm8SYuWaHgrVhci0GFVIjFaowNcFM8AKbqc5fd11yQlo59pMHEhgsKy
h3djKXLWMUHV0R4ctqVxiauTW3AavbT1fKpV98cv3PZOQeSFlbMTqQHbMmPSzOEg
YVIFhmOLl8zJWwPcnt1M45F34afu14Rp9AJo6QxZdzI/b5SFtBOpjg3hzco5Z8F1
xQR6uksUIjSUhFF2IPdr8ZKhfCijO6CduSmc/VrIgQMWvN+VlOAc98y1LbOSmsn0
Qhe3DKEN6qyY+d6UXnunafISkTTsVlxuaYkLJBxjD39d+/oE5c+BZlpiK3ORag/B
uBsFHEyLVB6xIh1QmUJEP93b1gpAt8JHrCM8KXt9W9mzqhYOhJ/5OqbG0jcnelun
Bb8xaqn7hPeYxkW96PDH7hcNY4SXI8GcvKTMsT4u2eLPPJTzURYvRsuprk+8TzM8
CVW3qq4iERPwzSPSY6s72WW7lQ+qsdBsKxeuBQ5GIqn7TXP2TT8ByUFfnMUk37PP
dqP9quIJR4fDrY+WRWoGJdDCWWDVbinKg/vdy23POhdWp6uMPlepOURgB9GScHIc
a70sOxuFH6uOccuvwnkyD8FYijE+YTIDw/h+phVKngpuxPSqY4z11RAFTip18QVd
Lg3ZLOrK5p/mOpry8D6kp+lGgEZPtNb6fdj5QgffM1pWM9JO7g9zclMJ9mPybxI9
vN8qcUxR4a9q2IluTCoCpalhf4hnbszQW88JGSSWXKzn+cTHiAQMkjHUnoHdlkt4
3ixa2XSCtEbLLDm22sN8tuUTmMC+7EE7VWCbGbIM1s78kwf+wlsrukIhJTP6Y1uZ
h42Ofrb+3UP5Y4lVTE+bFPCCNOrKvNVb280e2jRluul8Bs9XLXYzP8Oucq6BXL7a
ee8f8H9MEGsq6iUGfdHYV4KR/U02WiM5OXQRzXKyKrXovSIleWlPmDuIbWbOhdb6
KSAIuaE4RCONIWtpcSy2PR78OC/jzW8aX90gXF5QAxUenj0IkwhnKqxH+zXJwrna
oBKBNWCIukeNEp1ISF8SnFTxYsoDzXbbEJqeNLBR4bkgimmrCNjbVof1l+Xx7B1o
Z7s3FCM2YII431Wtb7THdonsKqB4lrPX2erXubBSHiKt6JTRYNoQJRw3o0mtt1yF
q1NHYyffUsRHy4XGua0l/fDB5G8kyF6nTmHg/88LrzNCJ+zvE93WRnoWTGMBrdoJ
qFrTqvJ5bK3VIwD2MyIIwS8IxiS09VWYOXwcd1nXxNM=
`pragma protect end_protected
