��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�����ՂF�1$�xU�	�.�g��z�!2�l�7��Qb�a��O`��:��p��kJ���`�>S��E�J����[g*4���҇����o�$��A�]?��硣�u��!YbּL��V�B;�ٽ�6P'�&��[�B*�Hk�
@
��DH����H�Jh���#h�j ��i�׊�M}���!�T��y��#TZcZj��\��L������1�Q�^�O.���������I�xc%ӺG?Mį������ȑ�c�0r/Vw���/�&(�yn����d܋i�r�yfәQ�D��/���[�4%>�,��F["�,ɭ5M���	g��.�^U<���b�1�[iZW
˵�9��W�3�����o-�����ݛ�� J:�vq�6�<�1^�K�D�o�;�G�+���ww���0�c8Q���ǿ$o���N
E*�ai!�rg�e�cY����
_`�;^����\ģWRDI6��O0��&�g���H��8%~��k���4�g0A�!maV�2�^���Τ���L�~:
��5x����d
�����jw_�H5:q�\�3���iئ�A�7�+O���U����Z��J��YE`r܁N����1>�e#����pU,[�K��c#Ϧ���Y0 B�9���H)��fY>t�Sŵԟ�A�'��q�Ĥ�E��0�!o!`��[��uz;f8���#3����ȉ�%)����J�b1��9]�K����g�0�$�G���ʦ�6{:ͪ߹o"ۋo3\no�#���Sf?��x4�x/����5�4������۷����|(�}�F����zd��<�?ݧT���{	��� :I���`�r���c8��F��.� #���+&�;��Y��2�oOR~���/oe���G�I:I�#R��t۝x_obY�E$&�"�K��4^����K����Ѳ�֞�o��±M�"Ὓ[9@'+�%�X�I��A��2}�����1�=L� ��F��^1a� �Sc��">cC��6�vDk�?���7�A�=qw�Ǒ��,�Ғzك^ۂs؟�Iy��Ww���������)8y�������x�����~W����������՞�eF8�h��=�aǽ!��YUm>�-Z��+�y�t�';{�2N�c��}(��zK�*��@��x���qܵ�e;as����=��}3��3z<UJPE`�ME�����ƞ���T۫�������jj��m\�n!-�]����*�����H������L���K�~q���+9WSL�^JECM��Di0̚0���U������Fzo����#�T4� �t0x@�2AD[�0��؁��DC��+L�c�";����*L�Hup1����s�K�o��evo�r��/�#��#g�6"q0'���#!�'�w%ß��\���U�;Kf���[@$T��l�̲�Al��^+=1�,"��*���}�鈎Ď׾�NW�Z��3'����� ��@
��:�)�X�H	��0��5S��n~����� 0LE����'�M��ׂ�[b��$��:5�r�j����c�1�nB��&��^��T hRMaͮ��YAW�e~�X:rD��hӴ�VR�ݥ��bL���6B����z0>;�5�o6"w�7�!#E�H�՗{�$�B��P~#�V�*}��d�[Ӊ�����#Y������UI0 ��F�.E�&GM�r��P9Ǹ��E��E�Wx��V,������FQb��kUR�H{=���$��KJ{���`�-��3�������j�;�ڞ$k0%�l��%��KJ*X�D����UI��ö���TX��J�ar�s�Ok�T����WQYA�>R��w[�/�R�Ԝ�T����e�v~M���!�0u&Z%�9�C7+�/7Z�
�DPKW��4'�_
�gD�Α��bK*?Yx#� �p���ytߨ��q�������G������x�n�$�-q�����	��_{��]���.~��(�ژ��*�T�	�ua��/��@u���x�8"����(~eV� {��V�Qm@C���1G��{ �.�os�+�K�0����u��~��[+���MPn�(x�5���S@����뉢��k���I}�Z���[h(�U�s#���`���筬17E���PQ�"S�_Y.�������=Z�yG7�����k�sAӌ�M��F?�*J��7�m��	��\�4��U�S[Ր�]�`�9��P�ݘ��3�|��'�E���ݩ�5�E�I�V�Ə�a4?"w�`_�0��(5���`�kYu�sg��`��_yƹ���zR�:~�fby�I�s.[;�@[���ԉ���Ĝ)FAW�n�]�/��Q&��$��ِ|�Nu<��)=��v�N`G�*��O�B��_#�5�|m��V���f� �
�J �1�㯣���h�m�u�oy�r^E��PX _�9r�"��!��!��Ğ!=����i�����y��JۻX��l�]'vZ���׹�r�;���Ł�p�`��������U��m��1ۻ`6�<Q�|�T���U{8���X������F��r�9�:���]���r�G�͘���J�.p@J��6�H-�Xd������Q��۪�%��3f_�j� V$V�O~���k`�n����qE?�m	0�����U�7���o����?��Z���%V���̸=��?L%N���b���$\!؄���Y^���Ѡ6ܜ�=��͝���&60fPF�j��^9M�;�W�߇}���骍Qx�9� �9�9.�L�iN�+읛m��t���]<� kj3xgj��f`�|۩:'��}`�F���j���L�������q��I~�h�~J|
CŮZ3�K��&C~P���䗪�v�� ��d����2wᭁ��%�N��� ��EcI.tI��������~\9�2|��p�팸�;��%Q<�Pl�P���w-x�ٌ� �3H��k�g�>.�`�'|]�&��&����p��F:g��I�F�]x]Ct��U�ٴ��|��tn��Lˊ�>�V��d�$�����˯b鼮������~�@).��GA{с���*��c��e�0=c� ^|t9�wC��*�x��J��X5.1_8|��L�\hΔ�nxy��f� � CG�����NvJ��2��)S6s� �he/�AgX�P��3G��QV"�P�ʶU��,�N�r�e�<(���\���bj�L�\�g-S�V��L��O��YcȜ���E̞��5D���@�K�@|�\ ���bI(��*�5��Z�;���o�S?Z�&�$������ ��WL���$��!�r:�Ȫ��z�ӗx���mU���C���	�> ����|��$��_C&"À~d�OWza9Xѱ�٫̜���i�c�}�&��m�H�P!�/0L���V�}8�Z@����N~�č�|�P �=��M�����F��\P����⸨34�X �J��� @LϞ.4R�>���ufݘ�B�p�� +�eA�� _�U���IgX�<�����Q�O���M&���8��4C�V��`S��VzPB��A��l���@,vs�$z�С��9A���Dv�����qS����K��jԺ!������M���
b�j|"���u��+~+�[���~0Ae�Td�р���|{/
"���T*pZ�K&g&��ʲ�]m|�&X��nC�y��XW9�0�1��k\)Y8�f��m�>����S��?le�/�F!�"
��ZO�oe���-TV��z�WzU�T�� �F��7��K�� {U��,И�����(b #Z�p�� �<����{�躥���]<���3PL�L-{�ܓ@Ú�X�᷷�cǖWF�q����],`�q�\�1�' �+���bo���\Q�^�^�4Y����`le�Z�3�:O���ǈ��ʢS�݁%k(��g�c����
G����t�y�Y�|_��~�\2{�z(�1.vRV�l���uu�c�#��\v1p�\N(��e�/:�8���В�7��(�ɻ�9(@@b�	u	m�q�ܾyk�49�'�I�7�����+Y���@L�Ect�}n?�ww�r0�6�Ǚ����(U�� �aʹIgu`�*�B�>s����&B��Ww����e�}�h2%M㸴S�Kw~֌m`��[-��Q<p������
X�b-��m��6�+)B/�]ezo):b�bgg1)-XL�Ҡ��Tc�ս�WY�փb+>;P�o�����[�����[o�ﯿ�+��f���[��r���[�ϱR�`�hl��ʬ�0�Kd��:,AA�2��e�~6�,\}��h+���y<_�b ��~̬��r���,B�?�y���
��msG8o�F���
���<����TYB�<}��91:5S���n�ﲲQ�!��&Ht6<-wV( �r�|D�_g�~J��Z����h+� �L0 �̳���6��-�6,3łt"���}����͓c�58*�!�ފ�.�����p|_|�׭��'�@��2��ӧ���[�Sr�YŎI�}�?���Wڋ�%��c��{U?z&Jݲ�L��L�)Y�>5��3�h�}��`�cP&�ў��3ߎ��s�BOŭf���l�cp���ҳ�X��	LMEj�X��S���rr�/�B�[�&�Q�l���B�Lξ _��o�}��2ҌV��T�!i�--��ZC�j��ܲJ�2՚��/Ȁ6�-�M���M���� h}��X��IB�9PB�eBJ[_
^��T��YG�<�M��E��)/B����w�r!��}�T�A�6�E`6RoJ�O�2��w.x��\���k��U3<"K�p�؉e3N��	ms.����P�G�6�;�/��� ��^�x��
��={K��n%l��=�������V0&έ�b���P5���S�+�E���ܠI3�v�xJЏ��F|�d��w�[��L�C��~|�1��/FqD�S%s�ns�'LU&�0�,8��=T�����E��e/7s�?��o co�,;ӲVB`GM<k�y`/T�.(W[��]W:*�>�AN[g���h�K��E.L9��
��̐/��Kv2�����(�o�d�C?���e1�G��%x��z�:�n4V���^��-�ؙ�<�6�K�)}����E�LƂ�/z�M��tk/1i;V.�	u$,ܴV�Ѽ�1�J����s�G����`h�B�C ?��	��$}or��R.d��������7Q�� �+7��IxR�ق��M���)t-�J�ؒ	�4&�L�@�w�ߪ�#ysS"��<�	R�o��2@�����o�L�XwH�z$%0�|PCSu�3�5]���m�k���R�� !��o��J5���S�|^��DyiB%���U8���Z�J����O�5������#��n'��_�!v��&��7m�"�3���β*�8�Md�lg�zfǐ��vI =�'���ѣm/�5�Pf8��GO�h!�#J ��r�����E��M�'�$r�/ʉ��/��, �����%ڙ����nC-�Ⱦ��x��Ax�����m� R�)L�g�0���|P�Z���X�����Ȭ�`����J�7�������.b�ҭ�H�_��/�'�H@V'���x[J���T��9
M��G�=(��,�$�l
l{�b��r�0��������T��叟�$�������+y�y�����\�^���u��؈�Q9�"{֎ȴ��3��w�tYXAޥZuNF>��8)ӮFK��k � #2�gv�.����U]шj7Z�p�,�Ǆ���p������\���"�����sx���,�{H�F��/�5uɣx
F3�s�N��ڽ���< �7��(����v�s���`B�]��!K��(�z��UEP�*�P ��O:<V�F,�$�0�ǜ5����F��`Ghc�F|H^����-�뎐�^Ew�8�w��������_
vv�����˧B�SL��R����,rr
L�����f�줲����� *^�����춹�6�zr������a�)l��ml�1��z�+�J
���6��������g^���F#��}�i%���u/"���h!�������Ȯ��9}��z�"��aS�����n�9
jN�,83��ą�s����f��]�8��� �ʠ/�+�2Z*;\w����]N���;W7f��ېU��qsgL���K��<S�G�5 �
X�`ƗLO�&��V�C܉��:(�Gy����ֺ�x��XjY�I"�(��9Q�J� +ۢ���ʶ��K�*�e@�>J���jb�;������dWt���.�R<�DE!�sn����:��*���� J�t	-7&.��n�N0=2�)�"Ī=�U־���v��46�8	����Z�k�Y���-����ґ�U�
|.��5���C�{��y��~Zi>i�O�Q���U�*�:�\=��	���?�6�Nj���v+��h-�:e%�f�g�wA���:O!���T�P�,��i�(�����X�v�͝�5�̰��|�/h������e?��nC51ï�z��@b�)m'����(������m��@z���n�8�����t�+=ODa[�ق#��K����z9���P"�g��i���_ţv��׌���Z�L�/o�+͑��`��g[z��޳3�H�7��PL�w5�07p�����5x�&�M���%��/#�3��8�Dȡ�;�Q S/��Ҏ9����c��T!D��]Gʲ
�/#�z����^6\����T�������y�Ԃ�heT��!<����~�wq�4J�-�_Wzd�;�O�n�(�:���m�à��ԫ����C���f��̔yE����F��&Q�fkì$��:P����"E	S�nkK��/-���B�K�b�����8˿��v���g��x��({���4Jc��П���ҫ6\D2��Dc����6���Y�_���U�b�*1���z�{���q�o���FL��V#�1p{/�b�J&D��"��3(����u4#!G�˿�U��t��|L����';����n31��, ���5� �f���͠!R�-Jݾ�����|���c����©����TF\_�Xw�� 2'��nBU-|ĵ&RǛ״����lbɕ����A)�\�sNSfm�$�^��y,c��d(�t�Y�=�+G�#]���r9�ן�WR��<�_sa�M��<�w�r@���D䞄Ԣśc��T�a����H�b=�ob޼���Ju�c����xhB��~�<E1�T��{ZJX1�b��b�J�Z��Bc�e��M�nJ'�p|�U���I<��jT�(ڠg�������!S,�3-D�����L�*�����0��Y�!�^�-W�#6d�	 �W�c��l�g����J�[��A�����u�ɂ�W���'����\	��H���)�n�d!H6S��x��XC�O\�6�7I���j�1س�^"e��Ze@i8x��Q�.	�_'�# ��ew!�+��V)u� ���y-��h�jAa���j��-�ۍW�ٌ���)eÔ1�gȠY4�Ãk�/0�K]&�8�6!>�3�)�"pw�sʮ��<�:k��Ā
)�Oʖ�cHz�F��+	��_��B��SM:{��=�����1��5(T�Kf����6�=%�K1��`K��!�7�ژb<�����=�@t.��A���>���|��j�O�]ks��F�������'N^($�����d� �+�]'Vo�	X�P�fvDL���b lʒ0oê���8�w���#����M���Q���������Ne�+�GR���w�)�0'�,�)��M���)8(����i���h�~��	e�a�[�2�];�QdY�f#}1蒃8�� ]#��o)�5O�����Ν�qc�[��o�PS�[����-���c��	n�Pnt�B3�jA��c���]������~>�G�'�l��|)'"��iZy�K����}�Q���ہ3�;ah���(d�69��y��ҕdF5�)a̦����h�#��s4A6���L��.���N��.�<-\,�����#u�;����l^�=�&Wv-����s��T�;�;a���](%�f��!�q@�Ob����2����YO�Y����;?��װu�[�[Ǟ����/�4�K�AO��˦��X�P����D>�Ϭ7�)܍��?Ê:v�v�z�Y��<?�fl8m&�n��9�B�	ɈI�`{�\�e������9�k�g��w?�C0@��,i$6�;$�-��NS����cX��%������I��w,�Gdp�l�+���*~>�D�khAǘ1v�	��7�/����H��C���{H��F�0c/���ǰ�;�Il�k�&J��-u�;}hĞ-ny5'0�4{+�7&�X�q��8�i����1���B���x��������Ψ�x;j������1���*�d�T��g�I��Yt%�5�V	��w��vн�.<��)';�2�%F��`./U)
��B��$����K�9�/�*�_��roG`mI#��w֏�@=���i� {�J�4O��X/c�3��Ao(�5�q��H�53�-pF�5�r�&pEo�/�C�a�J16s���ō�`d�ct�T"̊7ԀQ��Шb�Y5:�)=�SB�ELO*����W@��1��M[/�J1�;�Kͺ�4?G�Nۇ:�#��6=�
�fr*89��#�ڞ.wlg�`'��WZ��2WR���&\���~�>~e����}�h����6&�۞�]�4W�\��`ۧ$Q�̒7«3iϙf���A�Af�%*�أ͊oRY�kX�܍mBC�UƱ%F8\�T�����&�_i>�,��so�G�S��PT������~�dT�}gYU�`c�?��s++�m�uY�Z�zx��֕�������s� ��H���a��Gk���,�<�/o*<�ŲD�ї��^�����3&�p8���_���Jf�%�&��'���_}1�g	�Zӛ�*x��֌Q'�����0���O��k�أ�jQ�8�O>c�8h�N՗0��b��Ap.gS؀���<I����9x��2��߾��O���qd��S�|��A`�����Z������$��W�tP/B�z���κ9���8Ǔ�k�׈&OV{���y;��-�q�|x�-G�u�/Ǟ�vX�K�iFY�xA���ƴz���s
6�t؂{�ލ.>�n�N��ہ�ܺߌ��C�ltT\�%W1`�7�W�Lt��A
ߎ���(Ʒ9���7�l	�ɆߥU����ʍ�I  ���x��Er0O-�ɸ8�ַw��e��HܙX�«pA��YO^p�P ���2H�KH�z]��E�d ��f8�w�7�d-hc�q�j�����Z3�E(^/_zdag�^��2K�!��5�!��J/;�	��ϒ�*�����7$ִ?X2�H��]j= �"�v��tz~ȿ^�:�@�>!]�!�&�1Xp����)�M=V��-m��c��!��]��/fH�X��7'=�dg�O����L��ޑ�v}4��HZ`�,�O�k�R��?c�ej8󚨱`�iv�!؇��t���T����+h^�|��Y��q ��w�!��Y
�|��}� <�x��~0��T|X����SI)���&~��Z3Ye��Z�ݍ�R7h,������++H���°��{q���w�&�܆Jr�ĸK����t L����D3;ӥ"A[��b8@�z�;����R>�(|;�n�wa�D$���p0J>&���pi�>�[����������*�