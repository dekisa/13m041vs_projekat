--------------------------------------------------------------------------------
--! @file data_gen.vhd
--! @brief Simple component which generates data
--! @details In this file component is presented which generates data
--! periodically. Data is presented on register 0 of the component. When data is
--! generated an interrupt is triggered. Reading data from register clears
--! interrupt flag.
--! @date 09.11.2017.
--! @version 1.0
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--! @brief Entity declaration for data generation component
--! @details
--! Simple Avalon MM Slave with Interrupt
entity data_gen is
    port (
        clk             : in  std_logic                     := '0';
        reset           : in  std_logic                     := '0';
        bus_address     : in  std_logic_vector(7 downto 0)  := (others => '0');
        bus_read        : in  std_logic                     := '0';
        bus_readdata    : out std_logic_vector(31 downto 0);
        bus_write       : in  std_logic                     := '0';
        bus_writedata   : in  std_logic_vector(31 downto 0) := (others => '0');
        bus_waitrequest : out std_logic;
        irq             : out std_logic
    );
end entity data_gen;

--! @brief RTL architecture for LBUS interface
--! @details
--! Data is generated and presented on register with offset 0x0. After data is
--! read, interrupt flag is cleared.
architecture rtl of data_gen is
signal delay : integer;
signal data_index : integer range 0 to 255;

type sensor_data_t is array (0 to 255) of std_logic_vector(15 downto 0);
signal sin_data : sensor_data_t := (
"0000000000000000",
"0000000110010010",
"0000001100100100",
"0000010010110101",
"0000011001000110",
"0000011111010110",
"0000100101100100",
"0000101011110001",
"0000110001111100",
"0000111000000110",
"0000111110001101",
"0001000100010010",
"0001001010010100",
"0001010000010011",
"0001010110010000",
"0001011100001001",
"0001100001111110",
"0001100111101111",
"0001101101011101",
"0001110011000110",
"0001111000101011",
"0001111110001100",
"0010000011100111",
"0010001000111101",
"0010001110001110",
"0010010011011010",
"0010011000100000",
"0010011101100000",
"0010100010011010",
"0010100111001110",
"0010101011111011",
"0010110000100001",
"0010110101000001",
"0010111001011010",
"0010111101101100",
"0011000001110110",
"0011000101111001",
"0011001001110100",
"0011001101101000",
"0011010001010011",
"0011010100110111",
"0011011000010010",
"0011011011100101",
"0011011110110000",
"0011100001110001",
"0011100100101011",
"0011100111011011",
"0011101010000010",
"0011101100100001",
"0011101110110110",
"0011110001000010",
"0011110011000101",
"0011110100111111",
"0011110110101111",
"0011111000010101",
"0011111001110010",
"0011111011000101",
"0011111100001111",
"0011111101001111",
"0011111110000101",
"0011111110110001",
"0011111111010100",
"0011111111101100",
"0011111111111011",
"0100000000000000",
"0011111111111011",
"0011111111101100",
"0011111111010100",
"0011111110110001",
"0011111110000101",
"0011111101001111",
"0011111100001111",
"0011111011000101",
"0011111001110010",
"0011111000010101",
"0011110110101111",
"0011110100111111",
"0011110011000101",
"0011110001000010",
"0011101110110110",
"0011101100100001",
"0011101010000010",
"0011100111011011",
"0011100100101011",
"0011100001110001",
"0011011110110000",
"0011011011100101",
"0011011000010010",
"0011010100110111",
"0011010001010011",
"0011001101101000",
"0011001001110100",
"0011000101111001",
"0011000001110110",
"0010111101101100",
"0010111001011010",
"0010110101000001",
"0010110000100001",
"0010101011111011",
"0010100111001110",
"0010100010011010",
"0010011101100000",
"0010011000100000",
"0010010011011010",
"0010001110001110",
"0010001000111101",
"0010000011100111",
"0001111110001100",
"0001111000101011",
"0001110011000110",
"0001101101011101",
"0001100111101111",
"0001100001111110",
"0001011100001001",
"0001010110010000",
"0001010000010011",
"0001001010010100",
"0001000100010010",
"0000111110001101",
"0000111000000110",
"0000110001111100",
"0000101011110001",
"0000100101100100",
"0000011111010110",
"0000011001000110",
"0000010010110101",
"0000001100100100",
"0000000110010010",
"0000000000000000",
"1111111001101110",
"1111110011011100",
"1111101101001011",
"1111100110111010",
"1111100000101010",
"1111011010011100",
"1111010100001111",
"1111001110000100",
"1111000111111010",
"1111000001110011",
"1110111011101110",
"1110110101101100",
"1110101111101101",
"1110101001110000",
"1110100011110111",
"1110011110000010",
"1110011000010001",
"1110010010100011",
"1110001100111010",
"1110000111010101",
"1110000001110100",
"1101111100011001",
"1101110111000011",
"1101110001110010",
"1101101100100110",
"1101100111100000",
"1101100010100000",
"1101011101100110",
"1101011000110010",
"1101010100000101",
"1101001111011111",
"1101001010111111",
"1101000110100110",
"1101000010010100",
"1100111110001010",
"1100111010000111",
"1100110110001100",
"1100110010011000",
"1100101110101101",
"1100101011001001",
"1100100111101110",
"1100100100011011",
"1100100001010000",
"1100011110001111",
"1100011011010101",
"1100011000100101",
"1100010101111110",
"1100010011011111",
"1100010001001010",
"1100001110111110",
"1100001100111011",
"1100001011000001",
"1100001001010001",
"1100000111101011",
"1100000110001110",
"1100000100111011",
"1100000011110001",
"1100000010110001",
"1100000001111011",
"1100000001001111",
"1100000000101100",
"1100000000010100",
"1100000000000101",
"1100000000000000",
"1100000000000101",
"1100000000010100",
"1100000000101100",
"1100000001001111",
"1100000001111011",
"1100000010110001",
"1100000011110001",
"1100000100111011",
"1100000110001110",
"1100000111101011",
"1100001001010001",
"1100001011000001",
"1100001100111011",
"1100001110111110",
"1100010001001010",
"1100010011011111",
"1100010101111110",
"1100011000100101",
"1100011011010101",
"1100011110001111",
"1100100001010000",
"1100100100011011",
"1100100111101110",
"1100101011001001",
"1100101110101101",
"1100110010011000",
"1100110110001100",
"1100111010000111",
"1100111110001010",
"1101000010010100",
"1101000110100110",
"1101001010111111",
"1101001111011111",
"1101010100000101",
"1101011000110010",
"1101011101100110",
"1101100010100000",
"1101100111100000",
"1101101100100110",
"1101110001110010",
"1101110111000011",
"1101111100011001",
"1110000001110100",
"1110000111010101",
"1110001100111010",
"1110010010100011",
"1110011000010001",
"1110011110000010",
"1110100011110111",
"1110101001110000",
"1110101111101101",
"1110110101101100",
"1110111011101110",
"1111000001110011",
"1111000111111010",
"1111001110000100",
"1111010100001111",
"1111011010011100",
"1111100000101010",
"1111100110111010",
"1111101101001011",
"1111110011011100",
"1111111001101110"
);

signal cos_data : sensor_data_t := (
"0100000000000000",
"0011111111111011",
"0011111111101100",
"0011111111010100",
"0011111110110001",
"0011111110000101",
"0011111101001111",
"0011111100001111",
"0011111011000101",
"0011111001110010",
"0011111000010101",
"0011110110101111",
"0011110100111111",
"0011110011000101",
"0011110001000010",
"0011101110110110",
"0011101100100001",
"0011101010000010",
"0011100111011011",
"0011100100101011",
"0011100001110001",
"0011011110110000",
"0011011011100101",
"0011011000010010",
"0011010100110111",
"0011010001010011",
"0011001101101000",
"0011001001110100",
"0011000101111001",
"0011000001110110",
"0010111101101100",
"0010111001011010",
"0010110101000001",
"0010110000100001",
"0010101011111011",
"0010100111001110",
"0010100010011010",
"0010011101100000",
"0010011000100000",
"0010010011011010",
"0010001110001110",
"0010001000111101",
"0010000011100111",
"0001111110001100",
"0001111000101011",
"0001110011000110",
"0001101101011101",
"0001100111101111",
"0001100001111110",
"0001011100001001",
"0001010110010000",
"0001010000010011",
"0001001010010100",
"0001000100010010",
"0000111110001101",
"0000111000000110",
"0000110001111100",
"0000101011110001",
"0000100101100100",
"0000011111010110",
"0000011001000110",
"0000010010110101",
"0000001100100100",
"0000000110010010",
"0000000000000000",
"1111111001101110",
"1111110011011100",
"1111101101001011",
"1111100110111010",
"1111100000101010",
"1111011010011100",
"1111010100001111",
"1111001110000100",
"1111000111111010",
"1111000001110011",
"1110111011101110",
"1110110101101100",
"1110101111101101",
"1110101001110000",
"1110100011110111",
"1110011110000010",
"1110011000010001",
"1110010010100011",
"1110001100111010",
"1110000111010101",
"1110000001110100",
"1101111100011001",
"1101110111000011",
"1101110001110010",
"1101101100100110",
"1101100111100000",
"1101100010100000",
"1101011101100110",
"1101011000110010",
"1101010100000101",
"1101001111011111",
"1101001010111111",
"1101000110100110",
"1101000010010100",
"1100111110001010",
"1100111010000111",
"1100110110001100",
"1100110010011000",
"1100101110101101",
"1100101011001001",
"1100100111101110",
"1100100100011011",
"1100100001010000",
"1100011110001111",
"1100011011010101",
"1100011000100101",
"1100010101111110",
"1100010011011111",
"1100010001001010",
"1100001110111110",
"1100001100111011",
"1100001011000001",
"1100001001010001",
"1100000111101011",
"1100000110001110",
"1100000100111011",
"1100000011110001",
"1100000010110001",
"1100000001111011",
"1100000001001111",
"1100000000101100",
"1100000000010100",
"1100000000000101",
"1100000000000000",
"1100000000000101",
"1100000000010100",
"1100000000101100",
"1100000001001111",
"1100000001111011",
"1100000010110001",
"1100000011110001",
"1100000100111011",
"1100000110001110",
"1100000111101011",
"1100001001010001",
"1100001011000001",
"1100001100111011",
"1100001110111110",
"1100010001001010",
"1100010011011111",
"1100010101111110",
"1100011000100101",
"1100011011010101",
"1100011110001111",
"1100100001010000",
"1100100100011011",
"1100100111101110",
"1100101011001001",
"1100101110101101",
"1100110010011000",
"1100110110001100",
"1100111010000111",
"1100111110001010",
"1101000010010100",
"1101000110100110",
"1101001010111111",
"1101001111011111",
"1101010100000101",
"1101011000110010",
"1101011101100110",
"1101100010100000",
"1101100111100000",
"1101101100100110",
"1101110001110010",
"1101110111000011",
"1101111100011001",
"1110000001110100",
"1110000111010101",
"1110001100111010",
"1110010010100011",
"1110011000010001",
"1110011110000010",
"1110100011110111",
"1110101001110000",
"1110101111101101",
"1110110101101100",
"1110111011101110",
"1111000001110011",
"1111000111111010",
"1111001110000100",
"1111010100001111",
"1111011010011100",
"1111100000101010",
"1111100110111010",
"1111101101001011",
"1111110011011100",
"1111111001101110",
"0000000000000000",
"0000000110010010",
"0000001100100100",
"0000010010110101",
"0000011001000110",
"0000011111010110",
"0000100101100100",
"0000101011110001",
"0000110001111100",
"0000111000000110",
"0000111110001101",
"0001000100010010",
"0001001010010100",
"0001010000010011",
"0001010110010000",
"0001011100001001",
"0001100001111110",
"0001100111101111",
"0001101101011101",
"0001110011000110",
"0001111000101011",
"0001111110001100",
"0010000011100111",
"0010001000111101",
"0010001110001110",
"0010010011011010",
"0010011000100000",
"0010011101100000",
"0010100010011010",
"0010100111001110",
"0010101011111011",
"0010110000100001",
"0010110101000001",
"0010111001011010",
"0010111101101100",
"0011000001110110",
"0011000101111001",
"0011001001110100",
"0011001101101000",
"0011010001010011",
"0011010100110111",
"0011011000010010",
"0011011011100101",
"0011011110110000",
"0011100001110001",
"0011100100101011",
"0011100111011011",
"0011101010000010",
"0011101100100001",
"0011101110110110",
"0011110001000010",
"0011110011000101",
"0011110100111111",
"0011110110101111",
"0011111000010101",
"0011111001110010",
"0011111011000101",
"0011111100001111",
"0011111101001111",
"0011111110000101",
"0011111110110001",
"0011111111010100",
"0011111111101100",
"0011111111111011"
);

--! delayed bus_read value, in order to detect change
signal bus_read_d : std_logic;

begin

--! Performs read when register at offset 0x0 is read
read_proc: process(clk, reset)
begin
    if reset = '1' then
        bus_readdata <= (others => 'Z');
        data_index <= 0;
        bus_read_d <= '0';
    elsif rising_edge(clk) then
        if bus_read = '1' then
            if bus_address = x"00" then
                bus_readdata <= sin_data(data_index) & cos_data(data_index);
            end if;
        else
            bus_readdata <= (others => 'Z');
            if bus_read_d = '1' then
                if data_index = 255 then
                    data_index <= 0;
                else
                    data_index <= data_index + 1;
                end if;
            end if;
        end if;
        bus_read_d <= bus_read;
    end if;
end process;

--! No backpressure
bus_waitrequest <= '0';

--! Interrupt generation
irq <= '1' when delay = 0 else
       '0';

--! Delay process
trigger: process(clk, reset)
begin
    if reset = '1' then
        delay <= 10000000;
    elsif rising_edge(clk) then
        if delay = 0 then
            if (bus_read = '1') and (bus_address = x"00") then
                delay <= 10000000;
            end if;
        else
            delay <= delay - 1;
        end if;
    end if;
end process;

end architecture rtl;
