// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hYml/bvZBk4ZU4ALjfVT9DBvisB46+gXFw0RSQZwPwRHMCChoeCF5SEPBvtibWub
OMPjp6z5nQzlh+ARsgD3t2tP+OMr/5b6TdGBE9dpKDBd7n1is/OmthRcVHDuRrsU
au8NO4spQBHsuxduBqWt2lVI7KIhBbe46R77pjgfN64=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 77776)
tCNEPeONjV0hjnrgeG2aGcHui4SXYX2FcEF42ID7NRHKCwDLb/a9oR2269EpIXs2
4BGPnEFmueXf66zZhpvywIVqyaEFuIDsP8clBp/UwLY1MPJR1X/0Wo2Uz9bsVueX
Fjm16YGCiN7nkl0AseNA/1D3Gsbr74zaMTTPLWShM5s9vAdd5OIsEX3/uKdtF7PP
gzSAACSNHwdYs6IdZbwoMoBQmeu/a5+ve/9NRgRjgZjQRTJ/gowpkioqu+cz04wN
160I4agDNx9YOQOiRAzU82J+QqdIgDu2bI8I9JQcXHRHbdbeEgEZY3CnBzCbCJOm
gldZa8J/zV7yN0siTmbhjCKCcrZhQYzGZLdM0CYY70aXyxWYbSWveUe3W3YBde/1
unYCRp8n18Q4RG6fs6jEEGyonl6rV9MRpn7WRBGJ5l810q26MWkN/iMo6BgWqO48
PE2tu54HLHaElMsAlrbGAbX04/w6eW5dg4reLeAfnYcCmGn2e5ywFQKRfvA762l/
7eT3Uj9AIXBH6hI7KyUrNt846EjdmnSgcHSUuEOkbPYR/dtgRIiZWyXUfg13gV7s
Pb8Z7wY60o4HmZ+1iIfgHazs6u34TNvCjW33QU5U0qDL3gU+dDH5wwFNV2C4+89b
PkN0pBlu+vGu402Cl68kkF3BWqox6Apnzpu6mTm06Q+EOz9tZpy/tWuE14opZI9s
C6da/rt5kp0eaJgmsg3wKaLh3W7uELen6heLTlFP26rbq5f7ev+NBklRgcPQse5+
1pDBZwrCcczuf+sLrRbgDa1NOIpMbzydgWyIyGKh7uBxAzOX+IEJ64oCCdyo5RqG
+A6ltBFWIzP4Gz41Iy9zAJ7pfZtI387ICMBc+vCysIlhvy7rso8KP3ydHWS3BgXv
yOr82pXfn4A6kO/M2EWhyer3anxWyKC2xOHBmLdH/e9Euz4Qn9imRsIj0loYhE8r
EsQl67KgExNbpgxHHn8pC2KfU//wgU5EOqptDtIwt+JQ8JaQ72UdWyMXv11F3Zvm
8TTiMjcjMkstUnGIIzJ/eBWvueXMNG/MhEM6x4mNz7eufB3rdfWKRnrIOwI0Co1L
fLw4s1V+fMge3hSmJTFXpu6OPzoVYVO0jubqgPlXoduriiWVUzpusnRQ6vTw0BUs
uZX2HZCpg1hZBrSXQvveaEqetPRscTeIZE1rgtmM8Qjv3bUzYNT8fb/MqlUfZJf6
skKA88+f1r3EKdJlZvE/iAcaczZWPw9F5izZnXKbCRqZNDVKT0OAzQVh32FD6KCX
TvlcZiXTEQCEsGaSVIMAfE1f8NUfqmZk/vc6EE4NisoKn3FghdFPc/xtBKbeOQME
fbThp3AxzzR/s2xZUYta1EvlsyKvU7RJGXjRKzNB5pC4hNiu+rjoyQK6brBSxfhM
93ptiFVXsTKEEd6xEI4merZYL8sIYW/hPGZ9o5ULOr432e8yh+FesljJ0RTM69vc
SC7W2Sr59Rxq4QqB6aU45YEV0BpOi+ngYDCWPhWhDMFd2gszYY0Ag3HIn088zrXS
6Qa+om6rKgYfbqZkO7YNYFsknOQuEm+RCdQjwrYvDlRGTMGoffHfsnwyt6gsTvAN
JNAQdl13AtacjA7mD0D3NtkbaNFxmJFxn4uLl3fTmPrd4CIheA7Ko65odqZBRlkQ
BwGLhPmVxrdoGSaO0kT3FE7TkAZPdEHBop8sAKnTamgbZVZmfcFc+kZ9UoIcdFW1
BptIz//DTfEkgrAAmPMHuIiXJQea7nXyfdqlfmEiC5oaZYbvHU9KubFiZUJmP2DT
By0+RE6XMuQXoSX2aZcqbY9oX1eL6mfKBsUGD4bX4usw2RxVFZrXZqpueHfP9IxN
cBqT3p/XL3auSMAFxeKW6hrg0Q7bLP9Et453r5OhBh+yJZO64ssz19RJaVrvrRD7
fghrfjI+tdmlbGrZ5J14fgR9OU0Q3YMqf3K6zDNu2vwcwvKX4GugQK98vt1o0yGH
CDVGYyKnQo/ZYSSHL+xzPrLMN2rz3GPJpgOZYGDrgA0O7CNaN2wRCb1fASBDZKkB
C7B5uoHOm2bfKS2N96KcIoyxHa2MIvtl+rc6G2pGUmJ6q4DpwsxCOJdYn+g7XIww
7IqUpGFIJuuNQhCabksacWNGtJA+ypYaBB21rC6CnbHqVcqpelO9t5MydK6euq6J
CsGUXSEZC8LW5WzovlM9ZLVUenkczFfIgbUXYH2exk/Oeex503JCLOcTU9kY+D9W
PzBku3OSrUupAXvcJfXIN/v1CETt1jmRfI4gr/lGXdMr7aTrQjEojBeo7z6zEK1p
hzE9Wp7fGRos4IOdLzVh9HTl5WugkerhwhI42U4Jdbqk5A4fxnN6rVr7dlWuJ3EI
KIgyhuX51Zs1EgyBzFLlWzM89DmS9GzlZ7NZSqX/DhEEFGzO7Ima4NM5yOwWZv4E
dfCbUPbff3Tqcds+Ndv/FDYkHiZZjbE2BkQZeAv8AxAPp1KNh7tf4v50qfRgjD+R
YbPY9il0IlxsQMgd2lREX2jJMiLZaKtMKaPcqtzhWa6RgYe8INxXX5KnPTgcr+aK
etoWB41Th4iOdKc9yCDWDhMVOh28gQgUmXYstL4gaWudz950XVkVk/Z62mbBK2VS
uFrDdXPlhQa8ZW1S9xVv/Ibn7bvJO78x4pwtR0q+4ur4qS2ugKrlQ3a5O7+5Xc9z
vjWSevgukAdvExnO2jj9xZE3daLRDaGBmaEE0lKxWCb7fjigBQJQdFzVkFAjTqp5
ZJ3Rz4SZDeO0+9fW+5f7QpNT0lofCPfXySq9uhQCtJp4mzuN3LqM2FcSv7BvBhMF
a0loobKJWG3oaqdF3FO+lzrfho+gmxx4M89ZSCXQYtiUv5DLtwY1Zy054+dARJtA
Wkx0XCWCZBl19gaGIb8Ulvyo3YynwfqxOB9D2uTyDz72VeP8pzL++VEzMC00eafb
QRMxxZqTaOM2X5F9o65hWDukFHemBG7eTjhfWE8A7gZ6Cf4otSrIiJaVsGli4KRB
R18V5tTtB3V3mll8mdyWj+kD81RLoJ3yMDviso65iPgDTyKwXgn9W3aYyhp0Adw0
MXQsqAxthRMz36sg2wkSBcc7T62ikdaABYbkjnn0XTC6zPKuKoqoOrYAYsNjYPmF
3ptm89nMkUPdJ7q8UiXenVdRpImPoQVGlgfguWepKQ3LwY/rqrPBkelxey/BcPZv
gFCMq5va4RTG9SYPZHeJRIiF0BvpEXaTdpdOlPnzGb8gqmQP0TQziCXxDbVvc6DZ
cplKLuM0i2pq7Gf0LBJ6CZsKr183G24J2A+OXxGtVv4jRwrTaiVE3qQ+ObUWtHda
5WzfwX1AoxWirA/0YjHfNrMHwcCeqcR31VUtVegT5FpLBcOOjXApNtWYXQZXMZN9
2o2IeoZNPZ7X+hNRRsBCzTf2wHXT25g3ePTwUt1tTPKrQ8lchL+YGa+Y8J38WKhP
fKMVZMzFhLDxyQfYOtGTnbo1K17B2fMmmC9MCyzP+mUUdtaP/ouEJIIK3y99EEXY
REbjWr+2PwGFBCkLVOdRJ18N1dvhXrtJrIgizbw6qgIIPAztgnxvoWCFmUfZYVqg
4u09ib6Opjdg/xQ994Yl7lmd2upSp+LnXFSW6WM8YzA31t30SLdTFs5+FGzQe+vq
bIfEaxHyvaEuS3TsBPZvyBFXyMF4DXRJBqTawu9R1qvZPH4jBWo2u0zwjk37fjgo
isFC/aW/AHoSPMeekN3tFfxoXfRhik+rS1FLZUY9ajbFbhATduZ4rVPCqikxEA1f
KoXL/N071bvAbFo9kP5e6vo6ZbfTfLgFg+GbpZHQjmhwI4jADyWijYAsdCxrca94
dp5c2KDjTvfwZLFPqTps+X1AJMYRYGcS0MzybaxRWJ7/TNydiYGs/tP/y8OJmkGw
I1t+Tk/6dfpIlAp1kHqZB6S8uDFZ7wqRk/n9NZC80hOiaFWiHeedJuOv94SV7Ic+
ULaxudSUqMT5DApkIb1VYy5yTn9+kctSdqunydlxz12Ka3tQ/KGjn3o8r7y54v4z
LwxsHigL64Ucls9b/fEkw1Ut98H0UP3uKZgxxFwROvmREPKHjOndzi/olMQfTYlL
TyMNVEz6OU8u9YJyzxdi86bb1I+DFS4QgMB6X2R7x+G/1yh1duhxWkUFhHhuhnq8
zeICgR92PgQ5hHuMyGlBbQvJIk13hBXN191I6ecJLygIvobgMGbjygMEIXdrKxLS
AoIVEgYdUbjOYKuu3MEbqhQZXMURdWw+HXDoFB4D7obJ0snr8S1j6zVOhL5e64yb
Gyf0a1FL3RwM/LRTVkoHhXQyT9G7XJWLcpMrWq5ymGDpneEErpfeeWWd2X82nqGm
bQSuxq0DdXS8/dY5YluD7t9S2Jindk4/VkDytRZqQrer5Islgyf42buR9Z8BWVA9
cFafTP0IOlW6fTvK6qbv4bNuLBUsuvQf/1Y0SymNsKQb4MQfU5k7d1v1GjGEEbwV
9Aq3AT6J8HDVVkr/qi5arbY6+mU37OUnnGXOvl8Jo7FbJEdfD7hvW5yxez4jD4xY
OkU/3qB2WMTA+VHpxcqENT5LKmLsBVdIQ+KipqODx+8h5dyh5DYT/nUC+NK5tNtr
sv7pKPgdijSBKujK/p4b9D+PFJ88UTnZ9VuQvyomzTFhqSIpWrOn63qM5hWtF55C
9aoTFhQP+m/eIc0Uufx0eZ8/3+ExUihHwT7uJzvhV08MXoJ69dvj0WKAHx/52++C
NxO1UMa7wQdc+Pt9MKjWJJLQq5em69vSzBpcd4gqAaztIyoS9g8wn4bXMYVyVIQ3
zt32N7fO+TVClew4q7yPQNFQCqU4OyshCgd1wfiKXD6TZ8cgBiS93mozahAWrDdT
mv7JSpUcTiqaldO3OZvy/eowvUBQEGnB1+pNCc/7bJBwg73t7xAWpch9WOYcw0/Z
Ct/5wQVeBetwj6zBapKJ8uUnfGmISP72kcqRZA56WQ5pglw7xaRRkxQMFjKCxKQU
XU5xHtc4J4X8LXNLGcAMnsiP28XMSOGphAegd5iy2buEHScfW9rkxSYfamN0MZVe
/3l3TD/EauxCswJZlPTxeh1M4CTqkI00+0jj7GpYun16t1s11QPqVxhBkQ14d4Id
UUg/AA6hCzuyP8ETr2SdBAnNumleB+qXeqU8mB4TOP+4LYpQYqD/+IXDrA9b7WVb
aGTPwFWi8Qssba9ELLEjTh4/cfGvUxtni9MZFbeEYtKzPzd/xs2dx8IbxIU1s/p9
jnl/51fh1mE00cibB8QjHMizWscolaAtCnIBeVx+V/uvY944yIRihaQsf7/KW8ZY
BLHwdvdtjEnlJ5KOY7L7p/aVNqKI4PA4Oe8gri+TWsT3HSQ4pZIaiKUEc7AfXV1i
J3iZfq0J5TixU7XVDw2WyVc3DgCOzDqUzELVZsMxVZ1GCTjDDynCCYgnDQiEcbxS
BYZjqNJpDY610u6na58UBp2UHPH2eaallCMKdI/Ota1Aj83VxZABCldyb8imiTdM
RKNNMNY/n9qlkHMxutUCVaXUJxk/nLQD7D/IxIzjW1dkD+qoJh0kzLs01BJchla0
sMEvAfGHcruBMdmErUZK0Fu7asVxaEDGRAqazc4/OHMJnsMvtYaU2TTY6r68zBLN
66lH7qNgQo+GCNmpubC+a6pjK2PRWI1WOxHE7ZhsR3FPrcheHZHGbgjCE8OcPyzE
w6TvwuFJQQupSaPqC4X22d6FREe5Blk4rrLed947sxKUTqUxC/JXy6XE7MgyITVd
lpxYgWtcD7G/L99XFi/l/DjI6Gw83n7in3zYEONkaGEt6ORz2d3Uzb7pwazSliss
DX8tS64edu5papks6SlFkgAVEeAibBXX2WD0rYqb5bM6GQT+3ILmNg50h/H9wmls
MgJTM3usDoO8/PmJq4ua6H6bndF7nqmsFhFbso+8fkigqxwLlrCHhQrMbwcs9mwe
VLgB3hJiknOESWFjuqPRE/PpHuTpKe7TsncHS+6bLbSFiNNE1V36K10p2tSbiAK6
pkCezS4XVw1mSVCStT8i5jXm7i131SZvIvoy/H++Y9LJkubWUfCsETMj3NoBpyxE
Z99IctUl7jBKP42fYzEVLYcxYbVdlQVPVvaoV3+9TSPy8LqpI2558OkBprwB27RG
sJLC2RCozM6O5xccI4QzApF2cgvRFflwIL8ZGtHFSRrKOMdefNElW4NPo5kD+t4B
oCV2/m15icF/aeN98wlLvQb+RLyf0ruIZ9oG29i1sqxUwuOlFAsDm1bCAO/a0iR/
iiCvLLqesue7PUqDbjOQ2dCO38cV86NS63OAGUq3zjn986man1cWLMa6D8WF+/da
u+R/sdK7mS0KC+EU7WgoLca7rTJxuHACXFdZkxdO1fqw/eN0+ecx9FpqW6HFvn94
KHg470h357iDUFWRRQ325ljmvssSuq5Znc2wgkUzCJj0d23iy9ed4RoEYvVhO6+l
s30U+EwKo0ZOIJR3juTabx+vps7B4w/ahufv99ktfs9fk1cBX5GNH+xCCVovLJEF
VGsBAWewwCFlCwb+qvibnJpN261YPjtJ/Fby6OC6H6mCiRIJihEejNLuOb7ng4+R
UR6n6DknnopYnpbXMjrRlp5/0lg8ieP6QvBYTJ9PDqv1t0vKVgW/9yO+IbHXnP7i
XD1Zgj5sw//e0Hge7mejUZsH4uNJsTIs9bGtLZJklkbP1JUktuDe7jcKPUJ6JNK8
BwvY+KN2ERwdJaHrgik1vvWLW7cHY1hsXHy9Hv4wmtlyIe4BKqPBabldkK2O2ZXy
aBDz3W1WAtrIqtOv+vBWeEGQm6hLYdZBT4SjwepUD4b2wiYW1rW3kdFP2Qht+RbW
HD9RlbN9KS/7fexHEfl5Ls0bx6qs45thInCTlCvxaGcj2xFjdxngP+6c5SAkKFJF
dU/VQOs2sorgjRyUoeMwEai9q4nypiED0l/KV4Upp/4VUK6/PwX05s/l0sJPC8az
vQPQAidctVkV3+qNUV7noUd4HuhZSjoeIG4wnElHg2IisP/cV6sPDty/kctUVxXR
zvY1ic2ZhY+g0n2GXKio//FP0QQSIh4paYgjlnQKFArjwTssEd3dAgyqVVHa24DZ
bJ0qHG2x9dVwW/uLCGAbfsaPSG6FCQEeszkOUosro4feUCQUp0hyLgE+V9g1OLyj
H6p4UDuY2T+9zlVEztNqLuTE3O6GPFiUzKAnuaOIcwmarQS4mV1l8/3+3SaywB/j
ILxmk2wDr6UHzobFXXSE6dzKU1VGzE7f2I3uyTU2uT0OLy7yI/SGGseG/ytep6cb
lcr4nwI/XtJt8x3/RRzwpUiGCF6BsaPWkQZIWC2N0pzPdO5UlMYdBaK/+djbdAQq
q4es6N7NeXGc9ocYkoffItZ0ZrC828voq5RnA/hQM4Q8zbLgREwIsQvJ6YdWcQGN
IxgIHsJiDBdJ3aq/pHRuCjcx4UpbdztkJbK8VLk29ab51cZiB8GqoNKxQByAq7f9
zBqddPaZIy1nKOaDtKO9bnKYH90JjGBra7Dg4107RkQ6Kzu6RNaG0xOoxfJcfAQd
Ia7qmwUlfdA8/duxjon2FLlsX0+RQPEaSzrV2nvuyO9j9HsyG5hgojQsbc6vkc0d
/YSIJ99onddPOccIIoemT+mGkupFy48305GlpDFsb5Ga48j9VFzv97DBly2kDADz
LL11r/3gSSsrcEdJrvKDQIwwGpRmdT2NWhGdFcyjVi5e2H7Znhpax+PvAb0NKjdx
+YAIDJWPLONQJ67NrU7zfFM8aZQG0Dxnw7A+fTHEGnC5oYAp36jbm2qAVN8p4umn
CC9xqL0gb2ChwoHp1c48WsjFEeLn0w9GLg6b99zfDDmKIlbwRettKh6OB9hQNfo+
zZKVQp3n+s9UJgWNX9D1L/9gLtKyil1x8Q5noMhlklXQfTme7foVjFu702v7fIo3
SXOwtDt0/G3Rg6d3SZWqXWhSMO7wmTt3yrJItC0XHE96Y4lfDeX9woVD1PikUb8M
DsPc0oVbK6Kl9A89pfaote41iorG9PLAY+oS9fmEOALjILoGeWpph7xzyXjZy5vo
wueEimslmBiZ/tBnzg9vIPI5EdEITmouhijIpQvVz0zveAePoq2ipT7HvYfuLKgh
AheBepvzjZQN9zxV2Xr9mXLh0JPJmRx0zHgwLlJBSqMSf/1e/3cBcxE9oU4moajH
yf8NrxM3hSZfHCUnB+n/kCnewEPWz+aNx8sTvujl+MwFdXdFqWJjJgqjMCYdXYDE
8xBmX9vLDjqmHzrpIzsdxc0r6sdkWicRWOzGhTwfSanXArYQVy4DfMXce9e/q1rm
6nIzSCFq3IhYfYTyflL4m7bJgNkstBQmxVGl0sWGWptg5lKWVKpRXrhCC6imRnP7
iWEXeaFeUvaiGLAaIkocpIOEL9rMhckHWc3a2z9j6Lm62kgI4hX5IfDOYNaXmzVs
W8hGwQGfVbTf050gNnBjlr1lDGm3HWcCogK/PwG0jsDKF6qORq5g26l6jHV6mngt
7WPpv3gr2HpO0T5odGJ9jrFzWz5CjGBIU5Ys9L5YUyHB+eZ69ODRzGlLhsDqVxD3
OIxRsxnWheabNOAV9O+pNVTZNdEq1nmDaGOBMtIAJ6dGQc+kTaTB4YVe7WiKvzjR
qCHRFFTWpwhgeh0GESn43C2YQxHXT5mftp4kWwlQtSax3rMLob9hqgp0k/FEIt+h
YiTFm5pi4wpQHkRRtvWgnCG+SnuGJztWXPz/pD8bom5tBz706Uxv5a1AeKwqMmoO
++81bXb2AYpy1kzlOznmw/fH9UE/b5QlCl2qGB0K48eMn1X7vJKlwys21Sq/3tZA
PENjGOH1o89Wf9GSvzIzikl/rk1NiPCVa3X6JDltheaFnEz6lfSY0Nntjtlw8ZH7
fKrZcsl7TP7Eli/oOyUGC+Te2rS7mq9AwD9buzU5PdUbvSfduCwy9TNnh7kYoJVp
WUb88reWpFFEuGjo5HUyNz9TGXZDlZeDg+VdOvG75RvxEORlMmGxrKC7p85pNdDO
FA5+Cc2Q720KEC+9TWeG6rZj2Ibewz5OVJzLa0tgyTtuULY0DDGM4fHTG3o7cA1H
A2RuXHMbx2q3kIT28uq7/ztEJqvBpzjGcDMvgDu4MKK7P6Z8yDB2q6EJlTkdxgBp
g137MedHrROhi0I7MJPNYa/dkB3gjUhaXmjlv5DTDY3gttP2Cla3G+H7U+X071gI
0U6OiimR7p6SW4leOmBlPmmVdE6yF9T//xy/sJqVuPcyc7o6764NMph+T7m6ftXp
h/7s7iQPIFVJTqtkwwfv2NM6nwM15XVVKGtNQO9pfjszUs/2r9vxJxN87N/TMcsQ
wTeCndGp/PD8s1K455UTBwyofmFWdnJXLkIsZ/rUfGtyEK8ywWBgXpZSmESJkmN6
DIgxak3i5W5X0cLiQzidiObhKCixVcuFioHVqxH7xTm5kGbcmj3IoVJh6YXHx0RQ
Sh0g7H8JEJRbCEbp16ymEEuzVIjORpvmaeXL7HDm+5q2Nml72Dc0C3/A9Jrm8DsI
faqR20tuidofBx6HOrvn0sn1GJv1AfNcwTbf9eVPvQp1VKhNXEP1n7S0g3C5Up6E
5F+cIJMJoCUVw3w4bDtl2UO++uv3arsDd+JfaSj7B1RlffSJva6I+06Qm8NA+FQa
yLDlJwYIutJx/VkYg6ht5HxxN3m8ELig0wPWKb8VrGyljgeiVl6c8Ddxh40F1gO1
ph6ym6XyjHqdbO/0wckTTlWifKilb3VTiOu3SAm0INF5J8OSbigaksbXP/PrEWyk
cfD0BaZTY82GfyVPsoRUz4Pr4e62aXX5BM7bTRv4M/3qeqsP819F29JT8tLvvp2Q
2XTOmA6SDW/JJIgFvxTQLSLQVwpXjibaZ2neimbjrsIGiNFl2Tnkw3wmMk8f3Cvv
Kz6ZfqC7hERbFJbYHlkcVY6tOQJ+dxtQF7/39RTiISGmPveOzYcA+oYiaXElswNx
sYeNN5FC3jG4UhczSE0+TymifbjYpiyS653R9Y4Tb11ReIpE6Szh6eDfDfQKm/Io
Yq1pySbd7le2uyGC+5zM9RIA8waS1Itz7SVNxvoZmyp9P3Q3w6y1ArA4snoLDUv4
15eUwQhCcA/kxg/eWDis+8N41PCAydPFBr8uy1VeGVruOtecR3FTsPeEdBy+f7D6
9YRRPQv2zwwjY+CJjKu+AQWEKLBT9gvOw5Z/Zgrs4FgQCU8D6CW2dWEYXo6Xgdfx
6Sd6f/OXQv1qAm5Uiwr9dlbsZXYavhrLARtNk8OQMCd14IGBMS92Vvu/qGCZ4W4e
KTLM749BG3YjcOh/t/S6w3dJh6nnMvjNi+JSh+tIfLk343MdhXiWx0HcrT1bHIun
X39In2vsWRDHqW4Tr6YCFUbJuPb69dKXagRzZRarVmpTl4d9STKYd7pQ0Su4GcXY
CTj3HOcsXHNJpKk+2Fw/I4zi3g8yDBfFVnDhHzrg2UK4ItZgvDzOZUwi3Z6SuPIA
Sqkq/sTYwKMv98RkXtGFdlJ9EEJLQAyC9XlUCbWRzXtZMHFkTYIS3pFEQZHVurQy
7JIxSjqfHl1TIOTiHooWy7YgmYTfAeOFFia5e6sLuaGqoOdD2+1nDOZ0bZapqby/
I179eeltG6cj5bSnimFK1ah+zHWNgWKSVjrSDqvS0PEl9xFseZHZ4zLUyMI31/J7
5hBHBR2pnkTki1wXWpX5t1IE5jpaR9EzsQZPOYIM0C9Yz1+zXRoEz5wECYfMkNon
xMFQELW8l/L5otZnMB43p3p627j3Etgoo24NwwWoaSXNbHPnOnVIu90Os6/0V54s
nQh0wkSjNzD3UIaZFAx+F1sFZT2+XXBzF2nwOBsdnVPyc4CNkY2Ucsgo8sVrJpr8
p7mXLmBrU70eeZaOi7MJfuApCKrH8uY8nG61ZiweRpQlfVqnwR5DMrH26UgHfdlJ
yLCF3yghW++nZ1JQoz/fa15/xL6+DCRaHtXC36GtdsbtwXB1fise8uPJp/zJ2Efj
JJkXap0/4qhXmGfDKaGSureMS2WLJXU9lPKIMHn5kqc8JrBN4UaQf5bsgzYZTIu/
5juUFq9Tyd6sM7zABc9HlXcjpkoy3XiJB6qNcg7j04s3bCybftmCu3ij1DMvt6ab
xlGcGv63jKnoOPzHC6O++kZjbS5HnJTdqltkuCLfs84h1q1wZJBJYwV4pSX4VaJR
ckkMNzXerM77JVV7GmbJAs+TY30ZD3l7jTwGClpaBRBvQYXD0zne45rgShot12kK
geSqZ5JIq19aaqWWi8APohR3vM1C+Mh/9bDYTUtxAWhdh8rfjKLd9tGdEn8BjAmd
8GQJCuqg+tWKf247QPD7ftWfnAhK2vnQkLPAFgCkMNFi8fxEwbeCfaGSTmozvZGN
eRHqKbh3b34hdF3XAI5wXD+ApcLUJj9q6nqwunzEpP6mjr3sPie9J2h1BYAXGDX+
4HzrjMzosUPNbkFEBL3VzXJiTfa/0OMmajxekJeQb6PXAuwqecMUHZi4/V7N6K03
uDfmjLRkpMCFH5LYlS4k5UFWvNv4WiXC9ltk/wAzWRZ+2meZHQKtpELqYezs2tbW
qFtDXTHRXPFHsfBpo8uF/xwsZKKx5gb4Mha5xFeruAXR4AwAQyXVb1xb7z9lmJTl
Mj7p1zCosf3G4RjrCTSm/4gtfhb4D+YPIlTfaGf8mOtMoHx3ka7OycIZF8gUyOLN
hGzeLLsD++6iYZpO1xyEcGFYt1DWaLDiGG7ByWEYg94LrDfVhg4V23/AEDaL94fB
VyLUfdnmkcdLzNI0LQdkAxZ6CSTLd1ke4N/OhmJGhbHrepW7Rv8v6ZT078Oa/2YY
i3eSsfS+ZIGa8TlcpMjX8Oo/hFQ9YXrtxcONv3hkS8Li50pdIhOmQE7HzoPnHr33
R4SSH7vO4BZhPxJCFSwhMkH1H5Lg8LGnQSmRpJ+AJWcDK0rM8cHgw84n38UdSjsu
lyUFIl1hOa+nGUafeQzMSZ+jZVeZq71ySt+hHZFvH9JeLqbOnJQMHvtHcnRj9ow3
h5SZt7niT+XP97meALQPj1CEsPr0qah7q8u2uhevq3kxVvUGo4aFlub/Y7kkWC93
mUuMKDlj/5FbUOAywa05RWI5PHLFf80UdvEz6d6XnRB5Omv7/1X741JJcpjSu5IY
I63QxVta4LEL0AfkaUI894ljb7j1JposErhS85uCIFFj2B6z27vrQfoz3y0r1lll
Lorp/i8BzqQw3+A9vaiiT5pqhX8jSEggAFOF3Fp2f47maeecHmDeiRhL+FZ9OylQ
FL3CcPF2hBVqZMpRFJXbsMQhTDHTHcrVtmBYtJ/94lpX4ljYYDy9Dsbd0CzseIwW
QMJ4H+ygWeQzcwgfqaCy4L7pQSgGQuQdiYvPHFybQ8JCaazzUpcJZzwqJP3dr0LL
g+tO+WD87JdygSv58IlV86aOYhvAxcyBfPjw9PmxvEeZ80FCzNKWVnwhsDCrqVZn
zneWyoqVR59DzmzErHypimpmxD9z5lEFC/OP6lXFg8Yal+n7sLXvrLttOGxTMNEB
f7OWRnQuclQFIHoEL0EHQXI52rqA04rnx+Zim5tFS1HtlKawf2jwV9EZA0BRkAcd
+gQdQXnS1F3jSs/g0ldB7skPd6PU3OW6ob0aTYFPsc7EGxagthpAxwJ8rJz8iLmk
MYmGFx6z1oBC7t2QkOKDtMvaHyGPveGhNiE4YasoG1n4w45kvqYe/eMSVxX6m/0d
RHooT2IAogUf/L2bJQPEt9IVv65xZaD73agtMXneH9Ogan5p3wDvjZxc643buUYd
/LwKuCFTs5YAtRJtkRt485E8La8KPGhe/k4/bO2S2BBhLRGOozf1VKliYXD2KuU5
95QFvrzDUe5fXD+zMqx9DV/mrjZW2KO0zMRAcRLtBHA+AmXoKYiK/qzUNoekiwyv
JOy3UuBpBlpnZewdOxbEPGhQu76Zst6ra9n+0wFpNVhQtcR9Gr826z2+a+Qa8AaV
9gT8UW28LYdYgm6hXe6/UebAO82CQuSKPr9eIlQ3aIcHJ1d7v2IrN63i0DjhGjJa
DoFSSqVuVbevjFocEhaeX7thDgHRo6wO8ffuPTZJxI7wUHYXn9kfpNtZtjSIivY7
nIXWdkhI1LeIhFv2hSCJ4wFIlUdj37bJyxnCZ8nHp+Jfm8pvzLbbJaZ5x44ZtnYv
D+qn892mw2n7Obc9zgCbghwSb10OdEGaVlS7VhB1LMl+6ga0IqumsZlzZoH7mEdt
OiVEQGv3C6rBlvdlQcUQ5ZGYbp4lYKwkyZwEKbMnCWHjr7VpwDi+g/e3cwrXoHjB
qqM7/oyD086deFKEYjNNxJ5N1afVBUO8gcU5SnHxVP745BFXIMiu3zMGoeTnHTIh
unfwKLjwaX9B1+UF58BQp/0zpt+C9HDdT38X+3pf8S9ttshr9W/V70F7I81tFB9e
Zx4u/qq0AXgGT+JbzkUWBur3Wf9V1xALA3NXTamTO75xkc+hNKgrl16YpSgoOkNY
nkIjU1jpHuSkZWsN/gPV9HOivNnpaXORAutJaRfECgHRhyrGaHCMEmnzP4hj2VJ2
HTXJ+o9tHimnBPn5GdNe1+ip9oZd2ORaV709nincQrBulWUsBiFdJae87mMTuEq1
Y2m6TMoxC3jmYBlRpOh11igxoky+Dz1K5+3SdOKDT99FMyvSFnYbwhTBko17dm0e
JZ+sMaXMffqeM4mcbGP/mTRdcoeuBdd3jzKONhawET9y9mU40sjaP4iBfqUWquW1
e8X6PWM0sItYoXOF+v3nCZnUeU++LwubFL/1HC4FPmcJszxJColZvh/8ZlkUzJMi
xnQhDsZy/+M8YXxmFfjbsP7wjpYzDsk6hsDWLG0INXuM41hluGH1yf5ISp5hgnbk
oUIKXAMYelCaKnsEWOtjuBvJoyTvlmthRZ6IUdIW5oJYT2gm5UPBXzDkMs0ksK1a
R0XDmAqRm7dl17FzxZJKek6BZPwfgKoUE13cxiEH21R6+1bthf8BVgpYGGt+a/G6
EB2PgYHB43VKmmRDy3D0zxtF/OjKXaHuydXivN6hbYWl4tgijqEpvtY7yM3ijZor
5FVTEUatbuGAw3u+ZQEwCkMJIowxoyany1efXoG033g8K4SE34HZy8f4aAwg55xL
k7lPprmDkS1Szf+bVzl+DY5DfoS2PZDvQ+Hd1xFrUnr00qc/u3kKj7kP1/oN0gcw
VRM0xYo2RxlGooucLGIkdb7gIBhzD62TiOMwiMTtjD1UXWDgEJy+0jyQ5LXnEcpH
kHpeMm9+o/9RMcqC/HXOuSBHUh1xy6Cy52WOl503OuTQcWGaoKpCe1PcdJa5KFfi
eCivGd87T6X7o3xa6P++90UqU6XqTE51mOpfyA0jsVHGM26O5aPmDT5uPoAFteTi
etGCGdppi4SEs+2GaW6cpVWDSojAaH9r8WAu7hSvbGoKbaxyriUe5xK2bQ/SNNhW
v3j8iR591r/BLcLCS7ZKUgudU3rWoTwYZzLCjT/9nZuPVvzczPlbtLf71in0wvZH
bcvjwoHA1M4gTP0sdIQ+EkRW4ZivTR0jjPFoPcNadpyjuNY2efP9gJV0qnwAPoLJ
6nAB/ZcJPd+AIHMSgfDbh9ZYhtsX3TisNpBTUhCOklKNklp0D/g+j0jdULGCACcv
OcyJc3AjdN833xlEN288p0RA3hTFcbzsd44F2NBK5g+rAZmk7nSa6JlBt5cJn6Fn
R5JxGMb0fFU7X/QDNmzUoPpvS707pbXaY2vT8bfXhHa5x3xVz5KswVLh3DSozbAe
ZJhK0rDV5Nxygdv7ntMI6cFbY5T/cI1rZ9TTIWbBrgg3EhwcJAtDq2/0U2t3YPde
jkYnyHypoF8c9I5h2guwIgoZFuv98excsoiW3muY8pom/iLE6qxxAY3bBogJVjqM
+Yqie03qCJxvkXquU8dApD/tbUz4l55HGqYJNU0UpQZYibciNni32g/pO05+kLxt
x55NEUBEWTAU9PPN/H9ZHb5yoTHO+cnBn/hXNg9Q2hFSJMpYJ/acGx54azNKD5qN
AsoNLlT/Xo3Sxj9Y5pJd9mHWf/m1HeUqkQ019JKxEzCYLNCCGouhZwit+mRtyg1f
W+s3QPJQCrHiAP7mOy2DtoZwvrEgh//zRpOgxxPIVXhWlLQfLWQoiFIz3k3jCvNw
jynK4eZbGqjLKtyz95SaNqNysfIClNoQqQXIu+N9MPMMiPbxriP13wZo57V/LK0S
VX5AASrnCsXS/GFwUANsKsG4idwC+KBhLNOrFu2MeXTHPAZT1HYQz/KKcks9w4HM
u6UWaijLuOhXOPVnPUc1QOGCx7zMb01gJ/pXh5CzB7ehXaiJMGjyCqIL9OLkscaT
SmOL5j8xODIFHwvisKHnwAiY3mPaT//qJ3RYwbTjdZqTSSDwlc4osPS0tyFYtEdm
Y/1MGWnAhmFTU7gQ2UzAe7MPCi+l0sFIwyBIr1BFcOf5jHsNcadOjaA/pgxn36b9
YjD3RNRhZnTPYAXDo4qHLETYRumQykmPd9eySP4+IjJF8aOEKMVw/eYI/WiNEcIg
jWtPmwOv58WB+r4N3rqvt6tmVF/Ym8pvjfvdALp+HptCExdm6vB21qhVpYcp9NSf
0VQyK6G20ajSR6Ur8/TfbFmHoSJYuqnzgBFNJ4dmt80sfqsgr/S7gsi1wN+2+37/
AgfRYEp7XssE8JIWK2TptYEFFctIS/EeVQwjjAUr/QYhLmxHIK+mwszgD1+1MgmD
cmaCB9bHTwp6RjglRCW3BiJK5K0dQByPj5nhmvfvDC6kh5hYgfGoqB9g+fsFBkoF
qB8PprujbV2crMw/HjLe8ZFtvcOXBk79T5sdbbMdhzpbQQB6eNtjqZzvRFkGy685
1byd95Lw19NYb7omiXpA6NSsmvPpTxlEdDkuQcXH/HQ6TPFvrK2PuF02NPlvkhva
OyDetJIoh0UzofBf4Ii8UIMKXxqeBw8RiYC5wA2SYPA5UNuBpvXrlKDXpar2zAF/
CyS2uIEfexmS0PTk3kOFdXGgsaJd75VyAJdSzvCGJA4yt543/L6VQMHJ0XL0rGSX
snhWqWOCMgfx0uAYlVpiiUM+CZaWJGtg1hRA+hxUPNJhFRyLDZecRCF/rpPtAIph
3s80jXZK/GvYgqCDWJC2g1259KUDMwTsskBBnSC54FSd4wQlGpjvC1wYCclP5yCZ
J0G4ADUPDXeYnJbOSn5hrQd/v4VOtAEW1aGqOE6xBN4nHpQXSJ25TRvlgecjHzqU
zI90NVjqP1san8sIb9vSNKE/wZ2jWs6dIB4bfRDyqc5RrRnyMdr7qW8HQH6/diKv
YH/tpsdSkaoNHQETJt93giKdNSRAXQWMIh86EZKeK6pqzyCmuIKh/cCq9oe3MYxv
QmnHBokeBSNocPX4Rx36fJ9uMt7CiB1gxy7Ih5HwfdoJOYHk6NXCJhvs4CqGXhUq
DTCs+IJiRQRrenHf5m+OkHrkQ5f3A7cXmzUgR4NDv7ak6ZK9lk9s9w50JuTcl1K/
GtQC6zxznG5bJyhC8jqeE1Y48LfnFaXKxBQMvQtllAha+89tFi2cWnpsq3f5xBGT
dJ6eeJVDsrmAvq/jQnNdsnHU8x3J10bnlgnRBXSHE//Ry8clcR2fe75ntAeAYR4Q
JlGsYv1dSlNaqwkR7nrKRuj3zd+gWwTWTjK2zUTcNTKQgm0+3UhhTkDHDaSwa1+v
j5tGxwHe6V+iq7abFqLLQiR8jNvjjD8yFoPI914DDXK8KYtqzRJ7S1cKtsimCVfv
JfI3YHzZZKYgCV/5JnCfBVIdgc/0zUwhn/xoY/wkXga7W2RBLU7lEXX6XmeSVKYX
OtCbi9tfOKJzsovgDTVss2V1Mcum4gbKX1M5AJpIGg52uYgFwcBGLA+HdFV9XkGz
uRajpj/J3aORant7mXq0jibCN9AJxCipMnnQ1zaVg1Grhf9CdLVe8WK8tnMZUo1p
mYa6H/cnNhzGUTFqs+ej/veXQaVHGC0D1dNGJB9BdiNs1dW7Yt8uWHNi51LGAj4o
Cnv+c/Qq0r/qJZHF+312/OIzmiU16yM09Y/6z3larKSeFJckEyCvfOQCxbLt49sY
mll5gcn9DED0cbOVTxR2mJSBKlpVHcDVe7qfbTBS2EhTpMywvVou6kTC+pEs6ee2
OJKhWc5iPrOsM61ObPorzoDX9cnkIG/8jHzpOR6NQqrbYTKQdh/OwGIV6WZo5dmS
13KzVcAz7TzaBDD+ssO2CRtJ6OP585D7TOhCpVEv7CKbm0jht+Cs/5w2jHhiTI7W
Vm0nI9fdDEj5VWPYxRPCdwHtCU5Z4N++JHEIl9ylMbgNHzVaLEsytD1UWFnb4r8u
AloRTqI5GbX0/UlWde4fw1n28jbzujbDdagJDNB2SZl7Tl3Nd2ZnH23VI4w+3rcG
euzXCoHlaStVwnVHjMIQSCXciWODJxkgJ5J5LFg/UkCbFn4VY1/0sgppDwruF77+
hjipF+uco8FtjOfIP5SwY9fJBW5UDC0hVgp/GiLay5js1VVP94/sEea5d0TWMX2N
qnTqQxGwhyBOtxRNKml1dAC7kzrWR5uZhXMiv+hZmiQKiK/SDX/lTmU/UqqN7gUA
AxWgC3w9Ofx8JAq3eru2jvDRX67L7292Aa4tYS8Guj1uK5MnFB2G8Nq0jER28Wrr
9hFbgxo5usWbNLHNJ26dO2dkYZI20DUOtI+jcrYsNFyMmX9/zv75boSk9k+F+0mY
0qGsdioVsBjGR88emqmWZjhnqFOIBlSxKaXS/V2Vg6cpZAUIvtwcSmDkPjJp2aww
JCDJaQWJOSSStDOB/LS9+jFoB12ydgj+JGhItsRWfiXX4xR1izYJtQw0UvtjmvO0
7SAvrsj3pGKafQRi/1AZI1zf9p/lMVMapbHg574YN48xKUjOAlzPNMtt8VduZj1m
GRBzfKYbl31n0UgHtKUZ6Drv/Q8k0IX4b/aFp0+5jWbMQZEpQMJUT8j43TfcUm0a
28IiFce02i8tqxXimKCQ81tIgr55WMbZOe4IXZbsxZ/s/7+aTfyLfutOJUITnjys
xo2OnnVXXGQgodecQlwwsKoDj0LOCArqSzHJzl+8NVDw8rqieiEMFz24yVLO7L+g
HP5o7zBlwlVYU5/T21OY3+XVXw+YclE6q4ZX+kg4VkkweQ+rhqI8SzBFs2zQIHhD
sZ3id29qp8Dqb8o20vxhO6bc93jOCSd9aavwDWgKs4cuSP0IUyED+iXQWbNbN7+R
pqieszduwg5yGd5mZQ4QwglNiAthakxgf8eDuwmNxzVr/30qLQJWr0Kh6oSIJUR6
wTMLtErzpJ7ElWBIUggT95VUgoFf3KNvjyPVTEUphgD19tolYToegOfXBZPVI3nc
+tcq6AZIgOPZTXpF6qmBeIn7t8jLNyZ0LXp0D32uZbFqzhOLAvLH47gpgGUvF8/6
KD2vWly3R5VxPWbiZae0EgAxOj2MiuLJnq27LUJg/rwkd2tUSialOICA+Q7N8i0d
doX+o6Fdv1yrKl06RRExaudepklN0+yHVa+bbfh/TBYVfE2kOz8wjT5PbcjK4npU
Y/3VbpJ91U4fZ/4YCrqx8+lgQbNfZvC6ZlmCG9sLt3M5NV3YKxbryXxeVsbIql7K
d0VeZ1p96rzE/Xno5IWOS9Z/rEXtgrPn3W8xbmdlIdHounUbnvnuo81EWWyA3rPp
g0jlWgJZGoPgWtTFcSXQ3XdqvjABZfL2NQJ5Bd5WXpITBdnCGzehKRE8aUT+HTOT
OWymbe/mHzQl6Nkmc2ifkDgglSdfCY3PcIyeCbWBD9iHFVqrAhXZiFtuvhC8KiKS
vn0Xh1Fvj5aJsWxMHtN8ZkNv9uLKSziS4HJelCBrJgG9FEaKNxLSIQcqkEKz5Gcj
ta8Cao7rQvHL0mN53c2Fpu6lZzXlmhtNhKfLIOGqik9jCxAn2t48DtGf9r1U1KEk
Ua34z46ASuNNDVs2I7FKuv6ymUNvGt7toJhZ2SZsN6nWX+g1wjCxbpnVC9DxNqK5
et3tqJ6pV3uK/NqZCxdwtkgoFDnh2NlX2su1vpFnZs9SZCVZHmTF+hoYbXxo76Gt
CRHpwXkQD9OoH7CcZuB/zHndeX2hD5ynSLn7Dg2MmJd6uifUIPOvgmgyDdkEIoq/
vwY7eXNQXVLmBphR0mWSjJGw3dZgw63YKNp6yeTGc/bZsE1FdANzxsahg6+8t3Vi
Z+ljY8ZHwd4KrsHFWUfY0zLGQASvWAwtou6F2RlKqIy305k4Lle3z6MHQTsGHRNN
8NsrTqI+qoSEWBMz7h1K5da86dICnTNwdGjw6yHxmC9pF70gPLSinLMaFVPVa3E9
CJOZ9xOR7qzY8ty6NzUGria4Qiou4FAWblBmz0pmoMKYkGEhzA8hDTSO5EOwJoSt
OAltCSiEjGbWEdZn8gzQvTfxGvXsYfpVCKAqljeDCatkz06egUoWA4X3UOiqTpMM
TEuyWFvmFA9W5sbEE99kFsZqYvqAWc7k1Bkq06o/Us3/CNVYfvhgq5qn5I4IG0xQ
JGpQLizmo1MTVy3A1+vLzEjAw8efByFn1FmIT8tTwxVCo4iOtOt4xx3ksRoqyTF6
QW7nJxwTE3M4JGgsGY8L98j2wtx8xdO15y+ho5qPK5Y2FVuQGx1QszXx+g9oC7SX
dSLeT1RckLPdRWOfEWyK3T2blc9GsVc3d3xHMCvCWP9HF790t2BHcUjzfakt2qeS
qy9x0Et1bxzEOYEnonQLO5kAtxsEKPiBTLoRuiXlC9qHVgmbOm2tGpQFXCTOaPXb
ZOmRr5BT0bRGdng1/g0dL/yCCH4lg8GT2eYhcMtyINfl7aBNlNHoUPPqGGMaSRhL
OyZ0jWd88+kWfu8h+UPaJuj9X9YBGL4sH8dyTQK2baUBac8rB/+IFcqqTotkvG8k
O8y5He97hHNWcDasBBCM6TmT3cNUR6WUT/YRS+OZqfuy9yWD/MfG3li0uQmb5mQA
/oraWIcSk+HsabNBhpawPTJOLmyaj5ejrN4H3p3CHPOluzz1l0bSr9gYHlelekwa
kVii562HoXWNJYdm+C/fSjH0DFm74Rf7cO8hsE13dRP52rthrG9KBzFIXrfz2Hgh
ruYCb0Ev85xW7bHGnSoAnlHUkoxaJ1BYd4aKOJyKQJR6RAPrDYPYyprtaztBYSEd
m1oLJxftsG7OzjA8ap//Uwotu0GINO6CX3sDIN+xZTEASSj1+VgRoYPVaeJqryG+
/Ok65tixBEfmvTxdXFRqF9SMN+DmJdWWtrKJpMRFIWH2w/LvY9+DMs3RLE17M+Zh
8HEXM3kfWeg380Yb9YiRevcIdCAE3M3fX60QZbPaX1WA0cRmU7Oxh1C9WLx5WwID
GsvgHNr9Rx58pJs+sUfMG3lbfh2KGYQSRMwuIW3g6XQpcnJp+4uP4E3pRHO4gTur
SUT2qvGss3IISGjXqDZnjTLzaZrwWlK6918rJ9Q2JArRKxkmkAj4OBaObJDn3HuG
XhJyMuvzX9upUPoKdqZEFhjd+ArJCQsPrGIYlg2pOXNUrGbk6p3qaBkfRcSuk8ev
1MGmCZ1pQ3+bTVVYvJsAvHB3aYtMLzIXzAf0nUCw6l610OiCu/rWt/3xxQ8T+amg
KBeObHYA17kMLiiWZ+TpB0pcwR9udmfF2rJSG4/F4ABuepW17R3PyByMEmvBC64A
MpJnCzCq5C/US6COfQ+HTh94oha0aLKsnADzfRBDW49dY87KhMLZWgmDtF/LAtd7
R6GsQnoQYonEFuYHWHZjbA8rknQO5IFPU3TQtieFUt4+2hehK/NTVIW4FyVvO9f7
v0l33NT0Hc37M01p1GW54BFNI6FlnzGfB6jR2ugolGhj5KAhyuXly8tY5lD3w35O
JtycQgxDCYJa57eqC5vWSYnQewEQ7vBoGNV7oKCrwwkkw18JURrlr0m6rFEdg3Rq
/iEjj1rhHv98w1jIwIcQdEqiHhn1lMDCA1jbRL1oavkW6uWyEbLESxG04pkEcRx8
8WTy3/noBHocsxd0nn0Mmw+HSRWAbGn913EtKWhTvseJO7WtlRtfqKpnxAhX3d6d
jQozyLSjiQWCnXvkm+OfjjwzMyNVk96SCVRW1IZRGKQP8KpIoP6fMVP5e30NqHpE
EEob2T6D0ROEf/t02lAQQ9l77psyI6xeW7UFmPHvLJbXd2rdpZaj5mwjkDA83mnw
k+xNPjydfEwQnuUx7Rs3DCfA9hbcdMPqIWmVrJbKFre0nlyaoB7pdOwg56gvEpSF
Bsvoyy1yjgULXgzlRp/ehkJPlZwYH6cHBRzrfl5xVH/ZDyjruUimZRHdJnIscAWb
m2bcN5fKDHW0zK4k4r2r/jFPZ63nqWR+EN73WqJdMCQas5SR/F/5tJMtl1goxCnB
HiE6FsLEe2TzA3XNj2BnVexulyXoFNY1/kZBeaGBQJqTGz6dXL+QkMbDgI9KDB6W
g/Uy8tuDVEapSSD2CysVnH1DDfAtEAal3ExM3kOilbHpKiJRTNFxRgzVoX/js44v
WEWB8YRbqy3bqICMSvG6elXy24I6c0pLVCLrBjUwUSrZfreg3dz9ZHFzF6bkC+zb
vU1gL9XtZGEh/YOeDDPoVt8l7H0Nq/cRyJPeRJ3FutQBKW8USEX2qPt9FK4u1rWK
Bz/BhzDj6p8VjpIw+HOi0lLgyiXrISIsq2WAh2Fe3wnBr3WiwD4hE1Ph97todO/z
uURjQLl5mBh9cvEbsxNV2DHkqD6XnaEfMNNi0CCrpuIdBcqg4VexIF+JQ3o6fBwJ
OT6d+NcvJSbwq5zCfO57OiNuKTXYEkz6E3au8plg3NPy1+i9G8zsNmt9RMhPpNUf
gpxUOof+KWUQ8Ts7zuTj0NmovcYBgAZhrxLiWyoZ2bVl8ywIrFGxXLV+4EhREmhN
+uU9vAGg+zo9q2trEL59oCc3NYG87UBW7Nmm1mfgQ1iWy4qJul08lzxpZCx7L+sp
qyVe31QRq0Mu/+UuSI7c86hOuumahA1ALyZIXJ80qbCyN7fATzfekh4/E8SKKhIg
f/RPJTZzoJAgW8PSmM1Xw3duaXTBFyW4HsUn/aGm971BZhKfmGP35ITDxiR+TQXw
oKYZTEw8j1gVCgATpdslWzJ+LzYMU5pdgqCkSd/E62J0bJOjQTkHRkTFz0q97eCH
cLHOyTuPsgJiXnN9LeNdZbooLpMzZKT0rkJ3bZRdcrcJtds9UAcLrTXwcWTPKiU+
pJsZM5FV07LecB2vfD9+hE2AXvTWp/u01c1Gdcdd+BJeXWf3aEPn7abhYC7BHPrR
D2efpH1lYqaqlhS93aIJDTeFeuKtQ38VTKK2U6Bv0NaoxLBRQcb63HjQSyt0O1Hx
KYdrIkCPzKelc8ncIdLyT6ZzsiCYRf0aU6QLvsKCpjHKNz/U/kQUx/FUbXNfB+XO
kPhfiEcluhei+w07oZfPoXKkxzSy/uV6snYrcBo1TQ18AlZ+6J4ysE7Y6wblNftz
1/S29nIlAFp0Lkx6xelJc6CR5TBnRu6Vy8i9lBTVu2d4sQjP5Z9R5QmJ+PChbDe0
TRvGPmOaiUS0TaW31D7g0Q2c32+4UNH/KMq/L8RMLRlx6iko2s+C6vc24t3Phe88
8ZlMCPvI5MkLGkDKkCspWoQETuOh6xTT+KJSWK61G90BQlHPkcsmVgTPppWxz3GI
DPZQUwcdl4pP1+aB343qKOjGoQBkrMWGEb7hn0Er3JqwvnIXPKTOC7twLI+SaWoR
KefrdS8r+A+AtlzTwjH7JAu6BvOQYR5m1a2ODpxoPGod1mgBzW7PoinQzUBAKr7G
xsxP7PGU/kNKaW6UAOetT5iKAJA9XqgE3DaCS6h0Uq2fRahUx0fW5Do/NOKmOOjq
FRy3eX9e+LjhvdEt8XmLc4SxQ/Ygr6ht9sDay4ahYKulAYRE4k5Jnoz/E0vMvJ3/
ftLj/IMuqC+BTWzKGaoj4jIU344flvPYSakrVjucHI29uWMMyyf4gcXs58g7KhGA
dqrPct9VFYZnDPXtgRHqjba8iKDiJ9YX1nN78PpxFBJSOwy/k2djieq15QJ1FrM5
7aumXtqoqDX4xZAUslUdbd7+UFD2Su3ghKAMcRC98RF2vUUAn1kucgrNNl29A8jy
otI0xzhYNeXdhw0aR6Xdti4CS2xGjNzrKDrqCMQrfOHvdoyINq7WcEJqis7A57MN
xsFgbnzWQK/50hsB0ZfP4h1npV8T44mimH7ohdQ015VzLik+LUAG33r9K3g7zbZz
iMSR5G2wRUT9uAWmxaKWxFNlWlDcum8HMf+XAj/7jAz1DP4PNEswXqSy8zIyIlCT
ZYgw+Nwb7JqucStRlu0ospMYv/pbIpaiFCIPC0SwvxJirhJ0Zm31LRE+gm9eqa70
j+IzAEU83hiXXrKz5n3T+5157EXyMJt+Q0v10UInkkQ3m51CdZ0OeHbCLXE6iHut
HGaAHqkTT3U0ZtSBYNqHuV36aRFyNV6oA3pkO708T2KA/ZXcwj7nwnIfJs65JS3C
hhdanYxDE5U/roAMz6YPZPJc0yEb4DBSYiEc4IqZx5glRqFZpCAzxRTK6fp7nq+X
FopCyMBYsV/u0S+J/Yi1UufVH361LiPwVCWIWirY1rUjyIZ/56WIaPwbrbOXKlwG
me9NV2mqqRBwYGfsDIY1apSdXGn576NNrVSJqtCoGwjFd9yu1ZlJKCq2Hu1zDPac
OjlC4d5qAwTnznoz0hRu++V7Zb/bg4Cs+w9eCBMJrVVFZyond+u1XcGtTYYLmXCF
bjGmS3L/oHv1rHk9UZTT4yTDs8iN0ABOcPuoVUETxv07vTYuUMDuMOPBdj8aE+m4
bl1PiDEX94pajCj4pN5n2bpybs4OyLC78gGrQBAy/EIcpPpDfP15/mFNKrS4cbxD
+UtyK0Hrfc5fWNhK7NlotTeBfmsDhxyNx4612eQe6CfwzdL0dQXtLau2H+UHhjUn
GTy/wqPHqp81vO1V6gAJQbf6PihEV1JY1oY3eLJUSenCUBX614a20KAwY866n6n/
HX3YaOAWOb871GnuUSFocx/8HAPyl1n+Ahkc/KSRFbX714GMmEexlLrir4RpCAmJ
tJrwlH/NYo9XW45IyC5O7+yil71owbl3UHf5s+qiegu81zCmOlzywjs7adLQlTYC
8PJhLBn7lO5SGbq+1l78uSpavA8cPkjfedcbZUokqe6n69VCt9cS3QT2hSnO5G8n
H0y76Hbe7xIwWQZLM5L9p+kZ8NWANRoHFZ1StrGKJIC5/hl6o0ahOBsP8rHYQrUW
M/TbM/dl0loCa8GnXhqkYT8rzsWu+zoreGsxlDa6VAeeZ4ewFYJL6JDnl7XAFnC3
vpAUZwt60b1MZI8+wWjpcfoz04AQ7EmAsmbdx85THKINreGlqeOGQuDL2st1MarK
cc3t/KhovGiWw+U+L559blfFN4HSuP46Q1OcOoTe1XAF31yHipqq/M1HD8L6GqhB
3By6vWJovcGV27iiWfub+PzYe/ueQ28cwCwuXgtViuX1H/G53Wxn1JNg/rccmcFd
hpv7xxhU337uUk8W3wlt/hcQEG25HfrHFGTVgYaqyLWtjdwGdPlU/7xrCZO3Dg/q
3PeySYgS2zfGLnJEyFXJmV6q2YKeVbHoFBvVVzyXYQFN3ETi3foaE95zgdcoBkVl
q4RLV1NtHaO5VueoZ/dwAECdPfnfdqFE0RCUReT8c8CNcFp9F79vaW/+SYOJCVKd
+JDTKJ76q9m3OaOU7h6wSkWlSO3GkAx2dNk2ObLTyAy+AKGr37jAFRnLUzp/a1Ds
pXI9qPnXjvBvmvpoa5SauQ0jcs5K7ZbveidQdYJnTjXvFgu+qMMh/t94g17MDmdZ
iKv93CGVhOqjjPP2HyIRObiw/txu2TSybqHLQf1k8dy/M1yGk+1fnhRR1vqoXHQt
hhZK/u8dcw9g0PGpoxfax/IQ4Er5GVIZiRzpfVgLXmwJ0ZE1VZyF3zIbjCgMlg41
3Q/CnacwFV3FoVvNnYMVmsLdIk+bsJJ8/iD9P+akAVeAmRSWd8LDYQwomDRdC/u2
0OwBYuL8tNmJdpQpZP3jPyX9TmluFTFfCuhGxNJyfzq3mbLzDXTJekr3AskNA8Bm
luz866VWRM321gvXBWFkkpp13PvNUZzDsqwCKu18Oh0Xi5oeunQpTxicoxAepM7V
HTVgTVrWc+cGxZ8mn6ZIe402CqXF/w+PkIH7dpi19PvzYktaLwIN7x3tpAm9yU6l
ciDhb3xfcSWL10fhElaG2iVBgEao+vItAFlhh97ywlDhr/vjd0y81GUNeB2d3Iu6
8FV71KNA5Qv6xUy8OUl+9+M+Qib7CMzmNlyu9txpRE9602iAhkorYEASvW/Qrbta
MK/NNBSA2l5hTnmxOBeY2qJzG8RG6r2Zkt0Wma5Q7ACy1u+jpSB2DL3rPA/PAN90
n5wEXPusz6nE91AB1/oV6FCYF2DV0U0Z9ruQ6hAXyfmDTjyDNY0UbsoB5C8FWhJy
HbWVcVnTpmBqgPH7Zi4lqOL/6fIcrBwuoho0HU2sY/P4f9t7UbSPxnmadGQIUdRG
yTxGtlIWbCuo88fC81gSlwVFDKjOJfpWBxfvRXvHkNJFdkWiFYqbLyBv949o0uxd
fHsog6jePA+S6Woxx+JOV7hAihe+h3dhkfRlTG+hTtqNgisNtmGlXqEfpc2w/XX+
K8vBC9o5SbDZSmTsmoHcx8n/lwQ/2MGmKCMcskguIVZ8WnzSNpTukvjPWDmqEKdF
qG8lczEPhj3cXVp+8MASxXp4i9MHm0dE+TDMVGApgs2nkfQZI0uTmTlaTIp/qN1L
6tPl/4HIJu90stb+gxj/zDfLqOo8h8ALhO5cyMnxMXEISBoYK+ZtQvDOBOvN1xEL
tokfcxd04Dni0iK3tcsz8BSBnT53C6tPX2TS1+tw0ytSIDxt0v7++ANLko/97iVt
QUH6dAxqClTiYTHMNYrnAPXPDGAzQ4VYNK6Yq/af2j7AQHHLCHve5/RR6cGS0/d4
tv+Slx0G7fuTV/4SW4Eb0TyjWMOjVLPHjYTeSiDfca3jhJxdDeYPbEf6jQT08SAW
iNlMV6s8ef9LzHBTlMY/oWJD3Vp3iNHH/Z2coPCKjUhqK+rvB9pvRZ82SPSK4+vB
xKw5r7lxt83FbzPXH/MT7TC4w/BJE22EN8r2X17MnbjbO5e1vgzP6rEa0RwNIJH/
sfliyo0sHfopgRceesj9XctDvmObQGBWLUl1R1Aw+EUmIOGnc4bEZr0p+0qfldRx
89VX6VOK+4IlwHZ5qcxL4ruRqTCogOEJEhrQXyIdZ5jHTi/2pj9LhcAV0nuBM5Zt
8Ks8xsnj1CLsvydWuvLblflnA9v32WeZyCbggIDCAjy6C6iIe8ySf/rnknfr3EfA
tyBG0oxyXO3AT31isw3Jfs9pE0b6Fg58ZgPCsmOzDMzuG1+bvPFMfb+/VXmNYtxb
c9mf54yA71BPbBxeCVZw7w7WyPg6JCvJ0JBfittbpRxQd0vZnw4QHjl6+sz4CyIN
xI8z8z3zbL0NpOWRUOu4XHALM4e63lYgcYpLmzdgKlstrwpGQD7/U6pAc96fV47p
zRZoYrm6qz+JdEVsUawKeXacfEbfbY6CCue4EuFzYHvjyLMaI8/19nYFrmkF4kMz
IIDQO+WK7aVJCbBzFbF18BUJ37rvFckqNxDV3j1qmGh+idrLj5I4VjpcmUjCBndm
LmKBEQX+n9YWGEpYXdsU7InwmUKk6w91froegkoxohpulQZX2tVIZJwxzvFlgHqv
PtSiGYTe4BX9aYoREt5nRbC+5LxGennhfDDBJDBTqemSp0mCPesPwtoO27/Y/oza
tqN0X9i1SJMb/nl/5nzsLeNwYu4S7e3Ncb/cojv/i58wlrn/G1lwn5n1MNikoikb
46uEU15FK3OnhPb7/qHgrR5GIOkxQzDYrG13UtAsYEexdPTv2DxxFNOt5Cxn2P6S
esMyvDRyqdKcVlEI6hOtYClgVdog/72A0ODi6lBY3IgCnYBicdpOK7D45LuSUjQp
t1CcbBaQQ1uEZDrAm173+c/2K9kZ7B1740tEXwFjEJnUGe73goGBUBZHnLBhG6yY
ZtgZN2Q82laSoeQOhiol625htir1ADnmv7u338hTA4zsvk0rsBJMa6wXbWT4bdjn
p63pya6BrmUfsqSsq1jJ38/o1+M1Lfk158NENjIjVpo1jSKnkXDmQ0qIbYTbe5cH
krI9CNs1GErUshQyIaCf17nnV1nP6fIF/5ah9i/gi2ht6QQzJvdKezZHChCK0qHN
+OZeDyQQX0wQsKp4mUdY3VtGhD2uQrfCGl8/qJz71haXnpqbPj7PP4jYFIIKVBFu
CBUFPL5vTU9U/dWAY5mD6PcJ7qaP5iHOdTYEJi3sIDzG6Gh4Zk3eFYiDAYOw+3po
WEqH9U1SdJPP19ZZknSAvBf+6R2iLFDb3aUlMau8AXk8jFKx+TSu+FzwNKj2sKaa
JIHeGqfAHmg+zqi3sx0EZ/JM3eQhgJ8zw5h1tzFeeadYJQzB+n1BFYFxmwNC9AEG
xyA47xW/jwFAeL0bswxmg+LvNphNgeTDC/C6Io8ngK58jns/lidjBIvxWnRy8xXW
HiKAcCQzNSiRTM+F18XmijuvhnSGcnShmRqQi9zTaNGR6FluiKZBS6etxW6QWWyK
Rfdd7PICfuJRuTqwW5grDAp84UlHhk0ff1SjISW6MpADDmMN8yt/eopOstep76vk
4VS0LnpkLQBvVMMFVr443y2kBJi6CFgIXsk9B+ml1hwHR+o3e5FRpJinsjvI8M5+
XzXiNh4OcR2/51dFv2uqfeTxokqGPEbMTaW3HNkyCweCxwH0yNXMbJg4GXMgZgoB
PYkFNzb0M+ghSMMHzragLR7I6tLAK49MBq3P95RqbH1eGPx9e3nPiaDErciUHAyV
Bf5pt/4dTO3xedG5TIN6vSv5cIotVtwLFfhCxFtwfSf/IUCW3oSlzn+RbXhVwp5M
nJ4TlfsOM/G8erSzTG4xY+8PiEsJ/Gqh/6R3sWR0Gr6/U9joVcnaGI9J75/cOcXh
mqsSXXP5CsDGKIpGIRE/tUxda907kdtyQQP2Q7Uwq3/mdLM2zp4Wy0X1tJ9+KSy8
zAMpSVzsof92TxfhTSjVipR8pkCtf9Gnj4Vhd6TElRzYIgRtXyDTgsrfuNuhb1lt
ZJOTlvwda9dpV0qky3u4I5mWFJMqeZVfDPRCORg5QDiRKPLQLVtN+/h4HfU8sHgz
oON2uN1UCrrJXcRTcqRbnXID9x6VGHFycvKPkaeaNlX3hbhuRxlgoYn7FiwGkXIl
1G3rSbbOXLGHEk7R+e7bcP2CWJL0uPvAuj+AIQATnQxR0QIP+CQnm0w4SOhvwbDe
qiscJW10g0UnJVn1Y2xDC0r5krTnJX0peYN8Zu5WBPdCQiYZnCGnOkVlQXyqdyI8
ejxkNez0rsZbdOSBm4C8y1rXN5rCF4oqwmK4RMtOv2Duzm0Mg2u4ULLd7VYp2V/C
otMFEf5bVa+g+GnONDSagJS7brP3hAGVVYOYFJEQTu4so5HdVc0eLGoKk/Q8U4D8
DaVP416EkRH5OSegH1GKmKdoksyj7AvM5/08k+nEBZd0MMorxkJXH/hqk7UzFj6l
669AUe3a6PQhzZScFT3zegLky15EJc/Gwyvf1Iuse1SrcRZaAtEpFo9s1/yMEotu
8Ug1P7jD0GvLl06KIOQfrvKIo2UlyghbzwpmzNJGikL+hGFdQ7bGSzyJmV//Fv31
MNsfwjavx7pt9ZTCM9B1QXY4VOjq3KX1xwvqkVdu+g2NXVe/M0CYy2VCtuRN6dd3
5isWjXEv07W2733PHVB+ccLUL8Xy7tpnvvGY0vbDI/b2dFnx7oUGdTMIzjU3z1cr
OgDmjJlaeroVDVx3lnWi/DUk/MOuz/aU+aTjZMja9rzbe2h/NJVyfrDBBJwMhGqb
4IkAq7whfUZ5tFPHFYciyFT65wL6vobRu+HBEUrApm3TBI/2Kp7nnOzLUG7olK02
QdtX5GTcEdF4PJ+DvtoCFSWMOTh+YalK5GE8u8VWnCTlG7NfXgIAuiiuI4dGPzZ3
DseEx7ar8hU4iv6RzSQJfGWekM2dhtUXpPCObjhZcOD7g+GDCCCp4JfUTZ7AR5JR
vIC0ebzIhMaygqoRMiD9P/3o/T6gdQPZ+tXAIufvtub3WH6wLloKebcd7N8ufyZf
XdOGdAolieToYx0hqSPMpuleqPBNC/KYKuI+RTr1Qq5vDaZQbjw9oPwxMD65Bdpy
scrAuHLtL181fYyekg7Yx6u+uxW6D/zTUvmuLBNcZybRVpA5BD6HjxHPEdxa1kRo
Cb8qSApbm/MXUumfBDSY4OisHwIY1XAxd0P69gHz2+ZR22T+x1H3CE/6VrVHGHCd
4ojao01Up/iZ+f7qWl2JyFfXIBN2eQDb2H8YoHkLF2kt26TiDYGNbYkGnQDjiYa/
N0NkdIPoJtaqmFVDQRoiL0nBZCH8rNMT1c6b9vlLNJEsvcqbv79dG5IgFAlSJ3h1
pkdE43vonqMYQKDC5Gf8oytpvmehz2d04mVw7JtX2LYJ9Rlujfdp1PCPFMVZG/FU
FfGx0dXJsLeQ0Te5UtI9e7QD4w5FIlSMyP1iYzgeaHIVR/9qY4j2rWZ5Z6Lm0G0A
jCtFScEW/XByv8Nbo10nm8zFF6dGCwaD6Y2qR2vC/+s1fBUDueSruCVCeFt05MXg
3DzZnLszHXJ6stFDCUFtanbbqZFz62409DsZzAcxqVBrfxquRNHh5EOcmWOJz9NO
nnwqoh9WZCz7Yhxkwq5WKP7SwmmbDHS9/J5dvrHPSQGbTGC3UlYXX4Ip3PzN3WdB
nqANFSG8vDNLCCS0SoHROWTwO7rLAmc72PB6rk4l7PRMIUL40Kq8PDZGTSiMXwxI
CPOGnSsmPWp7WxizrWFG9wyGdKKuAzQ6v9DK26PIla8yt79nmTQrnru8dmg3wYe5
QLOO8magJMNbSkD/IeJs0x0noZOqhYdv9AI1SXAOlVkxXTMHd+e6jz6LLXTQW6bT
onTipfDAWIukTGPu2qq15NLcbWxovPEZh7hWeWnkPx088rHpvJ56HTfW0x/xYBjO
QXJE0pWZKWMVBJYc9r/MSh0zu1GOyHJu8VVEyWhU1Ufx79zkU88zrjUJacktOHUQ
dYAXZjnWV2qDLoJZTWAClfJqJzv9PGbVLKFOoegafmvhSeqSPdKD0QzJH/+TtkTl
c+q5saDb71S19ZKPv5nzEyukEPg/dxcZcpcaR6YBYKFEGY4+1k6ke8U2hal+jmfv
0uNc09N0947RtowvB46g9v58b636+Gehu9WInf4eADnH/ksuWeejXq+Nug6DSTez
4Glu4eeoIi24LLdbHg7MjcCXFw2Gz7+y4rRv9W62DPg7AR1P7ADVg5oBT9OD5bxh
b7jUDkCALJqau8h3SfGjD2ewJbCwEl1Q47nd8ero/BIvkfPdskRSs2tNF+k4Qbww
3IZiFtWO7kx5266hjZ4dE01U0gaTPbgeswpWn5tqLesBhAH6GfPpVS4kpY/34tTr
tVf8xQeyY1YQ1RhpN7biy2WMFQTBdlk4HU5u4J8fItdY1yUQ89cv1M4MZEP1wUV+
EPaL3ttCg05UymyLVRz7fNoo14uYmHdHFpEpML8y1tsrqu1Jho1/98P7mZ8Ui3zQ
q+Fc3v+GXWoMolUGJuhjc+yOzKDUtkUHGkFIJViOlafvheTgyWqGgVwi1h94OQfP
Zr3YqS9U4F+jcFfAkK7nJnc0lM4hOmnQVSeQ67gwge7492pzsZVDv9YNoc1Zk56u
+KLCDvHOK7md8qSSkrA0piE+WguaEYRBQgdquBt8OhQIUsvAux7fnC5gmd6K55H2
uk2/7ylfSiY7RJqyqdJfv/xIjHT3fchUn6RPW8uz90jvcTH1nRnL8HBI44M25/T6
HkWMYDQ2kKiU4cky3Ql2dazlvSci4HgAa9fdPrpISYYZEOxnSOGVmmEoMsYpnt5f
PtURc1oQ+H0U+CM0zIebxh8hK65Q7hQCOfbz5rclN7vi0vfqREoivqdKlRTX8EOs
tTOFeJl925XADSKtJSsQnFBRkccFs56jKNSfCwAYiEmw7uVICmsrF52Y4xteEOBZ
BCjc4cL0HhZBIFel8OaWRLGRIhHb3VChtsFVw0hNl1Ubc/1lLYzoCdVaWtS98mDz
DVZr0O70KcaPr4HuMHbG2kO3vStu9dbPm+tjYYwoXN643vWeEhjzorDXlDmIPdY0
xQVjoDV8XbyZ+r6cIXBoetdJWkQc3AsAdDul5asYhme5qhagSywxQWxgidKBH/8d
9fd3nMkUAvRW2HLjTUdoaFKpy8v8Xsi1VWydDxwgvlxaR3Px4gRaPnjbesrueqs2
wFJVOIa5/hOElwZp6WTUU8DoRnEHBmEez2VaLfXmDS3DtzFnGe419qLlAY03X1+z
XqdygMx7oKm/u96rf1MYA4P6Us6wbkLIbZi7DxsplEr0bmPTxoCXCx4Eo+cQyNKa
nBwc7NOfyjHBcG9ExSS98tOFyq+AqJ+3TuY/AcqxKzs5ddQSwG05aGoJidO7M8mJ
yaKI+rNFVGaaE0dGjBJjv6QnzBFepjCFw3Zl6pIB4HIEbknOBhqPxQAIPOPQ+nW/
UUWN1NxiPXkpgeSKD+i5K4VC7IfHmIYyJJ/Pyr73LDUPcFQUUaEwY8ubYn9c67yB
WUeEn6spZcCnh1iI36UylqrRkgzxaCd4oxS08h4OjNlplrXWEBWy6jmuY+IiA4U7
MSTnfQXgeAKgjr9l8R9si4Z1LKHMons+rO3+48JPJQJdzcZrOpW8rOmzXr/t00f+
MWkXy4dw9rWRL18vEz56feJnGeaJx8oPjpCSYiea7Di2k0U9gx+fP8IgdmQuD2PK
zmN1VtFCCNLp55TlsL1dmyrz+97j1NLc5qUhY2EBjRA2vMsoD6Ig+jGA1oSft83O
hPfFzbOo18qc8mjlSJyh4b3joYLZLPN42+DnvbcURt18gMyToS1is9Wq2+dWR/Gg
VL8F8+3gFC86GSkdMz0MK8Nw8qcNqM01kIZA3hLyosA7k6SoUwTsW1Vhf7C8yJt1
kX/rmH5FuQBQnEU39bRqE/Lo38aKNC9aGMWBs3XPdgYr/fJnFCIgmbCdKYoOKcLF
sRp7w5OjclXKt8EfQbvFKYn19mqnwu923O3Cp0PzN1RxuclxaMiKtIJ6NR+MRush
BFzFcokkBNDzYtZG9rZA2I1wpSFSZQQJeGl384RcYOOb3EplRG4I9M6+gveCj34/
GWpgzz2en4AJn9w0TeGIvPp/TYFotBzxn+1/cjPM+oPSG03aqfoiiL7ckI0yJL3Q
MjkPW0Zr1t6Yd5yxvE+6ZdTjN7X77sv886wzUnMvpV+7dB7gZzc0W9fVb4lzS6hD
GT9RLW2U3N5IZMhCM7Kc9sEZJEyZ8m+1Nm9pMR/5XIll5SzewBfv7YMiIPA4nIWM
nmAIjZVYS1OBP9nCVe8v9JksBpILJWyZdADk0a5Hz01Tb0D/QWmeV7DyFELIUal/
rZbrqGBTBZ25TeAPkCU9ZIDBx9GiiEdydJpx0qMamV6Aj46ULL9JUU/Nzpd7K51s
Z2ybhDOT2HI5dZdY80HtiPuDoDDGh38ye+Vorh7L53+dydj14SyzfkuzePG1UgR1
QEheO+9Tps+62IboaSjAgtsliFJKt98c8wELu04EPVxdtmTu3X+rHdw+nyXc49QY
neW4Ap4nl9pa7/hu38kRbR/LQj0vdv+2KPnh/Hx+Hvojd+0SX7eWZAU8N2UP0dhP
MKbxeCygbAnH0JpjNBsyPRMtWGM9l2bmc00PEvblvHL69RdXsfFmTd76wkxSKMdn
GK2YEu+kTLxcAvnBqbB4kAldmVzbi08V4L/286IWZWQ78K4dyIoplRb7cUX+Cnho
Y1ieq/tWwOIWwWWhPrB136YmBa74wJvQ0+6K/9E6MfVpv8txgiImPozg1ZYzu1Kv
fcvkMQI6uh6yUr50f/7RrZOswfyUVyP/gm7epfYyWKIO5ow7gazw2XC38xI251BO
GAX37EAZijnPGOSxKopVe3ugaASe+XdQh8Js9O6u7j0M/jaPM9/EEQ3RrsjDUeTx
NyeBkeaIfD+6ByCMpIhGhcnUGYyFTu6RfG2vAdPORzhS0ASSPdMhScFVQn5jKIIU
Btq2EoHLJJJMZnRFJTv4Lr/hcDc7pliMxeeurF3gvuPNb/4GRl3hTL3V6bk+NF/A
8j0skL8/55MUHVyD9fcKZewVr/Tf85FFAyD7gvwsfOCmqX+mx0VC/vpXPr4jJqsJ
EtkIMMUjf9jwVNxZrVb4MyWNk4ISU9pv3FuHyeJsdfOXS8xTDPiWyGtmP8+QhUhw
+76Zqeiu6RiLzNYDaKe7BhJdjF4Sw/BTBHoHEyK7Imw0rG/broYmbWlx02quq8H4
M25CjdpVeKCKLjHzEhOUjibBUSvg/H1hAJuCe07SQxrHd/aRxeKra774iej8Qm3Z
Rnb4OOu7qTF49f0Pyl1D3T3wNYHGjMtA+WUnlNBvVMJEYmTeVfuiHnKN3HHVu4ov
Agts/KCkv2OedNfVhXjS4FQ3G4pTn7q4825ZVo0X/exOgt/Yr/9Y68KZnyCbniv3
9/oG/xMtdDHJ+xDKlz4WIXcMx1tYfX6CRvi7ATM5SOcUyH0hBvQ2/QwD99EyYi2G
fZpOdu9JMqvF05nCzbwL8Vm1E10MmjaFrwMAcAVnrTVnu+dOoiBbmLxZHU/2ACcv
EDSpPuS+4+i42EtyOmw5neo+P9ui85lfvYp7vLz0v+wA+mTCAI3hJ0eFzXJDnyS9
G4aaBcIkKQHS6H+E6ttIMFPqwYYBdLHB6vehrW1QFTqOSjhDxfXzIMKSkQuMrxz5
D6ZI9BkMLbO/xKLkQze+LHf7n6nLkUKbb8z5x8KUC3Iov2Qv/TDCh8dzLQaQLvfC
OZJc9088YPeMIheucaK31W4dghPk9XG/+thGdHIqzl63uEhk9rbXoIG+V5hDTf0t
+pGp3Y4W5ROxHsjgI0drmoXcdDVQKWMfiLhhsMMUinAx//HAEknNsjy9Aac7io1E
QQsAS/GP+irTsfVwIMVHNYghQEtuk8raq+/WmtUhUxmE2TG8L0os0kTBIVe58CXv
aY54Hc13gQQmmtrHZEQQc6H+Aoo4WDSBqY0ie5aTElbyjoMD9g12wFok8Gbapxv3
teIQmqgCDDmo0axoWQpZt+BjnoO76f91DBfK4KCDG+1rJMnhww3ET8QYxITJkb0t
mrLwXRwaa4TMUhhHUSak6JPmZUCG5m8aEUj6pe3II8nsralizQ83bdKom07e3Ejx
GD94DIw0ny7E36o+qFQ7NVJWi7f7MlLXhdREi9BLVf3hTNOmHBsdu2P+duf3nL2b
G8rTUztSUcGPtS/r+0ssPnkw28gZUH6PSH+bPDxOb6jW/wZtFhz6MPXbJJkPre97
5Eia9whrN76IHKm0b7pBvRaVyJFq31vZd0EvLX8ogTQ04F2efb53/7hVxamou/Mp
hksBn9dcKGm92jWy2fNTkrgLaeD/RYL/O0T8gWHJ6cG14ylUm2/OiN8PPTAdu11I
JzUKiKhyncpH+dqBbo0rSVZD6GCnyKH6hSLcXJ4G0AvF2ZurmM9K5UEyuPUQHKp4
b4tlSjGHxhbqezDSpSdRwcKO2S+FjrGQC4+1M5xgDXGZx/qTQsLN+V7B9a72EU5i
722uRZKUKafnWJfo0BcTXYJuS8C4xvMxZJ7B1bbgG4O5MNkzwbdLqU+2GtBrug8m
JR3do7TZ4k6eFKrsg0Cem6sv0/xB6iqkZK3xvlSlAOTFakIELAKDtHzzeOlNKvJY
n7cA4FpGaQJTrul+tDXWhj8CKZ+Z1xRTccvdmOORqRn1uBqlG8ESC0bI5m1Dzs1y
e00z46CUKprVPmnGKyR1aM1i48LNGAfROrl6pcyTs7aEj1ytMVP7W11AwxceYcfL
9qDYg0yN0v1cLxUPndpsB5gNxjt/RagnrsAlbUpdypFeJJv2osOgnIrO9IQyXmA6
7U0VcPk55/zbrT/I0dhmW/1dJeIpBJXDJTYTP4mFTLaSyWAaZZ9AY8mWufVxtdnr
UqMITO4O2qrrL+6Zfifp4LKphTQpSOgXcGIt+jYlp0DxZrmZc3aKvYIiqICkWcdR
dXrrZPxkifjVUBLH/wbrDHIqYd4HjLPmrju/adSBmGVQLJTj3THg/mdeMGyweza2
fO6/CaJlsv+C9DenjUl7w7hAPCyfIFLw1vppqJfqnpmz3DfA9pHdtYaZ/qFeaotG
ysRyOCe024ZYE87rivpX7Kvjr1afNJTx4kiU0kY8smBwuUE5vVPOoR9fNnFJCXJt
CbyGJkgdkWcOEnAo9IsrVtBqEZegSWE+lv38JTSma9+kB+D/LzDefyNx5y8Zo4+O
ZCk8Tirl3RsWymKLwTNmPN8NuqBqpkKv7oF5FJAirYasgooJIHI60qdIte9S00Fm
86ds93jyQo1zJ8D1PhGB/T9r0jOvrsvh8OPPFKaKrHKphvkh6qV86N3FLEnZJ2D5
komdIq2NXIf0B1S/VPNgy3jdVSTROXWKRxBD0LevWwpTPIYdItYp0GFO8BGbfMN4
/ui43PqaabzMHQvlT5PYs8qQtCBel/7at7+gHDBQYaqViVNgFxTdO9lWP2+MePpl
uP4Y+pEpCnbq7hclIYwseI3HoZbTQAp3dQTHhmwW4yckAacR9pxomzHwD8fkO5U0
7ynlH8desUEsZjYtCLyrQ9/CeHXZbUqXkggg6FriCgHOlKdT0sDF9zBJuG2EUtBj
Qt/jf575uaf3gy/KOE9Lu2Hy7KpZuBG2LkcnRG+OS/z0UkYJrvLFDTE7qjrZjtpK
m93of9TdhjrM9/Z9/DDHdGtysjLt6vf5tEP5rKFAJkOhXa0aTctRKj09CeANfaiV
JuUM5TvxgShq3uGY+P0mJhky/uLQvh31KWlKND0sqorpJRxI+bAbJdplRbjr9SdL
yHX+mDy4MDWShma8ztUEJPn/Xt6BJc2Q6vDFcDghyGspmTvojkJJqb54p9jIr5hN
v2PqNf6O1HiWwe67+AX0xSJ89VCP7Lxz7T1vbJoRg2uXxgE6RUTVxdzl+J8TujwC
oa89Hxxvcvst93OWo8mM5Z5PPoCizZDPZkkcOsJzo909uDaIQdKDD1PLmeu1eUC7
9FeYX6TLIyKyXhQsT4Qvi7BN2rMLxcCHhNGgLIhrLzbKKjNqXItNvXjgHqxvRoda
/V3+ohITHrynCoguk4YghqUubK7YPo+u1pEKB+yRmVz+aqAyxGiEpx2fjLSO7EZ1
uW4p8DAvV89RHlprzCUu3m+4/UIleYrQUMZZ5zz9Oo5oavO1bPqlvAO8Y5fwzDuH
38ih0hZpFqIay09zs0V+XsEP99KBfRuwDz2gDjSWBnMffw/aK47lY3C2YYUZRqmk
C38QmbxhgoRYrVMhVncMXyvayWqHVx8pLHiT5Dq/RNq7UEu0XbPfC5lnZyASpgH9
YtncGck7CeD36Il3JwmdjryBGT6Jzs1Hg26etPJDDsF/lUU95Naax8fm3SKD1fP2
oeCUi7GR2ua3XtxVJP+j/CgXGIOmQxrb9CbT86EufZFD/NpjpWau7HsereR+IPZ1
AgklR61KkmjFbN5wfP6e5ElBuMCCWtwGk8G5C0NUQWn6EulrDMs4ayUPMYLaO3tf
tTaNpIhtXThwOtNR1hfF9qN+McHGYibUHP1DKWfmz+CdYE0TPsgTzlV3EuQYGWMV
5n7fj6/egRrNGENHT+2/gqQ+E7usJmQq8GqvO69D76362lh123IUs0n2+Sb+vY1B
JWQBNIuKkyF5fcTkCPq8uNvxeiGXsByea1mAMbCYSaDqDjsxoo9bV7I32yQ1lKUn
4QGjI+4ra6Qehd0P3ih6PznthnBK5FjvONOFb4yUdZFuYaXwfLfFqzNxEN4pntuc
7/UG/0Bre193qHK6CTJIOCCP2xk1pyXhBoRF5+eURU/UgXYT97LyWJnQ282Cled/
Xq2e6ShCTiYFOUodQJ6OwwL3qq+XmXERwku6Xx+gdQdw8GAHSXm96u3FHLD834nu
xCjK8hYkkeffEAWArBQSQIFS74eItIh5adQ6wn2m76z2R6fFHUj9TNms2bQIVmWQ
6XuOdT5skniswM9+Jzs92rug4Z+x0cx9Buyrt6f7DWT+PNpyxmRoydLN5xvisnAl
i6uebtgBgHmmWw2zYiJkt0RtiSGHPBcwxM5Drr2mir4nT8tjjeH8pekBaTD8Jao7
zkwgAH3mSJL5iEeJZPoFdt+DjoLnU+M8a1JkbFvxXvegchfDVIQEKzelNZRHfuI0
cBfYQ0m0Wgicb15hEJdYl2Qqs0s/ijd9L5O+YRLFOdPsnpPcD6UwDA16Jv2o4JAK
y9IeBkEW2rS/18P+YCsgBkK5fjO31v8+Vxqosh1qTV3+PpT+bFLsU0ZdhHhOuDv6
mKPx4dZovPooH7qng0qr6Ya5DaXlD4h/8vbwsy9a1wu0gMtP7M/JSc/evrWqvAfS
/y5UzfhPlS+9gHf/8zUensFT6gcOpY9RHybGQM2IS1eAbKj4rSh655uyT6/HbkxZ
ninIVq6h3CkyHA71UgnnSNoDnAhcS89zy30gzVxz/BJPX49ivNs0E4XaH1GqsF22
2b9q9dqNkodDyooQkR8gl2ss6znoLiMjEXi5foK+cg9ygf+12ZPCUstAR2VL/9Uq
WTlSzcb1YJoPY1Lo+7hFILawG74fPNo7Uy4dXuBS9lUyejc83mMgO1qlb+9qjnef
JQgnWQQSpNqoS0tp1ZeO2LM+nclOg2wyX55aU7dUIUBwFos3197KTfY81N+xpcvH
3NYoYSKjiAc49Hb+XJnJdiiKi3w43A/uTeSuf3VkJbOc+B2IhUhXfjRxc8b5X5jE
792QJ2mL+AZcHueyeJIM2bcqsGiLRSbsGAJZq33Nz1LHLzNOKVXICvxrLNqlRUhT
/7qxWxUVHRhBdh6xQ612Gd0emp0avrrMYA9niHgGe+NxRrrhFtpLmQrVoZftxXrB
eHPi7LYXKgNBNazRSPs1YEfiweZlTmcoTxrtfzGoxku7d/9Dspa/8CvU3R2ifNJI
hgnA8tsyLoCceMto2wMKwEGW8N38T5wwv9TxOX2TuDO0Mdx5iRFADxwXF2ac9AHG
QI6QTLCyVHIxrGJbYyTdqy/Nlzjt54QIpmrAnzaeBjTTLju1XUH6TpGmqnzXiQtP
gaaYj2mgLMfDiiBY0UDUIIAGwApSAauJJ97n9AhrKqFl9kvqhV/tlUxYhTB4LUmj
yomIlkbgjdp3ZUqXuS8jLA+KVDnoYDJOH9arO1nixBmy4JiK6GNq3gCv1gXcWSAT
P6Yhhh2oj959DBb5jPw7uOMGqFwFI0wSFlcB1fnWnh3MVgh+L/+AQa2P5hMjUigK
wQstzwJpHx5CH6qNuDfJC+kO2kTDgEh5PyN3bQILy53RUofkrZAStwt28GnxG8UK
iN4hWvmF0hnx0hyNEiesemWkvuCqZgDFiBsLALmWyA790BVxaCA7SJak137lQgaK
aoO1FBbJ2pVichuKZHXmTuWwIxnDmWizeG/gLsj/lP+TW3zwGQoJSsYIWGCgTVp1
c3rUxbHogj+WGwCVtcKxU3zMwC8179ZUfED55NQCy3Luw3Rz/GN6D4Am0r4nLN70
wC0s+dc5b1zmE8+am+h/RSc7UO2ZhEwkvtfXuZo3ClZ7IACSghQwvORspLfx6fFS
5j1wYCnTAgi06XqAHJspRU+WAIrKUO5y9tW+CnO5/j5YLdV5/ABLGUzvPM2Gy/Zt
MIILoKoTmqdd7QCFS3xvynX9OierMEA6Bj/5vuye0MbxZH27cN0vBbfbGOIKJpPS
j7/AiX7vyR3UmlaHG8PcmXUUr0ANmKzxBbQxlvpM6LTwrZk4spfocuxToIoC4jj+
/gezLOX+kAlgaCa7hOl0VnHW/C8VVsAaZku9Z1VZOokDgIgMVK+TWrJfhw+ki1jo
Xm74wY57SOI83gjr3FcYBWnFk/7/WvBlDx/ZKrv20q3EP0L625Ooe83o/Swn5tij
dVSCpnjSac7OFftEZkNHrsmGiTZIb5hYltTFhME0K5w07eUj06lQhvnirZM4BNq8
rSjw7oe9nPjHsNqP9qZfHTfbUvwZdcOpGVC/CCG5zp8FzLM2fTtQqJO08xaWQ813
UbshKnxv9RtuPeyRsrzH4Mq0i2HXUbdmEDwjDyn6YtsilWAKLFcei94R9eW2PdHs
YJ+OygzBgnjw6vxiw0nCE+Yw1F1hRI40Efrs/ZXoBif48rwV5H3HQcUtm/dypNVT
wq/ctaV2nl9SgJN5ZBbTMDRDCCLtWV6ksahhTiXbfAEyEQ0SbzLjDyQc9assXxDO
VPIfhADh3zZsXbyYUkiLT3yQzq7Qwx2CHvPhSVGUMIniYs/XjsvCQxa1XqE18KS1
WZJ/lRBLcXV6ic/9HEqkgVFDXCZWsDQ5tQCXhJ4dm1m6iKH3V7wkAdDxms9/HLJo
2Bt6f0uJgX5C5Rv7W5UGeqmFybt6HwqFTUfLRcS7Q93J7byXhhTU1AIR19cdWetL
bAyVKAObBrBsyPWOPoPfq2uV4qHVkoidLwpo3+CCYwA4sro0K5JC89GXIzSrWg9y
Q8Xgj469H87H5IEGdwfyg7hALuTeS6nA58Hesuis9H+dJKOBpGeISJrMdO5w348o
sAiPVOerm5mMPZOpltyJ21g9k2zxYH5ny/Y9xyNPBrjNXDxEQTmVXSRBOei4l2sX
gtwtJUNaG4CRD4l60JUeMgwYb3QhqpP3jLyfxJM745Owgt93qM9/orhS5M/VVRiT
Xh2KZcCihEhmE5bOChRdKpxFE0yAOw7sjUaakMyPBz7znxxdzdFjcfyWD3sy+Tc2
9XmdStowHDTwKD+GXd293E7bHuLJx7yGNlUCAsUqMGwlvnJquvlMN2ernOVbS+ye
DPw9EkoIqXEQ9/gInaF8hMEvcJmgvTtgic64KKdGRJpEk9yUPyleT7L4b0cqOp/s
I4WqbRcFAQye0cgFL+0SJVTWTdMX2jjt5IPcEdicIamXF3sbEWQHnIyxl4/6Fotf
dnhf1v4bGvOZ7wQOtrDDso/jy5yeD8IjKzIj28feD34iNof+LUU5nxAcSQOqw1TO
l3lmop//zYoHXPr+6tB78Uq7FhLwHMC4X4S/3O6ygPPq1iqeHHLRp/PUF8N4xjCk
AEaNWTav2R8EO51+fDFRJ7PAWG6hTf7VafWf8xt7jnAzdt5rFY8HgtxQKoriCrnc
gqbkpynsGTctIdDXhHKQWf4/tW0A9hrqT04vIvUOD/x1pZ8HI2VV9zHbNGff8pkK
kR2nJOnp1J8zQCNHf0DDf94opboFpOdXFZ7IlFxZ5DmAW2V8Kv0cRiafVm83zBsF
0TR5qEjT/E3JNfpVvHwsdYuv1BXUv2rzD6b4UvSJCmplPnt7RRNyBUj0uMVokG3M
0iaZYQKLiZL+XeBe27FHeglpnifOo6/cpbrQRT7TaXEQF+ffPdU0yitqi906SGuQ
Kh6YkPN7+G7F0Ok5TxT3aqwVL6tRRZP14HGrx3FloY0jSz+ud5Q5xzkyYpIY+e4a
3RPR0HGM0cri7xrZg95taaRn8wrp4GO/5AdzQY2Q9hmNWIzuYj3Ui19uqMpnO3FL
+hkBQ3sxW8+LHPqjfDy4TRkKJWrXtjHYW38u1PMc6PETvrgUuX8eN+yvrr9ts+0d
LDxWCXoElNFFEb2UU5q8kwl5nKL3kUUsuQZhNWTEgIv+H0/+YP7oDCzFg5vOCJdg
WQjXA+vXqcTrbHxtwfH6GmB6hCJVnq1PNNRQ8Dh6YadxlXL18Guwp4Ek916KGhci
mlJX54DNlS0ndy0JoHnCLYiYtNcPUPgVqb48hSEUUwyoKldskUP30ZoZbIHIyT9V
KMoN7WUSLWIJxGlq9PCAFTtk0qC87L8cfNcc24p7JXrGQZqWkNNzk19sqLGRXgWe
BtJuTe48VsziN69oQQkP343ca/259bEKrLUa4ZJaUIFEiHPdxYydtkKYDVr6orZ4
QwkN/ZcFGYEQfeLHmTT98XQ+SwWtoUjwWZkog0XazO0yWb1PsL/krAMABDt99xSj
lshe7MO5YDVuBv0slqfSHWIOJ/JWvAvbLhgdD1DN8Iq55Wm8rAjr+zYVEqS6Uy3K
M7EwOU3uPcMCSZy+xNU8C0m4MlVPTMPQKKMwD3iOgtgRd7cOs0tmvJUwn1M28MI3
jwZMoZvxCz5wLrdNyv4FfcHSRWiJhomI62emaOvhgR01UeZlUA5P5/4WArX6cFli
DgsKp3oJ6ZFa6FLJkY9rL6e8Wq9q672or6Gid7U1RIsRBgiOhHnKWtvww43U3tFO
BVgKDstaPwn65n1fM3YF7Y8sU7v8Jz4zPdeGeUyDnikIjAq1FpdsAwIHMoDik7qF
0Rd5pYX1aJB3JdvhY1vDo14hyrTC+LnOp3LudX3iggOoFHmkKUm+KuYHgqr/Uifl
Q2PXAZh6UdnsV8HMf1HC/g8vR7fLrQpiAPOuXJFGYtSRd/wqKUzk9OgztfROWQV+
qplmIJNTNaL6xUq8x82PHW9Bmb3DG3NSSlN7VWWJAAzjFWIZurX1r9Ue53F02Fgv
kep7Jz7AnQXvNtskvf5QgGMXs9VJ7Gh8EWXFFnobI5oIRiziujcBOPMXpEZ/TPpb
LXUMMxrjwcaHz9DfQ8m0KE6JaNyyGo0aCh/0j5ubiSFV1eBD6k95S0uMvozhlUc4
JwU0hTTv9OqlJjx8mUqUJnHEI2edS1VL9Q9oQ4Wr5UmXijd15y/4mF1hE6LlwjFx
nsp2T+BMWAVlg5+V5b2mF/uNi9RmFtr9+D9EvfXq1RDzAbzI8eM5sj8JrUHm8cfm
VkDVDHIk2Y2urAB6c4UP+dXcLQI1Kh+Ocgeacf3z4N2m3f7iYt21Pp2tkXVw5olX
3OC8zhK/cABg0aVGGmxncrdIoB1m2pv+xsPRlJFry9+/d8QygFihviG9XMX77TnJ
Y/4pc2zs/uunqhEzyuoSixiUiziSCW6UpZ2jlurEC2FuM4xnwN42Wa5wLFSzvxwN
tfdJPgX/cR0O8sK+5UtWjo4TLIEzGVTUAWGD6XJUH8wuKb7r3muuAh69cIhTk5Mm
VRHw1OVkG7c/nS5Tsu7l58/szHEwXcoF4E9GpQIhBPvYXi2BCYq2OfxXTyHFyE3n
F9JymHneqfr3mCBeLVgsawAqfX219SzhobWuY17fYiC7T9WCqIMf9H/6359IriC6
hyLkQ/gnqMTAao0wtXKPOkcgV2hkEQIsY932hcp8vnxH7BDXVRubJJTwSyOEBXUh
18W9woH4G6s+otkfIArGGeYiVzO2d97Frzux1D/xOd8p15iuS79zLbKFSlfZXT96
jZkfSDVkn4Uxu3DyaXdovRtB1XXvrgnoOZkegVR8D9u1DUloqUjUKwISBGl+twoo
opMUAhmYpuRnSBE12nE6iCvNd8FTF/nD5103OvfTwqhC/Wj/Uib4ZwjFXCoMglwg
1hnSF5O8Sb8q2o9Z0L6ftXDCUIng+qvBd8BJHxXrt8i9Wpx99x2wW3K+TUBXm6Ml
O7I7Bllb36CJyxx0iKiGVi/ilXaIy6ccfRsVw8GPG3F1AtD20od9axcggp6sKQSo
K9/Q0B8nds2VFm30dGYD1GZ/j2v8BblEnUXQY6hibiGpmMlXTDD2rr3pLHXz9UMH
FvmIPddinPa7eh3MfBvN+KsPc9DJ8j22Zuxzd+6ihtyoMwR9SARVzbfuc/CHz9z2
YohiDjF5AL93U4PdCyRrW/94uCUywtmVB7VsSz3M/Rob7F4WReLMH9wxXFdRZck5
+zNE6qtdAIWWWt6WifpbNKnHC7CXRgtyGRdiVTqLVFy7jhAXJBCy0ioUVj8ZksXC
Y4JFIXo35HRkQ56iwNnAHEK+17kMXE17++FqW1RwR7P3cwaIgvBugLn8blWtjPuy
z3muv9eEKzkWE5zzGFHwtFtcutWKjbv+VfEqxCyeezv1KxIy5FvOYbP9UImb6aJF
sweggs33SU0EcVr79NYTgLTKlbvtYbxnx9hdVBy2QHuMzBaQP3xObyuRL0YHujRv
/iirjbaW+wWLBoozPViY4hXuqfqAkrW0C1fhUAN2ZkOl5KEteFupOurn12w13rQV
YYGfrHAmZGfGRiAeP3RN/drxXt0CgjGvQmUB6UVNapByRaxnQNb+ejiVs0wtQU8M
o8+1A0v2V6RGjO8k5xvkdZY6a6pzbTOUWIjTYkpDxNiYeZt4rUvpde2pjQqd6pZG
WB5GG+Q9QrTR7OQEL2XjPQ0Vr0wdgO4/heEjWawRi/Vue6HlHukqPJHbSGQLHvDv
TR/+18z1U0yYlOAV+pdCFx+sfqyLPgDr3XnvQaSEUs9Drg0gEkhn3Iq0jwv+AokX
yXSqQ9DdGvy/dchpp5tC/teaz635DebbITSOvmZ3r+hZppzFuEr3EvgW2Se7xIFT
5Kcnr1oTFyCjUt9C7a9SWM1R2cQI5U5+/9L7RLA5KD3MusRo0GrtGtqZGGICZbI+
X+q4du7DFTv55KIWrVqLy264bwTkRx6APWZpgtogx25FawF3qiDEcx0j92Vn5Vfq
/x3ChmRbL78Ll+WjpLfAx5Lln7UBgIIEeEDR6D4cIyEMckNskaNZieezYz+cVBsO
xJX10gBBBxnCW7mfemB+XbRBEUZiY7fqZoJWQtvKWTQiHcffypgMuzoA1CbDFUQ9
he+324wiX+2wuqsiu31gzxfibCg/TXydfWV/O1E6NY+w8zRDddLtrUBwahmTQRS+
XoE7nbWLZGEffORU+zP3pmz4HX/SMbIKg440uqo16PHt5dP/p8qOSGTsEpAb99Gv
Io9zhe4yNYWtCKD0Uh2TkcTlk+LYlnnl3JIvvjEjQ+c8LbKcEe4SKpvMVqRR1hDm
op0psU1b3Ri0p7tdU//kYSqNwoF9PZZmr/tBp/KFNvaih7Vot/KOFPG0xZL36Z2+
SuIwOwThWEfmVq2lfyD6g8LPvu9nBWnzr+LDB7nzTetHcOmAzCb5cMtR5fa8pFOE
QCXe5nXUoCzQcUoGkpgyj/E+VOjWdlcl2x6KKz16t1bhWP6fulWVj62LHdzmsoLd
dkVl79dsLcHUK+x72jWREOgWYs/mbWKJy+UH+wvfb3nOp/uvqu8S1KZaF1Dv3Fmc
Gv+CjbTyM4y3OlGX3jmG2zJIew5VXlrp/SxxCK6Flkre+pDGe3/u/L6tyOpxHX09
boEflvYknEUPuR0BvYPd71LWTnb8Y+A2g4dAkC/gg03m2XESg4QaCIujovk91ao1
9lcoAd0dLXre9BJZeRBGEfm0BR69PsTHfBcRBXyQIMgSckK+TQ02UVKOLwdC0NLK
lepdOzohUqgXsm048AuU7x+bCn7pWjpWvRb1/6IKLynLVZDFn3BFj6pMYqw5Ww70
+vQxgb7yC6qJt0X95N6pz/lcGtV/TtAtzYRmJnl5CgrzNSyLPYepAfu3dS+/jxEB
vcWtU5c4A3VtpS1MrCaUNQepcZUz+Q/J1+Uaf2iOA9qRXxp3qa0fJCcV/dl146Ek
7RAUTnD7lNH1H8xWI8n/iyRLlZQacAKezbBOMKdfrqFyCPw+d81HunodS7bLfFxj
vpNB/UxXsFW0l4tFJoRZ/c77yagqx3MHkJ+dvPJ3qIVLn5WOP/5aMEKR091JcD1C
dhWCyo9DotK3ILN8HshUKeJrilmcxnh4NP8hpCM1m/AYxZG337e7SMLDXKuRL5kf
KqjblHdhCBsn0lM6ws9YeKm0YBXIZqJPrhWO85h/fipieoD6DlBO68hnqRMrG7mx
T/3jS6XckuvJNN/8XY/ICe1mF8R3tROc3uNaQvb2BGunRjFPMKN4QzmK2dA6rNon
1Aiee+gZQylBndkCtKYJzBAN/b1mqAJhvDUYYxyK3QVnFUJs7yWUmU3VgdQJqmh9
0ANuowlDXxNmKzLaLH8F/4+Lh12KIgE4WwRHfkHaPdLCmCiHG3uHtMx7jDfpTvjj
koqD/q2pQQyzILnZ/wZc00G3B3raAd/0laXwtHlIExNcLmut4HIaZs2T2qB+EB4r
6jfGmFxueanwFxqIJdiS4//CJVKXZ39bqA/1ok2fwduSLtnxWREy0rPEExYVp6lb
MMNJCpeFbnJ87zQA1YDnwD7mSthghVPEFh4AnJ00zCIA8saUeD0eiZNb87YOpVGg
pl53uI/8w83DJqhaRLKUuo4lht3qmkkOEOhNCGG4DCRUMUzQVciQX+utbuOCOPkr
wqc9uJN+rhnXAdU3+kqVBO1+66tfoDV3wZzDUZJnVlofe1V4LOJbXKnwEGJchyYo
/NzeLQEqTpF68AfFyR6GSJFS+X+elOo3ZgYPp00qQBiE0Nu+A/DXRLoySgZGZVgs
XV7EplI7BymJP5/8jWomsKLxbam1qvmGWr07UgysnSzCU05WVlA7TeYPFwRr6uXL
vpLAa+Tq3lWjKL9TNndTkFlsmYveXzwdgNTfxmFXbf8WH+U5PEYb/a/A9ketVBkE
DHT4gpi8ogcrjXCOhZ8NXWN/uTITiYMerlowroeP7d3mzGmwWeS8V+orans+Qaw/
fDhzBxVsRT9yyOH5uWVRkcs2KeLoBwvIABN5tjNYFkFL0gD/FxGETmuYMb7uJr/2
UXJqXmPUVW9hog2HoGVk2p3yGqeZ/dv7Y1e95o+PSgVK6xzQxYTBhWd16mafsh+2
TiiNz8XWDQKBOTAJxhfYvfmMBuToK+PujZ3mdWnnpdUTlCjUmf1YY2MAAFFNKy1b
Ca9Mw6/gr+XPC8DDCAhoP5waiWs+aj3PhS51xwOfuLGgZDdggPlM3LMMyw3zbj2f
jrZolHaWBElmJ29J6+ZX0A0j8SFQGV/xT5n2g6BiHBDNCE4HaC77UC6f0Yx4rALw
wfkWTWcLVonLseorfJKqT7UMpjn25KvNoadkhI8/wMu35P0kgnOH3+WcMfiFlFxM
pAZ8U0UhPtndfNjiYTIzwen3O4RaNxazV+Zko+GT1iXo5JNDtfm56TZPl09KrZfS
PMavd8yWvpU1/OEqISHcejELFmmMfmvBgFbv5ZB8BdEjmUTGqQe+V8TmzRDiI450
FOd6WGldfxNUCD8NJRypSwXiM4p6JkOWRfb0aLO9MStTJlJlg+apVrKtbeRUlKb5
noNFrbN/ZnDxzxZq+HMWoIBFNkSQsV4b9Eh7Aq5xFptYuskYGMRi9//JYMiy7M86
dwQUejDy34bGQVu7i6G5mIf0qyBm7swuJm+ARD0ZMIymjJ3HHnwALuC6x7cel6uZ
CT5J9g8owJGydrxtS0Km3J2lrGG1n0WvIckFUBK+z4UmcgHMRJmGNeiNTB7mMMOh
EpWhPq6OE6Ec4XnSpwt356bQRWbbWKR30w3+kLTo1lcwsC1azU1V/AzxYMQ/NKY+
8v97Z+ot4e1oFfPxEyFVuE2BSVMa7ZhjZ+V6/h/Dk+h4144BUhTJEtkdyRmngDZP
E8EGkgTU7o9U7XRxwQYjd6DHV8vtIDkAdFAbwJzH9S04hop+7RfkIMoNp1tTcxG4
TAal4AoT1u30n3kw+wWOfwOMyrj0MGcgsF1l3XUznCdsG9SG13oIJMQ0lbB5Vm2Q
z8attEr3nkekSPutwnDXForQ2STReoRW1wlEtjyyApX0H5DWsDSnZAMRHSLUXASU
gi7atDtHaZo54vFm876QzI9X+9gsbtpxv/udGSPO6NVu1nFoc3f1SmEag7nFw0/e
mEKnKu3tzZV13ycjo2HAAoujgtdTNH5QiFDVMLRCy1vhvZXNLP2GZZu11zwiwmxT
Sf/9OEC/hfKfhrX2132eF/C+0tNF6Zt2nwIKeee3DJa2ZyCy78Fsr2g4TfZYqlKu
+yzJlkkMSS1t2Jh0ZmKCn4jmZ0YcMMvMCw9ypxozDRkfl5nFSvFNqw7+QHwr9flp
BH3NAyBJ1xRjRyo0kes6HPMJwxcXC7qZptolp7fueYNvyxG1YeEwwxZWotihro/+
cBaLPEYH7mp4Iwf3KVrzOVVFO1no46PBk4AKHuU1az/rL/GgbAPdmE/1AfVUH6/q
kZk27OOCP7pE0fyrxzM0sAXK6ToePIsAZyEedRh9kXaWv3UmlcGHNswtBduO95fh
4LMd5/HTxoWdyZzhvO8v3W6u6qNfym5ffoLCqkYFXQPeLxs1518laN6IKgi0xStO
S5M2dxgb5/45wOWdAW/n0DLyohTlfXiIdikZ6TLEEJJQttQkznWUFRxOHq/USSj0
Blo1NwNGZesQ+qwfSrs7fYC5tuvrqe/jyChx+2AbgHxzbUbp7r0M64qGLdeEgg3j
zxFFfMTF+kr9KgeUkivY4CGd3LpsZqlaJue2tWQIAZKJWO2SzN064C7t6AqTc0sH
o08uMgi5oWpjdZ7kHAo64lU9ArSLBFuSHwC9oT3yj3BTjMpZ8GTE2bVKa1/wxRqo
d54Ot1xKMZUL9XJ0GbwglExp5liAWGViOg7x4aA96eqZr4eE0Xd+HZbRAlqJKAi7
9TUS+Y4GbP5WCQXkzf/t7NsbOIqNOTsV82b9Qn3c4B/rmKNIx3hFlABHhNHi7iUR
MMqp2lv+1z+dmtfc/2QXtHQ4qWxGDEByl47Khwh0ye+/h60jcYAQG7TwbIAvs6ko
jj48lLrri39aKifHDn2sQLXHsE/XdmJyptKUA085gQMBTUWgUSdtJ4lyIVGIPhmT
09TbVln461noKiyptoUSDRZKQo4a2kOhbbkvNjSmfs84BsFp7PfRWAABpTqt8/cM
LjiZCTXPcJD0Tilk2IVqRfHhnLT/2fXpA7qEmnfE0Hc6Ecy3RBq6YXARIl6W6FIi
Gch54+FLVzUl24JZavye7EESX9bJHgDz07zaHo/G0MJ/IzANqFtDWOnbZrAxLQps
s2vihcSsT7N4ruT2Yv24oIus4fN5SUc4bRrd/WJfg1iR1p8LXqAMtOA7IMs2YrIm
kFHwwKsrbSBq0EkbvJgcvjTC90z5pi68V8omoVlCS/GdImvO2fdzKz6AzRBGKTVo
s7cgG9mMXGshTluFBE+lqOoF0RTIfM7E+XgpMp0bLnu+pqENWw2fzB27FEILF+B8
3ExqCz+F/fz0uRmA59Ms52AJ5L/uesYOTVVFMb/DVBkSIPpM32joMfADI7Faq0CZ
Cg4+eOItsqLuJQCW2FMYgjkihC96LXqvMxQKdTC5du396eC7e0ZPswpMJWXUGK0M
En3wQ6U6voj1VW9pkoGtv23oJr0gXvYi/GfUf9jbojSVfB0iCXfBKTTouUM9X8fH
69+0qm7oT0KB/xN97IG8rgWaP+E1s6sz+/2BZg3zeYG/4ijGCelffVxTeJyhI2dD
bh0U4R7ixF8H7G8LzQdiZ0EkK385OgEkmSaMlU9+knOfJTkdUGU2FmIMysSCrXMM
lECBpVPzNFqJe0LNVtFW4665IRwxYhnALpF7p5Vd+/y/GF6QNfA7xYXEVFUJxALw
Z37AkGN5JFzCO20Q2xN+fBFaVslAPsz5ONPRDzSaiwwTuE9GRvmscggdP6qtgvpY
pOtTonmX53/CmpASq0zsT0aKxKVQr9/u4JJIjFMw4DhaGwgnrpX/lwAEL7o/kd9T
xem1JQZ8XUnZnQSPcfreNbgv6x+l9OQuFaCy9dHCyDZpzy+gwOsm/JOaXp73L3pp
hjn1oLY/2oTljSk6a98fTO7IsQCBx0+F76Zqrrrh5ezPDzlTo//DINN9SrRUQCeN
8W1MVWzHu+ISYNd79HpDOG4oo85U48DcsXnG4k5HWaIo0GGZ9aieztGaz0ghTPpG
9SISbosRAzp8phEUfGc0usgYixZp85Cu3BnFTdkgYUN4ovFiMT2m9HxolyDVxL1q
V7zqkWCAnyiVdIgQDb72cPYvjL4NoVf6WagGCvEtqTuzMFnE0QiDrZxW9AGM1e/F
YriXh20jrTta6Hfsk/JRPtpgH6Bb9yzo7LQwa/5g+/hyISpT/LQI3g8qQ1jYQeob
wOxHscF097ul8mkhOm2r/F2aYYNES8L6X2xag9/kYI6VwNiCS9LWKC4EflnznNG1
jmMCjITlU2XOdODK2xSGww7sWfG1XWR67xKhE4Ry7vhqLaU5Q541ci+9T9J320kV
WIHEjKBbeP+++KLQOVrxo7JSqpus4AR7uPtF9Dtqs4vCXqYJKU5NIn2MaP90kNeS
xmZVQ7RiMPlLPYA6EH27HlElam8nykkHSyMHThe7azevAC1tVp+4FpnvXtC/j8nk
ZMML/unxHwWn8fhxfXA8uCYLjFwmLtMuDLPeeg08N5GHUsS0IiF7GJv01Ar9dM4z
BuYTZkglZ6x0vl04Un8h2PnQUvsMKPL8J9Ktw7lq4Xva9lWxJyipRglFJGpCEbtn
+j/mFHsQpF1pOTxmjy8C9r+EuDZCV/JXvC5/uCKe3GMu/yj/VjcSkEojOVdUb2gG
BD+1og/k6QZ6FewgzzVKcKuia5pYZsKB0r91soef35ddoyzCEEVP0hZEQ1SovghN
oT4PZWGpomdz6xM3tGFa0ZJW89bwvZMdekkvZ8FOPdqkBzBIVic9BF1EMWKYsrwc
vEhKCKWTNVB6xnigGAXOUEfu/snMRsaxGR6vqh08F8trGRUwurJF0zXRIdQcc6Gc
Q2DzHgYR76oFe4LQ97hTpQFLRgMzoiqpvk/Hcbnp7OElPD2YOtPTE0kbaAySNXO0
pwL7BqmQfu7bq6ONGw4Nzn3Ubil5y8UXWtT8vByyHXeJRSElt+32grfChQcgo/FB
/gamyTv44aenGwKeg6qbqYKTeSk1EP5O0bEeOvBvywF0TvMNqqowphFLMasLhexz
0udXVxDO57nwBw+1R6R2aPX1s6c68PqLBp/4X4mPB7BBt+hZ424Xs5JZbx9zflTR
CTgLRBLJQ9zyw0tJyhUdDa9Wt2SQ4uwRR5zzTzXmgJ/OnSxWjvuQLFLzeOxUKjt8
PC5cYLSwMxOFxnvLNuV+hYAlDxb/gQSUfbmVrli0Y3O6OCSnUleRZTVp5T/UkOaM
1kGREpA7v8z4VHY53iZ8vsaqwJwZg+34qKl4xhQPmtG0Hl31DiNW7iJE+Rs/mQ8L
irU/vu68E31VvB4dFTOo9b3paWRvDKRpDRtJo0DLlj2FPX8372W86LfPAJm6sN0P
4ITxOUCZTwJ9LLf/bPivgCHQXbNeycm5PBmzCnpKzaM0j6yMdVo1ijLdpL+64SYd
B04XdWj51Ihmt7p+sgid3DFMgaWBC7eyoj2V8+X5WZ+DASRUNiRIEJkgPx0Kd3fq
O/8un8vPK4SGaGpq40tMLoSEAuWcBhK7TObRobX5oG9/JaddY189jnAmN2fJWhp1
HOsbL2TMmInaTiw9dWW6FJPhp/dkArSBT8dwwuudT8wO6x7ZOLE/IbdAwaIMlRQr
gLt2eyI7zvURqRcZ+qru/y1ca8hW6oj8lU1tLWEo01oOFNGjAdyLpr7utdL9MrtT
r3SGUud0uwsrZ4K1b/k3oRajPCSYKlNw3nD+lyKm6pTpw1ZTcfqVPuuAtvY5NSRL
RtQYac+Z2kx3C9L8R7Mt+nEN4KySsBHjwyBz711ZTqw0Y7Tr/TWmk2zg6874GrKz
5NNG8Cr4pqSxfx43xucQMvIhbA3SxercWI13/rMnlxzWsi8cIKxcafF685NaePlp
hvRMaUHMCKnKJHVNRVz391AektaP2p39zbBAmPxFgda5eAG1qd7t6MG0wky0VJcx
+CVWX7bCb60Y67Qrzaz0Hnqo10QRRRNYGSDfmewMpse4fpDrGxF7JjV83eD8RmlG
xyuoIN0CqAF5JWV24rOM0qm1KzGey/FSsWjf/xjZD4CAicRQxmuBzUgfogRE8mwT
iDiRCo6BdC76nyA4EI4q/Q9h0HHoeYxTRw2mZMHRaEV2qCzjQjCeNB7MU55YoefV
YAtDBTsnOR2lsQWx39XCRiFxHixyymH0COe85+Y+glWP3bN8MNYy3Rj/xjwanmv1
owvcimESJQC+tcztvuxgl+50cKQVWVCG/W3/oJCtpHvpvYdfJh19AW9v51YDnCdW
KtK/3oY743S+RQ0UPhFdC3K4odJc8Th5R61i1vkw4ZNdQqPMBAb7RGWlZxRdFz4D
sj3aZUqlzoeqXcZgBZwDJzzVnuy8GAh6irNWpz5DP997hBNlr5WTinC1hXNIq9aB
y8NVY0z1DhW84iUE5eUaQlUBoaLir/QIC6j5/BDC41CLC5yD2qt11jH8EJmA6pvy
Ukggmf1G2xP6kt6pLqgcWSE/uY+mO0NWm3+hYujflJSvYQGR73ZxZetc7VeBbNsF
foO4L9Yuef+MfLz4+xyJ8Vcv3x+c5WdhLYtbTctmR7jFWvpbe3ltFii/9zk+oOwy
XqR3qTKLN1NRit+Q+btRrEMZ07O0Iyay3lZ8DVRi3duGMQxzg/c+MRbHACKkgoI6
F/azb35TeDWyvc1Ol0niVXgu71EOsyP9ooCB9UdKx8hnl7YUuHhyjRYMIeZ4zXut
42X3OFxFmGPofhfotpdtnU007FZhuWXNdiEWG4tdxjM5dZB61jR0bZzHu10DC3uj
Z43rIVDttjY2zWwD5Wlc2fMbxNChhE5iI65EwkBViK05A1BhL0iFnuM76NfI5qq5
wC+GK7ehpslZWSPYrDDCU6IFmI3qc7LgwtvW9OOX55d1IKcdem45hu2yKr1AuV4P
ZMdGNJiRedM0PUNsh9rwZ3cl8x7phhWbNxlDB2zFXy9Wytix5Cofiq1iaRkx4Sg+
WWqbF33T1O0ZpJQZkEGw7l7Yu1m4d4aHmMLsCP+QesSiACBoQAf8vRvJdOg9e3I8
93fsbntLh6Ixn348zC88JlK5K5ai8rB6BLcfyceffD9dESwYLVBxFljDqT+KkJ1y
XALc+MQmAeq9Y7WM7bfwZnHVxvoLHR9rsc7YJBFXhz+Ui+zTWrA6jI1VLC1ak3qE
aW08R0kRnUcfiL5qKQu6gdtTqQV2GpEFh1i7Lq8BexZBDrYxtgI9+mv/3CIOSI1s
XiCelqK7XGi2K3wKX1BfiJ53ijmkfUdK3Dq7HnTyaWEHmxhIYeYVGQyjSY1a31XK
Yj/lnqGxsanOguZewv6LkeCd9iW0jjVrEBEprz6XQFvuc0lixMw6pseXGBs+MbVe
ESyhQUznT/60RAVdwCn9QGlIjkwmC/3WckxwWmFlVhEcUiKLmy2se99NbBN5Prqv
7Ocp+Zjilcr56MP6o+nueHIWbL0jUphfBvU5Uz5N/4tmgCByAglWCNKR3cMV525J
X+RA1xaKspRgwknEnuTyOEoyxx8jszcPrm4SAag4frDvPISDj7xe5CMr1Ffeg9iz
oZDJf3nFOMQlpT64CO8YZse9dT0YUb99VN1XvJMW4b7yBEGybpW22Bzm+LLgipoL
sCmsCx5AIcWVZGtSyhzIxCPLp2Kl2qX/j21YMMTqa302F1J9J4RZuazjvuIdChbg
cW+GrF2jPxdzr0ySLZDZUcY0OFriwKkPg21f+Dv5Ac1RddAaaSS65A6vcoUNfyW9
gd9gZyhggnQGNUg8OMhiNXc0K8IS51fgVBMorgtD0lNM3c8f2ro5nHF9KoFxpG5z
6GyAzhECV/o5pB6yTMCJ2sJHJVxrQgJ9eoPpDtepdMsKEfMnW9biK+U+EYsE9ykg
pfc4NSeY3yY2zgI00gI99mymP+pbY8kgZEBUNXy1wS2N64Sm2bfZBpt7E27CQxc2
PQxYZ7YB+SJ3AVXmkOz0XUXv8VINPq2XoTWmrnsef+U4lJqg9nZ/Y1nFTqYxMAfR
8nkClKC1h9k64ocUV2GK5nlHP3a+rwUN5HggEcpIqDKKrnYwAkTUn7TJc7mQxsRs
Br6J1Au0xWZZVBP+2c/zBfVPeAyH31fxU/CynTw/pklt/nxTGFhf1osg7rpj3n5W
cGb4PvC2pcMacCQHP7nvE2ICvRp0TrkZln3gLYLQFH965yd8Jgi2ZcYlGIxxoLWj
YvicHCxhP7tgX4jwVXtPs3seKEgk+gCESPUfHheGwd4Z8IXAiKeD2rN5rz3Ybo7u
2HKq5MPmbys/NU4Y2Q50/O08sTWXxqRBRimwAOkHG0WAnRU/wrh/98DICDMINkNR
GCJdjjrW+1FMIslZFHlPG1RxLVyqKx/GSeZ9gzL0+I6zRN585Vf1T4qJvvHqeqSc
yDMX68SwOh5Gp38Zy6gBEpLOZzQsY4kUj3CeqsNNsCygPK770cMOICZVfiGSbnTb
omWanp43QQltxKKG81k4BoJe7kjcD6TSU2homAuFV53SK2K+JoMOp8PPCaRcRX16
E8yx1+pyoFeMcjNCfqJwTlCdBvmwoop5k/9A24eh2uO15PE9x/fYO9JsO94oe/iF
onwTjtGX+hCrFnbrAv2bPS4kzc4p7EjqiDPR3L9d7PyimGG1ut+IgVwfNiLIdcnn
NHBQjsVm+gs+HlEM5UGqShPKlUl4se98BnfS0b1ssws1hpgcfbqeMpw2q0swmF/N
Yz+dy0JGjDFjBx33U90tJEh7z32V8iq2GhkPvtrPFAVmt2bFAL0iLmvmvXj+YLdF
RoS5Sw/65ZGa+aORRrZbrmz3WMPgxCFcvmRhg50DwW7R1Bjtutvy1+flWjkdW+71
UYNUDev+QswlZLdFgU7ggNSAuCn87ej1TH57H/IVu90GD4EpoI7dGobxDIl9N1xc
LXoObW2AXplhPm6whuUnv2blphC/YKjj6PjD1wvm6NuJKaM9sZxIzsegalJtZfMi
cg6/eLYE1MZTGguij2ZNHoN+oRihmEJQawkRr344voVEp71nrYtHMvjfFa47Xk9/
ZDF1ZB22sEGcf4JBBFGmBABkUuky+rwjKKqWJsw1WhbtcWRFJ5zvlcuIRsJRitsm
xg8g6454L21IGo9j67vraJm+yeXj+VAu0kU+ao4flhtr95BrX79sGSKyRJfZyqpE
kB/gm7pJXVM+2X3Ob620Nbkp8TAXKZud8+0Jq+VGoSnBOrWh3JdNFklG5EqNdD1+
kySiobyAX8U7MbI/fF6CCCY1kK/XHb7tfxGCwwua/2us1+HB3csknpwz6uK6G6oF
nTPQwNfU+vSFY7BHdmkA2wipe4kjYL3MNKxyQ7pLdh5ciVgQR1mMyyFHbfab+ZRz
+BBm0WiAx+H6HfPuxxVxUuY12frGxD5Xo2gozfW28kUnVrO8UTE5CRN2suW6hqJG
VU+lfa8S52ECxGcK9IibBPp+6KvVtaT9Ek4fv3SowhmoNqYB+RpoU0cNx7i/egHW
WV/orqUt1Iu+DaZzkhAnWt1KnubK9v/eNprk8PTjEfHcbsHxOip1EIblPRFmhrHU
k63qf33sy7UeT0EpEfTRvamGBPp3YZ7vRcSvZl1H7pVulwUwEXkrQ05zpFmiS+oT
AW1q1fzkPnnFwlFESxNzLHEcL85kCgp/n9eBhS3QloQl4VhHBnhpsGcavMH4pUdA
LxkzcodWxKXc59Dujy9mSQyNmboDoxDqGU0XdGIduXRrjC/l0is9pQEqzo8i4Htd
N5u5bnjudLd+5szUpjN6BesdKxNapvyahQ0cqqTiUUmJWQ3gRAi//epZI6omQQsm
MrZJ1GWutI/mnPtriVbYrRRJWScVthZEzBIfmETd3XSamX5V5dDd177dfmodt1Mg
TZKZtZsY5iiXEa+Sn0YKru3fQmuY9McCS1KrpBT0kF/D1U/+uVtPGuKBOEwBXtbT
WcbiCmNDgZ3amvdzIBH9aTzgwtfvG2TeW4cuxM9NPMvuijE1hVoGdnYMk3NBoMn/
H6ZSWiUTAAHiDL7HfTJ1TQgWSFMbJAruV5yXamUeSTxzJlixZFisU3h5/9fVG/xa
NehGZ5ZibNY1lJyu7fUW/pJWPh4JfM+9LUQsn0zLvtF5bmoE6KX3cOoFYh+IbgeP
2BlReLZp6iCEdc5Xi9E2xADOz6L/q3Bk5Z8uZPQNQNgw3z2dC7BmIMFRzhqrPlQQ
l/SqzVXw+QJSJx057KwepbXx0M3MQly+Xfew7qJ7bwBY0XaapyLTd+ZaKTYM+6CP
+bDE9MGmliKFpeTj3uwM7+hJAFAsZ85RRZpRXMdOe5VRelsiakJ0Bp689EbC7/I6
dtJ30x5SHwW/O7LvJR3U7NFxksXhqHb+SxSNru4fDh5ky262Pv5LYrMnJ/wsikRp
YXyy+ZFcOQJmQb9gmzLC+PzFlBH2B/aODgGeXYk/nxbWvkzbU4dWqnVQutiOc8Do
Eh5RTfNvx/V2Wi77LlsUuTdJdNlMAalZx6KN11iu1eKiDbfJdj1BSudssE7vEDX3
tVdX0uyFAL5o4IOGTaO/HpAhI6vIRdSfXpto5gFWGpYkn9Dtm4WPjZJ5TZQH+3kp
Dlhyyx99FnRlebXT6pq5oakoIm15EoOUHhi8tdC3PvbmvF/i61wgMPOpgtdltjoJ
abIl63PAxYQtJpW85e20wf0a4g0pWv3Z7T5ZTax7WkmBFqvaGuk6oQT2lUFfIGfd
4MkSbPVpCyJEjVgcXRB92/yYjtuq4hfMcFAXB5NF1EOU5DdI1MORb+aU8F0e4oTz
lM8BCXqBWURblj6TEgN6YIbbVFLOmYO2NW00aLmTNyrusOYWu/QVvh4d+7AZrMPJ
l4hZX65oDK4oErEXvyoxiKuyRM/CTx6oOD06I6/vgEOLu7FHZz7a5uHAgPrr1QHU
8iD1+M/DrZKIYG6c12HVH/VxIId9bCJNQ7FnMPvkHnsk13l4TPgrSwYnunUZchjL
DW1ivHIoQmctjmMtfr6VNkIpsrdkHZDX+V9H+vtB91jFEriSUYFG1Ol86woEV7gq
A+KeUSr83N275NmymXN3vHSUdwj+bwxuKx9r560nr0vyoJbD6GyvqYsEKFUVInsw
GL9oicBgE0K8bdfkGwpJP1Sr9dqWQWQlQLSj9veXJqtQJdPQu6wLwZLbodkVQZ63
hsR6VB7UPn8J3Hv5azgCizEGKuvWyrEf53aTcQzGKMstM6ev+7o/IsQ+4K++OmNX
RI0R2jE265QAfkJTsIxWf6eNClEj5Zg52qXlzi0dkZdVBNVpv2Ftio8ua6szq2cc
gB+Ibmje4uZweQWCv4b1VTEfXi9KTXAu86DhrmDIppAdEgzYsUteTkYTRpRIbw6c
hR9rOjpMBfOcZKMcRH3hVqK7xJqM8hjv81XOrVrnL38Zmsc/Vc2o3Pizeyny+HKq
C11gvXI5UvIYVRBTue+75zOB0HnqQE6UUJuzFfVB+HkJy9FBj0oyc3nkrrsJOAmz
uCzmZ4yRKe68dlrpebZnBAbDiCev6n4pp4TL1CeIei+1vRSWN+KZu1+xIEgfNKv7
0wB7jZwirzsAokgNUXVpVYtlbe592TSBS6fqH3WGJryd7/gLeY0elQJv12VPHx8r
gZQ9eHsN9YaX65QjwMsxRPFzgeff06OpBErKQJ1p5WKfJLJ5pyvfkRm3BXftNs9Z
yX8iQjqGpr6mhbzJ/oVNAUGn9dobhvlMhsh3fMMXp3q+V9iFe0zewwy7B9DYdToc
aqc2XsfJmT/Omv/Nt7KTQWhZuX3sQc2kY7h1JAn3WFBOLIko5L/4kihIDsb9Ezmh
GwWIiR+Ej2OlHmxx4vu7ftK5cKkbUJSylJHVr/2ao6/9QqWbQ9ktasdLL1kdX9ip
T4jEcmohsDEtxE5/nfqKbifcjV5DtHi4hDkOvSBW58/ZvkbrD8yQrOMf2kRWsEwP
tIBQkdMFQMTs/fK2s0FOrVjFdgcsVS0VCJEyo6czbbMEVq7QSPXpl+6wTJuEVpTl
ajh3HwbWEigc5yWru4HdPQZS6C+RAqq+L2539nsd6mtJyZKqcMCnx5VK1EmBgcoi
aSU7MoEoHJYQt3AOkSYxKvEBFQd0XjoJY/bvT/N/m7ymkX29ClZsJkuUIh40dOfI
bCo1YwWbYTUdN+p7kQPeIOXxlyg2yGSzuGiA7QtnYOfEURDckd/vxGb9eq9bWzIT
Vwa3oT9ShWyVlj0MarGLpNe7wuZRxNv6wIbkXR8v+7Dk7PcRzE5FEG878kMDcrGv
MgbPxM9oxftjeqDMyV2kbymSZ7v/rYhfILgd6b7wNe09nZ0u24pl9weGfijraNgO
uJvFIFvGWUfLFeWem4csaV3UTVb+BIW29m0t5RhB1v29TvZYmZ0CSXg7zp3hnnqt
8Z27pSn5FPCoPUrI6alnUkDJPqSvxRI1Tod2xRDlLFCJDkajwWujXDmZXz53o5xl
U++19NWnLiBvKgLqnkQrjlTUit5BLWymTC4dVGzEfiRloAmBdGoZquqhB1zAD/ie
OiUOPf4Frgt52z2CbQ+u0jeOfxGcV7Z9BosJEsbQQ6GpdIXJyIb3O6tGvNQFEHcn
3KBLMpsj8dmIvzWPoS35wNWSyogoIzo2yYr/De54V2CmGBYx8/7S0kC7o3dWzEZQ
SfcLFW9HubSX3o/S0iiwZnQl2o7BBXiSiu+sJH/O1oUQ2/88pm+VyuY5iioq2anv
1yzrl93ur0ZJSjBZ+92a1Ti/ZT3HA9XQ6ePGYXcrbNS3RMSWVQf1gyLqIjPBQkvO
5QJNYlrtoebHoZkIPlwlQ1kLI8Q4V2IVn35ACPMv507Fm4Q8o8hLYJF0GwqsbvAq
UJg9w+KifDuv9R+1bbMfzlE9mvq+CokZLd7kNqRy7BK0gcIuvkYXjkOfHclD3yFA
ku/vJZx+fJd8LxzYSPi9DMFg7w4o0VPeeT7y1E73yME8MbquaZ99fV/IzBM2tcZX
hVBrTApF3H2srQuxAXmd1egWJQ8drT9dki2XdnxBi0rqdJh7R9W7T6DQ4tX6jPVb
RksJGM1BU9yTvftP9Q8B1/8GhoSoq6mpqniKDKO4cFMTS3VzFX3fneo1Em5qaC1R
WhxK0g7gyLxFQFBqXLqStDRiYWqVbc5ssblzma3QSOjn6dm5wc5ax+dusCkyLp1J
hfeSIAQfbyLRiUP34P0RE6XiI76ruu8xNqsXXi9lKb2qblMYIL0kJ59h0g4EWKcj
40pGoarpbu5+cD5G8qS7u2JPvr7yESDYBSle9xRHT3wxu0/PeUf9zh4GpXkHMI4w
IJ5XYzYppcWNRio6zL4jCriaEtgPdp2PvKIjo3ZlX9ph/mqUyDHJfBa8DzRO4ARV
B9BiOqkwM5bbUWB5+rn5hukW1sZ7u5u/EqmkgTy2Q7GOnWFbYcc05XTyYuUJ/0gW
KCZf8bujTKcsYiqyO8EjSu74sB1NMZMx9vquAEHmOTYtirta9ws1h2BNDWQsq0sR
RLZiyWjPb5K6VAAJLgKKHa2kN6k494ORd50F/Pn55byEpResGRI32iv6YrtCjHh5
23+TnBZkNiRI9+XhUhkOiyOZpem1RJVZkgZz8dlYmsyOYX/ro8MjqRxiRuK+vwJx
Xulfb9WXHbJK1h7gtQtOj8lEk51vtEF3ot53ysbAvE5VEY5Ws3goX4AiQ9VI8FZP
ErYBiz+r9yokbRV6tSgpZ/9R/XWPcKU09XyZWFrCTtgkNeu0xWsS8j4gApoj4U8v
AK/T6Ik2jY5KWTlQgMzs6TclP7ZOJ8CUnUsSlEccM3d53y13ogaKCd0V7rnFWjJ2
DnhdUwFoMePtZsRNTjRIjIsTVdVxLnar0LO/FxflLfdDfZk92sXb+WFWwj4FEuO5
YA89qVJrmbaM8wVxOLwAFMlvXCTj9y36xRuzA074PLGVargJ9A04nAa5lPXrj2Zu
s/r2c7L/le9+gYACIlm4lBhGEgrgXTvW3Pgddk/VuwWf2gZouV0OtARvkGxZ7L7Z
Ec/ymqD21kmj9HsUCk80pp5A2QMbFubN6etF9AKizqPsPr5sNKl3tH0sZlANcqfw
y8dS2jdlKaGriIB2C9/zsZBz6VTY+ftOOmVq1EVPlz9KLvPI+xnHfu8HG/jRZhtR
QyIqP89YaI/GlQULJ++MGGKrSUkpbNOWtIJC0r3gzJko3cXAXeX3k4egQtXF6WhK
ic5umKGW5Ie/70HsRhc1kOTAwJ7CjVhYhulviMHOxrzrqSDVvXETlgNQQSBuu3ic
uEVtYwy3AYWZOPvAJQXJkOFkckzkJfDXGlpri8wGElAnsJEumejJq1DDcM2tq6OO
6vBzkdIjZu+it9p7GDDZSnN0p5EOu5A+8wTUZN4cB8iy6x6WzcNrXAa4jI12FjBQ
3J3C8sfu1S10me3VRrAGV+2nl28HRpM+WJba+G0OSzPuRWzoVij3wZjoJMsVSNK8
GtDuoEt6WmrpEcmggtgbnhFOLkBx8uznJr9c8wIibkimBB18pvXmHlQHnm/D9m7M
kTkbW0N6biQ2dGz2SGv4xJID9gD4v//RIY1PXIRa2D2CUcWKryeERVb5ePVCoC4P
SdQBu5HhYQvQ30mWVMYnvmH+FzVynqWUuHD5iq18w2KtNyeMPTzoiamNGoPw1AYb
HpxlQmFmE3+THnRlxkC3FuahU3/KHA45jOBK6tUBF7V8pOKxWC/+DuVL50i7isUZ
az/Xy2wQTPA2ZX+Cyj9Y2jWTKuDqFDA2weBJHXMASvPEeTFCy58FujgxIB7HLSlP
HFn2xTJDkGQk6jKxTY4sfv4NlqVm6/Tu4nRi4WSAsPIulNYGSF/GIV0o1WUybHU7
VZMaVxpx0hRLzJ/RH19r7zRMz0xgeIXiMnwpOcFE9DvzpZXoMapLMAO85yJfvKWW
lnBqCbZp0Vf+jiHDuvAgvCk0zOMPQqtnYvkj1Ns9F7ib3jdWQrGDA3tMftmwSLJT
e9p/6/7DT4qOzBD0GT+3GuxiAb3aOAmuLJdMQqLJGTOpxbo5Ldl74PERMARUbMFp
iKZPfvNUFU/I90xos0ThoJzBjGwbdM37xjHiNEr71tb7gAfLlCZIDek5cP4NrW6i
3x8azsl2n5WiYFh66K81WBbQSCyRdhvkClWuHt+4qAB0piTb13dRZvPbLnBqxsXO
wY1/jErQpOXV6IFvpRyO881cVzImpy57TJtZgNHHEMVY7jckjPSecnaKZJaExyio
va32qOHk7qeewJmdKky7X2OFlk0tIv1JkxzQ4dndbACkc9L3Giz9rNjDLvtz7IJO
8OeGsbYoVd47HYKMkZgs7Tk8upUT04/UTHamCvVT14b2qe5NDImjmcKgZwEMFhYi
SsYSb0pDAefCkJyYvNnTI4fAy0mbRaqRhZf5sDDh2rkWXEaUt6JkWqU2oq68mHEy
r2C5WrC5VCr2NbiDUZuLNtJNfarX4g3Ue9GyHpu0my8VWrYhmh+ej0uNKeepY/KG
RNfObBvsJ8BkyNbS0jIi03Dsyyg0/P0gjGMcKIvOEH3TyAcUU3kP8jbVu4nDrd8/
izOVrzI3ehR2dfWHcEnDBpc9zd2LAvEd96baIEJONu80qyeD2SOV5wD05RwCVlo6
M3BWmHtQShiihzHRSpULb++xGHRfnd6VJE5/o1UxltEiSq1xd7wnY15LxsZho1V2
kpizhVgSWO//b+3kkl+Hu1WgAdBO5e7Z4C9Oly2oz1t2alzdC1l+eaB/u/GgbuiT
//QQRkbkqH3bFjQ0VNLJGxccIZCSA7EHSg6mWVAJUbEghNBg7lucCrv5ODKm4CZS
0YigwjT4wDl39SIgAzSE40Po/fCWMSEfFxlzFHx+bb1KenRnw3J42pcxN8uig7o5
y3xglFxorR5wqYRqOY2qNmEdUToMeZAxkpKisissF2YZx0CuvFwMMOd6bCypv+Rd
C2BdJpkJjqshLZwfHICuIpofEHJelGi0M7LCORJi2YaT2ymTFSSKNidn6fYiCDxE
X8iSw759WOd6gActhrC1HyNGmicgNvmq/GnsRAGnZFoJ66ecAbBlNcsXfrczAThN
WLocVhY4uOaEzmKUMFjS7BfiNrdkwZMwBzXdNh9SQ1fZ8xJKDiXSoABG3HQZItAs
yPYjYhZAS84nmxHZA9PkmFHeQttLlFnMLdLg9q2928ndGTRv7l8itCmlTqsDubG8
ZMxNO8luGyzq5KUQUF5jR2ykyzcAeim8aUowBy7rNpVMXhEdpDpgbMG+X2Ca+Fla
VfL0bQip9hvvXawjTwAbYrc9NhunHcucvJeu0/vzadXy0fk43c7f/HT75aoXYz9n
8awSAQZuu4jssM4RJFMssx87swfM2tA/KQZ9T+D3I9nuIe1+gMVplbx0s5lKUZF2
YXm8dXwB050hjyPh719lzDnboXPTcod1+qv+FKX3SB4j7aodeeaEVudvvsHU59z8
lDllQ8a50KWaIhe+HZX4VlWlA3wxmqY1o44OgZk+2f11r5gY1whysf8axYUPmzA6
4efZUBFIeZWjK9FZlvsQ+QoeEUfgIXNRSOkkD7cL4xmhsVZ2jMf11nvNlv2Cr9Zu
Ba1pTVOS5/JcTOnpB2b84/9PWjW+6OeaioEjIJTqmPrfw5jHaq67YL0qXVCvQrWU
TtvK9xsVzEjJr6X8s4u+nk2VWu+cR/IVheQxrb6lpDfhcQHbOSfwWJPUihhAyTZ6
sx3/dF+XMLX2Nyg6jFQ67qoBTypaoXMEWI3xziL9nHbgJVElq668TdB9jCMYA0uP
vq3NnuIBjkO+3WcKek4v8o02qCrcyCSMtAGyp1PT59cvKYKTFJ5XDPbR7XvqQ5pA
iy5nfm0aq4oQ2bdgalYeLVrOj4exywCHTa8V8acMq69wY/XCRHkpykmGSvqRIv6/
+oLrO0mkGrmBEyqyKTE6Pv7t6zLuMB9HIiLObeqTNs52SqzgODgkgIcLmjUX3QfI
WK6azvUYY0E8W4fzF0XNroy07Z7Y5QWRk4sKa9jcqjKgsJJc+OHiwUeugEhaPNAi
TLzDNtn4vVsJQo5TxUDO6hzi4J9K6SU7y8W5pysdraT23kyZg6FaPKtnk/dnFZcN
qwCEGfmCZ+qkezc/cYUsav2oRwDWgem+mB94PvHnWeddgoIEo8uN93Bg7KDe+i70
8ZYOFVgdydkeps1B5D/ipQp4TiTKVTgDyTBV0bejUFp3k2Ko8Eg5wNSn0lJizd6Q
L4xp9omthvZqkaKqZomDF5v6AYauUk5NTZcA9cgo4avgyKfQUs2rYp1WzCZLmoTV
cS3tf4vsjcmSy6LC2THviHaisc0qGZzHcvK8+SQTvUDENba/ER33UpHwvxvj3WcN
SwXj/V5HO0AbaSRB5G9hTqmLdeBuna57uOPll0aAsWfIntCtx5nQGXuvS26DrJwb
xlV/8SjFZlx8w/ZGvA2b4STXUkwVrqhIxpca2G3i4yf2Z2mi9udnrnW42yLgqsKu
55Dz8QpPjzwYkPlTG8p9gbfd5G/9NNHjKtudIBmDNpDDB9hNywRzP1HZLsi9zI1b
VvEAPb/kwlaYlr+M5ctKWJSwsvpjRNjIwZtLdP/8bdbT7XMHXgbj3nK9I2SE3F08
43sDziIQpG/BHZHufWlcvFfk2a2QTN6R7ETt6kBW7UK20JbdV0EcC3f/Mi+gp98m
PMtP8W/Mr3X0RKf9BXvEntdnqdAyl9IDs2C0J+oqmdFILmWrQnrw8QhRzyH6Dqy9
cE38NKBathRqth0OUOUv168X3VkFSqYqKEcN0PpEk/3R+kvvVBuMbOGFLrprzWd5
kEwvDzx5Jqu6Csj3pFMqzxj6976sho9dOmUCcUUQnTWQqBMKoCZHDs8IZae1nI4J
WXvp93mjIrgLBkCTQJg5077eEzh9jKu6IZb9kCENDR2j3EFROpLawGgnXyEXgutV
zvZi5xY0udpXZcBHg58KIcGWGicqC7Rt/eCpW9m9RbfATBONH0d3c/A7QYlIaccK
jMO1oHVJh0Huwrh4XM/XF9/KTmAFmONA/P3M4Downq94e2aIm2yT7ftJRGKpvPIr
3dV21my+NZnQArqgW56g6KNNTfbSd8U9eOwHihOalnO6+yWI8/8CZDaV3Ny4WZ0Z
NBJRRl4wPlOr/K8XKghrRMccYKui4s/HEsOKZA7mA6bJxe6r+0RjZ+gc5cCo6xgP
JfQDaM7uX3fFLAkofHe7krae1Q2iuAD1dJrBVRhhvNxTz5pOhw+ZZTmSge5Ut7kD
/nvAqgRk2V/PYTV/FiIDwjH066ZXLmlxZgZVG6TqLBEe3aMIPEQcWJ6/Z9VDOCXJ
9IAUlpalbei4XyiK+w8RrzTvFzcv0PGD92HvIZfjHiwlosT4iRNAvKy4iJUIE7eu
KFM2Uxaivwwp+AJMGpdcYbtJ7WuRivEQ8ml4rWvm3d0hqGx6OsCXjA+4KobrWt76
tAlcySpq2SDOjN9We2kfmNiHnpo04Bow9nsSQZar0E+f8/6vps4xWVaM8YbfpPcG
/Sh008ug1h44Ejl3yjMSSK60O4g38jZmY9wiVDqN0ccaVvnlyAXbEuRMKhZfmUsm
YELkqL1NfHfIRI6aM7cuG+78rE102XUVi03b7zDnxcbN/U3oJAZ3V+E8WooUrfgb
wX0FhvbxFXCftPztxItIh2QNW//qJ6DD/0PDSzU/A0u2THQWyCMcXphOIJkEdi7z
HXUC3WaMsa2JCZOdDzxf//6Uwc07ULNytBn/tJoViu1mt61XhNY90jajfTTcLDYX
7K6V+5SXkoHUial2Pui5k2Cole+PnYpIHS9u/ZbqRwuG0I0UdHnfcJUliHw4dVa6
dWG7ewP8HBDpOCSdJdrEV9LZ67NYjeszyWX4McGO32YExVYG4QUZC8UsGPPaAUR4
Y6S8AbAQZqBbjMj5UmdHnXau1ZgK9+M4jN83D8D2qFpomicr0gKCGM/SUKr9U6Q3
zRNYKXpTOOd3eknITaDkzMifmHt9+HDQNtQsZalasLjTSOcoGOkRCvaGRBzKDHqy
5zHyaIVxi0B8SXfZt+S/9vLc4E2XbsYZaglr+jSHWr0TA9p+mCS+UE8bk20zJkG1
nTVWZ3uYJzzJk5qeyz43LgEZUN6iDQLDDSn0Hjh4w0683r5isYp/t6mjDg1Hhn4a
DZbrcSH6E5loekpSZCW8RB7PxsvlyhXS2rf3NrSu/pQ1c5TnUVdWVIXTvdwi3OWY
9++MHYFyJh9FZWkgGR3nEaiVwM1xydsL3ml7sAlu7kIK/7C6vvJKp6vm4EHZjC1o
kg+U1EzzCMcK+h9GDTfntMnjmwDp641BGSWdNy10rMqREISnlWIPrnGS5V9oUuQq
sOcH2tqw0AcEyFIhd/7oZSxlsXg+cWg+c5DsD0+SIVYayDhzrEMxByyH5iiwGpzu
en50OtmO49qF0K0XjGLhqAXmlhvk7uuxSDlau/wWEIobT0xerIyUicPOom1PrRUz
mgLnqHbLoM5bUWGIP7/XaGiQeOM+CiMgpXbuh+GL//wr/0bjYzgRi/TsxGm+LFdC
Trp5LW8GiN9GZf4F6hPYDY+/mJm/7JY6H9eO4KDPNQijoskki4RRy1Bxy7cvibbo
ilGi8gbZrR4TjVUKmpJhllQczVTz2RR+G6CmL1JCsoS3BzJ33cl6GwSzXbFEjeXT
+/fN5+EWQ9VvtxUFJ9Yq5yMcGT9Ac533oiPCBTVJxQRLf6TtJ+HiOx6mYu5zGEZB
M24NLDxATlbKMubla6xkLWr2lc9OpCPdUC+Sfa+fCC6Gyz4sN76zoW6jbPYJQtqm
K3w5ZbC+lUnQoxdKI6icaZT0W+tzCkOKMvpM9DIFO6tCW6BYnwOuS8+qyB5jrvPI
jUUUF8qi/qKePrNtnm3almr/6X7wgAuWBUbmEZlLRIYTzdLtuAFVlZYIdz3rBbWB
lDrmHLwFYBmHjstD49rva8q+gAot8PKvRUAWWaGeJtvXC+7oBfDqiMjsncb7GlxC
iz1U+JauUz2Q8xF/dQOmEitPmGAliSdIfLgk3YmdMkE981xwm27g6n0SoFXhxGeG
i2zs0HhrKmuZmlp9F7h6qX4aWHXEoqt659y/v9ARzhYp01PZipZYzIfJzvGThIRy
V0kfAuoSk5ZYH5EGIm6MjT52/OctVCj3GGIj5zvUP2ATaPhxwOheFphNGgHEvPa1
va2hLdI9t6UxmOP2eLkco8sXSdNiYk8kTCb/bLoRnem/wkcok09SfoJyMoiXbv+J
SHTKFjhcC/Y+1mA5DJzFYrO+n15PeRtsc7i/fJUnb9KRPTkxOjP+4VzPe9geeFMr
KyH2nrNWBabTHkxZl0DH+3GNlGd2FmuqnoQMtEkdo8XK9RCxgQj0qJNauLVjZQlq
d1ZgU707Bc3Um40BYmF96BehQSrNBjML/BB2ZcsIffWKxU8nJ6PcwiiVFAkRwKNn
SAaDCwa0iYQuXwDhVAtR08I/BcV5TKxIYTmjjQ+cJQSwJSCYo69a8syFJKUIxpzU
8WoNFvnACp5YCLeWH7gcsRg37NOmLHiSHHetvmBRVw/KBH/otHsbaCTbFfDOh2VI
1Ap32Bb9wvXjBxjd0x86VpKJlYwBcnNVM8hfLRH1eLnA+p8Uw2F3A4oaeJyq24B6
MNQBh3xuLPWwx62ZX2sInOCeQLn66hH60wjSB95o82BnS8QMd2orm9HkyeukGD0J
kFR6Roej1XwyXghDAwR5KtxPlCgmjwOmDVI2xl20K4/uOfaDxB8iHRJ7QjlTS2Ds
ymgGpgylwIY/3visKHW2Zd+L703O+hVq2NgtIG1I3pWHDRRUt+9mFnuwk5UlTe1v
2cCnpyiSxQcp8DE8giAJNTNGIGawmAJl/Izf2rEFvwTnE12fa5KuK0HB0tkA//3L
Uus/R5HuGC7YULVasJYtClgNedsK7JTq7EA4XRuZxD50JHWLH7O663O3kVz8uchN
/OXXRml7LkWdaLBqj8UJxIYNQvXbeBGB0VQtjQkvGeGkSeAkiwiI2MFqzs9UTwjZ
MTTxnm0ppHdhRxzOmTKOEOd6TGSG6kEnW65oerCwjLIT5NlJleFtdgbW+BcxRLVx
koDlCOrnPNteBcOUdDSNfvkgk1W4VzXyPP+Sc3HEYwwatU76JIiZ1lOzOwnU2gwQ
Te7KugleDI8qgD/QT18bc60CVNh6yotau/VJOdhkxuqeCCLb6BSi6RxNceA9KDzA
N6VUXoVoTqct0i0+Hn6FaTO/tE16Ej98b3FM4lpiNfybVTz7mQX0SxfSJQo69VqZ
yLE8DGKI0rnRurxm0ipAtA8dHcpVj9Ek1zkBzZaRY7MULFoxkuEVJvCu1mOlzAzj
VJ7FYmhmRATv+NLmUs+RE6y6ibUI44ZRCM8M9wWhhVFaUF8KE4MnKrbfocdJ61Zm
CMf5GTLnejunDnPqs55W6rWm8CqiVUgYEwiOsfU7M73JAXAL9Ic4PCIee1WmvdPo
MaObe5MEun0ATbfEW+mi+V7n0YcIpw8/gkWFA+Ot1lbWAIKMyBfCZ07dqa3Z+V+8
u8zR8g19671Id8z33Nk4BPOrTew16VH6i0+ILqcGCSxEcVn2fnHPqFfgIhA7KvXH
fr778wHlXuWfUBucfvygA2KpXWyanLTuYjB47croYa+sOALi8B1sGy4AYzFQYBO7
9Oi9AhRQueA4mb7wtcOKDcDkXSlKDzmoIYBviRACvAMC58IRanafBAVvJE0LXhSC
PqMSTGf6hVY0CdQFU2A/bZOD+1PlX5c0ekPaNOK3tMOLlOA0ljOPhzvsIrGG3b42
v6anuD+GRtZlP9CZ1R0qPFdesZhVtoakRWGCkRNyv0no9chGfBm0EF8PsA3641Cx
T5Mdl5Mbkvpu9JCrGS6mKgcVsonuMHbmS59pPiMeQYjCqOm9CUc086Tv00g7u12n
oYWfdS62UZqSRkP3g/bufNJtdHJHGCOqwYHoXe1+oulpSk9bU+ghgemS8QD0OTLE
mo95ekrYNpozEqzP1N11qf6OvxOeDMtR5GdLPBRYnCi7hTzOdgbkmIl0QuK366S5
ubSRA2ZENh6XikCcHM2hZjJYk6KJhtqXp+u0dBlMz9soP+ZyUEzmBcV2m2tkd2UI
TYTvb6gkyFy0wQ2E04Mraj14OPX/zxqKr7nWmWKUwAv9DDmfRhGc1rjOHR8us5LI
ODa/HXYshrtpwD9EZt2NwpbgTnyo39/kRP1BXfS+UoLzlS7v8bCwwxRvz6x90cXI
d2k1kqYtZgwYUwgpn2TelSUfc30gTZWMcWyjfs24jcQxK/8MRJhkng0IrhMSE4Ij
wPNhJRTtDPSEvazlumeUP83KQJj/wwUDmS9PNjDFPHf8OMQk0bL5YiW9OQtcvOn2
cQWEzs5f2mqgPZDFHqVr38wusj6ZLa5M6s+Em+AUWQYMriADfPz1NglLdRyuBo9h
tK0zbyKExNnChFstoyvM96iB96nqfa9lU9fekW0yCZ4FT3QL2f2Lw6ywZIxQxnfy
tpk4nYq1esc1GIy5pO1ZU8xv6PjQ2be+f1PO/MOyc5jA62oqhXkNm8zVZALsTWFx
LVyDOoqEvek9TJ5zOtZpSkIfQCvTofjVu2djkUOC4TFfkdUjLUi1bilzdEyjzPxd
MSujMaVky2pN7/pBg15z1m8SvRWioF0lkBzR5R2SZ3oq7C9ccMVLYMfCv8uLCZ48
ZA7Cm9QF7HBiSSUjGeeo6TDp8nHqq8ig+Wf8bdMdOzfUWySfJfsP1q/0cnlVqAL7
oNH0tZ1rdPCyAn4XuKxu/mDFQ0tJsF5VOM/iR6G48a0hB8av7hH0/5Y8QQfL9BHA
JVIh/MbHG52/mAKj4uhoisSn5z/yDbrIHWCUdQCLBFe1x888YbWdpzexiP3U0R0e
0NmE5CQ/kO3kfyKMNaBDXNafg20BmsjGI7tjuWS3e+XKvxC3NCijPt+T4LCte0WD
sQM2+RIxrD90I+CgZE+kHDX9llWCQA4/AjaFnEW1vyDwNXTDkWTXvPZ7z16R2gLd
254T+FPaMgaL4A5lEQq+bOUdqbR+kkNGLTmZXk8XXS3klv8ALBrY07z5ngfrvcjB
rMrGpmz+wZTlnWSYsj15FebCQ7upuHPvCyjZqL4Jl+3lWvojIC8gfVwZySp2RKfe
tRZ4Y3XgcZwaq+5fg1oFTRjJOG9uoxwRVlRdTcSJykrmSQLwH/JyfSR8Q5VbHKTi
nMCfmK/Y0rs1YiqVkuA3LzwKOewS36tzNUqkB2OaxfqSw3XLa/WzWWermD+xQJKP
UGNox0kgsKgfyGb0SX9L8vzQoagCzmaHMUtQ9v/cn7ytoh32HS9fZkmYIWwt4ZNV
AmUA2vC8FITHv3dp8i+A6NsTqo1s0ySFhl4L6v15NyMsLUVKn1WABnBxMgURFZpR
ckoZYx2Cn24I01sYCXO6Wz+UnRIfF9PxwSQCuK3GeAqJ5ZCV85HFLhZzoTVZB3sH
XjmxjExvRpvsQ09lfUrgF4aslP2X8dc9S/OLlD9hTnzEKfsrrV8zu51Vnc0Qpg/U
1D6kvQq0uyuKGYVyXlBsjUk5aUTDR86yQkKRV2oLUsbGg8q6+xxcHOnekxJnjEzV
WUJ6/GoRY9F/9ikUrwgLUktqBwCnzCYVe8s6eSqsNBLNTVnprUYrKmEjMWg8cIuO
iHLwgEp2JW6H2/XDM1OyjOtaTvjdRGv3qdag7vfbQ7leUGnCtFDverhCmJ9pBBhH
HTr7g0Tn7R7daUMwROmJp9Drqy5FH5ynTYp/WBCCi0b7/pojHD9MnUU9glRgnii0
BLuWCZR6swlalTm5vEaMX0mN9H+b7F/w3pX/Jk4qS7STTkCvAJ2TbcNPa97Jtl/+
2v7vfa/RKzfjB24xEEa5mW4YZluqUaiTEE/aDkT4SqXbl6tH5tvzVOI9ZhYL+50m
g+oQ6aPo49UmMbVd8sSddj5efm0vme4X3BZy1uuUxT+qrZMlvnsDMjjf7FV43SV9
soa6HbD/egYuqYwMWNz8wBQY0i7oGkK0lOyj1lOar87sNatwC28otEOLyFMchPN3
zpFlOterK2b/90nJHsfmPeN1VEEYoIxOzgxI0/MBS3niqswontjKJWSxhC3nPkW0
m2Wt23rOppAbZJKmSAzyARCScc2x9KqPzqkk8184mV0JhxQxAUP24hXZeq0qChmV
tzs8NK8RDkcAf5EQLhnsyWaRn6v3wUrQRXeT4Z7xFnEPqEFqcZ63c5CgPD1cVcik
BwKXsjf2Dtf32isJKmz5HsPZLCld/fgV4C1ZXXmLXXib3lpRNMbVzxxtli9dLPhb
Um08ubLPFYofqbiDo8rL/Teb+BfDbIgc6UqPMvFP5ym30RXO7QPy9xG8ViQ5HcNr
uHW+uZa4dRrW4UBL8FoVI4JJDq97J2cnRyVspGH1Q++ZQw4vMhipRcstYOHbcA91
HknGii5i/uTrFqo3fXnrvAAxUyTiOqH8tQcw3ZpwVQh3LeHY7hjzsOZQ7oxNA04I
UZiECDG4AMMYQeMfH88ROOdJDDs0cHfBJtbXUClKkWQASI7YDpxqKy+eMK/iikJf
Q+X4wRhfcMj+e+dPBMXuWtwdPQcDV+Gg1nDicPu4RuxYVfUabVmIGQaUkMvhrE0F
Isf+FXq4/921n1oM++irp77/JNYSI6mqhDF8VYwlD39Bdq5PVSL+wwx6Jm81PHhu
5D+RwfSaANrUS/ksE+Y6kvJ7ONGNtDJN2jabqS5op33PcJ7UaMzU1Z8yHyT+13Y4
wKHkaB5n5u5T6+zY7y57XfCPUo4s8srhT8XIIcKxPXcvx9SSNJfD+NZPPPOd3abH
/lL0n0zi29i/1LbruVjxGiOcfSaeMFl8WRCwppCvmPfB5XI4tvhzZFSs/9hhBULk
Wm1r6rCYsJwle9vKf9zFpe9wV+hVNVb2AKwM8iks3XmVsfeGcH/k4xhtylpk1i6J
CI5bRPF0t5zwyvyeUhYIHUuwk8LkfgoTABWsvGfVmYAJzl9zW2psru4nIsMCqtvY
xE1k29vH1sNKPIDavxYFHBnJwuShwdHI+O5AfNKtoZa9NEqy4lvSrbN5ixa+y+dY
LA45+mf4P7sgVZvWD2unWRIJvdORpg4ohBNqIQ4z+slsLWajX3p4cmAoMuKSfdio
D2aB4gVFChbjFBACjcryXMQV9+WFAYLvF/XrSneswOR8YUL7jD6hmB8ch7wYBwZf
Oloco/AsIB5z5P64ot84XIQR4upJGa+XfqhJx3WjqxreXuAK8YJv8xVoGcD3MiWR
17eGHPcCJ56i8nOxxcIpzFGFtc8Yq8GUHYClmZPd3JWpIFG7if1Y+dLL1i2nZEYy
c8HzxP0IRde6duEGhS4Vct44XU2NSN5lqtx15utwUhT15707OW2q2m0mtRN4bufn
QHPhNS53vbSc2tbwJTC5dgTsEQWOiLTxo19FFQOTLxYWmtAqXXPRny6Zx6AK75YQ
ANdqA8yJAh6ezf/6qOfs+NE/n17MToHshD2HJ32z2o/IIG/4iCgop+y/oAyb5abY
i5OvekZZtWB2TjjCC8yAJVKqkXQb67Z44P3X14wpFX4vuiOgzEBZfIfxgpj8+RF0
q/3oLut2IX1rfGGI1oWnTirEY+2fvSv45GJ51Luj8tjnEGnShCvuhm67mpgvjIxC
cB0C9DXvpoIJ1zfWld0Quo3zwrEvFSalfYayOHvB4gxydsr5GClr832BAfIbQVD5
dPOKiMXS1Sm+Bg/svWNW7ZT9W2fcEdq5Su3Yd22zJ0SgxmaphboV5671meZehlly
MxAnyGVoAj57cXTV7JQsw6eXTHn8FJecY8m1/FyLXvL7CxTMordo4C8u2Q2Q4Hwo
Qbz2EGtuewqZQcNWkybGFSf7owIMFeoebnZZUGlVN5IGI1aQKgX7YTXn9bM5va1p
9S8ChZdR2WJZr105JljoInwQLXxNyIHz3Cz+U1QZRgqm1ys6RarjlJFl7SOSkQ2K
DP6sqXuHFEgzRtqc/J2hHeClHyqEJ14uSi6f1RLP0pIZIbtN8rhhaFyqwo0IxrR1
UxFP9/7U1GVRpjqvoRFVVRCLh48eyUFP40jnx5th2pmDqfckxskl4nWuAT60xDY4
0Y2lDu5rup3Yc5nSQjiT11yIyYM2cm/7kEAnam0DhrqWXo3vEzEAVNHxLSRhKRwx
fv5ckpAwdnz78Bvql0ieJqJj26QknwU8SinXhCixuQ9baVGPsGquqEAicmRZAca4
dNthnaIisM/J0wKUljCjGfv1UHZrxC4fz2wE5yxq5kcuBcHsdI6UjHIPhbMS9MCJ
OG3XNLgEi525CxD8Q1aJloQl2zPsHJG59DUfNQrHlXLfRcyGvmhcYVYKekkkNwsH
GssZOZ1DPvTIWINTnQcafnI28XHxXbFFvuruYdIt/t9eNNACp7NfnrgveNNdgXKD
Ru1awi4lUZUplDgOiJn0s1nIuqm2Wg91bE36GJOqr1KEAvyZtswuSwVu9XBIlWJf
DNz/6DXE9rJdl7g/9AFE54pIbENf4jutXdu7B2hgWM0VjvEsKLF45Fft+7U3G5qe
R/ArGPhy8QDtZfv4LI7ZtgqXmzwqF3zP7lph9e6hZBDnorcGGBQBzVZg/06E+sfE
tl+ZjFycfKCUJsN7va5r6mweDOKUAt/o795A3VL8ZzXAdiHoSDsjsh0vrkeDCIOc
DKTRCEmqqM/EjGY2h8kANJCXxcDaJKsWMldpvjnTqG2iRHehEJc1EEnFcHYZRi7U
EP+p5yCfynMyefcDTZvPztJb8M/Xjlz68Bpir+REcGgzhOt0gGZqId4TmHYnWZkV
a5isRYGqoshYVYOs6A0xzrudoun+qognLQIwoDTiXUpNymUhKGZ4+9lNkOyvUT/C
osq4rGujeh5YUuQ9WzKPWmW+EqQebkWCHYh8fDJpSHNjwuXzKeZF1rFpHtS91FCB
zpXRWbnz6RwBhgKSAUsn1+wUclFh9CvCdflpLoDp7I0TP90BTWgOaqHxQP3X7uOO
dWGLgyieJM69qiwRwgxJVEaZ/HMB6ANWTsxDbLssAgX6hvS7bLHsp6ylfLv63gy+
s3xRfStPaXpHuvpOwN0CNLWYlaWAvLid5jQZjTazlpy4GmKEtfOdeVUEfZycrgev
T2kSlRp0JeamPE0HTbN5+Xskzk8HItcy4CVAx2Dm7/XeUiuKgFx0akd1q+EOhmtJ
0ReG5iLB/yHIcRoyVUBWCVN4Vlc8AVta9uXfbfYF9Jio8PWNBTacdl69qmpXuZ5f
bfHfkpoWyTlk+Tnx6pYznSCHwsDF1Q8+2LyiMDHn6C2efZekybmhlaluuGty2dZ5
DEtSdbB1bwgrADYVc4DRieTifJEdGapqDNuoWtJSs79jDC8qSgNcxvobhxodlQps
j9CZ04FAI5f49FxV1cm85u5ktplpfB0d0noMxkcimJc7TlW974E927s56uKaIo06
bmnQYRD2VteSLI2vQG7sBLLe7Ps81hpU4nvn66bKJTvJz0GVQAbiPbAZhXsr0gY2
rFi7TtaDuQThs7iIC45Ke1hnpJi/RKZKqdYbYHjWxhuLdnax4UooPTSjzv8Hz30z
/D97BK0iLFt5f3Y8AglS5uVBabci0HoWqNZjvJYk8D4SzsA4+140Uuw+Z33daPgD
LCswd+d3zLiPZZWbk4KEuFlBrgqA0QsMsSFrg0GwY8+xZbOdVkwYnCYWUpUaanUr
VTKs6rCNtznKIwQNT9m/FbLlH8YXQUeMeVJN+sr6QeJukUf+UdDGFrC+/WQYerd3
iNzOv8wq7OZexoji4JyUYVJ9DUDHpeUmkfIrJ8HOhsMOoF73+q+a2j6xqwha9Hmn
8281HgT8+UxS4w+NsDrwWesZzII29KoRtN/xKgfhvIQkhkBSK2L7iq/qZpFjIWUI
AVe6YOPACsRMcU3YRAzhnd19xbqz/eG7xcskfyz6xJ8H7MwJoWy36AUaoKTKeho3
ov1tCT5zB13fNgXVv+Q7g5XjBrCSR8w7TOInGRJ8KEyyuPHe+RRMzpkwWiTn3EfB
e8qKyE2O+MggytX80tikTTUSpTOdq2ohkZEF8/SwB3p5eptpIEoHc07D7yV8u5DU
Wg0c6HT71N2i7LXBD3yQ4vMPlzbMujSGewPTJ/p3p3aaulBjALS1U8z2WHnLcCCl
istFDltpNAXIoMcHlIVnndxE9b+KKQJUuYmCRZFKxyA0EQJtks6R5WKGGqemnrur
gwapQthVvNLcWR/KJgGIPiRGYEJkadatObZTJuMQgdmAsHkDIKHnQiQg1btAEzYY
gsPQ2lBSunaePkLHoluU7mdNXC6jUwT0Wx1fXFmiGrA3rg3s9TrkbXY83M7PGUYv
ev6MpLitRmD3M0mWeiNRQihTPnthjPW9JRfTgUHfmGkTd3GnNDommGY8X8sNZZw9
uLUlk2ERWuwO1ZtvAu4yEKiYCpEeDPZaRx51MQW2H+nwdYHsz0T2K5LQDlbJwxll
cNKqEH7C840ST5Rj8PsKlXu53QRH2p3OSyi+NO4tLs1mi74dEeY1XAlfwMzERntY
U3dbKwJOPE/nVzqx4E+Rtt7qoVkWMR7UZQOmnzejGBwT3FfqQM1nQVZCTE3YJKdH
9HvHOo1ZNWCd2q10fxGgTZ+hZDSodCxmbcwLBrpQMSixtmBBecIA8m9bnrylmsaE
H95wCLl3S5g2W2w9U5V8McFzffpg5hzjYwkBiViSHC0hAizIeKM6oiXffbbXaMeK
srYvzGSf6402JDEvrmhiGrFl2nn1Qc92Z7418Dti2f15iNXYk/dogOLkvIWZotjB
n/p5aZchSgGzSn4dqpwoghldys0DB9EtnUJj9oQqZUml++ajOJWNaMKpq2VEajTl
Ka6yErVs1DZw5Hw9CKQorw3T45XqSEQmdP+u+d+1u+cwaazuZwkYxNl4Vxq1cTcS
XTEGIf6KM58k+aIJWOwW3i6jy47RrJlXZkKzPYTXxp0RjMqoPbNZB41x13jl6kwC
2jC6D4pPI5NXqIfN2cZCS/cQF40Ok6Q1XKBHuDQ73P2g8qdDn5SW7LkeZK6IeYpu
P0g2YEz7sBoVROjzWXIdQWxQsQ0mm20o0OUyeN/x9WUX+SStxWMooFzvrRmZi1K1
ZrDBKOVX53xxsgh6jHtiAHhYbai1av8gj1Oc2iTEsyY20Gdg/33i3O877u75JXCB
MBp8HT0bd5y44ZDQxt8OiXG5D2GitnD2zvnG3QJzjBtfjcynfrMh4Thnaarr/VQo
Hc725qluvK8XH3DKtB7peQ8pvy5OlnS0MjNHN0/sIgHzbo9MKItteqsMvxdlNfr/
KRSq5LsAEzkvqAHeSQwncYgptIJV4dh0o8rSj+3RxiRFnQQO1DVKvR2juOd+CzIo
2bEo9uBPFl/m3g9Y94t9Y9k55jpoZUFgS2BLcyzdxaohpqde17ZCXMAD8cDW0tdc
/Mja6HmMJqO/x31xNzXEqGNos6nFogQdK9I2KQIE+24HmOvtN3PlHbXPNUo9dYU0
hMje7CdrHveiR38o/BqOS/zXQArVFYq4KeGShnhNnGimLaBmdNz1eSeLuruoD7vz
AqxDyWM7rTkgDRjAJIvxsjLqroru87Id6a6dob7yrhOcJ46+VFmyoZLf07uqiJX5
k2ZviJamXyYxeVSvZGuGWmEkg4uBi+kDQe0V6pTOVPJf4Trn/XEe4FSeIYUnWfW+
5pBuVbzijvb7tFmQek/N6/Hk2MDD7stKD15Tp6i1PsLMpcQWPzstisNm1tQ4b8cf
EZxicWf3Mopxq7wL7vb7OpS0Gn7lZdL1/ISHW4y2r09TWKCTdlHhDljtser48Pfk
Ga9lS4zV+HPjSFHi1KCh+Y4Z8oJVRl978u40CCSxKVF32wci4Iu653c1GwWzywYR
34AUUqk7pfSnd19bIveDJ9KbouhkcGBLfwywQ1p/jk0FtFTzJimqhexOz1rJMg57
AgaPNaWqb1ysQllGnqcVF/lTdsTGk5NkPuXQelbqvIwYYkFwIVRmbEJ26O3FXLJe
w0n/oDD6VcFLVMfSYa4x7mxldENUMWXndheUGDn9ikBxFYGltrGsmgGizjEd4JPi
5VqiXdTprywnUeY5eWQ+JljKm8nbc7wdkRlxjVATfthpCvkMRdxLBCltvBX/0CYf
XkbAVoB1ljzXcy3iXVczP4z9OJ8iVIPCliyNgp7U3zBXfwpPkv6LjpQml9/VyjPv
L7Ios99XnSOX0iH5/tEZ6XRk9APO2J2gnD0gvBnV6CvGVkh2wt9hqFA+MywSF1lj
K9X3/2ACxPX8lwARmoc+ALix1hdo1rGoJqeudV14OGs7Hv8TDIlLtehFOEbMIPKw
Dvsydi4UbPOUhUFKE3YIatMO0E7862VeKBXqt5ppjuGyrVuLWlg1e/t+b7d6pTm3
cUwSM49H225Elp4sscgvNXNLcpl/+Ql5yxrX45Yn2vjwdBocfa/Kr0T/TOLPTWew
FfP1u+J1HL6BsfEb6lt268KiJoi1ENvHJr0e4gOENEfbUrE/UCyPTBGcHFGfrd2q
NrD32J9TSo31lHhvBxKXQaloWI+3oJgCwqROrJQ1joljvwo01ExtltWH+tEuFdgW
7CFue9KcadAvxks6cl9Qr49+WBeEeT+Brf7K3hTeDyyGUeJQZY7rxWTi228RyW4m
4CYPHjzd9CVGvivG7iMUlH0rbuldDtNNL6dpky8Ot/Y8JZKzjQ0XbcPGma8j+CcF
oEp1IuEmsiSnEZ+VlEMkj8r+1U90Z+iyiRYNc1xlDS6lzhgwxooUi/iU6aaZaYgm
TNv/yauY27XUm+/jPquyzzdTsnUZ0hA0puGlJqclmZ8ZOEyYqaqxnomB5MYms3mF
nbpXcAIchp4EMuqWSWZu3DEPS6EFuKAtTV5aU4hXxraDWVN3jn8UNv1JDnsh674k
obQVHLxhyfdnHkljPvOxwExwiO1sKWBw5Tb63UcMKxFtx/Ds+GW4mb6PoE4asJoK
szQMJuS/aH55U3LxukroH0/Hkw9g30FnqkpwtoXqD37aa60jk+KgAVpgA4BdYhAP
5TswZJHBE8F8irUn637hv9DtgY7G3CRoZiuxCOq134Mi3FejHNCzrpgTH9TMZBB5
Ok835SOPIm8NnDy1BC615uSO7NwowPRKah1fNXxrOZdUyovtDhqRi7KaF/NaoOMz
3uQoHAyHdWBJiBtnlZTtRvSnV3pW37vgwvXgyQcJnuEw47yAE3UwnR8AwtZzy5Qg
aUlBrOYGjN31YaJPA7o8u8HC9TwLj1klzxuPL9jz4TW2qZ0bGhtmp0nLugLN3wzJ
0Z50vl8utfXRREPa6Z+rRE5HJIu3cakhhhfzHCHesNcAKdhuXBFXKpQGTfxGtdl/
hbbfoN+BxUObyJiCgUmdQBKgNp841KX9Kc3ViPjEdheJycov1Y9wArPjzgzu/q1I
pIfJcDGaqnGLKkSbukYL9H/i23mN9QhREmbltswDEhILBnwnWABlBgpsnyKc3aQJ
tK4xkGH2hFJv6XUK2y3Zmbwv1yeIiFvj5Opctp0xEjysFqtvDUqVLfqmN6azsYDp
AVH8vFid4AMHLPM7UbfYB9g3zkIijumZfPWDoP/rvbmFqju/sdRnLxuO2P8VYcL1
jSGfsGRqJxrSsyphVpskyksKQvM2LycAPyBnM8feVsH3W1gaU5O/LE0iVS0cdTjD
usLpqJ3MZRafanb1BhDarOGATnqgAhiZ83rcEZZG10u+np20D4j8fyWQGzYEOAZZ
7VpGe1F65eYMbJP2Nf2bR/WjgRbBN2vibcY91xLwnXP3F8tApIy9rLEOsGsmTw4r
Pm225cyUfuF6OviEzemYZAihknOFRmwPOoCXvK7w2hUdewf/aJKx4SwAuxE+rcq1
wABKlrs2pwnlOOMctk+ztzLiDH1p+P3fzFUzPeFPdbsr0AUIQUliZYQ6ltr7corJ
Fjt704C09ycWv3IiZw/Gw2AZ/FA4rWeOlMk1YD/QLVCS8qPF/+UMGCj6RpqecJrY
yWMHAyUaIYwbBONoH/bZ2twrMINSaq2L55KKQ0gXhQc3nMpywFJ4LRfta4jd8oAd
WQTrR0ZsEt+GgQcvnR4qYAruaXnLip6Cw+DvIa8JIEr/SCgkWdRlmi3eeFoik319
NvTvIw9k3Ym4yl0ER23vMTmm/n8wuVyRzNz26yJCMxBWZgUZeeXQ4RUii8xNIUJt
I+T59hQlxqt1FZOVGxVruHElJtRTzuRfKa92QGiYp5G2G4vjIpxWkSKndVYVnyzU
9iDwma+qnXshU0wwo5jUMoYBymJpxliTjOU2vN6UCmN3eXt7x1MlKLFgL/5dldwU
3BSxHlKxtiu1mwbUEqC8o8b02NxzWGbVyd6LqVmh1r7QBhIm1htqb3ebs/2D18IA
elBZi7jIwszNK9XlkRoz7z3atCRFN8ho4oKInRCmWa5+7ytyNauJqUKpog3WtvO4
Z0mY1uOVBbqO6pY8DQZP3m25yg2L5v2veeo6lbcKUeVEMZdtY5ASXLP8as1cgNXj
lwwKkOJv3d/VU1u8CgSGLM4k192i78a10wCduj286ZF/jWoP/Kl2d+efvuRD1Qz2
clooK4JmSuk4HvrFqE3MkEZqAZdR/SBzaBHLS8yKd0pQCI548fMC30pMomSi05Y1
ivfl4gKOuraq6Jw3c/8YjT8STHFnl7g195OAljTQR6hAMB/DW506hL11R0xL/GZX
E7fSkskRt1cDqvfrpM2M+wKqw7OcK2HEgkZle53nNEvfbluFpUOiErVe/PtOytLc
KR83pzIjxS3Ao1fo2235NoV58phCy8TF2lGfq8HQdK5lgV1Dm7an3MRxwsUBw4RW
uBtMh2+8l90Kpx55uTTDPtmmGEb6+n1T/IQjuNHmL3v0zlP27ermYwuDjI23lmX/
Kuy3qbcn/eCO+uYS8F+r8YDJXHiVJYOYOHABRtNnX7iKkLb+dFcPK0wupdmtVcCU
QeB2Xp9h1ZGLErHRix1q7qeZFbP3buH2q4XEQ1VCsGdPU8k8B7df4EKjNnkM1IVR
yVXxGk0asWkzkAILi9S/7TvrnPhDlBTCmmGMEBdPM86SOrlU7W89+mC4/J5hfrUv
Wo6rVlDsYcocICBHLnwjOwyU211uvFBbCFN1c+zyFcw76rr5pW/d8X4D4TVTDG/7
tyZXAOy7kL+dFxvAEXNKIUssMQqcnsP2WBhNElxo3pTezEiJ4P3zUXJoYsVJxuR0
01fgy71l4ylRkIji5SJE63Dvo0xZVgz93oMhFZO5nL89ZVSDxmGZgeEJy+RYCNMB
/b5BslWPvxURMkVNnXScszXIel0ChZeEeJY8I5/nBfchgSf0EDl7iJLApNv3cD9Z
bmfPiEVoUaHCcb/0ZGrz1OIXIucpl9vM9dqPG33mHyHNwqb2iTwSQk0oI4HUaW1g
JCiELfrEfWt1JVFVqgHLNFZtHywRnBxI2FpLgnGc8HPtQDvjN6G3Cpxd2ARHG8g/
PaFUrW0y6NGH84BeePsWGd/xfltRb3lxnI3leLeJg78scEMXTRnR3obSkbiAFYqV
XlAwSJd+SZ3IZIQHTFhFoCxI5lxdB/6jTqtO/+1g25Tw7mepEYsO+Vd8Y9s03fAi
cEmcsTrJhsho6AG05abnWK6fJBkkTsQcSkK3HI7YdoWb621kTIuGPsgNG86nf/uV
HG3EfrQWmplGd3X/jlUdHczG4NDMk1eayKvKfqs7RcQGJq2MyWvHzalcp+rkFMU4
exw0fziJewNwodFm4NgcsQJMFp4QgHZfy/ObBLh8kVfDaP8q1WA2VkOAeMT+nKow
asx+E5M+0RwWMcJ5cPuszisJDCp94qe3SwagEL4EthqA3gQhlUACrqKMlUMYGFvK
b4qiNhMWFFZ3tRFvmMM92bIrxjJRgIFXaTT8/9DOc9NxJzXu03agLSnX3uVTHZuS
QUBjmqwPW5t/aj2Hd9mFHkaD2GMLQqGmiEfvBb9u60POrIxaEsHxeUfqsONyBgQU
rGlfUuCg/Lx1ST8Dg7DoezJBQvnAdMDpXz/Fj49mHfx81r2NVpl/mGu04q1sDVvw
mJiUbpDZmvqjgayAl39ExyArHbZdADgnOI6pF/ByRfzyF+VPT4hk/qcCnGYZ+7Bv
Xhk6VPbYwAWlf/811VkLhiwghUadDE2+KLgNt9giu4e4gADXY47hz+iomSKJVdT/
QE3Tl5Zcz2uZO8E00NTkR+6a+Tz/hDxeZ28bGJNPic7ENraBAnttdAX7QLaaxDyN
enl0I/PBHOL5WsWCUyNqsEJ2W+7jCQUjy5RV2qQ0TD4PGmKURpIYopdyknEkRuY/
NXzzVU+2oHB4apwtzkJwBHg8AqIfmrnk9H5w4sLCWIZOuk/TdCpGqW0DCksTEy05
bPUil3yLwmSE4+Zi4xiVdgmd/K5/7oORsNAAzj0tB45pw+XPaUpHszL8d+/Tz6qT
6WUIC5lTawbHeBEyYEJLNBN8hO6xmoPCA04AFzQ7XaG3o6vA+8eocOc7WjLPa4Tl
+qauWsyKar/O2ZJ5HkYJY8rywDQp6mPZSDCerLVdx4WgDw5+DalblEeUs7uz5znK
cGtRF4e3g8PChA3jMZrpw29iyNAiGpKAr5ZOWEIpit/EZ/Qg7WLepyX8AxyySgJq
VdfB38xZkBvTWtqTET2sL21gzZeh0kcIBO/cboH4p5rLj3f2dTa+/0ORlYkGuGSl
4Hoq4BnbvTgpcFdeI3uAuwhZZ5y1JnjGVTD77Bx3V5ewJRcZ39xvUvXoCionwLaQ
dUCi+LCs07+dzLDT55LBeRdcCtnIh6AKtMj+Ws5gtl8RKRrpyPN4rbb8CP7II6Mz
RSrpDQs5VtQvjXqvZxa1EFZMFpMlEjy7HLqmr3t553KgAvbGy4Hz9Lelf9jgFito
yWFVLjyxSG123hF3cbRGZ+Txr1DPAD+jZqovO7E2HMGf+7iuEDXbDkF88DgtT7xz
INLRk+/wQGg8wMtKufP+Cfj2mkEWNPqVxIq+Ihq7mUN6qj0CaHK8zcdcJYYK9X1b
AihJSffBanZyC5U53qAsXmKeGYQOES8sZC0hNVEAZ1TMD7eXfstNfBUjmEgak5It
16Gj0rV3usFnMz8TwrzQiNTnmKc4jpzBcwGT0+4Y+H02BSk89DAHiWH9atB6kSjE
Gyo+vwFzYHXQb+QUeTLtYftls+bclcJ117zByaTdZ1aRH3T5XgbOxTTQlLC9vbFN
8IpgvkZ0kN2WKFIGMhNI/3PgONlGtqYBg6+5NsAZCzfQDFyFQX61nBx6rWoZH1Kt
QSz5lKKq6nOuTy+IbAkMWvvZfFh2S4ODqzJHi63IhNnE1AnbolUtV8xOvIwOIvCS
kZQsE4NmJT6a7ji48APIgOvekQ3nKakfO+ALazJJA30fD7as8/hOqAN34ZQs/8E/
BgS3hWbzkpUt3DcGmjSHeLncnIxOS4PpZBd+dz+nNTC7lN5x+YdNyaDheuxpnvh3
yw+hikR0lz3vG/3dkWAmmZLZ4XxSciBhwNfx5+4449Iwa/M5aeOtUyPoDMO6G3MR
FFLp2iijTOEmtoCD+YY2/qpy6k0aXje4cTHi4jjW1wD1yfuDbkPy796S1T/RATA/
e7f/as52qLEO7bnCm9qFic8FpoUd9nWh4krgBvfAzOfz+1yrIiTvy8ZzVdNT1ten
pGkijCjuRJwlZ410GjBy6/51tGR49GOYb1YNzKNScylynl0ZgRWYkdPIuuYChdHb
+M61Y+sRBarQWPCbgoPlUTfgFtQLOUEVVoa5HCzoGQwO/ZvtXJjj+k6PXOxalmcy
PbDIFfPxCDIuobEyyBgXrTujZ6kMt90xYbWtQ88onKzomKEvuDgi0UF4fDfio5v0
axKI6YvlnMPU4dcrODCJU/6X2YCpOjNmYTPcfvfwQ4aYu1yVYonJTQQdoDyardBV
FaBFpBBrUFSQOKYDHO39l7ftvB54ZoHXXEsuYO357/BMWiDLoa85PYJr9AZpmtv9
hle7MHqwtYub2bAXTtlaLiYVngJ/6U9wABK4cM1FCcJApGRWh7cQ96UTUNSvy8x/
AyKWV5xSFCIE1TeppnHyTy5Dgt/qjHHJAxvkGrVr/ULvHyWkWV366pVwKjFljFir
b/fZA4oVXipIRw/lotEihfwGfi4IXTwOtmOoxV+9xlhwI74X4bQElgLDeWR5plry
PUy6MeOrnqT2rOkMHrUcEWx9j9dOCIG2C63dinK8j11QX/bFeY6CI+VnFjhCvpiQ
ath5wusSACdCgEt6r9iEfqO/1iQJbDQYa9xkcdcwJK0P3tsgcQOk6WhORyM3ox16
X+X1V1WrMemxKFc6ITNgNHq6r5qnvSIGQdw+r1TAY0pjTiYBUFHNfJR9wcUUlG5b
6kDW0DinUpTRc3Tc+Jwh+0tTA/EQRlC9oBw0TnQDGwmQl5ax7MoFUvHggnchah+H
PJzmZobWmbbuv2uKp+ir6xxssUaXPq0pcR6VOCLlM06acXeXDMmK334MYlWWS0Re
oLDx1DZ7Pcw/JyUNI+yxTwf2mtRUbY3FzKoP7kvGxHPx/5VAry/+XuEo6ouXk5T7
xQO2CQE1KE/Hz6B2qltILA5PY9iqlOX8H+7CFMG3HNJO9i7L0HIBS0Jgpbo7JSkt
/kzxVoyecpr8V8srJZKdch4xV/Sp7vKWCgtYcXB/Hkojw3TeJHmq+UZLFPmdM0+y
7KEAe0okBRkbNhtKw3TrOG3k56Adw+yxV3J8uaxlM7mt7OUEZaimxwg4CN3f2ZTv
mi7Pb8RDNsCITZGpndy0J7Rz5J8QQUFR+A1E9TYMcf/MTA5ZlBRKMVpv9nHYfn2q
dS2CGuYPFwkfZN1HrEhuPw3RVK4Ng88BmVdN2gQrLAmnvL6wfA3733xEYFsTfOaI
ERynUXe0GU8JX9kjqcvyi2tMO6bItfBG7cpz5LxcGzG+bKa0JQ120eFw0nr3nM1o
1CACl0BecuAyTOLpjYXt1VNehXFKMx0wvqaLktuT0SVrELJqbclpAZqDY/+l+rRx
C8iS3+oOcw8zYz0CVZFpWnAlz1r7H4zoJfsYXGIOkym4ISRARxjR7+8LggU3Boyd
u48s0BeV5+QnAPgcagnloW//UDWneNiQA35Qr0vAZWQ9UvpPzEIZt+n7yX9ugPhP
cF3TOXu8AYCkRvMLV24RaaDwg+3haYu1TkHcu4ADTaBczbUpQ1R/v1SsHTEBuDP4
xfC0MYfxzNMS1Bx0VWtoBlH3q2jZ/7nhcvsqxWuliHW1tsbA7i0pGbuac9qMsshs
pQEsv7E6PWvk/E++fZ5aYTP60CcoYs4Rr+MrPZM/YY7awPkwrhM7X8mg2UFCzSW6
bzPseLrRIzhuk/w1lDf6I9Ef/Sl5SD+MRs1LvuJUHoIgxTL02CWd+MdwAwoE9ov4
cB7Uo0xy3i4ChS4M5VtUVHo14zJxBX66BGn5Zr1axIMlErkV6kNrtcQuPdH0D7l5
D4m9tELWSfSaX2stLr74mf13+gRYnj2/iRwDW/mlA70OAffzkkFTkhaj6bPPcKk2
YoxXDSlLA+g7TEg4OYyLaFvgcqU1y/BBkd1Vd0EafE5BMz6HqjwHgka51szEA+Y3
55jm5MZ4E75igddYINjraW2f0CN70pOZPzDKiETkwGomoDYNrLlg13MaGf46DIUO
fxUQBD3Fm3WGC80iNEcWGB5vkJBy0unRFMseWKqsWYD+QwzJ8lpRR8HOjWoJHrXK
IkD9o7rQxosYY7b7IWjY0XPZVeY6gLdW07N80Skzdp3JC9R1QxP4+r8bhSna5zmV
c4Q17of7PwDPuEotK70v5REUpTmAus21G4MJaOgUCJ1mI6oYvZ8gzVgvoCyxr8ss
9lr5lsPVbqziEnOS6Y5yhttqChrGs2IJTjyWSingCsZfIlLMosWtYWKjXmO8TM+3
hnnWOLqdx0cjdD1wbi8HDyQgmiwIx8dwkn0GdDQCNOyMGJe8tUhx8ZV5IrpS86Yw
4Z8RtJxlVw3+5A2TEkHoUcFt4ye37kEvYM9wZzx/vmI8nGkZkblQeH4EhrWm4ChK
KmQGhH/vqBbV2L8GSXWh4tIPfWZ7IOsBS0DmuwgMsQIkZIyc9lZ8QCkyPGfVFiLD
kqOyOkAJYcsjR3gkUOvdvRtnr2nhGmaeJxEmOPWSNCVmxD2mrkPggwrbJE0v5O6O
+P1V0rOpmy7QTWZ9CgLVb3FJ3BIYq4zhU2KGRtABovPj8Yp36oOPTsVVieJ1BldX
Y06BnEjJr3dKB8En96iYzs/WPBROwsDDskUtQ/rsPR3JG/7ktvQACOfS0GeOYvlH
UfdPEeR8U2C2jFPFqa1Q07aXIyGMVLLq/FcDF7XlHYml6ve8EhngookuIlAXrITg
BUQERXBd9Fvza7nMhMKi6AWfdBBMsyH94KQ0Kdc1oiKxW4U9h22Qj+7AsWodW7Xf
F2aghNoIZYbZGGcbiol2SL05Mw63MCcZRF7AykTtci2aTnp8V5DH90ong7w/Sx84
R+EzNzqtvVxoU5FwcM/hsSwOsX+VphEw46OxoWK+497zN/SplimvTd7W5lAOK2/J
pmzXyGBSF+bN5sXK03hN5HQhLTFK5ALfHv7Lue8An/ARDYz+nUahiXf2mvVpYW+j
Q3UZAH/R2HifYZHAOM+shyBhduC+C/zoRfZXsPQ7Iuk2U/+00fpKEMFLFZNqQO6t
hxGZkENzwW6GB+fUur3AIYDeKECQaiUbKhCOVvovDSVf1bs/oqExL3vSSaaES8gX
iHW8Chu7Upq4F6esJzBFmX9/lRocmBliDd0GfD5fhFE3Z9saK6DgNwWHE3HRJtZW
RYtKQ00PjAUmKO77XIY7oBtGrMBSils8R1VkDEbGXh6oSwV7Dg8IDDPwU1lAgSSG
jOlsWkNBrmu4SgIBsEYuMJcZbEhKvA3G/W2H2knOrh7fPcN0f8DMlTm3GYVzymLZ
vmWdgL2CjU/4oY2vbNxLD0zInTEz7vACt8dlGC8A5rQLHxrsxa9kvNH8u/zBlf72
YrVmkXRQdSBOjcUj+RTbRLo2gpvadkxKuDz/RfS3nlPH+9pccCo9QIDKD6v9/A7k
Us6aohcUCsZ7aj5remSrLn46ohJ7pi7Qd3WAoidBmkVVJz/KGf7gDv3wQIeLF8Po
I6taU5NsWfrZDIBXDWWQqPVmqu3tg9zSFyUJiWMzjXsSAAeDNKsUOiHulw3J/4x7
SF46G51RGYRdPY9nYPQhlBvNgRXSfE1Ts12q25LJK6x/5I4MbUh5EjM2YfQEcXn+
nwGN6qqu0ehtEXguf/5bU9KckLbMyISjFlK+1F9O1Lv5ZDNFfDYx2FeZG2LN6pSZ
8T3IYFxqFO1APmcDt3P/k8mi4mVoEEtO6a+s2+e26c6KJcN7BqB/XbKA2njOaMK2
TcW1SaRdMoM8Vrr16CsoMov8BGSwqJLM/iWiGXNOj+ekBMKHtENIIq5kihg8ixOJ
6Hgc+r26r3+RodwBnscGoii3nnjVEYoG5x0oPyH+QkPyuXNOU3fXfkv1ki2uCxuh
g8gPu9wDbJkqpJAG2cbA1UgllbuVgtcmEZxbcyZBbL5tYqpx2jFrZoqN+D6bUv7d
ly1myP/ENvEVdnIhpcr5GK7WWo4f7dCcI5gyxysr2MtqgLrfuumHoWL2oat2Fe0t
MMn7CggaAM3zXcnNUeeMXSMRDd5uwZtqVj2Atd0EJ9FapzhF/YOLsqyLjpjTYJeA
+EUB6hrhNdNZ0O4G2MF/0Vmvi9IbBPXqPuT+jKOAIHkL9ivnFsJkDMPQlzj67KCK
apYPx/RfhhflKl9WIl05ADFSXS8CN/0oMS9enF3gY3TqQCsQzvWlQ+rfKEjJMznY
CtbLpbO2uUrEX3cCEpyLqB+Bs2ZmNZJT+9gHDxTpUQySrOXJ/m529s+cgt1Za77D
mdovwacjFRUDyOLAm6x7MUsr0GR/vHC/0fgFRvlFKUdizzpHQZSZNj2gTzLDGda+
LSP+hAdWefwf4Fu02KCPoM1KrsT6ugAJsfwKEcdOZoTEln/e6HyhmU1Sm0bNCycT
6SyHkKHcMdVJWE04YBI+WGBLig2vemXHsJyi0XTaCmbG2oykLzZQ6bQZyFEdeEyr
F6ISQ/YcEPDmRWySC7VhRh/CDYH9bUQzs5eASM9Iy8om/nbPaM/qRB6prBhPF1ey
Lz0n4QgKcnss8ZItP4OiqghQyVh+QgzES8tTBjyhl6FKKGabyuWyO1pFNjBWdybl
wq445t/s30dgktQNptqtFmJLoOl96GDFn/4znI2rs+Q9e26nSPefZsydn9vnR9Y8
dNYIQCBTLYCQdKBbvkmz3b9bQnY2OzC+8D3V7llrlpoWxxyGEs/c8rDR6zstBPbB
p3D3w8t8jwBsg0MEKyqnyE0lVHD567yMzYxcsNM0CG5V0QDG1sJzO2vANoyhb99g
R8xW3hilNX6M3D9/hvZigZ5YTSvnfCiJ5VCaGU5ze0bwTOPshGP8XNp2U1zq6Pnk
R1GD/YCm7szZfr6aXqp4enrAFa6uTB25Y8PoAlcN6/gSg3BONV2RX3H5eXJLl4KF
CfqvRZ8QdoECs72UeC5ynO4rE43ywj6vVPekxEjwfu5F7FAloCNcyGc0vYBD1pro
sBu1qEYDXPdH/76pjTrKno6idueDdUQJoudCh4ZiKC44W6pksEFuyfsIJXlCiYkr
G9WFr/bFJxQ4tOfqELs8UvFhaDxXLYmcq9e+iEqZcYh0DIFuMcj2huhND1gnaj6w
vLMEViKOqMkWJp2427pWh8SfcphO28fNTTjr5xwYOdYZY9Iv/rbcU9TUnbN/3vDA
eQ5jK1wvITkV81V9V7qT1oasjvcWvE7OqdcuVkQKgU/2hPECgIoKDIP7OhsfLOWw
UxbkUf/YdzH2TgwxjRwX3lFGajbOXf+bkcNArGza3vmlZOapLSkVdao6rdK0AYFL
maw2RVv0hmqCMXjCteY7IGX91HzuNiXNA8235o3wSxBiwrGt3iSLZd7v8U93ab6W
zBTLx8lY9F8Y2aKhx3SVkyUEmz2220KOR4GuzqIhP3Sb3RU2MqpLseqo67/wBvp/
ixFOUim9JDZlTY9litq4X2gVDppgYkdVFmy6d6FZj7KGOsyIPLuvQS4nMcAW8b7x
j16Ne50CGO3R/0HzMVJPgQuYmScKi571GW96M9iqj1i2ndYSJu4WR5LuzauZEFw3
rrrceSkp97+tGWb26xQwO7w/vnkGoKZrqURO3k36AoRy1vq57gMNPF3OtJrhLmcc
w8LESI8Ap1cIXLYt8MtrcKPYaX57mzVT2G/MsjMUQ9KzDYWyMIySTHbsIPfBEUDm
hE/MCKo6fX8NwbsP6tvIvMLVjIaLSB5UX10YrNGW3/khcnAlFBpajdLAbbbKWjUi
W95PWgZnn+C5VUUAdF79/CCGHchEk71DKK5aZ0WkgD6hwOXCwLqRYBCZiCfX2PxS
DegTsMUrD1GfgeQAVkgB6s4MvIPM43oqVu9IQzMakEGABtzLWBKr5dMVI9hu+tq1
ZkppX7AV78nJqUTkyIXj/jTDcX28nnVDMv5evwjHga7x4Ns1VN9aFfTEz8Cd9dFX
TjnfD1Ikl6w811lfqqWqrfgEOfypZ4ALmuHrECwyNje4EcugkFLb3HLsOOYbtd9V
D3JeZRUKenQiBivvcOfxuoRjvcIE8++ZffKKG3LhMsvE8qvnUhUs3y/zU6cL6NNt
6athSyGFdjCC2wTcloAvCm3cOHQXVhEOBqsE3EV3aFTwrrj+Tc4WQ70sfDcz8Eh3
rN4uyX8VeRKbngJ2DFFSjkBAuFrFYVS1rfhvCRpP4TG3iFT3LcdB59EoRfPOozv3
3lKWPTan1Kwh4l/vfY1t6azAla7aeqmNSZbazEKMTSHD/o6fxxRARgx0vxnoReQN
aCO6TueAxXnlU9aDUHOcmtoFT3usyGSdG/vSzY5fTsDro5QskCRQ2dIDMZBPWcmy
wXE3y8dU6nmdkX6XsTMU0t/0CSwsmEL2M15uyuFjOcQVwUjRVCq4RQ9TUdkqX3nG
hS/4ZalEzx4LhNber6t4/r/ect31X4fnADYS4xKYGjxdpn4B0Wt5wi9WnyTpqKwp
DfhxVFXLRLpjAvAkfgCIfO3OtRxuIyAJY2ep6UuVQ+BtRtCgRUV1HHEFU4nSQcQq
6TbBlbJ0lyCFLTjgwzprBWroHwIHorRMU8DdKq8wJQZ1ZnCCUSoqIeGGQQHGHMBs
LsbUJZ2JTOa4EGG2lIUth2EKs2Ae8+2qNG8X75y4E7CrLqQAPJl0nMUnizMj1JPF
HZ+96EZ07zVarIi7SnHt77ltWvu4k1B9PvXCcP4smLQxyoYOQGKyX3Sc1RZw6Nyr
RMjYF86nnOzSrnxk4ATsXhW3ka1GYmSl+oXPG2RqL2slQDHuxIsLmvo41Sey/gMi
ny6FKoOv+UYK7xPLp3SAl7w9skXs0DNzkxLT6IixD+vzqDelEErYiHhiUwP0y/jo
wSH7yTWzOASPpqUrPDqGvJWgirvXu5PMTsRMtYA1j6cWaFK5gUKQu+P27t70cEfF
UZuo5ALmSNGa3WeIyjUFFeduMYX6Bwz0B4TjKsugSR0jW1TlBAd423O1IkzUZtqp
WbED+CZqcdjCjlKcsgt+aD1dNqmtCXuRSDSIsHkQH/AkJUlA4P/fwCkuIzmbECEH
ewSRqTEco2AvPrnkeaLnKT59jvC7JILWGW+U0nv8uWAopTZfRrPY1QdHAtxgnEU/
SCEzhzCKpnxiQm5GhkJB1cZS/lBAAhQxFFUpVuWpnLD5eN3YYc2UoPBZRTpV+C6E
5ysg4n5+okKwWCM18eH/L4Wy2Pp8xr2O66VqzayCgLhPCUpFOfpZYuwKx8n9D6XS
/SI+M5nfycHwaSLPQoBFvo/hiIhyOiMKnv2xRiX1GYI27NKXqB5f9msB4e22QcU1
BvNWoenQPHCMAlXXaGRkKfi5SP5KfA/Yb+ifWbfsf5xYuEREd/0qZjeJTIwSzmEo
IMUMceXOpRvjAXNbdrkPY99tz0UmcCkxgebygai7X807nUgEkP4r5xCXu8z1tFj7
tMlPKhB/pBt6o5iVBfhCUDe3RDTe+Fh+bxapnIX/TL7KKKW7iDUpGcgkQnSvsMZj
tMAQk91+fo+1lsj3QwvOZsUA8vvRDtC3Kr6PhohKRaMKo1RVQNxeOr31XpThanug
R5UVBkK/TtMHoB0jvuBDLC+J3zbN+/rNuwqCJP0ZxvgY/5ZkqFPlnum9qzJuBoeH
SJEfRGHU548yUCRlPNmIEl2VxaCvMgPR159vmxMz1lxrvUEyFxSLUbzHIfUrIelv
9AoRHkYbPCaKt8hQuHwWNYfs7yckGamrX4doei6ieA/wqQ0/NyYKlN242TH3NNov
duHn+6iAzJivb0kpGgVgeLCZLwFfcgpR6atm++Dnw3KaW8zNyOvTMlK92xbc3WUP
2Fg4OmHr5Ab3aAv1Mw3q5YElU9Olr8EKT+WceaEAc2QKA5SElGgSJLtilmFipUWj
00einlhHZSXrj+qjMIPTaN70JLebafEyEaPeIiSg4D7lMaQZnbS0Xn/pqFJB4W95
5XPhDQv9BOriOsfOMX9/z7H0lsthzR7Z6tHhNwu5UCbSO3Wq1R5a/ds+reaSQPnu
fVcA/cJJ1tuusPkbzDVYl2RCkuxiqjeyK66B1TOpFbVM8ANEdPvaBwrdO+SKmiev
/HADICKjSxWscgacBt4b64BUhBRniWdx1nqgrgyqdNt7BOsVscyV4kcI4cUy0RDB
tsMiyhoZ2aD8S3ldGhAmAl8Inw1h6r1I2MX4TES/1FGp9GjcG/L7MRAqU4pOzX3v
K6oDRx6BTsW58bQ8tUYWCmm75xWBILLFM8esz+8NGJ8CceomiIlQRJGj6Oai1FPa
JUZ/rOK5oo8sq0Ss+DhYQqmQS1g9HCPwwW38DNd4nHF1I1sMradcXYLZ425oNhIs
gyalr+amzs2b0mlDu0ExSSdvkKBAUHluxW+hssWAF7WJ0V7u0NUuHMBwokw4nVIy
48DBkQZNu+ZKrV4iJAjjppDk8O0xe3tx8cUVmBFxKlzm+eLih81ZpskMfRIrxcQl
ql7yNR/DDJ4D9K77E+Ru9+ABttfH/oHLxXKjE5hj/Lwpiq4LsSBMWtWgaXEdB2iZ
xtbD778ivS/TvRV5m66/T3CDKaFZPJjbeZckUslnlFa7hX8bUhJ9YwIzu1pRPx2+
z3mkEs+KVUdb857qSkIQQp44fH7DiJJnMUsx5RCn3Jxwij83GTy3DM13mSTEG234
+DrZPmt/R0XslpwE2fB2PEFVf5lFB4fmNBAzVrG1+GY8gmD18nO+BOWIao8d5Ae5
dLDZ6eZuaUXKQiaPharLS03UyENEhflrnZOVzBJryEC4IuY7W/A+/JneJSBc1h9H
KI6GB1MhxbjgJo4PiZ2XdY46UakrFo/bqW/JGYaciFjI+qs5a4uGRJgLXF3lsaXZ
/5IQiDdLovRJ1i75O4tWAYThAGEUKmIhv9lnlldO8vQsj2/9q8XBhVTYjCd30uB6
V6RuGqQP7SW+shtXWqHhhjMAMVL3VdN7UDuTLZYlLFNQIB+BVJvHlLq44FPXC2Z3
OklTxG1IOc7Sk5WDIZ5LcLxd0lmnc2kc7jEow9jK0YSc8Dwuos/CJRsqNTFLNKW+
qCBnNtBS4kLjIAu+2L+SlxPagreH7eWDM4pi1ahD2rE/qPAVgw0Nphg/Mbeca5cU
02xmBWZV4OM1/HbUJtc1uQPt8Cy6jGcvUpPDHXb700LVoafyumW5UQvTNMhnION3
Knj4QN8/tZXlsmtMlMfsOUc/25+OUguVIww3AMHNZtsVC6eNfTEKVZvWyvnzQ5Oy
CeyFwBblE1NcZip4WMiEE8v8vMWBgKSmA1IDyP8koAC2wdMc4BnpC3qjUlUAdLyF
Rq6QgpUMdCT8EW6R+pzVJVAizycfhiMTmzdv/6PaXo7DyvrPfD4hObhaka9sGGPD
6NO9/wsnpG7Zq3pJFhWBPmCobsaHV6dr6w8UIbsj5ZLw+C8eXjOwNJ+R/MRuopCC
OonmBnufEX3Yw75gQwiDlqkSri1eIcTi+bD0JExIzYBV2FyOZnj27TVx3lradRSW
vNAtzLhPAmTL5eJ/D2JOdsmyPkKTmiBBu3bHPFXaVGBin0rXWDkhOITSfvvVuToA
4mDsDv65d5+SIT+XW0077iIjEbCS31Qqox2sPoOY4Uke6b5uy2eKoWlw/eGjjnYS
tA2Yh+A8T0As2OcsnmtWpV7wolsisuc3v7/oU7E7jZpUnE9zJPZGAOig0vufiV/N
tvEIyPV5lU9ld7QY0Eus7FsiZWc6HuqDOBWNVkZmXibTQYsEOpegiIZi0/gDjEaR
Yz80cxrZHKJX0Aj06q7RSogt5DO657VRWX5t9Rzsm2z6m9GF2ikv+Dyc2qWwq86g
8lPVTIhxKeCdMQXZmLoS9SRk1Dgeer077RKpWfnYXXM4SboN5PEwQkw2Xws7aBTg
DMr0BEB7sA/xRANRU2YdcSBLhsdE6wrGGLCql4wmeJF8htPdSdeQHtgkqL7a+5rp
DiFhmdnsXavtqJzXWlr4gGXP9jJW6E3/1A0xuAXLKGY0BEKXfNltgXcbV41D+c7Z
ZsxS2WLdnYx2xMihv4382l/1bhD/eiBj+X0ItcSSDHXixPEA8zlOTYDxXzbTAhSx
yZIi+3luDCWCWMV0LJcRODw6Yoy7YpVtPHszgkZQAb6Brjrm/REaBuCzLXv6mwlb
Zn5spvgPdFODDZFGLxWxAwp761mndMrxmGjZPJZaIIKgQeMCEXz7GshsQ91+xpTb
nuRJmObD7PPlQWz08ySRsP2ag4gylw2lTM9AmNcku3mSpPuRfF+Ofz9aUortLRMV
jSNqPbMGa7uR0YoLUQeDmsUbyYK+xsTtTKMBeOmqBPWQwFKx3LgksMLACGtFHdHY
rxh6tkBIM4ZmoKPRk2MuuS2d/WCuiP7BidS7fnQ5zhzdjWUf0AehKyIcA4AMkcJd
qSihuFuoYiKd6M+hQMT7Twq4V6Ngpa578akvrq1f1FjWCMm88yeWC0wL6ivHaPju
aGD2gFSbB1HafZR1ncZtUZdWa7qja4wHs8r+4/Emq05Si8MQ0tKuQ3iuck4KBEOJ
PBVcbmFWZ24yHFqGhRUhYNt+Ulz6Q6B10qTRauOcoCwkTZ6j3XCtOjh6GZBm+CQk
CFub5itiasVTaTTeIXS5MCy99wR9h1ExZm06NSeSCpbeclorYmdyTPwj1FNmpcQr
NjfXcW+qJzM+AsjaV6wK3e3xoA/O4hokZMj4A/+MBbGBTaZS67sbFPkUGegADt+I
iyuJOlXMI1fMy5DluIBfWCIFgQQwY1w5Az8UGgjEtj4kvxsfHzTaVTvEzstFL+HD
oULaj4otTuxEM4quucX5x/CxRfGc0aB9GBSYHnyanFt2JtSr72chQivPCtd3gF/T
W/fpc+ZCOzVM68MS9Pm7lKxLHYgv5Rgo1w2la5LhkgHlVOca5GW1vRm6BYKXPsGZ
fl0iKJeGcpoB73B413AxEZWEv3JLxhlgoMa6jCz7X9GOVP+zsjSl5l2ztbDq61Cc
WPEARTjaVcFx3B2LgcWKQ7JS2PoNKY4FYb3/QuBChVmPhR/GlmivZ2ESwbAMwMmm
3MoLZbact1ZvAOF+NqBVpCFatx4G1eI7wtEJVYjTijc5cMLw4UOtyV2YOUW1/emN
BrfAePo4ssnQ1Xs++0jRZFzvRkdeZICLj99h1zaOs8gyHxSsNCnCjEnNNfMayanj
QA6uqt0i7OxjTERyK6qUI4Y6V+tK3R1dFJ9+zqYi6ihEVW0SligeA2+kgmarl1KM
w8xhDVPFlt3D2ggChcAdLLP1KyBxfo3Fs9VgqfpZZqyxwFVTaZ9/yEm8Pd5+H4Su
iii+sec1BBmxyPORg3pnv2+adw3VznxRxxyQ0H4jD1VMTAf3D7hA4/T+T7naWy6r
z0Xcf1JH0Rt4y1DthSdjFRzVTzR/e+4YI0+XjPAOBuvFJayge8gG7nqb3jclKWgi
pLhsqbvGKt6NSPGbDDnq9PShng9jNzjF2NjVameq2psUpe7NrosHw4p7FyvSBZNQ
fNZxIk2a9nt106kLaHv8Q016SNcC5TxqN+dWfPSf1lZlfxtF6XOKgNpGCBNFb2IF
pvE+LLp3CbCe7aHCcMSix4yur0HMP3I9larHi8ZQK28WH//55OKB6HKLvv6HbSn+
neo2CllNC+pVxmGcuvmDhrhuXrqLiMhxjY0k3MpMcjD+s0KXJtZ2PKFE9MhZ3l45
FeianiO1bH7v8GdVkgUD63YArbyu8AGTC5cHpihVaoUPlu39+SDfUIaqhUiQICYj
STvPCpTn6szOfj/tTi0bnhynxztML3kXhGRVHj7Fh/FTEMnqynWgqzsmSU70QRK+
yYssAC0lHHArxof5Qnc/LeYfyUlD6x7IdAg7WCMh5txVKXfFNbQ9GdJAruawH32X
9bgHHEObnbNkdZEGQt8Y5yLc3HqcIA8FHJiTT/mbmMlftJ6NsgiEtuYMvz8aR4ab
bV74ozIG9ONbkc0bUcEUm3LOZDVTYg6e+5DS8icovkoOGRkKWrrdCLTF6V0Q1gm2
ZbjrT84ZG17pBqHBPMGOaf7sa2idw9diaEQLFeyvhn1Q/3PzYSseY55SLfdRPE6L
OGOAYwP/zQN4zixHKeu6KM6Jt5zfFdboiYeRvUUL/8cdAmWqKXVMYMqtDxp9RTX5
xcv5iWul8Nf1yBVpeCR+gWU+J6yNeBCX6doOv2+ttTw/A4aKUswMLgMOPstV1CYw
lSijOutadC7Bs4/Z4KRkiu/T4bV/vtPfi62KM8zE7E27FgBGfJe0oBkzkLj4+6bG
a19FOQCzgLKH9Y8jdqBk8m2H3tx4hXiuovtmUhmXvPkGVvIZmG64rQjxcO8XNSsl
9QQC2fn2OaV8+6M/NhlnIvma5yJWq36z6fj3LeGvy4Ktbi830dDSKE5if8HgVNKj
tEnULIPvNlSmdRZXYGlinS4ZrDt5i3fnJPyC/CoXOvev0ljmLxvFcjD/OGCZgPBk
s/31CZysPTo0KiCQXT2TILQGOqksbTL/AJSK70SGztpafgMwn48Ijsp6U+vZFWdX
xGi8O03yL28AJeMUXOGZlzmbz0LsOHXLBcBFn+HaShH8/bILIS2BjNfmajqlgOlS
GinwKBwVDa6Dbl1ncpanI4TLLuxoHkuLidFt1BkBPng1BBoa6BwCpYdTwI1Zf5dK
pt3BI1z0VAjrRj4S/I0NqOU+te9yz+TBewjs0S3fGXXg8qZ7Z1I3kFPR5BnW2Bzi
rc74+xbYLc2NzK52HKDUpSLuSD1aMC2Z74fFzm4WINBDdyWSOhp0k2Zf69pHo9TA
jxARJ/9OcsMKd3Fl48CaH86W/elkPBinrSyu53Rkue2+QDrICOQs7rcxTKWQtimY
sWE0Z3AxRpX3dBvsHMaxK7gYfv8tHAwoNksKKmbAYejTB04NDl3z5ysvRbSjjLLb
GdkQBi2kl3AJR+xNWIKE/kh7JSHMrUV/nKViGl/mc7p/AUHKRb/bgoyyi3zMG5pm
zCqC+l5O85c0FlFG8yUt7dVOHrgcTZ04dU+QslM3E9Bdb9uq3Jpb/ihGMT+TN9Gt
9qBt/I9KQuL1S8ykGWRL4xWdcXIkGHWFrevCCU5iVoPvH/L84pGf7RYuzNOj/I3n
Qs+kmM3c/SQCW7shMrNAL5TnTWzpKg5kQlrtUGmURVhRTnO6q09nGc559GeWd2yZ
BXEYdnw+zo6Z+SSJOITfJEyjmBNsugXL69quofiv4+fz477e6HdnMnzFlfmGu0LJ
g3Oei+d0bwGwg46xw+RjPZABMDnEOSqKRWvhVFYgC39l+T9enMtk6P2SiKniefTq
Nz7vBwppxWxfrNgMxlBwT7bV7w5Th2Qw8OuO7UhHWBt97BnlAkcm/L6ghgWzRlX1
ezVhgsx9n0kWxnK4ZW7+uWZyKCj2CjX/KE3QLx4Y1maJDumydxLHfhxbEEyeLwsM
LVdMVVZX51wgAKEOqfCvtYeY5YFA0hGTdx914IKMSjLgnt74taG0nmJOlZtfK9d5
nbzqykTYafACsImzv643Mou+8fcgS8QuYhhtqBn2ypN+frzN1Vx5/4WiBs0m7NBq
+g00hFupJO9DSQCw1MfrpEyBYw8tVHt5WSNDIDMw24UvP07qiDOJFJ6YBwmcqcDm
WB7i7ujnQ/mg7vueWJ6FTSD3n26bp5izhteJMntYZRLcrso6XmpIt3zy3sw1Ay0T
c/UmlLlsSFOUQikwO7IdnWCkJNdThs1y+OMBg5p71O0gv+AGfOj1PtG8kTt2Ud9Y
d4JlpKLD7nGWtPK/ITvYe9EBwbsVT1vOqhTDeWpbLMnF3GYNvxj9OOG04F/h7GGX
Tk1RFW9xhTkPvqKGyiYqTR3WUSNbrI3dRdeG7mQTt/R53rW5FSFx7UVpinpqz5br
TGccJg+bvwJ2LXLQXH9DVUbtRPkP5HiQkLWuzadO/SKb5tyHiA4YuyxSPaRvYFC3
d6pmmOZEpHn9o8dLU5SAFItxaHWCP4b/aP8hUgswP43DqQCOQzhTByHa2Asohg+p
F7a2sbw3dniCtOLmE4jDQmtBUuicvbDEqOJ4Z70Wk3H04hLVNKNRAMV5t1fF0Oo2
9Au/Mfvdc1wSVuQYtz1Xgk2TsKOybg1BLVvQPzrOMKz12C4YGLDe7LJv4TOWoilH
qRaqkILrDJPDa0+6vlfJSEuCk/PS0ay/yJ1pj0o7T2uqhWVL+J2VIHOZ9gXALQel
TNQX+srgUDPI930JmCRFjSOPBOHSHnnr4F7Miw9ZR2YxeXezaS3PvZiq4j3tch3G
/i1VXdBw6KnPUIPGoAq1RbgqaUk5VyJvnUetC0MoNgoyxNutOrQYx1cM71Vmc7Rc
DG0aMTzc03lNb+1WW0aIh5CmJtcWHvOtGnNQMw3nI8+CE/1dky++FL4U9QVqr2Az
pGodhUzZcHlBJaKztl5ftsQu69M3y66aOXjEa1W+3KS9osw7CR+Ee/Seh5Im9HuK
43OIKAcEe3dJdirGfZXjLAJSUT2vnVXje1CsMfBmGApkPIkFmYWukMjL9yLnkqRt
6C/FdzYzXIlNT+jhuOTeNk1ha+VmFQjK0uWlh2k3w6+9/Gm1MWvwc2Bq0udvkeLd
HZO9gS3NAZATE5AOLWTBj99THP6NgX/4R0zyOrCMlm0XMqGB088Fbq17d01gmsGL
3v2GHunNpm7/aXENHyGLNrXmKdXvk7FjpVAxFO7aRxKx5Vn/JgJFtMcoA5S+qKwG
k6Zxy9ozc+Ge8ZWLGWMOnPyJBuUGsPk6gM8W3DRUpkNh2u6+/axd04GVzu0gyi/P
ROcKkvsle/DspLGSNpURtuxKuvJaRrVEaAuLd8urMzALyUSj2jUfomUML9ddcwk5
uytXoUw4fEGWF5wb/3faEwe506kkbtBJ9tnB9L4cPB7MEER3lZ1gy7IEvFyp1g61
25E3XJrgei3oUHX8ajRCdpvEiHdMzYFRepiiVxvYeeLcZaSPsAjfDxahpvFRYeub
l+yjnktFs+gn+IJ1GPxzAXB/Nhc9MhzHwC8r6ZgorNcQ96fBGwYb4OZyCQ9We3jR
YX3ThGwLt9gJVRX2ygymEoSYqZXl4UGJ8a/JYqlZQ3+4sAUm0i37tykrAr2zaeI4
656qBvXfJ3AsIoKevdroBxPBoUESGg/xVZHUuL6umnyYGfhjy2zGYfZj5CxpbTlu
HT4XkumRW+Xe2xCAJd6unrM+ExDBzfy7aelCyfk9v5XdXRNjViafeEAF2v1r1itS
V9MYGilXX5+rhZ0mU2ol6UhhRIea5jsEa9Fb6q4yWp+s5uoDQ8O4vPsRpVMAi5Lw
G6U+Nti0UbE13UmDj/gIRt/DamXjQaKF0lar1L3jCS/BM9sCeYDNZqkwQVB068Hn
LYfGMtnXPjTXM+40S+FRRMlFqFYsfKUKS10mbxQG/8dncQkon+66Vlb2g5nPUBfG
lJPoGf2vW0j4PVwvmO6oq9d3E0URNYdBlqLhsQwQQZoU+F0uOvrzj0I2AGR37LU0
FIcNOx/BD3B+H3vtoPHMfdp0H6umvauHVnF8P4cAfun3oVLtI4PHH+XNCJM2q0UH
aQi/OH3uzearQLt6d++wh+SCQlYeBB/8TZH/8HdPaH0jAXe/0BXZeidQtf9glHJy
9nJYVR0dOS9qPVyC2X5dzWSfDuYCbchVPSFwl/vDgFT1qt9e4dRzyJ4bVdj+HgZB
y29losJOAPIgLtPrKwER9y1QU2zJB9DvXVv0HWTOQCPzx/C5RL4OzD1ybQ8MWKID
r1hno+nYf9EaVnF7l7t9usNeRLyGchdL42hCuwCzieq/p2zACn2WS2qDrSgsQH57
NugafqMlzgsde9cAW98GH7o1AGVDAUhkN3y1EGjkJ24VEbgM1rd+VQ3JvXupgBF1
Gdn3xHNt/Mm33hUwOmegw3oW718giMvoS0Nq+6zA2eZhNYq0nE+KOvjgDh2kB1qW
SCUwH+gOpC4ddZsvc4tcGiPX2EYy4iWKcvsJDILUhGWgXMYzqv/dFTHvuB71v8BF
r2RIVA5IhyJhkg0B2lX3HGW6FcvvPA3VmoDaDqtpbadEYY55i2QHwbo4u/yXoLzM
0HhuxQzY3/GhqWA1oJ+thSGqlagaZRW9Vtb+TYpgO2+olnQEQF34er8Xo/bO236P
zojyUAV5kjtf3/bwP+CfRT/PhDG9t30caVuxl3qNFykiII0aXqbzmA87jMd7E1KB
d4fn8zIvycuKh4SZoakdkC90RQrmNAuZdMdDykyaIsk9yh5PnsgbUwndG8gxL+9c
WLav0kd+N2WQmFXJ8n4s9FAzo6PG0m1lxRSuRQ3gvoNe//0SGb7Jk1/4eQFqUCYA
bipJ6dk0rhTl6f/xgZO5ngzb2OUIhG5rPNFU+brAuPTLbevpR0Ua+K4tZATOssgO
QdOHwxrhMW0CXj6X8kTaAopoDPEEqy/zfv0/zgVNOq2Bsr0WNDEDlrLxdB4iRDu5
C4g3IsfeR3XA+FFDFPzMQtHnYzmz1YZwsPeS8BvUuH1ADq6j/3oFLMEVAtYZCsBF
S19d8p7mVjHhXJIdcJv8yw/Nx0OB0qJfzEhKpGYDiwG+07U2z9vpGBxjgY/bI8lU
rkMor/YFVxXBU/JzJbPsXrLslDoon8wS2KfJMZMS7DORyiGNNg3xRLKm2dDaIGho
m+LuTEdaivfa3PZRDVqR3uNP/TIFDDAMllCwhUDdzE5xqcupj3Fsh6VYpK34DKGj
AUARErOk4Ju82xiGWbYYBhBPoShOl2etj+tktAIE9yaQv9+5CTxKX3AKy27RtTd3
dEMC5Ab6hpyMRZXIlWpCQZmJq9qFK09GcgsPQ7yCNNM3BX2dtO+IiCqAqvbx9TdN
DWRWgztg6Cr9WkHIfy6p4dtd2DpoDTZKN0yjRPDiQjCxfK31ShzE1zqwSRKkX0TN
GbTf5xr919NgtGUkMs2rT49KJQ1tkBOIs17hLDmCRTSKYEjvmM7t0cuavgiO9KFL
mucO8GCfI9kkP+rDNxCfKX8H8Mtw2Zb7avP+/yuEEi0Ik54Cc+JJZbZgoUzfkrXp
4f+Y9NMe0/CxVVTLTrIgYGSxnKEPBLVuTmRA2RJv9FVW0CyG3DRwj7PofuYIEXo6
eoCjjvN923CE6MRwbLb3UxfDzoWZ6sQj7q42rINj/cm9H+7BhqtFH5o7F3CFu96e
+/WZ5GesOxgsSx00CypH4uI3Um2dzEYvwUEds3RblToGjtYC6J5FokkqVVbJCSga
jXuHhlKtnKmyJ7213Hxz43jlyuZSzbGa0BCLO5AVlNP2ERRROZEAUjXEbRAV1Ghw
F1r/4xcQv+4sjkV7JNe3/2Uqnwlf9lijGuvWtmDSPe1W6CA0lhh3omO4kR+q68Yf
wZ1SfN8XE8x4rgt36WcuDP66hBZkDrR2t2IKJXc7gZHJOd252eUsY57oBjtiCkjT
Xo15w/URjd0myGaV9fEeQpLzqQgNInzEDsmy51UYY1I1OvgUyeP0tfHiwYv9LXsv
ee6ULVx70HV+DE95zNADxeu4wr+QBZiDaBkHT+QHAPz5tUMbmYjDAg/ruWTEALyb
PL21uJT1bb+OwWESlZV3Y3m8vLcQqRUYDxMRcFvicsu/3ErD3Re2TDeEsyyivKT4
q7+hvDPdOFNPdda3A1SicAm6e6mxF1/+4PFoQYixgkWiy2Pgil3TrYrRqJzhsAM6
XSWmRMoAFAjo92SkIbdO8FPp2LuEigW4zMSmzVfCANfsLhHAmquSrE9AsBWRf2mY
O39BDVEBkgTJc1NuLeCH4Nx2QLjPivurLGa2STml2G5ECcCZjNISEUpKdGYyEW2G
HDQYoKosnVAo+IQMbl1XFaDMvJpfPfsD2z0ClXh7T30mDJ9FOJojCzP6R6rLThkT
YiKdnaywjm5AFVinr6LEe8saHRutpxeB2wN8p6Pb92w7d7oB2jpKVfJiO4IgJzIp
uj65WdxF+aNwPEM7DZQvVQQaa2fWzOcfqMfN2tCIu/HuwWubo3TccYcrjhZy8VAf
YXPX5TeXi+/j2/SluxN+K6J+0LdaPxJfUbBsy5Q+3b8qkQjaIOc2uMIBa4ju8dU8
0lrzr5oFn8mfoylBZyRssGpkUz4QP4nbW+7SVE/iAs/fgq5PVralG6Sl8YycU7g4
FPiWJ0JdV6S5SXEwqMG2WOu7D5/yzdomatNWQQ+txKcatixiWQUNHZGjbJ+KrmGu
LhiAnr6s+sSckNAwIPO3dwpyzzFJxCNO99v+d2xdb8PfdBLJ92D9xyTLWBkeOtg6
psMcB8qm3OT2XX8XLmDqzspEfvBzY5476k9m9BBSdSEFZVTjGvcpjY91g7hUTkjB
OMYUZe7Ltu52jfMQrpROSjOQzorFArc+8bbX/EVdoypilqGiUaFqKWsnkkbyeNZQ
IhpIawhSreBVSHFNtiYrbFUfaNKrabfwbiVQ0uYndiJQOCNwcOD678MtOt+BXmjb
9xHp3gwfCKv4cJPv79SKjiQbuS0mRvv39ewI0bIKBcmPuJ7dcTd9E+sACTYAWqGl
SMce4csAn3j4zIbqRBnRTizXMR5dCVcexex7kCu7SJ9KkZatbmnPmJe+J7XStr9P
0jURwWbO8Nr5OE6FyYdaZyX4NOhhotllxbCIBHJubcuevy4NngbiNzG2bg+6ruFG
keS1SpGuaPIM3uRVlJwFjEHOJ4qhxFQ/Slm3AnZWH4DyrIWcXzeNbwZWRaxw75aG
+1moSsDbt7HnTRFZUyboqZPgtG8+fRvMY+uZxZYsBkEVJzg6ZLRDytetuWT8o88y
rWwgxNevNq9BlKX+8ZJzBMGLSyt3jSilJ+bjQLTILGwhQGKIT+87aeSWgI0qLxpq
1UCRdWIi8EnfRC3yrqx0CNMIdcxXFrSPZpCDez3go9YIv/pJ48fbThKqhLZ2dGCO
ozPKx123iPJxq/6sSdnK9yYMu5vnV8/3iuUQgM+nSuJ2fowVVZRnbjGq59nGdHLw
cbzX7syfD+c+6cl/hdgCfE3t8H4IqkJPPcj7HewlQjc8IW6vcfhx+eAlSQW4nDic
N6QDlF5xDkjXOZHDt2UPx9lQ4eiyzkfamLwVpDh7jZQQAESobx+WGub52iaBUj9Z
3xdcnwfXmOvqN39v45oWpNKRMXgqQKC7JVpORquiG0GwME1UoWoUZPLHn+u50d1+
TzGP0Vl2OzJmLKgS1GteEY4+YI+QrICvhHLiPW+zh8DgHXBcRDJbUYTdIF0rTyuB
SaPyJH9VTqVIgAVcSj6CU0HdCPKlu2UhSf1E02uXXAU6aWbyyI34bJgjR129mEYU
ryOuef2See9IYKitS785NkaOuDOuRJsAtxWZnDnqSPPyVnSWtoZQQg3rBDIJbJH5
7xoQ3f2r6OSBtLeaHG9JpzvA5tU35n9wxT/vfAAYchMd8j+LBSC0UvgMt4pdrubj
4J+aLszhcNWO9yLE56SutTB9daLXqL7E9sXa/IqQw1/HniJhntEWG2hdfjMCIy76
KB+TNXGW4Pzp6/eWbwWQHbwQWYX5siQ4ZWx6TNsP1iLuth4aafO39GAHOJxW/Epq
vpbr8GoqP6NgrdoJJnVIo7Hu5YRO/iG04pVubPe2UpEFN/EepAWifUbNhML7o6BN
jHDpOOvNMRUHoNuYCKnY/8Wb8Ziu/ZGyNB4tLLe8LQbYp8V7CPTm10BLRy3ScJxk
N5W1oK32ma+769pB8r54JbT/PKRi702o2apd3CMwPwGp3QFw3wvbvDJLLxg9qged
HLN3DbDiUDhr7bvs5DtuKslbLNZkr1lkfni/N3f9zLXbyi6roMsW9HQtpqaXoIvj
adZeVTVwD3mmUkIGh25SurQZNkfwwq/n8SHhwvNayjeLQnMXSpDfZkeq5Ljh7Cwe
kvFxe2ig+0ATxYy90A7/vMcUqmyIkj2QdwKZyBN/e1V4fD/ceecAmgVEKKEw83fe
f7k8yM+nld9ArdLT91wzFZY4ewckzHowI7Kni/1sMoGaijlxp1ChRWYRdrV54nSu
Qifu393eluExUFuSS6dl7rvh1yZ5OrIHGzw6+qmrIhfpxSzA8zv6XDr5vSLPT/Pn
etU0v9kYbIF0hlndSZQtGhZ8azwi3bm/VvkNFufjhOttYFn57xB+j569cD8RmJfm
HgZFTSQhV+kc3R2ZZVILAiLpHqBStft5JKedcW952c8n0CQJKrp0Vlu9/uQpc1w1
6eWQ81NfO1VLhjRCUmydNtB5LeVdRdbSgHBAXgb4fwFU1UVSUaHUx2aof/lGsS5a
/XamepeNS4IuAaTChCzIP7vIZ0A1NHt5QONahTuh82bkzOeAK76vDj9FsSMqQIYm
n3NNeW8jBt6cSyIiDIdtvwkAO8shd/AwPhaXRjwl1w4MnHfR5LRVTY9xH8GfGhew
CUcISgx4owRdjUULOYNdSdAp7MlwIPlZm9r41Pw1qCNvF1RNAlR9rEB+nyQC1uw+
YZPqCsJwU6gTEnaVTOMgSuzbBfg8neeJG+SyPenj4JDgxgKp90jz1diQ6NLt5r+A
uimvKcvmxbjWDifwuF8iSCFOFfMD/EZH1GXlvAR6927TruMc7Q/jmc0Zgi41bD52
SgDd/1a2EMCt5AWjdFArTXyr16bgm8j/gWzj3KGnDiHYLdRRT+3pFTIgh0X1HSZO
URztRB0LW6CiaLxJmsHpxo9hYsXbC7LSyHk+BECkqXAN/eMOYvMn3oahi9vyQVNC
TQYgyaoFgA+kOGJaipEIVopexWBPE1BhvjoY15Fl59UNhIa3tJvqkPO9ds8RjxOS
ZcDUvtkEqd7OUSNcaav8F6W4Vyw9+f8qsb9gyHkV+FzInVDK3YuafV9tIUYOwxct
xVOIrNIaa8lHazLQ0TC2iU9YIZysnyrIreunblP/d0IiuQL+ygqwOGLxwD//Fj4V
WaogUVnreMVxO/+gU8bLTBnn0dadMEXeM/nhsWWlhNYbwKO1WqBJkirUX0VGDzrv
xMeunleMb+pD+BdGg+xqbk/s5eImYDUgDUM2u6YAkhAab0EVWJp7x7FjB20moDId
qMhi3s0dOjzsXDuOTJq9xY/pcd5h3rKo3U6FUjk0GqAFraF5QpbjUx/WOiqlM8Lu
RZ1sdflbj5O05c8zw5vJolTaEUTamQKYX8nxoXmPQAjdDUbhSoapNbKT8B/pm1JX
i+wrdjXbajWFtFqf1NfTAbwYxAXbXKEp1AjelEjZbyclb+B+hJ4sqzlEfEPPVbGR
RIQWSr7q3LaCuqiIZGw7k5zvPXsMd5azrGzVoY5g92rbOVrpocXyxROVs0xwSVCG
ZP3fDI8fc/R0RmKm5/xphb8LisVWhxGeY2CBZI41qDhDhDLoFiIiu9+fRU2ZvArq
wFm+n3Q5V7twkR2sKyOnQoAF4+cAbBNJpVITWnDoizgL8RNS3EmwXpMEtBVlzGIi
cJtKF0FaYtbt34s3l+KBpqirkA+5l6pshlGDiCc2OQCMWFBV2+vo2KWNGyfZEdsX
Z/oRnuFsNUZIPdUoEWQyZD7IPTzTtxvzrxtkDLDKamyRdX5F/dPn52P7DAgkrWS8
KyDbAc1i/+0phZrVPPvHDFOnw0XH56td3cfZ4Tf4Cd0zX/9CzsUl9OtMY5HyQmV4
G6KmsxSxbTDxEkKEB/zVkqResTkqT2mcp8dfDaWF4+LxvwVdBpSjt683bQPVW9RK
OW5m1h2cEwtvI7KdTZCh2RMjMHTn8PHKmAKVr/gd+sShmSt+UxpCCk4IIKwsxm6Q
S/TQjrAXFEWkV9pF+3j00iM2eaJKm2xfTmqJbmRS36nwYJfRKQOsIMDTBHws6H2Z
EJRz7C/1a02kPl/rTBHSKvP7iFyvjSg50UPzHCLGoAZ+h3WIUEw3Ssv7kKVNqR5q
h8RSOjju3xaFBspvyFonvVjkbzB+lQ/mo/riNCMds+FJnvWpknIfqI/7H2fXhLiP
Ar/0f7Nx8s3QeuCadYwR923eCZVVr7nBlVQTaOnOKSQNI1gfoJqQi9JltZM01blu
v0J3u3e7v6885OKRS2NnwL6R3EGKyjQxOchTFg9RAc2vR7GT290Q+zlfGIDKtsJe
sXZzmHvokYYkxZK2eIeWhyDvJyW22OpwMceB2zevTyNUOFqpm3b2WtdFmn0akPNC
73NbL2LlKuOQHc+XMq1XAfaTKYGx6WMA/Ofik08vrBsOaFqCri1c889lSv7F5Usf
ssfW+gDWFXktBZ5Xo0qN7V6RsgUJn4n8dwlGxjlC+92h9yxEplvii5r4R61vlefr
Sbz9y9u08ueTcUUpv4FGp5ccwIMy0DJdNXgMwJqbx7jhI7jgl8DPr/1UcihadNPr
MJAcbIMh5p5de+saqK6MoXpUY1gtPiiuf822VtPoG6SRBKtCY80uJUoj7F5KfKuE
p2YWSjBBg0kLqt/s7+GNK9Nj8zD5bmPhuEcwBkUDkqiTZ/yrRYb3nWR5xmJib50u
jddTpZ6XKwi4UlVghG89jM8y4A17JG/mjoTG5yUdmD3m6Yyxg4AXfjDHWs+Aa7RU
yFZO7jDLFfFRImu/i0cBnzvI9GTcxqSLvLqVENYUg0XP4Cfv/xPkA+tN8mb884dp
jorGtkblqjM+6OJndp/nZu8RsfoLYTeb9rBZBRHpEK94Yx8xDUrv2Y5PjtWIVyVp
OlwZaM3fDi3T+LKBAcOLbIpKFMoMIO7UEfIF02Ass0FlWrffgMfFsFRNL5lUzM+c
UBuEpccOQZA0v7QyeQVQzCr0zDuBS4TUcVhV7N1VBwERaCQkTiRmwo0CuQcbiiuL
nICeTHyMmrOI56GPHeXn2F665jW3VnbZMf/YqLeKFqLY4hASLgf9GKSRCr3jbUru
E6RdnLkL/wfd9n0f3g6krwmnypNQaroCCVtaXy0XeHCzgHSYV2nEZ8BayPYSIEjn
FQI0m52M5XfnDPDstsn57Dnu2BH7RFnVf5Fcv8CR0B+1xM9JOaF4Pg/BZ7zeKgdJ
ogLh6j5Ikevt9RCImi1DGDrjT8cVCrUTYKpywrwjTRLxlpGomXu/6oyoAYNtW5Cc
AePE9f9C+bNURpIAlD2DUQgt4HV73ocpoDsFwjBc9yCua8O8M6KilIRfQqaKVFzb
3hI9wdBkb5LBtmaXfSJrLwYfXTBV/IcHQAM9aHBXlAOy2E0m1SW0ioFZOLXIS8ez
+Y0UDLkK6UDtYyDGwV3MK2LEJKD/GkbOpM1VN2xsH8M6mr/hXuIvayUoDqwxCWLv
FSNrMKAXRXCgva/tmpQjFrmIm3410obnoWURgIVnENuzQZN9bWd6ECDcA4osqYjh
DmVIW2PEAKxjzYdkcqJhuKTBXaFP2xb1AFvp7g5GUSOUFamuKqs6mY9kcG+GDHlq
03vDeHt6osYeR+hKGze7G1f+t65e1ZqG+pSeevRFruXAIjRFaoOvTKLPyBR9g5Wf
qBxpxyljStjWf98YKRQsZ2QBx/tdo5Eiea4Cf738jKDr3IJ6lWYHe/AIjVp+gd8S
MpaBqF6sgHQtHltf0zTDwRJzb4blGEz6XR3Az7nIdknREsYv51pn6T9wZablxjre
cKziYmXHJQ+luT2HpncVWfpvlynAUwHFL8WAxHK7qwwiJkRF2WmyjGKgpE0+oEYY
yX/UOQ7UoVlWbQg5vxwwfg==
`pragma protect end_protected
