// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rpi9xcU4NzHAfMer3vxEJBvnuVDjo2WWqxsRlINWkqJDC7YJ+pn+7l9fymOFy8oYF3/l0TOlLpZe
WmNZ/b3gO7zEoR9c3SZQ7qLjiJO0ToaQOYdiOT+6aQL0BZIyyMR8HaWugt73moCCtuToWoXjfVyQ
DUMhTyDgrnmk6ZHkyHsGLXbR3nhHXS1UHvsKV4j9Go4pG1nGjvQlxHejYytncsZYyno5SvPYiu3u
Moqj4j2bnffk7uBpL32oZ7QzliT3KR3X7Gv7vNWiSIJq/KmGYkPsVsKMQUwf/qnri8AdtO6Kj2FH
xlds2v2XtGdIBWuuUUBNrtr+RmcMop6rtA/RPw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14352)
ZPzXBl005VETMljCWcPolBSSidCMUNr+FUlufMFfO5l4il5yQomG2B8eswvwEPT7iKUgFO1+698/
6wVRqXWFyAOJ8mPbtc+VeZvUL+JphtkKJK1A8JMrYnBxkZZpblccunX8aYEIvpkZ4wYQwdpEN7xw
f4XYE2tkVfxLvaD7ioQIfT9o7qKSsYRKFhct2KGmCaymYW7NckwFx8RsaAWK+0ltwCAWOtUGv33P
a2jF1k1VRCcDJ0OViJm7HUj9oAY9oz0uKCD3WhPnBlMcESmIV+LbyTRcKwpGAS8hqGeK8Rc1eMju
vejlGb2o40cvFxoKZQZvTxO679QoFiWhRaotD5V3PCojaKpiqgGjIocDglZkPdEele5vJuappLBU
SnTss7UVkHfG4fx6cgZj+L1xTHVPR7mY9YzKNDbHQOpX8NIR62+unRwbCQcxkZs2Lac47zd60kvw
5aycwZndlRq8FFjmUejdK4nz6HCRWRgHVVKbFyNShPosJi6y0QmmzaZqpLy+fBAAZKOM2F+Pr5Lu
rcsSB6Cb3qm56QCGJN3JS1HQH7FpJHD6toUhC9tgNUiPwwxEKoowuIQAqGHQfeIKkUWzMHmsqzF4
c4r4roGTuJVp9TnbnLAxT7Hll32AvWgYSMcZ1Wt1zjARXLzLHrrE3L3nINcX9FQiNr241FkXMiAD
tuEGtoaO9NQevMThz0fNPDgks/GBCj0/rTBY9cEU+aCh7mXg3BfOJ1RSSSpircaeHUAYeaLyAacg
nX1YYJte2M+hTMx5zvFyajv0gmC1HUtnhBEIZ7uzMSBjKvLuMvekXJpqmsigs+iU0Kkq2xyqVcy4
LB3tIWoQZp1fj/j1I8vLOxH9UyrSj3VmAIeN/5LE4XuEJ0loEErkjaGoIFwTJym4k3RGU5yVGVz4
CPiMGIKHZhgaIJbo/7xSM76RgRBJ6uDsLDpzWGtf/Ptxc8HsTkZgUPZg4mgBsAitli9bmiUh6+m0
kOZWR15WbsGy8MkB5BtuwXVZLjbNccgZhjaO7j+ktBhOLa9VbrFxzxiYOwj/gT6MQjOHpE9KvXKa
0UEfSIxOyOY1m0ivH5VylFT9nM6/PqSLDLSSx4bqDs6czV7eWe1MXq9QGizbHM4lpbrxr4JkxcC9
NX+njbhjyyEPP2oCr3EG+fspoP2EqVmqmi4J8ZRKg8wpOsk4g+pX0GrWcvbAO6TRELLCBA15Z8/f
8CBFdbGi3b8ma4w1/VV6vBDQEOskhYXpHqAB78fc8NkLrNYYuGy/o3etp4y1/3Vu4GlT0vjnXYNG
WABd3QcF8rdDhLsVj3MBUWIvrgInKxeh+dA1+Fg9I+/xCseut+7pUSyGBB2pk9SCGNn9icii8yPI
L7qd5TjQHIIre2QLns33tGnn9mhu68QToiJ6mELNeym0Vgh/ld9lQkO0G+fgFbimzoN5yL+d/OKz
kkDT0qrHkjRkFqJxkMlv3LO0QaP0vrBAQ5J+YxTIzeOnLPQYpT46QtKEOVQQAXO2omQ+iIJQtYE9
UepBFjThT1wc3X0oCbKKFiga1mDWEhIsHzrB1YBpgCM3FLljIlbacypd90RrcUKCNeE87bZ4ICRX
XHsvrGWXQrqE/0zTXCZakvBUPc7NbBtc5pvDm/Oxl1/cdkh/pnWGteuh/ozdiCRwb33vCvO+Q0He
I2VPjm1vEXIkKxf9H8eRG6/opMjWvELyo9SYIyp+kgL/Rl+N37hun+0X8AAWs+lFQs5urTjdJboy
SlFOhPBiGqVVGVeWILj74RYSq6vgtqUrXgDlMAywX6fyX/24AfkZEpsWciKrIxXJL5MIsJh65nUx
E47YG1zu48fkj2KeVtl0g4ji/eWGOKFLtLc0wC11ZBib0/74SRI1gR5xsbUQd6EpDJ1vGrd0IR7b
mQu+XXTfKcWvdgO4hnQnuquoGy4hJ0PDPp1M5yAu/zwGCfNow0GHnCcHn9ss4YHi7yAv4kP65EXr
RHu8bazqbaEQXWgUjRCAI5iyXtPqVjZmEkGUDwuBE7EATzgKTV6eg+hjk/s1i64L/aDuNt+gwdQ7
jKhn/WRgbw17icFJ42Y42O8Dde7M2VQSbiAAAPDBJJcRqDQalt+p6z/q2B1MaebCXolduRGlvDYo
Mm5A9EPaLWCO94PXjFsv8AvTllyNWy0oPCjgIN71WcYmxAy82H748B42OhMP1f06Kp9ukPraBgt4
zuEfxrAAvmn6jcom8N8njBW+Eo0blvTi+0NULMjkSAUS2nGfL3qwH0ETcOLJGMTKOUkgsF02Twju
tDteBkhvoigPgE7CjnNdg9aEz8P/dQw/pHizcz5EPa8wt6zQ5zvOOOUQEbrEb+VjGw6qXhz+NMD0
8UKf+Eyzvrz63Qt19XyVFDQ4Zu0OWOsxKijlte4q8RzHVz7Og5KmVizn++WyqZuebnR6mqeBD6Iq
jqOZUrKpYH/7u608f1FdzwTYww/Kvht8vQfv32vcFsyvTFeIS4QSR95YNIPfIWbsCIS6diWgTfTg
PS4eFirQnJGT4kSYSGlyZ6obDfupfwyrVu9LorYndQyq9rF2qqXpkKGe23Q1+OPOTsvpBgBFANW9
x3hfOIlQG/qt4+tJ05sIZEyBeC52FnTW46nqNQgozKQ3fA4RSGkQfZWUFX2hMvNIYe8Qb8C+5xkh
+ausYlaMqBv8vh3k04uZl5s9GIOH8E2EPYZRzJ8uIcrNbRV/KbBDpXOIOys/W/DwbiavmmOBrTqB
Z0jlVUzkMe8U8KQpHbhVx6gz03bGaxTF1ZcxbGDi+sPH9/pYFUXvyHk6WZnGdABE2gQy7hdCe7Rj
G28P8ot38Fsh77/WhmV3MBJI8BwEDwCc+SuzY9NCCU3lzoo63zTPALnTyH4rJ7KXpA0Ca1+L7+qZ
H9aUjtzYt02MGYO271xksLRU1VfRbw70Ou5otndLmi22Vo4S0e4Nucop+fwUzIryTNArpk3wRRcJ
g/58kIzcYIaCO1CxHcI+wtC/bNpYPhRlPNRYa9laVGEcmSB83qCuq53W59HpdVFgfxeBrbcU1PF8
/6PMxnxP5R1WPrjKHvcF0moVmwsFEh3OYEvwDj57KeSWhJtdfmvt4LcXmNlnMaxdOAFsFW+waWSi
Wgtrv7AQUVAyRre7kazw1mUH/6pvKf00Fydzl0ONvJctjsG+nxEDsx2/amI1KUPIGMNdsQsCMwS1
tik7paYpDes+UEcnOCUQmeVGWjLYGVYei5jKiVc92jc6eiWQz6hWndjx1iI5FxtzH45J8fY7f9j4
2nN1Aj8ranBFqiK0O3ZxxWRBrZ/rLxgLO/ojhNN/2ZxD7ia0Suj4mzWKsT9oIvEmvkY9ScAlnWKU
5EjjLSHl7sUDDCRsiR1cOLd+xK9h9dMM9vyNi3QdlgOhPcroNbV3bI9UbRBD+9ChTfYLLU3/+2tf
17RWA9V/NIJHU7+gyP5Bk59/rDogAMVrqP/vOLZ/pmx9Qr9edD/pEBOD5jzoNNfbFzmwi8nQZI1v
42tskqbwnsSfhYFuuJLy2RmqebMXULmgv5wfIlYva0uh0znaeGVcdAPL6RzfaF1mdXclY1pS+eWa
H9iArwOei0lD2ZJieZQClafSuppahDrg5NEHN31Yrdw8m5JRSJlqFcYraEoaOHD4JlVboIvSMe/2
umpTIwaqxGC124bfWk1QJkv0EVZ/e7Q03G5x0SX9K4npRluk4d+9jv5DY4Utp079KAlCzXmVVq1H
3fo2zBHDfTJCyz42PCoZascifnRLw39usH87C30LLBxypIpZtdwmjSii2F+DbFsa4fh4cNJ0OX7l
NPYkJfIyR+tfEB+TnqCUOUl0FSsIiD2CPe5MDzECrFsfpMpnpN21XH1IY1T+H3fBGMUyQLUsw8k9
Y7Bq1PlT+ngErI8vqEUxT6yMZZnyX6SWWjjuNmEShv9yKYn5gVK3rSDcPhhmo5JjUVvORFrmcN8m
1Gm/i5LfUsp9cIL+tPR2WyHqkQbAMYnX2rHdv6KYG2n7V+igSxJg1rHNlyJEe1FTsZlJEs6B36+T
Ar/h80xMNhfUxNcu1HKHAa1x+pcffWIqoJ6jloUrDfyZhdlZXCqiwqpPQDsn/RlbFg1G4YMWe7YP
Rmk5Y65l6DOWcqw6XRpTPAhf3x1Pcc9KYKgVvx6QuERe2SySjrq/iFl42yX/qpUe8JNKJHDygKSV
rKsJ505l/5W/9Kn2oc57NMeGnscDZOtz93ymSFv26vXHpC0tpPkD4JxX038vCRknDoH6Wyhy7bja
h1v1IkAidw5RpFu8iS4W5Y2UwBKc+NuQoL7MGusWPtueb5EhaUfYoTpqM8XXo1gPXlZAgDbBTbT9
JXTJT7q9DFNjWMxY9XcsV++MbuAe0bD7eajsYMWZnRTY6eVKemJ+nwQwfO5DuSgPGqGVIptRfnEp
H3sRfAwj12JhOiV8qyXmA6kI9V8Fii0liDOiFIGtqSpJG4OyQxXg1uYkZCC4EOL1d/VzSziW74bs
12EqD1hO9FZsdD2n1G0jiYn1qBnVXLbN05ZkEXEx2p7uQU7UueijhofqxnbVhsDW9W4DoCPxGalP
tPrXtdB/7KaQOvpEQkMr1eBafjH2YU+e3T0hEWSnbkoZLL8LGVKlDLXhsFsqvTb6hgaadudW1fmF
Im6t1eOg84jcU8qbR8EAmfw1YzAlJmWkPavf06x9p3/vko/vwCSLsUPJXub1UvqI7+kLWH7i5Yl2
XuDtk8IFnpj4y6x61Uw6MHMEAs+adc9hBuhxziHdknGxg3JePzjm7CsYGcsyFXBnOQ8G3US4n9jk
slCyK+w4i+7dSUuW5JEsobPsI+DG8D5U32vmPRB5xu5fdyX6XJI+z9MIhRUpdHIzyXXNADh7kVjx
IvdE+uJpTJScGlNXmVpCUsAYG18sCvVD1w/JV2SvzjDD54v+WVLfktTcwsi14gNQwkKPHMJMlFHM
3eNPRke0E8W9fRH5KxadzXU5YlZOg5DkIU/qzcJlL4kFEZ8YFkW0YE+M9WsCjvLtvIfTLB6pgS8f
ejUn1ykRerBXWuPVC0BDb8Jbo4dlslZm83pkW01aTi1fAf9/QxSL/nyPyHwSJ/B8B5/2a5RjeXfJ
/MsnepdckhaaMvegpjBdFUhd46MjJYSGbT8xAVkVOOI9nCs6KS01Gswis8qvj8IcGSwK1IpwavAy
2t/H/eDbfbTXQtri3o/PhEMKr48aGokEcJfxwqfIz8+sCenI5RcWoIn4hpdAJJG+0C2dHa2juGUx
P8MnBhc9pLRn9uk9flBgZsoOGCeTwSooyYR6dveS/p24Zx8EM62H9oreLyLAgDBGepA+Mlqv5G7s
06DvPe5ARVpaSih6S34lz835VYS+q8JOZIW/6BOtKEjs2E7rLmC/XQ2nW7HeJwbBEP8DVku8mX96
7kAL0QE1+FTrgjF9LFanfWwIwZqEOWBF8uCgpr+Pr+ek3aBDmm7KEDmp7DnZi65zPjlBGvlwXmnA
f2ippcHv/TDylUEz2p1U89YTmoDtUp1EbBLGZGbc2BUnVYezSandIIzpgya8Zy6pQG47ZoywRUdI
aZHkbrPPh0AP5qk/GrOti2PBNAGOZoX6ewvESIXWbuWlWdEcLKuolU5m5yuk2yaKWSmeTmKci8s2
X83kb2bdADaDIXLqFKeGeFseiI4dzX06lso+WVTqy4QBWB5bA8Jyg/3ozSNzz5IvHeQo5Z03ni4E
lg0noSgxmAtpLVTRVKAvhvKEiH9Ty7Kz66CEMIoHdZ+mhCSQDIrwlfKIzf25rhlxbyCIneZwJxkY
/5WCBsFhFlHrwAEJGubISrdf9YLC+/owwroeUBeUvr0zo4qZGAnP3GqqJ0sbZFD53j487Z9iwoAT
Ni47V5funZwY4opTwMT5+dHd3r9q7BouzLBdva688YewXHkVnRY2WTBogyEK8WUmEoF5SYEPZ6S7
fTLd+d+Fa7fUAyPB05ay5Hv55MQMHHLfssghqsya8nyzIZLR1pXW13hDooIs/HjplKtKPyTLlKRf
ACRAEkHpmUiDoB6hLiZ08n6OHLc0v/O8uA8issni3cuAKNdSRRalQrOqxNjnuZtK0O9cr6Ofpcg9
J1BVMeI7Hw9V2FKuTsqBYsyX8JRaG7/OgGPYaNa188o3jxaWgA3o7Xft3vpv/zmT2W37djzWyMCm
sOB/0sbAtlgzwMM5Bd3gHQ08wP3cQBrvFKPh3d0t0RKBAbgB8RJIB67xhxBim49R9oTUOg+z4pKC
qnuHHn/nZ8wY6+NiwBKHrhxtr1IUFD7zcSxi2OcILocquVbb9ngjAYcOEE77xjuQu3x3v5PKxagE
YWREWO14O3Hw4AFofI5ClA2GJClvXZzpoVrbNF9qnJk+FmncHxQvuRyotor2igLQsj6n7oCB4tDe
Ub6ucUGvk/yze4SchfyGQ5QkvCgkj4ae1xP0sVo1MsMRz+5L7k2GWOx9lQdpnAWFAYmnHpZVg8oy
6mWg8VxGgE55NjeutNyQbLEXvL5J5+tFuKy4UliVOO4mqyxA9ucArVLh9HY3E0spz0nK332y7Zny
y5+BfrbJPSwsv0GBDHtLNPnXr//GzMDOo9bD0zlJJ3h0BWFNvQJxM0HBnbLZtZTtUDNHMc222EDz
77DW39l3FJC381tJWyAiJPLRPGXvdYo5IpDcaz61udIfYJKOJqyUb0NiygzzfkodwmZZmM38U1ZV
C/bl8iPpIJTCtG0skwHrUlbKW7PxZe3YoJrDBnYIMXVSFIaybeo1DxzFuJV7izOqeLdu74pGznqG
kfA8nQkB0FA5dhcZmPL4w1nhff2C0UJUaO42NMAwjCRwN1g82eKHuH7AdMehlEuCyV+anLteVj2m
KUIHKQHfqaZpNC5ZG0zkq9ORE+sy7fXsLhvyQ2+lSTTCmnxTUNCyb9WTv50RSnBadlsK6sv8hwDG
Xg+XvdBN+ZrRRofdMBo7U5ziPtAYNSziQSb0wwfivgD/bzf8ZYDgQKMwpbgJfNkzs89bu/hV/UeX
72Qm4jsTRkgXXyF60QLMuKL7Mi4WdQzUyZIwNyphAWHZJWoj+sAp4/L9WdbTbLStiD8TQbk9JUcN
iRRSaZ9jxXz15vjC9AhbAcngWeI4eA32UFHi33pcsqG6d86q8gOnNCMQMY8GR9NXGTA8A+FgT3q6
+Zy5UGd1wtheUNKGkVALiIaw+hNGJTy1Fl//brlfqklaL0DyxdvVUiTWzTTF2+67NPPbrtAETBAy
/CSmQ+BJIgEd6IV8x0hbiC8Gxih4fq1KVyNa5IzMt6qIs0yLLM65BWYWSFqd6GBn4WU1e7UM0+V4
A+lYSzh4r6JaMIWP3z42RLpwd6CpunnJLE13pbKXY/A1LqWUTmeV7VVRp6SXj+1A4HZaPU4fQbFZ
5h07/dDQ0E97Itl0zf9cC5bLCxtD0lDYhNs8Jz6aP4xP7NrxMswo9Yd1TB8KYxpaYYwSsUS6tn5j
uw8AyyUXsjMTzJF7PsMXNm8TvR5EruciKcTcWCd80/f0IcvTztqnUe/ZxQ4Hr47YA/B1i0kEm5kO
R7qwHXErk6zHWjxQ+T679FCXx71jAn80darhLwJrk063hlS5XuaoYpAp1kfRTXPiFavzcR5RCbrb
yXpxRtv+h+7UvINGGyXdUoR/KhVFmLLLbfh9McaMQ68RkwNjpiLtDoFbtn8dvt70yD/i8ToI+jT+
zTrClO2ySibTc8CpInNhEVuG5geCN2SXbLGf5eE6iy32CAdJphxrPm/4dJMuv8pxp8rOnUraFUMg
in+GfZJwnA7mdEIhF/ud8XoFLfvuJmodHZgQpBQeCIK5Jnymu17iLLPb1hlbAEUis4EUNQVFr2VN
nk5oJnRlAsUht3TjOdeg2Hm+boumId6R4w7i7Wik2EohTGWZ7LROzDLXSe0AfcLCcWHvoPBF3Dy8
bHorImyNdsfSU5wKv/wa+be2VkIKrJz2YSEK1ZAtPW2mEJVvLB6M0hwcLiZrfevTK0+FQ8nlODew
Vt6jJ7/j5ufHsSAre85T5VU5CiBZvs7u0a5GGOLmgXXH/xaQogV3yvzy7yo47kRtAV8iI822TSuK
mm2elQ6BBFBGuLk7AHRoTEdzFJtB6aBOXhu9r41G28ukkt7e2K1cgM/zAfWJbYGqeDw2kQUiz02b
Gvt+8kT2likrKm7w6kmneVbdfD9j8Q9np+R38OBvA/Lh0SzwNg3EvwSToBsves4GPJwFsWVHYqyq
dILUa+CbDQWocy2DAuElvHEhmHggr50KR7yYl7yTarwinwwedGeBTkx89UzlknO77sKZ+QjgPwNM
02hkPBYyw6nbO8XK5gaUHvZBscVGwram977lZc3U9Q6ycIdu6oxR+Qn4m+bTsr6nX9OdOrLPagb/
f8cosRvcjIipvOXtKIqq4hlmIcUSmVtccauISn18nOptSStkV/XFM8P+kbDoYMmKkL97zpdzO+1h
BhO3aNZUU0HGvtUX4hbjcWIIMeEUcjkCP9VjIoyvYPKlMXCyJCx82AQaE3zdpg/u9E6rSYlDNpO9
haRzoRH6xLQBkbXjxNSZOm5oelZxYcf6VO9cWBEgmCFPP4XGifY/RcVPOXiBTBzCxqnOT4UdRbRP
cE9EyBAmiKsnah646e6aDaktJedH2dfuYCS1KI2HJJDwWiGw34Z4ZzK9ItWkTvZUJnUnRD6v1o6q
Y5UtkWuz6cSAWmXcjdGU2vX0NaNTpnjELKswBJ2ANMKRhuUw44BN6qMQB10NOo3TtYlFhz9Ign/P
AOySf5/hURgN5wNAnoXePpkHMr9KNpdGgVEU7DIh+JOPUzJkuZ99Ye7rzXjMzzA4vtynFIYaisxA
zkPJRQoyMj+x6a/iD+b2gU7MaxnBCUTxBS233C7N9fepYtcXoN8OK7JASVLFpIdD2iepQ0KA6r+5
/WUg8bfsnjRhY8xKQL4II2zj6Rf9bWsFKnIuA8Nzl3mufhZAirdMFAzx+BrkJt8FpPSK3cvdjRCe
fTU0VqRGT+b7d/4OQlEH1sN7P+KoYZ27/iCXtFsDei7dUviKQmQLKr3CL8yu6W/DylfgDyVJC76I
XljsjIvCWwGx/SH6d7ht6gqsmx/rbJC/qwsqlQInEyi6MxN+LbxqLA9GdMqJPw9xVTjVpcB2Olwe
iG3R5B3QAeYEtLYbN5xku9J0rLxliG0TSVHe5gXLGxpG+C8ULjSonzuDsWDKPo3T8OZCZ88EqN0E
D3f0JK9Q8k9nPgZK7D0lVc8IX4G/0GB1OOPQYW4ZqnVNhkALyCUh0HdKT/ZXYgxwgdBcsGMJD0xN
pgOukVc6tlzaTejFpFKyAtS5mpnaw2sjoqUj08NZV6fzqOoJFGimJE8aZgWigXH5HSg9OWhi3LQn
HNdA11m58YtCD0+go2oE0HOGT7rhjDxZ/5IGXYzFZp0fRD8tCchpIZcVzLOQHhwYW82tRg93DGpk
cr4GmFlfPfau1zlJp2FdX7y9p81nWLB/MGTS6wGi13LFBppDrUqKYu/u5EDgMypEme5o+1IdK7B/
nYLNOJMBCr6SysHQoqP5GD61E2YLgLUuEY9WE3szzUTwkoGVRhOz01yWhPGaMOPtjyEE0G4yG7l9
Bbob1jrfJR0w/owggF6oGI8gn9fj2yq4kkxZAKNRxBfd3OEIv1r5jIL5pNlfAVYAaf67LCa96Ysp
egV/lKyFt+KcvYUHbwzyH5FkR9QqGXcAQvWzeVJkCL6AdR8dlNOsBGBSfdEF+WEAbIcsRVHdR0Pb
uymHdHTnLBhVgk7lJ+3V/Bewca/BAFeB5lajBWHddTMU9Kn+3cCxk6mtC9X+mqtcqXAojKjMJ7/g
jsJ6ucD8RewkRl8hUb+kk76WD1Uw9i2fnO1s8ynLyK8+TtqW6oNtNN0qb172HdHb5ZY248a26h1j
ScMo0FgzDoK8OHBUEiSl7eFsvJj0FVJuqLKOdDhqws2cNZbE6G+SYnjzCCFWs4Q6gg9apa8tdn6c
yFtbqUX7/3BztWf3QXuoYPh44ponsLYhHh77Csi/cwBWhZnULFdC4z6IDBDpp1etfJjUjCuLM155
hgQiXLlnmmt6yi0ZZldDTjpNXQfVy5c0Wl41qSFStq5ZqeDpLaFhUDGL5FuXklHAxw1jHbvp0lZF
mWr+TX/2pR+862yjoSdZ41P2rDUrm/U45qR7iM5Qi5FJ0wTOlAt8tqJ8oMLB5JQQ6Cr6qZPZ+55r
vtHeBw9ZWUhGWI4wzz+3TbIyTg4ZFNB7qLu3vZTEU/946QSEbRhiC9rsNn8n88qBe4jdD35+lOye
ZmuPJkap8ZzfKjd+ydEaSnolvFLbXIHXetjdJOUUcoLOppoTtP+WUbhupddLEtW2xRdQ4XkGo/lF
xnR5Mb7GB+BaY2pTCa5PsFcL0ekhQYlrsS+z6If93/wnBNyXRYCAGcYWYQojzHFHYiBusXNj8wmy
W0ylSI7cBqwd7+5Mo6CNAk38SGdigJOo6CGoQoTQ7wJLxWHrKXCI+b8KilmzzGHXs3p92SyyJiYs
QsPACR8rHxD8Djr2VW3M7BVAOvKZDFSzsR+6m2XSJ2PKo0BfSF7+izYnpz7RPgvuZpmWWGuQozEP
vSE7GVbwlUGvwfjs2PYLZU1LKtc8wPA33KX89voWuGU9S4cqVnlXbLA14RUh5h/n0kY1yp5SyPDu
JJDxtub5J0t8lbhDQ4KBUx8jbSQadZifvU+F/CqyrEDSam3k30nCra4zIETfg/OGqwAN8fvxt/7r
P3HqpYKp639cuYK/jiEY5wgVy7WmDamlpt4k0iKUmn5YS269Ls4WuebQRsGVUqtDDrnKaC0nOR85
ME+XoQp+u6IVVSy1DVwwY5+0L7VUgevKxzD4FJs1dR76YrzE9mPeK3h67Ejlp7gTXBoxrxhNpMyn
AmC9qne+H2fckT9IbRIwdbAML+4jAdBMjIjZBxpS3uOi/WhWvpjFBj1/BUB3gKHUH2/lprUMCHYM
FDHfsYuzH7N4T9HFFaBimuFNfUR8Crt23nUBmesJrEU4M7ch5hHOhwC/lMnWWIG+/jxEftaESBCa
CJ+lerjhqMva49UDDjGc+RYRbxAJkV9YicbN5bB3vP7ADvBKTpnNME53qzDv3UYDGQAEylKzpOna
1vb5dlrtWdi2DBYNLhvmqqcZBJep5c3NERy5KALf3Fmq0yJe78IcoU57nvKxAr/lJ1vHrLFRr5cS
NED2x+v0KVspb4Q7t6mJsstGzSHHka0TQuZ1fq0TT67rWegBj6ZQ54wSiludTURXDx3y6fBV+VAU
oItf4evFm6uTne76+cHOhJ935wOwugiajDRKJ0PoASzL7sumEiP+wcKqq4cDWqxbA+el6sUv98eN
Eg3jmgaUkbxqLi9lqhdREn0Xe6t4n7wAxSmsHhZc7e53u9/Rk4Xr/oob+AC+lRkbDMwrtCgmMcgG
z9LX/F4Y7KBABRGiFT+yAzfahO8MGAsxM5OLL9SqhSD2hF0OJJZ4LOrORA30TeeoYUdOFH9OIE+m
+Pko/qLsLoPdvOIo1QypU7Oa1Hn44G0rKMQQZk/yrHI0Tfc7DFr8XDpnTJ4W8yLajuHDga5C3UbO
4ak0O0xFfIwa0v7jPHa5XO8kIy2R2v2Le7vw/qP8+306GVtelYWoeBfH1NaYaWx40wRdGOOI7IZq
eMiXF/eloqrPzB71wFf4VNW+4Iq+L7t1XnrQXfweZiH+d/1UzXlc/f4elW0HCweCgy77+/Podsph
IvYAOeVGLAKh8vNaFWaocx2ZG39WEQlDWjmtFZPF72cvPi6ZLC9iRA92BPsr3+u1IstU187YXTDM
15hjXbbKc6w+XtrfEjXAJaQW70J8jamSa/VF+f447CXbxj0xv7HkZiEYLPoZmKCPpwHbQvcagjFx
LkdzgxZnlwQeM3xTe+siGT6qngYAy9xr1iPdzvh6AlQKkJjqFudvBS/hkmQRQ3E1e6gMrI+D0BAu
KI1y7aIcCp1SFrSSflpQqNmYe4o3MiNEeFtpTN+TPk138xaTHHDj7lpGaXWdfuwYEcCcwvtlWZlO
d2MSWHE6M+fVjLBheOzGiG9a34KOZeh8wgtp2qvy3xZWG8fYf7sXqcuCBefLkLkCL132MjllQ2hP
k2FhGkGCBp3M0JIPaxT8keqbneLSYortQDqy0hjxkFB5xIHkgRSlAKWKHPRPuXaCLK/ZsW7CdKJc
hKoEZ15F4HuKFWF0LmKr+rjsnAol6On4DgY7cZll0i3zddM4U3T9RHF7F/YXM17PQQHs5H+5rOfa
Fet8rLYSb77mgPKricPajRVjzdOLUvpIhCbuZgZP0p0wZLOB/kbZeZ5uZdR0xc/qZ5W0Di0HFdj/
F0IZKnLfN8FcAe0LwbdFLi213Y++J+XrYO86fXRV2oC/kfqM8nP6F/We2hj0AfLFiQbOM1wiTUof
64AUMWkIwnZtBPDgI1QB5p77bTLCa0A9vvSHfVXbQKawOU8E9L1i5U/S73rGa3sbz8IcUAVN9Orz
z8FM9oC3mVT2o9DUNH1IzhWjhpfKYBhW6do+YuVJap/vp3d43t04DhTLkq8OrbKobauygjNI/yL5
y1MGNqAM5mAgro52MaUhapgdng4RYZMlobYspuyk+qB7Vpdz9G29wzk7/IH8rlLRd6MlielZiLE2
p6eCMEPOpFQoXDCPKu0xeAnKs1t2SZQn/bJJYH2a8sk4G69UT+knymMNZ+xGlGmKn7ZFaO7Uwu8h
7igXq4+01zt+Dw3VYB0Fc9KvgMc6XCa/ACSOUruvxZy9adA2GAFADoNq8MmfapV1IY6hA6/7T5mZ
us2iqCcHVXwmfwRxFPj5y9ouBNHk9QpoIBTStss8Ufo3IC19LuARLpEL1QiKnFwvuJMTS0a/cEXo
u48ZARJbh9T/Fjg1TbR9Zt1dSnGiPy98qwR/QXmR4e05CQf1EDKySfIdD15vjbM5LGcH1NWpn5l2
6SQd5krfL+PaEyltx8Qs5EzOpM6RHhzro+cZJCDuWhPABCLPvbpgDElPYJ4nH5nakoGZ4Nbimhs0
QQF0k3Gn3iWRxdlTLCM46DhPOKyiaWyhmqAlKJ9oLM2325+TtPpz5RNVonBRP/XiaJTQyutPTvH/
dA1VfGyCLcmWCwSDMlba0vrL+1pYR3CYBMnyt+EJjn282UtPtWIu/wBaKADD3/5wh8RY2ob2B/IS
7R+f3Hln6m8e5xSr9GM9P4SUb24NTyEz+6AlRwm18SZHh3qVcpTF8CQapOt61c0bBFK4H6YHjz5h
tcBaG2T4Ktep8N+erm8VMlVp/jTQ4RMNd1rwfr0Z9PMOsrl7RqXh15KyiPCpUE6lN7RuFr6K49n4
/IV1E14K9HrNUGGgPPmdAg86+FFQzSUaswJnOkDC2O8RnrZSyJQnzeP2TrMlRbEeLnepV/i6QtNN
mZ+PYS3JKUbk2z855eVLWmbx8L/KUSyTbmQC1Tv7oKLwag5N+D9iEkf1ZvZdIopq6nE/sRkEay67
FI6Rvavyjm0DVqvsu1Eq94N0i2TNlqBCm+L4iH0CopVByu8n6bcjSOLV4fAbOZRoyDGdMCi0YzX7
1+kx7EI1S0QGEtR4KrY8rThRYzsM3KyydOj6UjEUosZYLdzum+LHEBHwITdtHwwK6pLBYaoSrzq3
VxDYuIIOFdNOiL4CFh63MdJvhktWdFKgDU7lll8gs1V5WplfpAQ+X/zf9WBaPtUhWaP571RYIEJH
FeF17ciM9b8sz1MJK1A5BA+bCXMZQLmqypU8GrlDb6F4e8m8xirZpxDD1d8LN9bVcqazNa0mxSpz
2NVoiloBqI1CEnQ+dkoW74On7q0DkfgPf51hLqbmmk5aOlTcljWxLUyk9JlFkPqliwV3nREqVq2v
3sUn/bdhTiNPjTU1ak45B1F4UeGK4GO8BJ6Hh4XK8Rq8ikt/VOf+o8EQd4QALo27Wz7jaC7tN74k
i9FYAaMW2j1/p69RzMY75oV4kXKQ1mBq0lMwEfKcvUpdoWLQWklMGN+cdIfKQTim4Vp0lsVU2COa
8nEXPJBUraTiwET6l+YJboPWL6tzWWDe6PrIKFhS5Zk0Zg3AjprvSsF0xh038zDm0dmmds/FQTrn
a+OWLWcYZ0Svp9GxjiG3UeXUhTwLa/pd3iYegA3XIcniC+o0dWmtsyrMRIUYO7KWnqNXhvQrxz2y
rE8GFK+fQBwQmwuLyQz44ERChRCWP4bGwXcV0O7K4QCnupTY18mIEpnB2MAEoX96V6D9ogbnRnK1
Z1BvtvQXsmnLH7+eSRg0mGGKeExlYyY4xqeoZFeoU1XNLBWwxqZ8KSLBg1a7dkSnwuIl2UI2SB9U
YyplVB+Z7sG+HGjsLoMOWkLoy2z/nEbn2rJ5eE8dJr8qyoUuRYdILGORyx2lKjquCy90CG5HS2E6
x4ROubfEUOzmxoHXFIJ5ld/BF6trhbsLp/oE+/0EXlCIot3Z1aypi34ZoeE+jjNC4MoxXhxUVkRp
65fh/nh3Kn/mpVXRfcouRX8iGE+3fxbCtVaPizStmxxBsDikIt035jjTWuTC3sWtRDbXqSXgbUcT
Vmgqp5wuF5/NDOrsGSHNk1xv1boXLv9fHyxdu9OSQE3kG7sekp1iMii5KUmrjEslYIjURdpIA8i2
Sx8pyfuBXMFvovvtOcWgwSG0/YJenXJQxfe1+m+ymVbSGsk+smZs44fnKrEUTDicQgnFGPW7A6ew
vz5Y8lf+frigFuThrCSJ8B9Eocmk9LwuVVUOeP7OZhiH1w+l+mLj11ek00QkPrZD7bqPzLbLmUuB
At4Tc7xt82bUUR4peIa3JrFOx8V9nVzlyuL2oTWS5+ma+vpBj1VgUcZS7/fDZzX73R7CykAO7utm
SXONs2MblLaZNCLXcjqU6XLpldpbzwHSdi5q3VcLqMAnL4/PW3TBKijMYV9v9fJsruAmZHFP9UYf
VaCTSnV6fRHPMAiR0JcyFLAMZ3cmVT4lYFOFmucBbfw6O1nnk/s1Rd4Kbkfl/vtovRxyr01YIEnG
y1YqRRCn4shJGlIngfq0rl322UpK3iGysQRAVpzJAWCaLsctrSUZ6LFhCCu18Fp9GpUNiDRchPJz
Lx5bluiN5p8JlWud39iftAtFf+aIMNgwAuewXpC31YXqEn1ylTtDNdgQqvi0i9PKOyYWXH483sMo
fDtPNkzbLYScWsXDmOPgfhcuZh9AgllB1CsbKO3IMuqUypIMpAomQwHC+/dqErXrFVmNKocqypbm
HVR5d+WI0hUP7y+QrvN0sZz1JpnWI+kuZWBloOCwRPO7RkvhmtwR1qb66vDyRLJJ6iiOhkkyoqZE
BSmmiWrkkSO+0fPl18tZuHEmemMwlPt07ezEgJNcQiJwt9cLsmq3XGgg4pSMM0i5/ocYSow5x4at
1ueFMPXPlRfBbvt1qozXCow0g+PtUW+y71QL/RlnHoWYW0HJIkYhpsMk81kfwDQTq4BYJUCluOsA
RNjaUtlv3bKPyXpVpU7ndwTP6Oo5v0By07t+e0iYMaqobaASMi6EiexCihm2QxaEVoYoc5L4H0lA
NyU0Tpop5iZ/LaElTgd8SWJWMnb0soMH6dhHEn5kMnROzzezD1j4tqAaMHqoe0u5pUw7E5W2GnVS
IWoO5gJJ0bGp4ephe9T5IQ4bBr9lGGamLjXtw/d2eyCVVHtRPyjENE43Uy7WxfS0c0jVCqOwhxJU
MBVc/OUbYWF3ArDjmTXrkQJEYHN25oH/kvJXw5JUhfRGMMS/Kq5MIHWgQH4JPMwnzK882MEAu0pi
Xaiygx9OH0zfPK8MbAPd5kIqb8eY4vDO81UMvPmpIB7QrE5qAE1ZFAFSt17PZNQPFJhpL0g8RD7y
dt8qdx/o3ewbdtGU9F45f5poM4SxSk2PXHTqblU5j5chdTM+2FEFrl6Zhifb+JkH2/3A3qBz3aMW
j4dbrObozx8EzuVowcX4RjX4623i9r2ov9S1Go163u6kgVW2NCl4jXs1MQEFBlDsvXX0PPqNtxvg
kwii3zLFD0aYoN41NDBCqSXdCB6QrqnIG47IPJrg+znnNWBhvGiX+GhDPrlvS6s/4hpxXBu7da21
qNd6cBLvRZwD4tZKonh1sxj6CX2eKYiBrMzkGyo8pSPonSJWjknlH6AZu4ioIbtGQV+j3ysAnfne
ljl5VQ9i4pKXIw+25s+3IlGBgfzWNuFbw+Xk57atqIu3G7QiSSoPihZoTwqtA0OFWlAB4av6Fs4o
kC/xuCjE69TbYp14U6luCpbNrK6muzVOjqm9usut0uV2gUSi+bAJWtN/DVoxDtD2MRXRpu2oC9xB
3MRL8GMqeZXjvsGFXHMM5ywB0YV/ENIDIubQjYc0Ig5ZbMLRAVv2Us27NzoN/sG95HJUIozqmyiU
sTCnowDurOfWodvs3ODIwaMmf5gJToxQGekdsvK+hVk0j0DOjFQV6nDHQSnsYKRjvAESuW0E5cAe
eTUwJPAzQHCvA2miGrsNUhYvW3+5rDr46Sen+6urWz39cq5wBStHRHeqDqmSqFW4hhi56ejPBRBk
r5C/ZueDKhxT82KBkqyWtxjUcvNJBuaufR/PcXxgiIPoY2AukINDRcAJGAJruMFpjDdNJuC8mtmN
qqINGlx27JNwBmP0r4rWiJcY3XRv3h+PwjHVCwapLHa9+a7TnnMr9DxkVtZuGLgUkcoQWni9a0F+
okFb51iQ/4f1Ib/TEP5GC5l+u//aT5pVPBRlt5yHaRdsUgbWuYIrz40qN+5G5RtB+W7kfQ77NsKc
H3xW/yG6I09F3zFDJVf7NVCaht5TncB9YjmqivW1U2nMt8eAbT2Vz/Na0iHjCIyU6niitmsFsg0X
2uiLydywROlGWcT1ZQXr2bb2BHnf6TtQGaX/pLESlpE3IjeSuBtJS5yfG0BruxwXTNb7brE2+oyH
JhIHSq5m481TFHcnUFyzihbg0JOjPFEFzn5vQP2g66E98jZ1SaxB8Jr5Hz6DL6YaDZMQGKwOGlna
Q5uyOSuVLK39PRNpVuUlqWDFFSYOAAYNQ7gsXoXM+fdGlKGOmR2H4WLna+vK1a2/yVNxlSAQXMVU
2g0h7Km0P0TZSnTlexN6pYg6+D7m+vxStpyE3PbaSeJSkwauX3vrfqRr4sBtF/0OAY3V+DeLz8Yo
Y78EmRmeZjvgXHLdP8SzUGNB7Uql8PbZBqjB626scaXz/fXhtzgzlIvlG7zZlTe7K5oGNFwZLQmi
PX0uTmNTefuEwNHU2tcgjz3ARfaNA/snbOmGNX9XutyiimWHhU7kn7/oNGU2nM9i9xxET9NOozvt
omyA5BMOScmEQwqlMallGqUCAE9IfZ+2Aw7C+DXGKmL3Sapnpd82uVdSg4/sIrD4y0Qz6J2BKvps
VaHcQz+KyfjCUcpovbS2vzjklv8ZGLMzaUMOcMBzljCsYtVc6IsQ1UHLVx4fhNiK8uDTNp72NOxw
pwQjvkRKtuEKvStPwS6bRDrcIHGNylykW/1KClkB0Rn4H1cizOw8rFFZ0H30Ns4riRdB+MAmZBUU
YwOggbtBzUAW2DrdWo3oR/zLoydV0XatnpNGt4WGKBpE+puVxNDCZCdiLO1bHsS3sIVZZISmQKHz
oDGpOFKW+dcU+MroT4YTU7AJLEWeVTfTkG7857CBx/7cxgTrZ8dO8+CJnCdmdJj9ISZQovprFm8w
HPMMX0xfau4+ms5WKVVhCv3yFUnPpK0bWnWh86Axipb+8rsmL+6JC7F/VbpgsEjQdcIYpFixtbY4
HJ330FELxRBOLw022w3W5jFpGYw0HRxl6mzitjxp+c/ewMKCmIvr8iBHMBXubv4vRjiFPkocfCpC
kxKdGNFOC5T/uNVaP4SJEXk5j1R1Ni9At13ITDZ4oupfcFFwP2x4vAnB4ZID94W4qQGEO/71Pa5W
jIx/pCpHaS6+dm0TDenWVGnPoYL7nbSer+7rfLpvQSZAox4RcuCRp51ZVD7UEMFzhzUFUFZYvCvh
LaMoTUqLgigPxL534x16Yw1B3u5ZY4oJZ9QEkx0bC0lm2E5bdGsUFXTY+FY40LB7sjww4+8AuWiR
Elj8evXu8i6xXX9N+5WELQ89zyu2dtUqmi/OEA/MSU2spucdh5Ad24xCitAllvHXntBrUA501J9l
aWW76elKDdKEEIroyKjnoHkHaqkiTYNqfJH0JG5CRr3Uo6ug1WQFDmlXnkdI3DkLbaxUS3looQtM
zuFbS0ySqops7qsjlc9GOV1RMnzkyHa2SSjCE1yYWJES7x7fd2OAN2Xwm+7UBok+SQK/8i1DhTlF
BnY67GbDpM0V4gA8lpQT/HU4ZXuk2IHWF0lJCA0D5JY3HUyRc1UyXOSHcpLMhgrUqT0QWma85Bo7
xvRSJBkqn7p1YVKPxATcA7fohXMYA2efZSkSF6KPN6i4dvb2nwsP5EeQWcol0PX1uyclGzP833PN
KNqAd5lZ4Zioiy3wWQ+APwRvIrOC2I2xmgLZNjCSJg3KuxIdyJxPcXTxVdsoM8RzujfkBsm6SfW3
eGWDPrhSccRIIc2BLRNkxYfsVGPcrNCdN/v8KKxQrWjsVxIlF+ATdIt3LKCK09FlO9Zggm4xWrzP
oNUODKlVAEAA9fuqUXhgZU0+BKpDVyWPwgb6hKSIFTogJHCwxtg5hx17QFqkapXc4CX74XEoiNt/
u2pLWFKf4VrHvaKo1adWQJYfUlT5W7dC5ACfNRn6DTRYwHwRapnaWMBTKgbIC9OHq0R1oflvvUxk
kB46JMq90avTVcI4UA3nKK5fKnHmYZVFAqjJtdnsZw3HPPV14ZFv6sF2Rm5QktwODqRJ2xNyWgpS
z20no5FhO3qRjiHAI6zTFwzso/Ud2cL0ZrCvIW76oM6yZPdai9TjeNgXRYdb0CJdB2g3jsq9YiRL
olg7LsEh6iiANvcSkSpOdsJbdm2FtPWU7K6L0QkRrgLjW+TmmM1atROvig7nlqgVDJMsj6CuWZoO
Iqxp3XhbKznOv7bQ1wNPumTto4io+RlEU8MShrzuAy6SWSjK2R1+cNHu3C3nIZ14nqUya0uvUUg2
C/oBTOkqoE7FcZXy4s6hHBSAR3ALIx8nI/SRteBvii+p95sj+Ivda0ulBuh47g9gSpZt7f9X5SJL
fUv21YkmsaKxpeTzY4wPS/m9rVcIPuf3gJ1nee+4WG8Us0jSh4htA9zPEFYu
`pragma protect end_protected
