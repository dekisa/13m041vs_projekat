// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
PGZvPdJxvHqkAAJVNRs3Zsx6zjUFPq/f27jXve/JnU4h89duRHPRdJ4HI8QqQHOTEqQtvuUBI3MP
qczjEygCHUg0RInMqhW+hVLJE4Chuk+qhDkJ9DQJrbJAyHAAQZnq/pfQuCM92y3Y0eCMcpwWC1X2
vcXP/NtAgWGycNZEytKKY8pbFENwCPZbAsFrNhufg+MO8vd5FzF8mBhAH8wfs2qzGx/btZBzfhgA
IZOH1vjkOlLTwpIhIuTRuA0DhBW6UGpnl2Op3ZzZFN6DK74trsifoZOn+RYS9VfxMXC6KXLpD+mh
dhN/L1B2kTAWXQCJwNg2rNtSde7kZarqWptxxQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 124688)
Av3+ilRAAGuhODXYvnUPXSYVqIyyCpNk7EQWEobPF/bVLEdryQhzzHJuf6QKdRUOtbpQeYGQtAOw
nv8FzNmtEmB1NemUakqk/99pe8eT/KnD7Bj380kKTEN0xb/K4/wZOo2crgy4f3vaymTJ/Lwnjgjb
AY09uchWt1ukQiOOoPzfFqhnITCNBQ9SAEvMJj68B4M0GM1quryLuHpJyoyIHkBqNgOsfp2LjyLq
b1jZbH/7GD759Ke3bCaOgODWf0/q+befDdOBuPiAtWHRXyJhvlwPpvisGqWUL+z05Ld4+NEdw9EI
1WNOwssMVc5mneNL6x0e50Kfok+wPl2rNSl8tSnH42jeqQ1i4W3XhkSBjqryWIpu3A8a3cOSML1P
fyA9YkyTUVEMHcW9roA69Jw0SEdxjwQmuW/dcjSedB1DIymJw/6FZtWzp1/g6/9AUbEyVfzevHj0
Lj805XshddGyenudcBVHNZ7WSQ9IY+N3xILW7fdSHYkzSzrQX9eeWvnkAI/DCU7FE4FcavBuSbkk
HmRFqtJUw3xTJPnZQ9EipG+6iUVkL7q7UhG6eL3jnjTBHXqEVRM6/ZnVFT0Be/UUj+X3xPPvHjRe
aq3aG1R8KLoAxUPgENmH1CFL7fITfuaDT8RykqSkKF4/gx4GllUALWVlAHLVlDBNWqvmJYWyWznd
mtZk0kNs8+1jK+p1IoaiJEyPZHEI1jBhrjL1nTfzGotQ9lfzt0QvFWAoPosmdSzjTYsMnnF0Xonw
nQFUMJKan8KT38cmy6eviG46yjumWnvpXFHQODBz8o8ZAspi6M2kjM7sAckhg9dvl2bsDpASQ6x+
J3FubrRHRNjv9raDb7EGwRg/b/K/HgXu9D49zbrDa007s40KlObYQlJHyCjIeu2bfD8rGmlOnyJ2
jio7Z81bpQclQYqTMSoeVDjFcqW1Ic2+AliFfHGMNNDORUxKV+QvYkc69QBirhXENcHSmXmSIQrR
TW9f9ylXAMXvcggr+GtLcEi4V3lSu7XLbUClUNsZtWHkptABaWHjlrY/+Dgwsucp9uAHFt+yTQ6n
4yOjyf5XxJZI7mbC3hmEl05n/Qz0Ma20mJ0J6gDJpugkcUgL8eFa9e6J1rPdzS/8u7ib6EVj7hQS
q++hekXLREyhksDezfdSYUz4+Wy63H5G/fL8M2+BIcjAOaBJju0004cgQ3Hc7eBEuN1qFDy7lC8I
uOjGyrsSz/gPaPpyCjztQP6442xb0RXWpR/kxauTAk/eDl+T2C2yuazmrbfvbwqJ6FeToSjwONAe
bkhdE8hng0mqwmTfYVlsVVjM/I3DA1hPGYQI1LcI6AIp7TQr0uu5SpWzfh2IkoEHG1cZ5AFujT7N
axCqYg30LtVL72LAKUHbxZu1Jx4JjPmFmpjlwrTgkphmCgWDjn5lsbdIeRLUwRfaF3WcGMyHRXGS
/MCZKQwhU6XbrBMvcwgR9+j7wi1Rtel4UM+8l6q6VgcuoEiDo4+ys0wtq4kK0p7pmSBFeuQxs3FD
rrtx/kW/awiOsQT91Xj95M7skUDF5ZC2stXgbk0XCCx69u1uQLoJ/qfUXb8tF39zy8VizNn+C1Cw
+DoOKdatwWUveq6MMOD0uAA9pkXYtbkEeRzv7EkIrEgfQGGSt/RzwB3zbkH/QW9b8OsygyEiAvGw
dDV3iBIB2eAHCFtUJrsJQSiFqlBCVbpAG/9VnUn1uNkXxkMkTPaZTMbvS+qMSzyhkBuTMf6Lg7Jf
bcsi/1RxM3vHCGe2akwkonKj5Z9lkQ+dFZLPxQRwd2irmtH8IAGQA3RKr+TLzMnTsxu4aUHRdhvP
h9GJpvenGxV0qHZWuPLTMhCbHu8FIrMDbGTOHWpEuLFBdFrc92m+3BwdLmRRnhZhdkVi9EZkVP4B
El+85hGorJ6NY2hTngWQw7cfISIRJPjhGNkFFpzunB1bDPEnbqrs+EIhdp5rmf1fpULy9MGQILvM
Vrx0G8IEKCRPb+yQJGoEmXHU9zc7dDjA29Eh+MFbjeNSJAKW+ua+r4xMOAPzra+8qr+OH7S5wq8l
+IJ5XC/0LM8Di6reN2p+fbOrz+5qA6uIz9nuYxaKW84wwjtOHdeAAEfM6Iid6We0w44dhPsoWIQg
/uzQFC/u02PgSIPNLapWw8XJt6iSVxQTRfx+JiMkNSdMJWrZWzImqKpMCHe20YiIcf6mT7x37Hg3
zSuBHm9mrPbcnoNxUyJKLW60Jy3KkmYVzmq1zrgv1Bl22hP6nGIBX7FnCfqIjHo6ghdYj72VlV/d
h9iLQ0s+a0GQe5/Nu+g2m2GJ0Ur/yx5u+CgmLZE/S715eeVbUH6oW+zdMqH6gLJBRMewDJTZuglk
m2BQVjXV/mtzX4QBTNaUZbiCANSENvZsB18MIaYa956ixsfJzePrDj/I/DoDqW5W+5QH2VoA4U8W
YjzFdhzBnZ5cdPy1sPDbXb0a5OfYrnGMgDFx+QXP0HtZDtkarZuyLEy+zB0qGUaTCYZehFSVoR0R
V4khgLQOYBcXPJciPWL+dVlgdTE29JVuhck9/mx41vkc5ny8Ca3SBUKX+qOJJ+4VlE7BxDSydCnR
6022HSHDIqRpvdqoHjJODfxVYqiegycJolfzCp8PA7mLMJnQvNnP/dY1qk6Pk5eSC5eMXzAwmcjw
FWH+aeI+tTHEJ5OOYj3oik7chKrF7a8jolh6qeZ13d+O19BuoYF3oN8IBWxCzDXtvPHEMNhtlptZ
zzdXGw2BxZrsqIWeBhA2aolgisEh5tg6RMBIl3XQIcRDcLO+x3wbZNfZ9DdfcpcPU4JxEEK35vd9
zOvliPPtlugz4vTrxyM+nKk3dMojfxZKUy1nXxmPv3r8RoBw54CQa7CLX0rEe9IecaHMuES94MIs
Rco5iB9otflPKKXGM9BKhjTamLNOAN2lPl6VU0Wvny9+cotW/gPYUxW4z30gd1p3baiS/kZ4OSfV
zF0NJ6E2N3TUBCXc9FB+ZSDeywAdkh0JZDY5UhFL1GihGpXUIYfvBbNtzlDpXaLU4wHKwsSdFbsq
+Pq2EPkcLo3L934guOfgcHyqKmLi4qJqDMoxYEODQkZfNuZ1+HYc5Ab1djGawsL1+h4Gc1XAMrKx
I3CuezrUNf81HxybB6JSk2i5GKslyz2VaE1aeqOcP+IW0MNhx9nLRkBCwLYB7J7vPUoEWaB91Z7C
Uli8CMQOq0N3EMTp5OXCVvj7xdmdU1m8QqIctsd+Wwwl0rJJcD0AJg8lKbNftxRnDdXMKDXwDWsF
IKRlhsov9F9zuk3GKLeBYVTco0wvR4o2hpZz8hHstAXy6veEbav4L5GQD/0EUBAaE43b2TMpFbMr
wLGc6t/XHYEv4Lyl9vAR7ktoZiabndXGXO4OXZkA2nkNuN6g/T2lt3R5v1qeyaVQL+6Dsj2BTGvS
Cn8uQ8fSeScey+Bz9qLUaepr2h03DrBS9avyqv2a/pp9QyCuOVH+kZS6qAiUsoQBYKE+WolnXIqM
OONDc5GFwU/G0D/YZTOyeLDDNxCkHaO/y7SylM24fBDseIZisojcncCqM6oliDk2C2a6rM5BdJZJ
UmzmrHcSntLhzIvKgG21Bdae37MqVtisg+Hrv0lZh/WkSx1WiLGRTO+9qAZXU6IQhL/jVyk+lWog
ByG3+QxIj983e2YCmzsjz2aDcwCP5BzryKD/XMzDM29yFb/TL3fYZWSJIUjtKaDDyTpy3zq/VR9X
tB4suncXAAHQiiEBZx9xIIRkfaqpbONEaF+1n+IJrOU0W3zJew4hIxyRIMNBrRITjtjbIrSiHp33
/HzAM73zVsp4jhwxzDpngB3BVwabn1eji2x6+XgBXVPXOHEz3GriiLrsgRIsmmybf2Wq1VcCqaBY
XBOdlNp/ma4rK8kZvh4wySrG9LQalxph5l4fJCOl7qhWZAo2SaBC9msNHn6xw9oQc1wkMLNpnAEL
cnYy9ycvmRbHOlhIdYuFmyJ+v90fp7k0CLCYYhKaH9pWLQIX530jPmrgWAEzRXDBbLZuKqOIsdxM
2S0hO0Cx1S5SCpFT104ct9SYrtwGyTrHBvoC97c74cEorViH5BnOPC8zPrKSkjeyGqPMLPALbXoW
UqGyTwrBzjAiOKA0kNqw079HpE3rrZzNG5UyCi+cfEHVqad+tz2NhUuarffY9Kvck5OxHqgpZuhg
t5+ri8EE9T6w5NNqv2T7h0WY2ngF82MIVBSIreXDIpSmr5Ii50kODb+iiok3hhXvUbofixKNnRGf
yJiRoPM3PsQAzxINDwdNYdf1PtriLxKdjwyLE9O1kZrD+VbnANoKd64csEYoH0sfJzXkuJLBJUSS
GMShZ+DTzs2RVu9GOMk13mfgcJXcOAhvxQnk7EwWDmEa/bXS3EEAihwNPTMYRsTu7xS0Ts8wX632
f5nyCV8EyRbIDVgZ9JqYAVPia1J4vR0BNgATVkRw934ZQQIKLmrjAImrBMLyXgAqRTeXt7p95atT
R/RE02SbMxqJJeAjk8xjdLjIAdwuh/WbxmkJNJE9/ObdDM0Ktxbim7B7k/D4C+H/Q0Esk5CpryW3
MGq6gcD/xt5Pbjo0TSU86SDU6u0AWgB9NRTCvgmXBG8X/fi4uprmXPuM7PErPzYEE3BeOoGNmY3N
5JH+D+iVPQLdTe2WZqvbL2fz6Xb6Lu+ShGewEIh9bmBrA9k84Yd3JXr4QEZcSSO74fmWjcF5I+8C
DGmGmZyswS2ekSGWPZR725SSvFVWvD9gXmG++xoTUQkj+mYXWkEUiK/oGbxEEY43KT05TCmuDdW3
Ou7C7rQOmw1m0FKtSHSTG+l/oo4YraFWmc0XXKlJqfIF8IO5clO5/+XEDA/X8hIURZFt2/3i4RmN
ii+xgzvwPngxleeQVbcIvR0qnrNKd9P9Gud9SrJ1nAonmZQEDVFNCDY41GBwT9tbixwgqjhO/Ihj
VwP4M1MJPVFVisnbsPcYvJsbfXdkiGtZFTaZQnxVuMcKX7wMwMBmPxt047H5d99K+op66hdGXOJu
tedym5rWPGnvMl2mQBrTY+tzxDqHoJsWeLkSN/WvaIZVFLxAHfdfgBiyH2YhfYMdMYvuYdVps37Y
uP0xG7YLAQ9yPdZi/s/PRiq+MF9VlhwF35yHPlGQagLv0QmqIPsp4ZZ8MsEk9gqpw4+HlWFLojNe
Ch7kNu4q2W6SqqPiEhZXJls1jdUv2JY4Wzk+8fQNYzvNeDNx3gULIZXuSZHem9vhAkNpDEmxJBgN
p/P7C+nyujXnzKcNs54vpNfm0DoR6B/Joc1R3l+THaGuD3B5RXMq/pd1E9Jn+SuhZzCvSxLEJxbf
lhTqPwANjXdL5wPWsHj2WVJWZt67g+tPF2IRE4ju2YML9Aw/7ZqEgNr6VN9BsLAzuezunsMXEFyW
Wnus2J5Lq8XE+v8jtk6QIHvS0aqFWyg18Br9uTiKmT4AYo6ylcg4jfjLwnAQWSNuK3NGf5z/AV+x
NwTNGelyAMPtrPHoteQez5X42U+MGcXvKtdktwkEqJlWRvPazkUbKs3kWoBdSaFkFxjm9bLH5foa
LGP8T9QD9f9YzAilOSIKJIXFIW0GehAJf1b3SoVmZmYfUcLMD8xsmkR5vP+H2k4yWazXSrZDYxkU
4IMUNLQizEzr6Elg59q6zJb1wJW/fow8brNPRAUSMj9keOgPGEyuAY0lzsLU2fAHCeIQOLC3xTzY
NoEylP5KgKU7bHLpFoPBHz6fSSPe1laQpJjCRnlN+YJRxSUp1Fa4w9NN4Gu2BhkkF1AHPGa6lGJG
csq4hnTHSbLXsnKmBLCo+7GooAVCUVpdSfyBgrUZBsBoLkC1poi/wOh6tDGWK4tlaqLFbP811Fpw
+ep70T7J/dDdr/I/LwmD11JekbG1HP/fsCUvT1J25IlCWEcbHruiNsK8jz6BfQniq800ujVD/CMv
xxjYPdsBeAHRk+a5M4Do7oNsNBFqaiB5Lo5FxYrn3oUIp8B7+olqQx+W/FnoGXgXFJKbgdTQE9vE
oYJ5ZteLvCNIzpfYVpLsa0qQ+8Y4Ju3bt4Byv3Raj96OHeTUF8ljmqVUtw0r7iziXjOh9b9TQdlh
DIcIfNnDjG4fGsqOY/9GuEB6ipjnQqneLBIEuLLd4yKU6p96Xwj8AIoGGlMbjQbgYXYdFilBC8Z7
Tr4Mph47SCPtSF4S/CRdSY7VJUdg8akBVUqODr1F230Xoqct8E2OSugoxfS9SHUk+1XGyCF3ZynU
GuiL6D56u4w0F9+OQ4C+z+j1g6bWKeU1eGd833hh4K0l4WKkDYCxBYSKlqP/VPzbZVLzLmBrKmBH
O0Cu5gKS3qbFMI1NCi9qY2AlGIwIig1L31OKDYEpgZDxNyutyKZXS7eTdvchoiC78DY4du+U3ahw
7ZWbpu6HsGbpQ8vwnooHUACPemDvaGHUXkDDoOYG3jTKdQ7sHXm9lnrlh2M0HJFRj0PQCGSKd6ow
VeImueSWL2cO+nBl8p1Bkcg4g47UdWG0s3JHrmEVEjSmKTIExjvYpf1dbQ92k2ksx475XTm6EBv1
WdbMe+rA+A1i0J4My2CmDgYxPLgJFVStjbl2wsbwgUiE2Hb+/YBgN/k0pHKNVouzEFNFKkSsHYO3
89ef30KBu8Ip/8D3x3s9YumN8DtrBawKYEX9Sk/6qVaaSxJJIdrEF672U6h7pgehAy5zX0HKqJAt
K1XNAJxof3v2q0bD/mhR4mRfdk4xBDb6pr+pl0pvUpmAE1SsRDhESfpe/4WaNuf/jXyjykbtwQp2
nOA9lay+tFTkk1JA9R5UP8phUY0gRe1JxxC1uYoUzEssWTnzsOx5v5xl1qGaGttUPwVJoDxDRMk0
BDNFs1Z67vtd4bHw43B0CpedR8CeCZIlm/EU01re5nZx5oKhs+muYdqwxJEw4Jvewm3ojn5z4E+T
dYY3D2ClCwPmKIMrPkl/9mdfaYDz+0T/CIUtemgAZtyiCKlUe6Izz64yzInIZwZ9AhMAsMZLWrr5
Ilaow7Z4t7TTdOX/avA7XxXBVEWFO2WsqIYzwllXLOEs/+OyFWxF8ud1lVfU8CS8ONPXmk2t1shE
cbwZAHKdbESAVo0lLN3qQQdWeCMN63+TDLpBb5umUTwnxrxuxk5Fwb/5ieeDYQ/+hRy54FlaxIej
7an1OrVFRSn5hx0XvuwLu0IQRqhVney2bDy6Mga/rdNmlRl7l2lWu8VjRdPRH8Vq3yNlgHTsTYde
DgWHb2EEwXGVsxbJOU0/jfQql0CgOBasNwjF8wMZlP1dmFPCRanFOjJYzEdskF3pqXrMQZAGreBd
AB7d/v0LfGVoLowp/FXmvcTAhZTyDauMH7I+hZvLheMnwmn7ZuRPeb2DMAsoCLe04w571NTKulUe
QPoT6vPOLJmaBP4od4OZ+Qo/+Rdg67mEJ+jVZmpndGmsRDs2Y0aw3BxmQwSSMaO+ETXpPa8dbwRq
sDwSkN3VjTP0g66t1S6x3kkwRFfgOsSEAnSrS4nc1GocjMuqzM2TrCqRiv2yCpAqtDIrPfX1UAyX
oWms+4TpS410W7gPxepPFruNFVx57cDKe6EMwKzrzGyDHJdEGKmOoqofTz5/viGFObj1Z5pxisr4
u17wbEhlifWgBQKgMMaWGBkrBcEVrNgKrcwTDsyNnnoDw5kLZtkVb6F8rIB8fcy4bX0sIdCfJTnz
ysAMZBstUJsaRhApNX0MvewxViJPg2sdS6MOaHsVkWSrZq61b/dEy1bP72MBLy8/u8V/yK4onEdj
Fma5049k0DHNwMo2j3Ybolr6y2Ol4zPwFaxjzm6c6vMI1nWUTmgSkF3jaFl67Jms1nMNA59Nm/cF
6JxGDu18ZWf7V2X9BMjNBlpu1Hq+LrS4tpC/flEgmG304b+/fdAj/7K7j7PSoXkU5kxHoty3D4gG
fJqn4raFo1MHbtx5C2o1izpWkWD4jFLViLfcfk2Jx7/lpZNE6+jFrDVxD6XxtGakVtpOb3lfAzka
/id2CDKI/eaPA/qyZLMOInF4/LEH3FWhBvqwSTZvWtrXhB/v2UqEGgznCDJ9wzyJDwiisghvhf4U
U7Pp4xAR7wg4zqBeRFgkoqI/KtjmtjFN9IX/bP8zH1Cxg173l5yqozE553WWk5PyxO2NsZNiJiq/
u6FVp7JvTPQIg1EiW5xk6xqARv8fob+TxVEO5AkAbZusicMS/jUvU7WJ6i4tYvJRgYZbf8kpjZlt
o03lWXBg77tZRutkpwYBg9KyjBljF4wUhGX/iloBAncFAn55CnDVgurI04a4NKA4J5gvpR9KwHWa
2cUothKad/dbTwQ4QglSTX1gjZ87YbAadd1zLFbc0ixOaDX9gIYHsvse04hIeX5iASLfHSrJmn/X
a1H19YNroqr6fMHhZ1sipaKVzycSwG7qbkBBMNw/k0jrjgy+6KnSj7oWy16RwOrznr42yKsjSLJN
YZtHb+rM/N2lajuYCPtluEWimGq0Cozf4LzsQjtjqsWxltNyxJfTgjbHku4KUaF4YoQCBHiUk0xu
TVf3B2wdBwu8oAULMd/Nuk9HilygyfwXW7cPkW09BJ6b7jPp0sfeNltg6MoNjArbLxobUKfRW2yz
ExVqcGOUd1Xx6HauNK2/sk9wDwMd0OkcQTzKfBcQVI6uzytdbi+bmDMwlt0CQw+oYzQQMzYWxR5t
IxIyHYRWRPWYwlmcCUJy/PguSW9QOh8T9EXD4YlumLKyTgNzBBXIkFORBoheqDGEkzyR9uW1923y
b6nAUT9BakCbgbnuZm5+ZRvDQQsN4axcMdtzmJ8G6WZXDCfb7EGl3xIfp0hpODx2UZpo5xyf6+Ux
pnn16Wupcsbw8j5VzlaPKE1uqhJsv0nnZBc5uTNIH6sWlOI+cO+Pf1xXrkpC1az3HOi9JDPYPpO1
xqRS4bF2TiFvPNKDegHYpegi87oefWNOu99ciY2zlz9/S8rzGHBeGqbfEWFYLwbpH91wMzqQWTc8
k+cTNqpnUYvNmxmQ1x4JNbz6lCLVVfhY3L5wfZKmOZAtjDaTGDA08Iq/qShxYgx9KDVv5cxACCux
BG9wg41lhygOHK3CS+/i7V8bXEjrJQMzldGPaJPX1t/FH1ICjsUxfDCzg8JCFgUV31P6IXMr5BrT
NOcX7Ji3Rj47/20mQZsB2WK2/52MWR54u6089sm+n6u0Q3Dsz7E7F/JloDgPnAASwcZ9S8rf90p6
trsYTvnAffXQmFvhWxSUzz/2JNNYDWJC+ri4BzRhNXtYFErITx0DQuaoCEw7kYnecFJ8rFOpetEc
jiPVPG9pROgF4dFwgNpksYGDatPqrQoiAY5CN1aAEsO1fvgqGInZPgr2GsAY4N0/PB6QmB9nB1TA
IoUVEypBLBknQgojN5mwgKyBo88aQikntvDO6KaNYvE8xnAtj5esAAXVUDH5NtCPvaQfNsZ4RQMB
kBjIRfaEp972eoJCV3ShyMWD+slBLbTm9xEC6ngSYqaANqnJuXWN8zmGo33r2lHPzu6/Ej8+niwt
EQTZDJlpp3h1mdccgAAbu4E7qadl/0Bc6Ivi3fkF4vaZoLTu8pVS7rl2AJtBzogty1c8wDplBXE8
gZaglwiqtVHXgsD2t0++wvfOLDR+z6r+QGKBOP6Ae0z/s4qwBz0pKNROiI33BINWxy6tdyRpRQWN
U8QKtAliCwTXCVNHdninmcfSaGl20CwX6AoYdM9tfPK+sJUQi7Vp3phXY+3mhKaxWhg4OSJbT+H6
phLrKJnPKGUBDQM8K3QKvXKhWD2tmUYxftDUbAONbhxsISUohAatE7OU3U/Jc2o66CxpOlPbANeu
4Jh/U0LHXzP+lO/3uI6puy+l7LjN8/oS1wmnheB/gQ+xJcE75nSvhsTI0w/GO0UzqUf713awKjJL
PhFRw9jP+SzrrTsQfNI/+ngkqzYjgVgrHKf08pDH/qkrQrFQ1MX2Ta5J+kBdUPTr9bqvlEPD8vAj
tJJ36wOSmeWLJ0Uzo84EQ5glJ9UGVMfl3bKyeQSgS4ztmPO67qJn/nF1qRLbgDnyA5whnncd8iUI
xLGQGz2Y1setAPXsBJHm2S1hX34wpa93DhBN7OKXVe+thlUZXxJlCNxyv3BdkRkL+6oCvlT008d8
bDNTRnRkKZg78aTR7ekapWkTlsBUWAh0BwZAxLYhcp0cnN1Ty7izb5SrJfZzdTPSjQ4zqSEELVxg
abi+joyFGZx3mwRB27bFxvGSDoUQ43Opkazl1bQA6/k1DX8jWrT9E2u+3n4GVI/hRjeXxQ8AfOxu
O9qbPE5nc2+0jdxixFq2jmC54SzObI52gXqOe5ewphEQFC/x5zApFt/1QqfiC+RPhGBCe4eG0Zut
oyIMnoefDYjv4u6pTeFCtJiNrQwgqKB8XDU0d/yKr3z+BV+SsW+hm/5iOUQjz3tHiLywMpcVQLdV
+OsyVQ2gUSsc2QxqtPXw6USeXRh12lAYC/PxD5zLpAUuT3BFBpX6Lsz137CpznyCjxFcs4x0upPO
gDhJDodRPoA3iFSenCw7wf2blVwd3CMvddducZBKdLzDVhZlU6q4rQxgtqCVrI0Wzg+uR6RNWxOi
x/Qs0u6N75gW0VVauFuz4Cz+/rwR8ydFPAoYfV1AeEhJ2d0xKprBPrtg00C4rhEF+clNiNFys9id
HwdHCK1g/JktuuodN4aRvOPkZWPV2T9meBAqVV9pkJo91cgC9i32301iqWGsD8d/Z8hQR+VZ6CK3
+6Jdp+AxrOIpIPAN3HEwITX7cCDBSXX9E4A2ix7tBuUwqmk8rUJa6nstJ4Xx4Cd/IWpy0V97kFiY
b7EkKHL9N8xGjImcxn2A2JAFQMrdfH68KtxwIl3FK+2WW4O6vBcWkrVdkJ73ptIS8yY1QjGI2rSe
1AaZN7x5vcUWxAtXGYIqTsnmXb+7cFAWw2KJjxcRSqMdoAdI8hHumOvNawzxuLaFbMBoy+1E4PBz
51yOcuJmP8eWRwp2nXq7H4kG0kx6Z3NIlRflQqWd3Mctno7pwE2xJrcC2yH4NthcrUzjDzoSHyS2
5dR0WaLVyyScHm5wyZ9j91ZuP6EzMmZRwMFrJlqUGL1MzQ/+Je5psuvm0BqcD1C9IkDLwRAh0iFI
TtVFxcWNHEjHetHlN68H5inh2+qWO4ppL5b0PDTinVv/THP2Zs7UT2DET2Nli3o7HfK6i8T3mOLM
SSAL9UhV9qBpxLkyhsOb4QYl50Hxa8F3sq+KC+CbrOB2t4cLqzWTIITcNbcxDiW7GJEQud167U4N
JD0qA3ZAoH8AJqyTe25UNdar7P2A+pt6Wkovea/SeFIkGoz4eOp0b74C4e/hME0UEZQGS/2JY8DH
2QWrPo3Tq8q00PR62YbxdpSAdIYUqn9P5zt75MH0Clf6/nn1Diz/NPcEQebMDZ9feXzgM8iNVHyO
6Gbs/v4FxI9J4a+78vNwG99qJeDuJKiB8EAYJhp10FnXj8XsyLkjjQuNZI8dWjEwaTsrHm0FkJuC
1+ask3EXN9Tr+7lQ1iNY9Ak2fSMNpXWL6ycDlN4sb19kugNtxVbKYD4EFaUbIEZvlUNGo87ikFo+
qAsrVrMPnuzV9LMmVB++s+ORH+w1pzgggG3AbuZGVAMqPeZoBKRwfAPpOfki9OuaIZ+AAvSXGda7
nDjUyhgQWBlNkmJ5jzkDNYAA7rP/jYNzGo+GIqVt0pkiXgIlt+z6rZxTdJd1wq/5jkMWS3mg1Xvn
jAAGdx8LlGylmuAaxjRCHb7uIEuN8wjzh5/QNCKg9GeUlwvw5x2cp75AQHzeebpftAmVhgWHQfJB
KEw/nrVDwvMEsufoYLNaqgvv+QO1Ott64Z5m9iMQpUJ8LR7Wwvs/kpET7xqqdqmpSxiaQNcaLuYZ
ZWXnNqBcfDOohUKNSRag22gOTn07cpvlkjZBc6foFCqZVx75l/WwUUZ9Gtsn0Fdlt8C2h42AE3QN
m1TLFrOJIFPC3fGt9hPqWwuQYqI0NRuODwGinPgI6D4f//7yyGbzJshK076doiJ5cJ3G9kFoZr1P
jCj0m/6MR2FxkpLFRZKW+8RuO0VufZ7WAbIJo40yhnkT/qTvdEhQhWzQLEd/7nMpXTza7LcBnBjo
B4TlChz3FllhjxI+bTUjuxu7AZenfPAdXKg6z0bG+oHHxXrwrHCvTOZSQS2dq/sb33jthHehHGgw
4+0yHRAQaS8264hgfpY+mRLhxP5a1Ah+FVyPJFzPkk0zIpuqdmYnLvyDKkiVW3WFkYpNDsJsvnD4
/tEWpTd0fwbFD6rKMFI6otMq4Dxf/Ww2v0ktYvXUR2lANgoLYC9z2UFc0nHM7eCdNhftmVQ8omYh
glpsmQQJlYT5qvdBIckiEQ8IzC3K4xEpDXZONVXDPdIfhYe2L040JZTekK36JKG4OLt+itdrLsZk
0Hr0q818woVunbN7NxMUGFF45FII5zo6nsn2GQ+y2Af3f4jZHw9AGKjXBSYqcIHmqtzi42R+tVbC
kleTCIYcOkjexSMzIw0DGUIqV5AeaEnDzx2Hnu1BSeUbR31BspSaqiWKKQqByuzGUDcsDINdkOYj
pyZfnDJz93ZPAweNt+SDpD946iwCvFiOYkOwK5c+i1tL43n62j2H8YBQPeDx3ynMfkPYk7rfj6om
tSJ/0WAx/rc6rtkQodG3mlQhKxoA6XVA1fn9ZvarEwf1OSiZ9b1dhh+z0h3twSpQ+u3pkPjGjGbr
nMB7L04FQqtjEvgk5R1y6xjGlvf80f9v1OLzRZUM6VLybCuleJA4EbbAiaGcZdsDKhUTpTNIATPL
n75F09O7eTqPCuVTrpaoYIU694xR2VlVnkKo9XekgTlkp0w41tXIN0Vp5QNh++3LYr6+QsL2A44K
Fp8Jht4IhW6KT/q0GwReYhRSJxyVW1GI+ClVYSGizPantuIt4S8lmgMnEZvOb2JNvCCjWmlCGOT/
t6JM1e62xciAQdTTYcAd6iShZbfxggCYtfIUJo4rWAQdcKxIY2GvBjlAB28AltMH59PaxrUgT+Yh
788HsLLGFgtg0UtZ01OjqVgKwh2LA4W0zThIc6yZlkhJo2ohbJt0LheBPF87VS5Q+0tJcXnwAboU
UoywRm+Q4kVImCAYXngH9SVkMkdBoyyUh62m/yQgP7yIH1ugRW7tBCMUcVCy5X0EJ0//OUoh9Tee
cqX3EEP4WrmEJmdtDei9hfzX/q1wHIjUJLQoNsEH7kSnd6N5CbLsMJAB0xh52hqVL9fyUHlCaelq
kgY/7nTfHA23dSS0D2W2LFPBKoGjDIHky35+5Cmp5zWC96gpkfnHI9liUtGWaU9DevZM1GNae4A+
S+qKerPYQPgQb2Fj7A3EMiLcMEOTECR4B5+Q678kb6LqhED6pbcxZRepLQOYOB5N5gPsWfgSu9zh
LUgk1ZHV2ISHHknbsmM0XUgCP+1uU0rdsZgTMYh36MArueWcKxaJSnAqCL0I+Df0yL4DwWN5B5B6
CMsWNaRrTsTOiaV8FMMFKpZfLps5bjShhX3yrJPOSOz6DP1TkoW1mOfIeEYjgYP0yCI1cJ5OPpjq
+yZC3AWNlpN0/mRHZdFfY9eW50agxUIRsA2S0APlCKj3O5gkYZ7T/G7vyg2bsnGZBfOAftA92PMh
wZqFiHhbf6mV7Lib019iqSO33Tn9PhEOJtziUjvr68wqtUJzHmkP5C4X21ydVO+Erwv9U5TZ0F/Z
fSLZ2lNLiXsuDNHMEmuY3ktcU5pnoMlwx8s08yQSBI45oKQ4eexZW5nKX5ai06wW25BhP3fE5wjH
1pGQ91RlfutjRCOojRiSOwpwwwr9ugIvjQpifurI5kSvf11nQ7GWPjtkDQ2O0szVkjhwn87C4I/y
AbvqLTeBoi7B5Q/rvODMjbVFnlMBlTLFyas3IORufDl653dQveJCmJd8hvE7cSA3ccGUPpZJJLYR
Fcp+pF1GWc5Wofd2tvmVIftZUmiaMZqIjtxKhH8ukjTB50wVhxthybHIqcPItXsQ38ncJ/rGqGUC
r7VdkIP6VCv15fOT12YIMfvrMKNYSnQthVRlK0I/dc8kwM8C3aIYNF8i/S1I2zygphVMhQuU+Qqd
vT6ItPugoIUB9Tk9VrW9hLKWCismzRvQWmUxlcN62A/wo/tpwuvcXuM11e7k8ePtzevfwhinZYbD
0F6PMEwcI2gjLBWzDJjS2ZwAlIBlpJ3JlxVgGkxE++i1o968vHw8o0uXlzEFoeTTdex0DdlA588Z
alqZDHydRzvPki0cdhjzm7YYH7rXYyShjxZHJVGO3zUjfGGx8bOgDvtLgu2pxZF/Tt2coO8WJwSa
bigCt+v2sTrjyEqBLDIsXa5g9ULF9LnAJ4Xt+MI7jBEouJdTgD2lp0DC/HWWyRVjw8QqwLdKkO4B
5Ha6W6bWEZVkbQeJlBEpseNBwCuY3Y41yqBfazXJID4Jmz3CNV3S44q48mvVW3r/plAtcWqgQBpc
9KxKJZHklFUPAu0GKVIULwoHE4dFrzRQXTacm6D/bk0rzUwNywTLefjLFUoIyEsBJLhV10V4Z6av
HtyHxw2f5xzLHr/6drUbg/0fRkiJm0aqgtMDqPBosIKocfuBHHTqlhzWtpG9yTTS5D6+fTvSzQw5
23e5U5IkSfDfJQPo4uQoeJfYWBEEJYjlVGuGU2hFeGN7qxFzyQNhTZuaGIuWNyvbb5rtL4B8LOFP
R6CHbk3+OGglc+J5EUcZ6x6UgezGFhj2t8XWah7ZNPNydaIcfacyLVc8g3KVmhph6u2fda0vXN9z
X2duhRbwJnXVIXX/j2M3jPJsDfw7LBThLry7A4EYm606kExwSM9smXzV6WLeb+t1tH7szQKBVz8v
dvC4UVl8eyMQxTA1Yetzf3u9qfZTixpx/Z56w0HrE385fW0hmyEF9hkxqfjpkUKiDPybjIlqE/Vc
Bvzrc0MouwsNBi2DmizKdIGA8fSDn87YlhYYQlYPycCJGXFLLJM2AMB4ZzLe+oPE9x1+FXTjPvCi
/RPOVnkw5Ud0rpdjCIUeOhp6ZLAbW+skU7cytRxDeeVupLhqx1fRjURCjZLylsgesqsPI3emohow
S97TokVlgLF4DZm1EUm+czmYXzfNgnAyRd1uoBOXcofSKsVVmplHmmF4CGmkTNnczDk69UfRSTyW
u0PG6E/UO37EHdqXaUuVrqoBjGSNP37xhIoHMUufF6mBgZZifY2ZAw8hAAzmP3QpmjGKVGbOrk/A
3P7WE1yLTnCig5NyeHFBgLYDKa/eKW1pfUFgunOyd4eprhtrrPSBbWEBgggWTEpo7O48puj0tjnL
0JZSmcjfJGnECErsUejAsS3ONotGxs7DI73XFtBw9NdvSBzkjOsw1yYEuJY0KcslkWtLVveKR9fi
wmk9lqHs4PV3PMs2P7TRKY4Rpq8t1wEreeX5hx10tu8Jfn7ceCYUYKCoTkQf1yad05Yv2xDMUM85
L+NbxS/83+E0D4LCDcQaFFYpjyy+rbgXZsF/PllYsPOi/tolaBfTGg2VTgsfX0D9vpl/Ued1TupH
AlifH7sqKANbirohzb8j9Oyp2OEeHER9M1wTqtDbyGnoBeyCNf0h+LXu3S/PQFtEr2yS56LXI08E
FYbDc9M3rHW4wvkNJD5RWQafUMKUfdEgRIoEEzTgbnsO66tKnrbeGHpNp6qMGoDoZRet457PrzFo
S4z8m+PvE0T1iG2U3hbrcjrPrdqneN6f2J5ummSY3fPWYFvjg6wVaxTulqxwLbeJP7KEHNSO3R/o
iqqpnkLcljm89p0LA+3beYfgfyhjzkDZ9jO+YQjrR0XLU3rEdiIqLNfM/i/In+oJfMRzB8jmZfQC
U1kXbazWkodpVHN35J7zuE6wIeJHSHXbQ5pczUxIU+WYiKoNaoLSQd0oG90M4nuuNqZPuekQJiZ6
9ypU0GGcn6igzekYx+Ao1dBGKrmXFwFNJdFIKKoQbJhnj7lB1dhFdXIry91KCDEGUbjv5G1Ahre9
6t1Sv7maoAur8EYZ3L7KoDRIEHA02dPSb9833ylOWqxr4oLVIb0FEZGJWLSqJtQRkkuYceMLE0FZ
bfwWpmwkXwHUot9sNaxu9zFou5MGbjus6Lxy+dx5hjnJKi0oOuXRR/X2lohYAKJRN2N+LPVFAN+d
w/dK3kvv1pKdPaPrgJ6A91D+IoCzxBfHxha6LO/LcLup1AVVkc+th8AZAwpu2cj2th9B3grx4G0Z
uKvz/LkJJKx7d5Zs5E4DE8Cb30voGSlkYqrl8lhdDGUQ0Azvxf7atkZVrC70T+U1lOXEPwSi77zU
v/cIH8DfNFmueL9lpBO8yhFK+uafkOi3OXD/GqGvI8kbhOlAxFJA9L/GkITm7NSI5hzeUJB3dUsv
03/Ta4/Kuq/KTk/wQSym2Sf7mzr4s3VbABOl7UbtViiGxZwDUzJD42ceqV1H2pzvBx8IK2x+Jt2Y
5t9q8hA7UWk5U8qwX+D1uALvHIoPVZUSWA5jufMeyRshjLzFoblnVYqmRvJT+MQU0qV5X0dlP51W
unU6dj33+ssna3irY3ukMUjxDF0Bm7/0ZKUysjeQtYp0Z2O4D0pIxump6FQMEugTdpw0gg/iNcso
hT6yg2+AOy/tzFtFJK9DPBR+wL6jrcp1jPaHjHHRoTtdRj0VwET+YvDjl9HhjzUAPuWdyHk4Fd+V
y3mrBYxcgECSHKOboTZwXIhEBudTjEcuJryZqRQC4KEtcy7dYEQdEMozoVJk5GI1jyUZaC/dWdOc
dkvKg5Jw51aAQi8pNE6D4frlqqwIjA2QK/RN+nP/j0ilRzVckeEU3YfMh/fsTPTLgd9nmTFb444W
YjENYzrFmbFIaro2iO9blYizp3G7pdQ8AzclBPQ/CSAZxjpGsEUsnoXC9EDZOmg0tiDJ+6V6E4zk
HL8dM1L3qpSwzZsQfqutCDZn5pHAiA8JUzhxjgBU6cQ1YxCy6ZQJwQDyBWu1jhxxsjnItAh+vxR8
jrRxpU5uIFSFxIkIu4ck3fpUawV8RIWVq40LhJuPOqNzAarQGe9JEfoH4xxDYfoj/z4U4XST1rIS
u6cllibpqDhB+nvQ+5kYsqfiFLr0Z/TxWdjG1Htld0IJWmck9vL7iAK5Gll/yWT/n6q94KFBSkjd
4lMvcZJKYpOVIrQJCTFC45AwoPf+CBqPb9zslta4lCWusfsBCvn/UQytrpvoQRxW6hYKH1SMOhTf
2lOw9sgrLmbCIWrQKz6YiPVVVJaTkZhZY8k4/1Asj+CBXwZUIOhDeMWfwSD++ZDqCZ1+tI85yl0t
ojlsFIhCkEkTNGBVlLHhF+VrbiPhZhh1ml/JeHnA6xgi3YCz9dvW6DPaxMigDEMIjxmUMg/pWhA3
VLNsxU9yrhtxIVwjierLgMXs60ED9yhsmlT93/EyDyn7XGqt40/vdXKuo5sJ6Wp0Kk0Z4bsP3Y6k
zk/NmjBoN0/Y3kY4mzGzvBpAbrNTQqGT6aJ/XWaeXn5kjLVq0osH0Kw3VHg0mf6Je6H18FQNeb3e
GV1nYCifk80/58qOzboPN68KyNPWROupOY7rdWFd41YLWFsy+I1eJJpcmxSoyCrmK7ZMQZwD25vo
bSzZ+zw4gLruMF0hITH/4peZ95g1fa6EZRi7vK2GX69BRzs8zwgzwXd7+vxFwEyOysIvGlcqCqHJ
H5b8msz7wy7P/q5LLrGmBszR8WGB7TIaGyWv5ZnQKHbLm+BeUZkKgjcp1V+LrF6gylMf+yJv184p
pnplRwC4KN739gWMQ2I6Yfi0tjeOdUv+Nm7iwDHbmP7jAzvaCJfVLbz+Od1ucflQeUWwDtkJLtLw
92Ll+HZXOu0jlVFGdFOVFyF2+GrZgjssSJ8jntRvIOENWLx2S1Jctk2mS+TM/tUZ/RQymHIKbmxm
CTCSVDSu/VmlX4GtinoCknnL/ryw9mFNeaX66Ac1aoDsGtHiLDBdTcxBDchJ3Oo4GUkWTfvBg4n4
1zFoiJmZkGlYq2YXHoXC05ZC+yn4wY/nIizHWM+jk4a65JwGTnLFsmIRyRWFL1A4YCJWj/dS+BP1
rXknmvA+XACoMcj5ouc0eFBJXx3k5xphoQcL1FC9CuLaiH6pp+CwofCJ/xdV0eaq5pQXXSYjB0Pg
oNPnojEqp//5ut94DLvw3vykGdwZI8e6uQ9YqrKrI1G3UuEP5fP8OdXdqVb0psNEOrR9iFro72M2
LYRMHnnvttcSDThwxw+uvTwKPVJgtl71iXxOdGep6N0fnjH/qzgHqJ7VB3qMcKemZZ8V4Ql2GoNe
c1PkfBXi+3XX7l90+PlbgahyeRM1gZxefoLs0HMk6K85bueZ7NxRggDR2BgVIqNxKYNTni8cu+ik
6hy60OjLF2tHLBhHQTqmG3yXabO4OTP0yCKvYyA27Q6KD3rtnmk7d/muCFlV2PIJAyBH4iASwGZ6
38zCphp9wGkXhLj++Y08Flu6mMl9PWqQ6WcWV4GV0/EdGkYMK973i+EuNmmvXE5CXcKhkL/5BE5Z
05yDJ6WqmIpMVGkGXTeE89geu+Tq58sTaq+SKWT8AKcyZCumwK1Ylnwd7hIbYvFbfc1rxDF6npzo
k3kDswK3U0+s7L1NN2xj+T3RfltQ7O2Su2wPI0+cBSZMZ6oz+3bbHZuVb3f98nCI2hoUZRdSTrk3
dHayMRUtnVq0g6Q6iKRMzX/pwUkTtz5uuUeF+UMxeHhOUw5NcsTJiLs+9lyTPhbv+eNwEayamhHs
GGiD/emfy6VLJlLXevWuMnwuOxkCT9u6wv3eFSL7Q4p+m+lD9lP3YZ0M2dPxNfou+a2nvaJz6Pfg
0DQwpWgi0Dxi+D6wM3q+8Eh9HzBvRSMYEaOHgtsa8/TAXNED+xTEWi/4UG+Jhuw3IWXahsMtPW71
yFA46UZtcwqdZaE+oBnapvhDIr/KzLy3ltVVqdjBkgKWxo46yKlsZoRRebPnMcugwptHC06IaEsL
sg2Jy2HTfGByi6RlHonEz2VhCkoUX+xtYWJslkKnG3pXWCl1l77k4NpPQTKGZjF9Vmxu7DAIakbY
dVzH2jX1y/f+yfR/d/vCh2Zfrq0hQpLRTz2Li8JAZvy0LkIN2f0gzPY77jCn/ZEPkXu1fgExgLAB
hR5vHlJF0K7zqKf13BW3Exs6C7Y9df0zAh8zpt7oUp2F8yxBm+Z8Vfo20QVCDgbt4HN2Wdrctyc+
gIs4e7quAFi3X6gGRUTRfwQgfU3hajBJ4SK8yPwQScQzzHYJmOu1b59IDlbv2F9bhT3/IWalh3JF
BYo6TRDaIQaRW/8JJ0i/3M5URBt+OkmtZJ7BQwTPxs8ABBJadI12gOynipdIfQsQe+6KJoUSCjLr
pLubabDYdA9rdl9tSy7mjyfrtsyA+AdEFmWYQ6zc0Pmtn9PZnNjyyA1M+zyQI+gMQ6F6roqnYWbN
H8MbFDActW3Zss7vSYckFrY6I2cKDy3SOdrW1Tx+XzcLjSm7KRrtoCxv6/WLRjTzDdh8lXtxuGuT
ewbhKUogKs+Gn4/HSh97riFM1FJkdSUkz33V+Gp4D1rE0W64RWok6aoXKU1Aw0nxLedoW1QcvJT8
78rN5gN+llQywamLkVN2vB9MahSRKVUBiZtUQV1yk04JMDbchLnE+fEXVhTE97y9lgjKym3iOMu6
yNmmN+3OEJI46ponpUHT0J/mN+LA5JDHYN9WAuUiYMEp/y+PSTfc0waSdaF1MwCaaprYZH+XwCVU
eupBRGamyw/wFz+9u34Ps9M7VS9moWp/Jv7K6RYnU/V6noeV4EaEtSrdBYmsnNEJAjfbEKiAzJbq
G4GDN/nhLTxLkZhIPh6ugaA40YnMns2xGj6S4lgsx1Z2kPxIG2GwUjGfW2r33YgHYdP/yyyiI6hL
I4NnjconqIh1QIeZd5fziUIi1Cbqoz55cVVsa6vSGE6Ojad9s8JZWJKnFjPAtiIeD8dxRryHThMo
dOun+Z2S2u4ehfN6AlVww4PLer6NEmiYPLNJuf9SGduMjmihFXbmtI/3WMS67C1wG2JUIa84vgSM
YNaITbayRA0Pc3BfPs0E1q1jHiNEE0y/PZZPwBz47zKZBb27A+hqVrqFATJonLmT++u58sRrtwpm
mHSjMl09KeE/8KNtwquh3GAYTgbHWmX6BsaRlaz67603RTTSM7ZdZ629Ah0UgPjGpXqpgW/LujFU
NaYKxhfOmP60AyPFdVpDTgtNlH1WvrxV59+sMxElKZjyVTgIXezzgnmZ2ipfIN3b7fP4bB25l0zJ
d+Gun8bkkTVjeeUd+H5glpGcIaSfsT91n4tb52RLho6t8f3I0p+K68G33zleUoAv87TIgv+i3osZ
tJ2rZhSii3AeXm+21jl+zaEacPpL1rD0tw+saCbGDIx6jPzH044fL3ia2X3cH0Sd+si4E+q/oF5Q
7HCNqBiq4QWTAWsaj5bFVWNZWzpQp+DS8r9gIk/vyRvJe/KJ8HFjp/P/03kniULzUprY1vjKB1QW
i4WMTiJPUcLizH6zorwSjdhBls9gXdYvMjDWLu3d8WeYXynQBsTQQVDpRYLYufuLW/2vC3aj3V8s
G3GzSNJfAKxcUNmSBdsPMuKNl6fu9ACV8sdMTJExzruVTuPQQGYUY1+R4B5BAduL3F2GlWaEfPHA
VnRpj4ZTdga4j5g7XFg1rnce1uvRXGwpj8K/JknG2huCgtzMu+K/R29ugi9NUcTtCiuJsJmTkOJx
WRCMdzu0fKEHAcUgob/g2Hwy1p4JjPnPqIP0j3EltIPMchsytat0J+Yx0cWHO1lQp4NmwWxDt9B0
iALksUTWk+dEJFVV0ZWDcyBnFmvvNInzu7sFZHzhC7uc+12tt9MdM7SLcX9BJrwdLt3Bk3BhMhdB
CfKfAS595L20GIlEaITFfKHISt7n47cXeppitrIG77pupVC6XFksSJ6c3HCcfZo8sj7kdIijtjyX
ONugTbSu3QxodAlbeLNp1YP9P8Ut0x9KMPcGzwcW34ktNEZJlvnC6kwcVRARTKDpaMc95CnnL6nZ
JPIXYanDWCisBVnF+s5oIA6tXXtIQhoNZagYCh//VOvJzS1nsC2T379rUMy/C1kjtNlKdz/XHaLO
3BS0YtIPKfAwhxgHP5zryp8+wOSLFyU2QAuFUZUbjRNoE++6v8FroKoGayp31Qt5uJTQTpzSb7YG
fxipHxl1OIybgPWonvcdoNIEK3naNrnmHJ2Uvqtce13FslUiVhw24qQGLzRsnfKyaOhe6r3PZh8l
Ly6a/hgOwLt5WdUYfAvD/DvULPcIpxjoOpq5dERkkoQIjfIxAZmLxcCCz2QtnYnwFiSfaTKBuw8S
DpGKmJuYP+0uZlAuNvxQuoNmA7RDMc6nFiH0Kas8qTXkLzm7PlinY9rXpCDtVwJMXPi80OtFGZ8E
fxAJBaY/bifD+gyqdlPgqMDDLfTKoFfDx1qD2xVsnivKLUgYWcHRw9+4WB0H5Wh+uEz5qy4LgFS5
6N85pBQYfFXGX5+wFRJDUPXlJLuUiAJjHa5tEa7aS97Bw6abUA6xoUzZNcaD7wzv6PbvoLolSn/d
xL6o9Ae+sU4ICc4EW56LD18CRRCYEgFYV3QAEK4xfQeXDhFjhB3Q4oQV5kwq3CV960tZilGnchjO
3cJPX8eDMCkkSr3pL+VvFGqA6Z89wG+QNtzNmdh3ni4xCKddE6w/WQ0uK83qznakzLSIb+uiuYWL
NF0wY7ZFhO9eNAf1xxvISJ/+NfHud2d29E+JCeSu4ST1gvrxpPDlcVxQ2SPriepO5OLrwsLG5C//
pDn2i80Q7vMiSnXbFg53MbbPLOxPEj/lS1oKsOD0Gvw2UoHKe6v8YFVBD3GKyjJgB5JQtlQW/BKS
xXl0MyuUEf11CJK7uhL5Pba1fwG8wrwGHyNdxkTqaIkTQyLrlvLeZaYoHxoX1ERr6LbHmjmcr4BT
ih9m3MWZuXtIF/uOYYPjhcspGtgGSfgshGZGnLdvgRNyQhWnXJKCxrdEAoqhDPvrdGawx1hkaAWU
KgrVKkB4BaLI0JsWd7z70ykCbD9SceWE70yT+05V0u1GFd/6nQKoDodAB0a/lWMYCdDxOxBoMp4B
ihTy60bq6ABfOiCsUqx1q3mLPA4ptLr2K0mp73xTKY/1At3GFoHCqZ55oX1xT5iDklHubt3sOqR8
kyp7IxiEY5AAdfZmBODFEVegvDxtklTua5XSv4hJ1TcZJWVAblVVLbbLaKNhK5zMu7rNAfO+DjHv
wCCapgSQEkZ43de3WnS/HV2Z9MjitVeCufhG4mtlwf593kNW5Udvhw4u30YW4/knJGgFyAHTAOu8
r00k0R7WeNvAIjm32aYnNTp1D/K6R2jD2IN+AztOUoOJbx0ARkslV4yuGce9H5NUadvDo+BsgO3K
l8y9icgHpI4KMBs1XjNhJbgGeF3Vdu+FHafwk8naxD8FcxAUEYbpAZW4xFktgbxyOgfVpA7DThlV
/KYaUNfxfVffc2GUXns59nUjgwqEd/PxxiQboGfaZKDMGCj4NinYDlg1w56FItapb5oGjFjqOsZV
nG/IYVNJn3t8zVwkU75/2+eKqAHmKGncoUzewx+aKgkJmBaiqYufwhHQl+tnxSU4BLiUewv0HVTt
T+5NgiF02qAuKvq2J+6lwr5R7WIWgTRxcylZnDDajVQWmjGsWp597eezN/W+ctJcR1KSFEVAs1Ex
fwmUX7yzcyjE+AYqnhHqrB1OQFxvib4zp/8spTmp9C9F1pfzeTK+OU/S2D3gxawZl/f8VjgMbQwT
J6ei2f1k6aodweKP7EXMvbAQgmM97kc7bgsXr2Yn/UxNti2aDRFmvJ31sUu/LJz3a2XyS7VswBjG
8Tp+VBGysHiJ9cJlJVjI6BZVN11oDy3CjwCk1B8wKqAhJestqtnJOKjApP9BEOg+c6TyW5d8PJVg
b8ooukI8Z7qIkAz8gKWSMr5U/fxwZ0yg4924bLi4+qnasdsjlZmSRIhl+eAoJcxMIQNxrkk41Kci
vUYY+jprAcBho430Wi6tfpFZ0TA47S58N0Z+moEpxyP4SjOpkQJE0aQ9Xj6sIi55m1ITLmIG4+FU
TQ18iGBOKoP2825mSnoOnQEnuULb0nBnGc9dOkyJatyqVKgSuwbXxhblLq1nnV4Z/VqRVVHppyCL
1dEMl7GVmdTLBIMTMzNdmcGcWwLiPj6dIupM2KO99J86bS6U1H7tHKsBoIkYorqEIP6Me0NuRne6
l/4KPF9+0QfabVO8DnIvlqQqFN8K4cRVnVeyZC/8jMI27ExPG7AGx2kS/OqKsGVO1z1dlzkBdXuF
JxArXcL7AMoj7fcOMtXKbIv13CojQ48dA8wlqsC/jQC3z5hjwbvxCcNUlP4g7CP+931Ky4DtegFO
8J/EjE/QMOh+3Y3i6TQiHZ53Q6Uxre3PM1kA9QNbOi9/QfnxQHMCEvzcOOrrrAqYnhQ6vE/w6rC2
6YXOPzqKce1rpYzfgx3jnZkcfzW6zxvot/zIEF98cObBCt9uqIpwT6tt8MHcuFzM8CXTv6jNQ3Ya
zr9oU39E1Neq0KHU3PXkMt/s+yp1Rc37Pt9HxDaz6LnjmSNwU6MQ5Paxa7ZdmgLLwvZiesG3LklA
6LUWfARzmlKNwFej+sEbM7KUaA3lopDUURN2BAt3A8iyuPZWLU0TVBAkzK8XCDEd3LFx8SExmbtm
1vpnwpwFmXKyaAf7ndxjDsdcwlIduUMw4CmfuVPFRcOwtIKF3eGpW49dwNcQTV3FIyUE4/1OTI4n
uCno303t2EprLuG67C7RQ4pnmxjAYARV5hYAy1Brpr2KJaUyTKk8JM/6Ptnj0dzLogr1VyorHx1Y
/vMfrzEROHx5VosYdckrOv2LzoaS/UJegBgtLEo65/RXNC/qvWHEU0QfVZ3H+Hm5NnPKLuXZ2yVR
m1DXno+RZnYZDswsuF3Y0fa+hERWH+O1Ybnc5qxUSfZo7Zj8ZE36ORhc0vNtw/jyDrOsjnftu6r8
1zwE1ZrkT9CMlDuf+j1ADypZhQqVHSK9WJR7d6XDxCw1lMKcJ11o1jLfh8M7e7ETq51kX3n7URw9
l0y0tE1DzYCrM4TUBc1H9uDCRRzgEUZ+e1LXVlyoTuOveUmRX6zlzEw9ra8S/ZpIbOKQTeq/WR7l
ppw2EEeLsGL/hUI4k4Urs7DKh1Hh2Q9zcFMWrpG3Nzcha79k+RFP5l7D/VTJVqZckFWOs0CM4cFS
CWaQZF7bUgkCEwUmOeCGKlBu0P0z7nxT3M2yCZKM+Av/ypy9KzToTxrjxUforJS4cOaCpL3pZqMm
JvZr+FHrUFxo+KaJ+Pw3bpkfq0wDiR3inOcmFcFPRERHpoU/qe3Uw6gK4NabBOOh/ZUta40teQN+
GOeGGZ/uIJIpFynOR1eyhq+B2yMVrmSvUmnPotYZAdCp6B6TlQuQ0dZoLhihgR4IxKOGn7TpUROU
YFyRH/vyl3L+lY4laT21f3RyKtFEFGMLquJN+YqKp/U4Sf8BCMrNn6S2c0dsQJHvighrUxTzJknQ
DYTg85onLSCWGiuELimrxznrYNXy1WM7N5Pu3LhOoWXpvG62PjKj4m09bm+XgHlMwdFI0pilIycX
mos3wQe0/ZZh1KB1kMAD4rhBRXjdk0JQPg8LIQO52TSJlJZ+rPGgcuCBez0r+q0LzekO/mPIHZYz
ehFwJqAk1VFIxqzT6TZSGHSZhPGX86u8eOGA1JHjDhpaikv/FYGhVIF9zlFaCzL/FLmg9gLz46oA
TTmkWu/oPC/1rIRmns+4Sv4YuJpqYlKtUuBdzzxqjogfBTUN/7iaJypyY30Oa/FeKOtpMvQDhqci
bXSyC2eG5xh4jJm5eXwxezNLWranHq02hbbrxiSwkuzct9T1sLeNxv9tU/ddv9NilGV7oZ0bGkV4
zxeK8kweXG/YDpvHCTlyG93y6IsvEhF6/eln1krLg5vsWWvCtA0GDvcix0xwiPtOJ+wtXut3R5g8
pSzyPjMmR2ROtQG/vEINlOx2UD6EoAj1nj7GWUQ1a+/wbnc6tdywyzHTGk/YskVye2Bwj+k7f77R
yx3Z7QwnPHdoIsPti6FNOIidCOph1lPsdCDrrYGeSOCbxhbA2ZMwhuoveyNv0QmBMmz2r30S01D4
yuZyNO5ZO65smXM0zjcHjzV6KL3FuoGK/fhVZG2VyCJggYt0ezPAB2OBBenYfl6LQYG1HdHLRbWj
FzqBDWcAIzoogowSeY4RmR6Olxi/RB8kMcT+0iMoJRg4IbGCWkH4Dgm/g0bHT7eRnIwnNcRn0ih7
2jujFh08Mfh+/YOPIeacGdvkxBuyA0xmnGWv+iAZpYA0uzuUphM0PdyVbulEdtOLGMjk4ZzS6mQZ
L4jZZroGLbwOQFBsdlbMynb5RqbWZkamGfhtLPJige1PeIeF0W8TRdisa7wTXhrkuMAgSi6KgW/I
jT9DpXSFaFfcpgGBLb/yXazf+JMUI+4cpufr6DoKAK6Y/jwMcGFaGBIitZide2PiDlhDvIJZDiEe
zMbRrMVRrn60O9Qxb5vR2PwALb8P7qVORJCwcJHVONKSjx62mG0c2VdOlNRkwMVuvJ80h6DoUf6X
S1a7fk0aL3iZ0bJ7doHbfcZ0L+F+zHzWgIvRAu7NV/3byAucehQGFkrCvaiDbrFad9G21uUlgWRi
VbSFkOhRBm2+mzvao3u3mDtRZzQn4lHpwVwMGJ9gPPtGUAPJLr4I/Zus0K8Y0KWAtxs27catxIcL
OPUKVAOJTk1O58WqQb29kcjhUp2t847H0efB6f3+MQkuld5rlcCOc3HKRVfcs7pd8ncslITAV+rT
9HxMaz4mSt031I6PqSeAvjGGrRBC0VdfeEtLe2ZuNej0EMUYuVCupvzq9ah0qyOOuj8ZLmcnWuWz
fTht2VIcuHAibt2DQX/cJXKsJQRK8J5SkYrSUXVaGfI1iu4l4rjxuoPd0pRA6uSS00oiiumTlpPJ
hCY7T98Wc3pMArdzLYZ2e+nbrBV88GsuMU1PWkcq4SiM1lV5tLfSyxNLP57L0Cx8z92yxgnvJ41u
d4uiDiqnnxKTT0zW1gJMgv4VR38xOa4Ux/frmXyj+YZEGBJrJCWs/k1wQRoe8HoC+eordYdp4HvX
wDzNB0BgpsyfAIfZSnviAOTF0K4zEoIXuZaXpGy7D+mphmgWVZuNNcQNiMzjRjSXRo03LSoq52PE
9Bk07B0IAlEy1hHIshe0hLUV9QiJXO4VnQRf1CI/7MWJh8y4f9/cbMsO2z0nVVKOEXKBL/0LvxRf
SRfsRw9Tlxp4S3NegrkBEGBPnfutWNWeBoOwLfzY8QAqZg5xPxXWY/dn2v+IGvk3l8CWYxsX+hiT
EgkUxxiswToAJqY12Un4QDvlHLM1JKD3Qf8J21llE6exi3KZJ/invSe5GljmZeEaUpJ9l07oRQWx
ho65QR0NroeaGKh4X4K/IGaM780E2GVpV/o/agN6UQvhZOZ26B4RZGe0fo11TYYg8d2QeiLI7MOU
d+ctX7opLVo/MBVxZgGc1UtfeNKt+PoDh3dRV1D2JXhgfAw3C/TdC92JvPgL9CmZ0gxsuU4cdCKe
J2Nm6eix5kOEGNJxohQ3uj19KaG2salsnZT2qo0Id7BFbgQlUun0coOWYzmhkn9IIvDeo04AHdi/
dR3camlGZgjBqNF6zkZwYHs9rd842823v+W0rM0F0+4//KAgzKMPPtfKp79OiaZ5gzbvW9DkLGzA
KvKaQKzzgzhLscL/BoHrbXSncEHrp25QRn13z0iu8tM5JTzgoZ628/+7H3g/E9xP9f/pMVsRdRcG
ZAyFRkyTfnvax0Q/W4i8+R2cgaXPBhtJnK6/gs6/uWmdicqnLqiC3nACfqltjIN0+aR4WM9iT0k/
rXG3CRcuMVeWfwMQMED2Aq7yu7+eGrwwrF3ytW4Fi5ftyvWTsQ4kE+PddhRLXCPAAITh/Ohfv/eD
1rAYyAo1PDhbgBy4OklXG27SWUOvPyPdFnSEsYt6nCZ+G8QLb3c42Z3ZzP+JzqwCs5b1thHrKGcm
89eCFWRwUzIpm4rmo5a5RiprIKmfiP3e4R7njSGhfifot9RUUQcOtb0CCxZXdRCGGEaI3OIZtTCO
p3bXulEY4redbEUEqZHnwL/GLf6zVOgHM9AwdcKlPdQFhsQtlTfICLdr+JhkeaYnJOSk6wirTNSE
3ntj2tL11tuy6WQVcki8j9gr+UXKah0j4HYxBjkCuqPeBKAQfzh6opodqxdFFXu+TT5+7qHqby5M
+PefcsFyTgivnRoUoQz56U8kiyZxq0/+Zan1z85ePT5EC9yak6/rDNq9uHjjXSEXzAtQ9O4rCN3m
OjLQVpH43f6uUzEVxJYyWlUZHrDi5Cifu4wBNg6VU4wvw3/fevHz+AoFJLcjthRdo1b+pmojfMDQ
wRqJDrgeqJ/HqmvrOwg0STrATvXAy13KPhMNMwS3xiMRkkTL2/AdqSmQ1nRdIH21GPvxeQp0S4z+
HjPiaUh2ibDkwXMdQ049Ie5Ubz2l/eJdXnkm0rm8CC2Ftw5TR5NE1SGbSidadFGVcU3OASz2ggMS
yBu/z9O1r3gzvKvdWfXyvoaxoonQTryDp/0pzyDDBtFAgfSXm18tqFgE2Abe1fOR/hMGRSbKzhtf
KenYvp320874ViSf0ki9USViw6P+ZXUQPQw75QkYF46+RIamVFHQJoEq/kQjHtUxzZNCz71fzHjb
/T34kfKea0e09BgTAmyCzhZDx3jGzZStOfQY3LXuruPB2EzOlwyIuG6S9MLZndDf/UgIOXWRzqvz
WGm6v3FcROmRnxMeFgF3HQBzcjS3zYwBlY7Kp0CxqR99QKHTycKpfogguoaMajFnhygjZt/UCF+7
hONuJmiSfv1r8zDnolfAxk4cKLjF0T0wMwaxauyPc1Zjr1HvAa5WocQlFtYPK1OOkcM0dNaXzfna
LvBjoC7Z6921jQl2RFt4h+abSqanTiU64qCPc888Oq1SGBn70hqgICvp//iMtYZyuL0l5AVh7iWu
kkYgoRIHM5J7tiSYEEIVGc7M/SRUOazKZt/cQX0rFT/VGzRU1pCDZRtoiRFr2gpyB/OvO/n7XEnI
0ptHgKpPQwS6njFr3/ot902jWkHg7ClwYyXRkkHPh7lvhR1JrU27CaCVzEaWcColChFDM76MCLeN
++gYNnsyxzY4cNMOwnajkSoRLsg63vLBJ4PICO//PiYEvOYpLsxMk5AVCteDdBxCcrCS8I0zdu+M
oZpF7CZzSaGCqVSaDhk/N0NFi0gviYakPLfj0BhCJfeXdBBRAwjrfVB0VZrnywRLQJ5w+b+oNenA
4Xz9+Pzn8UKxskfbVf91LaXm5v+8jzfTWvk0gdIts8jl0bjvVYehIqvydiVQZWrzJqkSAH4f9NIO
JxkRNu62ae+qUPIRyHLGfhC7tdpn8uxwaIzjyP8XJG/r3I+5liP24VpxQduDXNAMYWrVX1xQefAn
Ur90Q3DMnBRYhLUmPmhUt0YfC5Eh6sHQZb4PTYMtW7OeDzKfr/LmyyL4mpmVCu/NXlGSa4wgzvDz
ktxZf6sMKQDpwHBzUBWGtguwgH1Nyr2Si1OkZesvJe/RUg8fRPY8cNZHSSMyIe9EmUwPXNMuZgel
VR3E8+IJ9pal1fjWhtUtDTHuaR7sym+Wi5Xk4nXZU5KfsKovQeUw3mytVAve5ufkIzQlAaIYaZZA
4luH+x0Di1n56gF1bB0Ccrw0BanHXFxBPpbp7XXZyhdcYtHMBDdOfrc2Hm9aHYX7KX31/rBiYixn
fn+A8+KmAZ3vO8ra/9dVShmTbxxLyQ4pmlu3qAKz9DWRr5ITr3v/n3AaBB+kkQR24hJWYeOY4elf
UtceZ1bI+LgLwdiu4yktk17QUCMr4ZJKcs5vJYCj+cczydxNi/4ykrW8NETlcbmpoO03eaCQvkql
iV/Gbjk8y31AJmXww8CuJ6O7LyvcICUFKWipKKadnmS10otzqsRxxlkBBggBtwXu16Me0xxzz+wC
8ebezyGXJX/0LzhuTut+Cj9MRLUR6iSAAam/2xz2Pbz3nytzh6mN33KUGY/5jpVmvpvdGPc9YpLn
MerRE30Dg/B6zZGQzk954AzYRN25Ov2YMCIfztPNyjMnaENTdpdsPJ10fN1Q5n0PXtVi//KsxYD4
AxSHTz/aCnbIXPLSWzsFxtWXSFzUfPdg1xOE2A9QIc6tYLN79pOrEaV/6wusSKlGV+kUaB4HOCxb
1rxslCXiXqqD2Q4bxx5jAKKuikitsdpu2pugcoYrneda1KJyMKVecvRuEAa5u9yc+6ED0RvtEIdx
002NGErhqFiUaWnPmEzkM0YMt9Ukx8peqaannW8CoMJ4fIhec5AcDTx8eXKsLcBJhhwAVRyMJRWg
OhKpu2pE2qQtPpZzdr+Gt7tTXCuctVqPhwhn+mo7wzZM1GxyZmyKtWU5tm2qO+U0y2tlQNBfThjq
FE6TXeAxah9U/2EYtsaprnCb/yVD1nZLdN8GPfO95QIXHCtpH+kCu7apUvm14MEahLpl1ptrab5o
HEgrs51usnz1jB3A6zlEUnKgJqHqAAbnKApv7zLN7XXwJ5amlgPMFWQ457igmVOIPVPQVEmSsrZ1
XAzE/MdWJJlI3BYwUDhmlk2o0dB7hq9tcZCRC82RHL/Tu59O6IeJLExfEQ/kLzLO6tr0gp/nkOe5
hzevQtXIc8p6PB4aR/GLUCNdl1gnP3tGk6p4Bt9kPcgH/ust8P7FBOfjCAl3RqYdXLI/TIyrPEGu
mTNl+UqFrALCJoDsziJgXJ1UwHWIl9GYjrisbXgzgwj5OcPQxxGD+pDBxbJPCz6D/djQvLTrKL3y
zE3FQBXKPQJcfVamgziWmF/Kh0MDyM5S9qjTC2973AS25r59gHkytFJLAzVDLUN9cxJo07dLYT9k
54IMNrzzAFdwHaCDTJ8xS4LPzIuC7QyAPF5tZPCRCQ/JHLUIARGjVSk8KvlOnEVS/4wSGofbOrNB
UrkMieLqx1ytV0pp5zJV9QXBtFU6RLafQAKvEt4mkiYn0QfdYpz7o4x3Fw4uA6zmZ7LcdGTvjaoa
rdnGPTHYnWvyY9PmvBqk/7WqNpD70sfGQprGVdX8VvQfUW/t8vIHvVKrvZr4S0GVtxAUwCKlGrSX
lTF41g01ReTOLQHaMjuLnmIOncgpHJjgZEbp5RCcxndkv60pG5HY2IQE2rNUOngIChaya3Fnfml8
jN1SPR6DDm+fk4cPdZ+aDMkAIGqy1uqvB+uKSwau8Lhu8OwciCYd/GbpIJ0TeTXxiw13zZTvcidS
JxxWgTK48vxYkNqM7z8f2r5KWVQz8ZieXdMzA81nG7pq4vyplvPpObZ4TXjqFP1rl+7ek7xmm3Op
1qq3npfj/a0kuZ1b5poI7ERR0QcPMze0bgBfCoIpDjZd8v6RAhcab1NaeZVN9wo6arOdd0aliCfx
CO1L/c20tEDBvVQD9RlgGZqYlb4HCfVX4JZrzY/5YGkQYwaWDh8qzZc7UyUfpSK2MOGeeYXlAPKC
TAHxXGXbGYa9H1r6tV0c5Xo0TC+StSOJ/dF0kg0lbsBdLOf8YI9ImPYd4dpq4ldC2ji2cp+SRpib
PjAZUdnMRFCzBWActMH1swuhi7XdXWFG5mF0/OBhCYfjrlclOyqmyoBPE+3+O7FyY4O3jmvWjq++
RX6u6nDbh8/QutbGk1Tz2/gLvpcJT0b+0rlHCyUJWiTrPvHZchduZUagLEQbNY6OrexbidytIqVA
TqcmiiGmqJXeqFI38lIqv3x7M62fZzj2uQrrPVbTdmVz9isIKezpsXizXEv+eHh6i8TzxBPrhrqs
V1n+/TyCagRzQInhHJnyMbc/CyX0ObuOH3JJnrfCRMQ50Iqk64ZP8AMudxjsJplwMqevG1qVZ3SE
bSXKQTM3An7AzGZiNqWjvXWoyE2rrdxzwBj2aCg1Y+CTK0PESRkL2N3jn0SGy7G7LCUGHm+Ayc9n
XM7eHAcnBtk+VA7IRHxUKd86RxNzuhP4dvsbg+HsEvCfAahbsnqASqq7wqjBnWRc/B9KBZpoyRI5
3H0zIQh2YJwe+9r84faYfkbqGZwjh3sXQH1Jlpk/x8Hj3tWG0ex4GBJcJXt7f1Oz3/U+DyeIV3dJ
BWwnwcCN5eCG8pIcTJUboAxpduIsgxnCS5PEIgReRLPw5PPwIqHUoaHbsoFqO3BprdbFjuimxCLd
z9bVUnWh0ajVpv0Nudi6uroIkhgJsrr5+aEjAeHaYrwMOXewamlkGmUjYnuedl01NtTNakd4H146
bUOWDZLTNIUdZOJFcquydtR0ZfPz9qdxbdxsCK3xpLlt44MglMAIyghDqD2wGkqZwO3x2zNBLVL/
wvuXpR54Dhg7P1n94MsDx5MAzfoqG2QX3hEhZvVc6JdDUr3AR8Q++qePFPcvrduN7rM8ZdbD1gxD
0nBi1hIONGav34oMQMVPmbEG+wItsGGgm/lkoBNYssBbM4iDmrUuBFctu1u6HSG8WtHZIzWpd8Zk
WQJLdHtXrhsKBugPx1brQOC16dJU8IKrrIyBaJBd66LIaCEz6J8Sl8MdwbmOogkyVAB7NHRMQ8Mr
asJhtUetEeacxJSgAkwCF1yjvMZTAKHP4SYWcTVUgHiGwc/2lnBMOwyRz8JOZBxb2A6nOoAoPBZ1
ZdQSUtsF+E09XdMUL/CFRX6Xj2lAPJaB5FTavl1X9cgXqlmUMLud0uQ9sXWBn8EIRHjKm0QGahM8
t7ni5DGmXmsRtFwdb4fFebD1VShqvtlbf0gYtrtT4/Fdyz0D686BkcAbZja2i6TcbXp47A6jRwI0
MiXRTiQrwRWEmHpXUFLizWVaAnSApytVi7Op7ZgI+c9UPoqONtc9AcO+goAbZPowOWv3P4ieffzo
FKC5gUUGj/UYET+N5abgBPm5mWvThpxcaIsKGhzn6ntzYp5XX1E1h6q+KWvqIzmZtspqBGWLZHVd
PWKapyzFUl/OSFaHajwAk4WnNWoXRiRBHTSQBdv065zL2RhR/j6bTY8cUxMSeVaXl6tMBsfl05L0
Ey18IGqEhcdEhwFVrb3nw0MIiSkTZB8ktruBLL7uZeyynkW4m3Sqz1PDei7fekMVDS+oDH5M4Fez
RXEPvSLePXPWVQvpcOZb9tyVuRDJ+L2E+qpKtSR2HuQzB3ExP3KfirSDB62EWdi8C7Aw3H0r04RA
IoxMgsfejF4VoRzdpTVtA1h6CzhbsuOgpIdcgxOgMagYsPbZaIsSktjPTxud853DCuIkPdanLn4U
svYxnVF2m9/ECFgRGZ5gGP6tQFHz7VabCvrRXnGkBJnBPkvei+hiwVWFZaGn/PixYx5+3ZFtU/pX
O+2dCxkNcEizzyp698fy4Kc31nS3h8CH8ZCqHPbwBbtHy6yKGsDufhNJliX+4KOhOPPrrHWxXKnT
5nKkwLAylqIyQDW1s+tV6+xomvrqn3+7SPtrPmo4VSzc3NHpJtU+JtCg594iK3za+EPIBGmWgrEt
ScW2GZCqRKJ1u9wgN7RVrOyOAtd/UlbO7OFG03eXjkelQBdLpK5nxhOOb0sBgyjwDltMAIua4tsF
FWouSpnQISYXqOb5F24ra2fdIQ3d41Sd0nMTe3tGfdxql7TlN+yj1a7KB1hOl95g6gQyseArUuKd
NSWJiUU3hHWzVrufNe92HgcJHOWG5+MVdvjlPQGM0sJFsT75yOQiCPrwEaM6LCDJ8n2NZInv/wn9
A1y9ypaNFiecDjbd1gwBI5r9Ro8MZVAbXtD4wk/lkPvBKTvCOUTtnZalOuvb/jtmS6h4dUjSe+4m
nGYTiYAZbQrAGET8tYWS44IynIySuyDHZwzjb6D82cyEQnX3gQVlYD1S5oNyqeKZr7eokQFtNS6q
Pq1U1G/4aKAamzupPzypK9JnISJnpURuwKE+K5a/AGm0LRbG9SNDAohQ6eLD9yWwd88g9PWMJOUv
mDmBAPg79gBhC86KPIjD0HWLZXaxg4V/puKpVv+Pzfcs73alICwYT5y4V8+eftm9wfR8N5QTKb8f
YFpmtRjiSqzEe4mMf9EZVid4TYBKBN4x3AVje6GQ11eegdmfdLsEQKgJyE90UWXBI1BUiwd2pZot
XogYRtwnIBUWeOiJfN3+WMrKTFTEDQ3rvO47ia5SDQARyG+5d9RwZq7WrdgL2rl2vO67oAHRPRVw
mpMa9m3u7jZI8lVpgLUi+eUl12JuVZEADhdUMuoUGrWO9HtaNFkxiRqeZKMTJDUo/t6qHRNn83f4
oxkrsHXVMFs4SM5/J5wenOg+MHuf7Un7szeo0mmW1VCGKYOC4r8mIyMuh9uhRYQYHBDvtAS6O4EJ
+2SBvMB5gDIg9Mp5+O9sNe8kAkxTAoVJzAnBxjRdz7rawmUO5M2diFKDw9ltvYTxGboCji3lnkuJ
AdzBwuIYyxz4bHrqUgkmz3K+4No64YG8YZyqdJD9qAXnBS1K75BDQ7ZYDQoH/wkVoEbnHvJKz9s4
enASdT70VKfVhs888jtLWc7nTLfKu2XyZ/ACOOAucZk9Xq+GO0qAFjqvKp61jU9AYCCzjaHY2LIi
r+8nTcsqNLPYvDF71eslKDA6b/SRl8vXd3dHjYTTxGVD+spj2Xl61u5QrzbLecTT5mtLbKCP+fic
Q0FShwG1i7c78Gjcg7yAeIGiztknDHSS9HQrwxjwWmho0drrsz39w6RZZ9sa+NpoDo9frHIG1noF
jYQfe+YOTCh+HQK46cak4aueouQf1J02ErEGT31uJ0BNVUWEDeQp/lh+SS0D1H7n4CwNamEI62mR
lRgY4pO7vvPJybsnjBFUtf1H+cST3m9xcKi1mBpQ/giD5wIdy4ZI83vNuxDfPbuaTETE1HeT7SMy
4xgDinJK++mKAGs9XNMIzty5jxdK2+gRLnCFJPNZ5oFrSS6qIYjeIltMaTEVljzTjMOStK2ghvxL
K0Djd2yH/uPYwAnSmP7uHvghw6cPbjZMPFUIIxqL7+BGSrwOPZ9c1bEetkNi47ajVUwoFHtRWhbX
UVC8DoLskTVssVAJtG57JZx+S1W5e6KO6b/A4f3bmoDciKM3l9XM7u+BCvfz22XowCgVwUOLF7KE
gEocKMrJHhqHrdFmNmXNZBJDlHlGU1eduu3xVPdc5hR5zQvSh8vubVrhL3lrLdNU80kzN2FGw18f
LC5XNfEv2OKSJ/B9eOaNkx8vohilzt3coOP2WAnvYx5/Qg8Mcj2an5HTsNCZ1Ye1BOIMob5wzYLF
TMPSFxQ68xfM8rCtn9LZruiMYRcfEwtWxFX7RU2d6UFK5wBqEhTP4mIKm7/UICYb6bMWJqsNRrzL
R+GziMiiuXFKAlTk9uGy4NBPdsR9qHE8FXJ4+ko+ozrqI8evymnhxQaQLTSL45jZMA/o9ebwnvJY
h4FDUyzqkMNgohcREau22QGg8h7e9FK/pqvN83kiGEJetWYw9KNbSpo0s91/lkYuBU7JsKtkUPAh
mxmNbEyk1egF0Cl/+tv2wV/bTAnUKADUIqRaiAw65vfaJ9xQnacm4XqXo3qBggEEbm/2dBBF3Pl2
/LIc3AzotSR7s39YGwowYUX8kDJJZUTL0eBX/A4d5Xc6W3J4l9GdPP92m8YL1zOLNB6WXFKrN0je
feeQ6K4uuVA/zVYrH3O/whGRsl2OJhgvKTKIRtuDv1mSjfp73nF3qBrYRYoCrFK52Ji3DA4vOTh1
Oet7R4YQlmJFxkTI2/pb6fPqQoJKQjDSZ9FHnyr9CgBk22IaMIfrEI9siCqWoh61fOD/a3pN4WfQ
j+0yI7dTvgd+wHBHyMUH/z15t5asNOQTSClrpmVV1BGb4VTpS9tyDmYPykX0IWHCiIr95NVuPUDc
fxSv+WA+ErMNQRfTNBELfX5f3ABoWfnvAekDeijbFYMfFSHW26KqF8h7Dbma/A/KoJJoI7e2EUlO
m+jseEtSaQzJGhPRUa3MutqKxKEjTaqSj5i/6JNp0Aokgtu7fcc6/rBXnuVvSn3EfYI0jq0efN82
EQWrCh0mmbe3JdlcMU5jdfMpHwS392gBuW9jCoqnO1zJtwMyIEsVDI9jyUIo3lblC/F/tPqRKLHL
Hr+g7y5+seAlERFMTBMG4foCKqYp/wU3HSSgpe0KqoQm/cPEwtvfsSW9cbQ87pkhfct8fyy/K3vE
lr57sjLUjU8sYIvazDNhSHSD3wN2izwUFWDbY/wBx7pvwxG5bfsZRC4ksxykdytQuSEMrt4QuTZB
Iwy0R7sDYvK+9UZ22ZmjmD2+4xbLIqMqZS5xcQFSzyolpCHHC5YCCWvXfqHJ0YU8NTBOfoIjJgl0
/D+DBb0R3OutCutKpjmaGo8X8DrU+NPkt5oTXHBnfYafpJFhqX5rjh1lLS+vcj7K3RdhwpJkrp2I
3WlTqyiZZwSJfj41UeujSqdtJEy7ZTazsK6usi8hjLHSBSgM9hLMxW1FCnlNLCb0oYFAnM76oTH4
mvyz23n0Z6NDWBCWcCXXGrFeOEZNvqy4QLYYF4DaFzugcOglEpevI0qXcMPwI7xpP27nmgNLRXg9
4CRG26siaimNSAOObuG/gsFDr9gI/oAa+nVNk3B/ogea5shFUAjGR9bT1gy+Tr0rzRt35bQOdrSz
tNji6ImFNDJrfKgo6glRer7G2kuEoY3Ea5/UOF3B9eDtuAlpLPEv/UdHJt8kQ9hBwvBdk8WWzs+k
KTIzdIkDhj8QR6EGXkvo87UGaUymhGbZ7bocCjs4o5Iq9Z91OPPgVll/Zs7tl8sXDwaodrPvnIWx
72PB5ibqWpFP/E/s6/Y2Gu6WJdLu2ZB5fgEt5kWNJ76UrrhePOWEBnXmMwjRxbiRIHpg/eQ7049+
wNcNd0w/NC6+Xbm2Q5Ru7MurKnainZHNRZUlDvWcXnzk6ch2hHoYn5UjlHbVBMe9G3MHv3A9at07
wS1jav5J4WGsyoeDwX5Bn646YeZ2MuhqXOFr0eFmmLrReHo23sL+iQWn2W1rwdkkCo3fvR7wvSBy
R4QEtQKxvhyHqb8/PXavgbQwE1yQu7OA/nZjYrhAky/zniNbfIrvrqHrxMJsPXZXIY1LGORn0Dqy
rjeui3OR2vEKtKEF3ixcpwAOHmzMkqr8cSDHV3EPDSjW2UJNowPSM7OB97fE34yFEYvFhh0ale8F
eNdFn8juaCL7GQIrMIEuEfBns9DjpvvCEWZkMiYic312fYIZnMJUBCfh/LuPwyv0bNlGIyvRZjzX
yTyxUhAcN9FqMP9526nZHIHaOLnVRSUokbRzG/SgC407kGLNagRrRw2vv4ch/Uhh3pm5XixXFbFQ
tH4YViBnvbVyguQTTabiB+4L13ZH3hoLqjxt7r4+bj2arVgmEw/3c2EHhzyeYQDW8MXllfKc9TKV
Rzro1TvX7+PXZ16YS2QylLAaDnB5Mqv5wQyNxKc8ZbiBXAkIn2lC/6U2VYZDVZcpiclOoPpMUOZ0
U2qgWUaoXjWNjypFnteHBfntGIATm2cxzt/W504xY40VuI3d2LgRESlL+2qF0DGyWF+qgc6GqTtz
DpyfOk9IGyax6yCeDIEGrXIVtTG1hf6uX0MDG3BqfLqXYKiVeVpIySGAT0MYtX0zZvHQOSHU5Nm0
jTWoB+/Umx+HPKItJr50aXdZfzbADrHDne6lJv6IaSRfuMhWGLadkn5foZJWtSMAehRdnz2ukoOK
4H+dAasGQ/hwEdVkexgSkpI1IOpsXIc0RSFZT1JeXICJD7Izmu2ze5Kwdas+guqYyxEf0iM5HLdG
z+PxJrJry+5VF/tMVib10n6LP4UjJWlEy3oSpOlbU18Jel+2LSNX4NkPR495Z0oQXnHhFtPFwHvm
HGLeZFfu4sgdrlRNuQEGazgdrtyHfhznccm73GRqmwbD6MGFFCnkXiToLtZT3LQdD41DG9FkFxdj
+EBbSVhlNE3N9fZWE2HYazLDCqWqL5tHkdDVNzU9e0UZG5PvVo30/dHf1s8/aSjHNe20QI9/R8kq
7tFZX0bDgDflsVADdWlVixnUQ6If0+3/2PDQYThYNW3Gzk2RtXEYrvvGB9hkbEdCkLkpHO6Ayjip
AnIaG6LRo+JeB7PzWdmCpTODnYt6dFhmhiGXeOhROujLeKMxipe1RCRCHqUaFyYn+06Z7wkeVB7E
rRwpKkYdCbR92nMeBmCKNQGAQFQ4n2lbo8pQWDIkkL/sI4zW8jZ/eQDMsgAqLVwdUpIWQB199oY/
qjQlke4M2D0/kgb3a8YnvN3R9mOlVraF2NTV66VnlnQgGRZnravFp9rMt3Crjz1CUX8aGWgodaBy
ZQYi2/9Q3kV/Nus7iedbeWMhn4Mtm86h61JjHd4utlqFA02eR/TcIIG++KjNc44CENrr0QHKBdUm
XQ0VqWyuqLYDxdbMiFaNp1j/KwgsSxtzac9mbmgNiD+DlYzCeboMw3LE/M25r5fX4KfNMKr6z5fB
0rw4ngc/Eb/QVKTICbXckU/YkkbieAbwQPisrNZtKSe6kdwP75dp7H1HBlGrSuQIPv3HlLNP7VJ+
ZaauqYvW85AuRy8L37diNQi0DUq3ynioavxHQsxGjocdjiVfCDfw9V05ttXKiMP51nIPX7p12UKX
wWFBdMN9PNzTVhcwUFOx0yvD3KwxmnZUWUDy1QRyjWDpzAYTE9yp2gz7lAasGvMkoA98M/w7nUGK
09mBqDxQtljtZW/g99jbUscaGtKP0LdxG+IB1wsRJfw1GW8EeRZYVWin8zBWVDgh4tS+M/WYsf2j
u3KOUM5qPP7D+WxpVDgRCweIcjnlLY/OJb8cWQt8I6UmtcJi2ScQDvDwZK8vUIl+ilCuIqIHW05j
+yIcKlVG/7t5DcuX86V6lHEfxqdnVar4Kqa4W6CtzfcCrecg9rxm1cnfopobuh57fXWHbAR/juqj
BBdK1Rr2uNMuPUJ3EPOBKzRGuN7kskqTVnz31bWOx48sf9O285JYDBtFwTvJoey9NZ4CSDgKPWna
9OCKg+IgYBbgWhxiWQ6R/vXwMoHJQHfYsbXyvO+Oq5LEtT8L3vjeSkZ+TIeFVZuvmBW38o9wC9af
KD7qXCzBP+h72M+1aG2JF+GD8xg8GbhJ8+Jn6ONnwskvlN1BLpNOCfQI2CDFX2dQYc3MYJheC+Xd
khMGFK2pGt+UJd7mVdgws/o5iMEdeK4uVQXExyAPVMuJUeAY5SfLw20j2ahv54ABWVGLG0qQdIJ0
EUXy/GlwVvXl6tmaQHGffuLcv33kyEQFPNr624IGQWBR38IyF42RQXXq7Xvoyvs1vhlBtjhYiBeU
XebOB0L2o/Db3ASRgIoOssVuasTpvJ5mbn4x4DOuEEnPthSnlTxiJWeKzEgPd8iROTnBz3J/ZMXO
Js2qnaetN3heRA8EH6/5xwXcqk6j3EcPpb+RJlcxoUsOCg6L1qAu7DLXfK4M43GlSEfAi4DvFBmw
wqZVfl7ZBexgpEvrlRN1XhYjp2oP2u6ZI1nljGj/Jiyrlw6e9BxOX8GYw3v7/nkYC7sXEwfN2HRB
CHjiN3FaREfcpgAD6o4Z5pXZSnkDhvMWIx1SkJX9pmOv4kgEIo9ST8vsAbPl+LUMKKN6/nEsSv24
MGl7pCWgEOlNhlMztRcSCNK70xmU0ixJuz9BuqG8vlCU2MoXUig2TkzFwf1Jepsgwq/IrMe1GYZC
GB0BQBJQY0c4CcfPTnrzGX75FBec607U3VyiauGjywJbtvBikXGZGgHdCUyA/tsGOaFEfTA1pw0j
2MlDtGZkN3s2keQ9PVcLDK0cqbhkvUNx8vwmKGZRGZYKIbuP5YirkiUsuqMAI5IFQYo0dzebqBua
YSLJC6SLu+Vt7NEYifLUz30rvm1TJmeVf5hUyBWL4JQ99CUCTeFpFFvvpsPDcotH+h+LvXypU8jP
Y/5UI7XhgzRAuzjHpP/CYCGXBu9cBE2Glc1w8wZDXbpgEZnxiZhDmL0Y8cqStMBIKbeI2s1Av1FJ
cEU46zt4s8TsWnJreixlsMYvaDCdc00LDkMTKhNrzwUiAi/NXt4WHzaeJEOh/nHToSULJqcD10Q+
kHeJpmvyX7sGQB2eSgYX5ZMvP/SXMbk4G4d2f9bdlc2QZpcSF4q1uJ3v2QAc4Eh1wdftajrvUYIf
1C5STAXqjoCu4RUk7UY55XymlFNpIGnU3M98SzJc5ctqI730e2pzsr7g7B+DKFVo5XzULvAwvuVH
D6JU2xICRsdoqm9IXWXR51sY7WC579bUSMrp/xT5ZdAPLzeNVKaXFAy6EiO3iWXLcl3LdC5Ul19+
INoAXDhfXaHLH3O20Ks3mVA4NNPrBO9SpyMRn4EIqNJ4L8H71ccjrTQ5mAGONDvyfvVVShFc8XOd
Ptz71l9H4JjQLeutHSL6PCFgMe7CLSr/dHLkX6mYcz/F0m6YYowhpmjXVwDKR8G6CVPWyboVobcH
tHsZileOzRL4e667cy2DSQYHCycQvNAysAoMRDSs9N+Dtr7Lcj2ES00UPPv1ptJBnBamqk0WLby9
WrJKwnxAsOX3ScPHfwJGFqGz8/yz+aGu+V29vVDszMFDfSTnxlVjbMAbFA9uAsUX6jDTCEzuaCUE
Id6P7YDDd3QkbfA9r5/0T5breO8ZJeQAEUPjNYZ4FBFbalC96fwko5vFjWlPWJcj/YzxmxbK6Lbi
poPjOOFhfTHGw/a0XsQiGuAzuAtOsUoGkh6/FQWbaXS2bYmKVLjG6+XP9nyB7qElLgiOZiwY0s/F
ShgDYFLU2NJWcBjz3MdS/bjtFi7+w2/BaFYc074hZM/Fdqzhw0n4mFiBWbSw8l7AvKU0rzSyi1xZ
Edq/uC+KVUd6zMHU+ITyLgH9zXHEiJOqAAoIwgaOBLCHUw0wwrvh+PBm/jHq7YyOHR/chkJBopXu
xecLXSmsYSi1lWK7CXjRQUAKAdKTPuh7dKFTn+bh4FboSZGo+3xfgTySexwIyUeOv9VGqVuUPOZI
7ZVdSnAkrmmX5FmuX3Q3oatXvXWTQIg1DHm6gTIEHF3KsT8R/dBC/ZrVv73Xi3LYiGkXy+ZoTdT6
45cKo8bm8aSczSxgYakWVd9oswuCDbZChrKoaMJKKW9eSJT7DrFoP56tXi7F9jybIAK8O41NfryR
PJgpJQQEA+jTiq2R2ao8oSYQ33WPEAshtOcXvGGwWTaSX1cvjQpkAljMvYT4rgPnIhA+o1ARZ3sO
WVvSfWuKMUBVL9g6msv99ybP1YimKQgIp3T8PoiWxi3DObxbe3iYxA8GhbNerNpz1kOB7itBo5+Y
OlcM3wdAbN//SBDERqbuE1952yg6SAYMW5HfDlvymdtzeESQZzb3sXEDV+tNXuXZZIpzPLidKt+l
2NCdwL3GBiL0DS81JQ/s6k3j6BBDIUhg7gG59wtZOMjezr0MxkLVH4fC7Y5u/+mCDZnGez+Kypoy
6fsAzJiU3O7cbqnEwQDi015TAI3/6anuoDGuNNJXJlTidVl3Z3LCOjmEmBZp3nsBMJuBHFOMK9m0
RysgUoEGJQluTNQjj7L2Jn70BOh3KTNAeFK71Rngx1TDc8rGflW6ulRVfp8SX/jRtNhzm0EVkHk1
e0gc4J/EB8UstZQu97RAJVLb+Sc88Z1EfUb5aA3PcL9j1QTOLvIIvD7nIrULsaI3CzWIX8UPPBHI
4ymZ7xz2g5Vokr3NmaOBV9O6+jfXKGwdRoEid82+K27e1QyYFt+vitYskZ8kEtcfo1OlBDt7Poxf
2dI1hEUh7H0NFQZNGfWjYMkLJrcLpjkt2hWZsVP3V0oq45jCQGrTrjYSi6KlNVZtpMAONiQsSEtP
e9tzYsybbWxdAdjZTxiQkg6Tw8kcIIOj9QppO94R9d3epm+nTh1mXfZtNq7FCI3ZEOeUsqNUXqyy
9F+ghg0VG4KvJWBbhPhDjaa6VDIhK/CFB3l5m5DnZL44RbbO8C0xCJDtBq2cTYMPjdAckuQGRA71
qCwk2TISZf7Y3f4F4fGr4Nj6QT7OhJAP0WWMmPj6CZikpWcqsS9GvOXHh6Jgv+wBaqN9pxfDDCGY
omgE90NqZvKzh2PXcTEI2NJUwpUxr6KzMHVAJeTA8vlTsd/kWsie08XOV1tU6BRzhzbSSIUdMjYT
G0hCP+EtBI+qAI527ZX6m0w/pJWMs60lz2+eXZPy5vl/jY9LgYTrpGFk/HWQfzXnkCcIMjHKbhGk
z5vz1fgtuTEbVh5xH9+0/ioV+bMqCNgSLjqb59flTzg3HCH5h+tCjH3kb3g9wP2TEmtIfMuUhHSe
QunxeiEm8L85lVADzQ5Du+rt1aNGhITafnoN1l3duHnTgXuKVtFX/n+LTwQSVtNP35qUW7ABy+xz
9a0Htu0nHKU+wlSEvy6H/GNdeaZuxMPFfCqtyYOlA5p1D34nQ8MC7ooH6NpTYY45qwkrkVSHc+CW
bQxyTY+KUdujFVjWf2O114Wi1+ayFHBTDI9U9t6qsetT7mUONOmAKgaRgR8tUp6xE07wA6osBqgs
rdVnWqa7FVdkMIvvzQ+6HsNh8iD4za5oFksCLjM8NsSISUFmHKd+CWrsPjw8Yfw2RYTHgPkMXdIp
OH8OvEKPS9I9EFuxZQdWEYDfPnvQk8rTfx+1L0FamQ1HR48q57EaLHtFL3EUqtDt0eaBYDOda2UN
sdRYyxSazTr95JH3PoTkIyVVJesNLVQrWBvZXmK+eUekqdJXw9+KJKJyBvhgE2UdzBiee1VhDOU2
M3Mctfy2LCB/VcjthYTBdifgfK0s15Y5QkEHn9bSAihN4phBKbOS4km8eoTbipFpSKPrkaWoEdKG
zt1DfRx7NlUbXh6yxBKgSJ5l0HdScr54jslGHpqJVzjEpTBwvSU4SJu9s1f7xCWGAbtyG18wwzNi
/Wfeo22rCujIUGFTWtiZGWZLt4M0CVYYug/D5Sduas6OIAjLuPuqeI3KXKSaYsLIo2Vl+NBe1x4/
yy9WJ3YOQsl0TIDTAJtpW3CxS7JCovYr/sn0lbRqyHOKR7KVAAutmZWXIDsiR4OD7xsn5rYOmCYV
ESaxTwcjxzOgepw3n08KwRAmP/WgIDYkMPv+c4X0SW1tESeOJPlYw1Vj8AmB1pQwY/fSLk0q+4R8
YTVbPlJo5SGuRBe5TxadAbpgpScIdAZHG2rfW5UCPnQDLD7js7RZEAKBvb0H2dxuCJKvDT9waCuE
70Cv1l7QEJpIyNjP3TSufUVMKBfRWAXI5WW8Wqb28dUhj1UotgXiBICVNfQ+M8naO4PF0pvxPcSC
JRT6kflJjNm91ksIKjDlIY0wYemnVXPTWzLavizDxO8ZVjcLxe/ZWJnNXNp+va/jaMXvM5L8EquV
p82NAnSq5fKh3hJBIa1UWQVb4BzdwBFcObDAvPAowgG6yyuXTpjzCbk43NN07k1nz91bhMPwcdF/
6ae/aQ28YihdIBEHtsVJ8myZyNcJGzHrkJv9qtx5cFFIwGXulPNzEoVk8xbqFowAhAqKsIsixEJR
N6gzpydZ+nU8avwO7p8iF6YgZrAdc2xeqEna8qr++9wrOTN2cFLEqfMvIWhncNA3JPmGIeHrCcWG
RqHYrGwjJAO7OXjfdr1aMekISVblywrjcrzesDYpKCGmYuxXR4dYOUEAtLozN55ilUdkM5oHU0e7
IwFXOE3o3lTlbt3rnbM4yaUJusSVmOgtBV5yDhR2oO2s0oWprtsa3O4zvl/Uc5DBzU210jXz0sA7
oTgbefKW1pbrp4Ivl1m3AHjrMI9fw/uPO+nt6ZIoL1mrsWr6VJAKsWoWfJzx8qIBEfmJT0oAhyDi
JsFN//hNNvwfOf6H2IPtN9x4BkzZVmcImIGyOWlyHq9rg6g843Pbko45lcDl1PYk73EeulNmfBdP
XEJEvqj08KGigIW1HZyh8LYyEjrIKR/RNglFRsuvu089zh6Vg6jVCsEhadUcRjLrw4l5BzEu1CvN
obf1foeW8Yw9wmlhmzpCiyWtWd3erfQRsesy4Dcj+8jbCwKW+4/bdO87C+be2MYT8B1qh2FVYcrD
1SHW0yihWfrqvuH6mU4j+cfccrrPXDOBzNLSuT+ZKftscqtzLTGyiUnI2DMeiSwCnitFHCR6QNJ2
U8vzulfXJBFATKqdoJI6h/On97wzLMX3qQAIXtDDouQqHQOvidYpUC2uenp1O0Y7yERZ028JwYUL
2duwFvLgy4IqJVXsYAoMhjs0Gn0+trUEsFF3RmFcCSgJe9+8VufzsUM7vqkzoVRj7xucrOjQfJTt
6b+88VqjE6Lc6krutg+zxt9NQ3OUZ17GPreKVvnqBHPfVBWKLkijbqRV4OOIJSaU8jnxnmqz2EAI
3YIYHBmMnZC8mFUjpr5Mswu1l5B+CbCQKLzPe+/W8dkxkhS3eMjcGpdeU9zswHzx6ZiS9KJF8Hu+
IA3q3b/hIyH1YfuJdIVaItop0TXk6mD9uaQ6Zhq1Zckdo1+5z63rr/zx5khE650p0GF5iBgOkQ7k
K+PnNLir39/uZaG/EueooQROrTnPBOpp5JixTMfhX+XigxFQWE5jChWCGYQNrkfU7BAlDPGhm3sI
SJYoJBEiKKRsuPw5yWXcSKCExW04S6pYfwm4n23sHEPuLz3jzIM7aPjj808znBE2aylHiI1ek6zF
qFmb7oDrS82D26T1v/8zWP5+CRr8TRDuMTE2l3+1SjrRJuqMITqAG9ve/7lMVbexjg0D4/8U6dpO
q7iqyI3eohhBTvpF4Ip2E0kqbARZvxR8uXhVchRN7x9fIxB9zDOCL49qg49ac3LzUiCyui78eLPX
gaRp1boWbS45gp8zpOB4KW9jwiVPKydSCNQQdCNtD9qcXpDwYBgHFPItkgM9H2Uc0OFkGorDK6qt
tV6VyyUbZS11PiciyIJJ7g8IomPPPOOtzjuhpmsUwDRU0uo52yyGBg+1sPy279aUquje6PZnTjYb
x7Yd9iI1S7rGZpip51PmprNaUzPlrLHt6TOFCmOkPxg1k7tnzGUH1ex4qRXgtR9viHm/lZFgA2lw
BNisNhq1vGNoRcJ4CKZaeTUHlTwgq0Q5TdNt1zbbc1mTSO3zP1FLL0tPPCMQgGdQaQZtZ2PAethr
QXa2HRmQK4otW69oYWfr9obdZoBZ+6vBVRA6R0NtKkkSKBUhY/1bT0it8583/iC14QFRkyGUFrRb
931V3L0qxR8JvN37cHLYQZulUCeFXGHc/G7d1lqqiSsXbEWIQvUQH6epTqO7m5X7p0x+p3y2dg1Y
Z3cJJciuNdqV/Vz48rjTTXnL1Sg6+HnCIoCjtU9BCYmYaf5krBU1BmGqJ7hFKgxtp3e0TUISc5ky
HFt/K5ik1MOWkht6Jo5TEUybZYeQHwhq2t23RurYrbDmpt3xulVDJZR0isJ35+A+Y/8MfhkHi7Ga
V9lv2C6NulI+/ydsdkGEY580UowhsMqlBdokmWxxw5xcbYlx5OGOQsHNEINoZ+1RGli9xJYVxcv0
9IDl7+LSzzEqJ/rsBLPW7Pm4nyo2zN4vDgAXbFQSlU9WegHptHqJHyrFVsB1L56kxIsUb27PpZJQ
HcCiJ7UxU+8xbZ5cye9kS671Iea1GXA1eAql6KTIJwiFuoniSPLm9R3Baq1S/tRCdHLZhFDxJ6E1
CKhv0s+OlZln51FJBm3B/jzKsGAgc/1/qu21H1KbrfnfGBo1bZ13+WGi7QmZVo8Uu4XN+l7vEY1G
W0d/ZTsznkwZuSJdotqt1i36vQDTt20V5xVPgWNOgsAkp5BgPCG43eIaP8soTkUm1rmALJQPNq6Q
j5zokx0z5Gk81bPkMRRc3v3bBqJr3MSoOULee6njkOGhX5pgpb3xGEyp8bQoCdjrg8lhAO6l9meR
4b4Nr60iKnGBTu2ybQVXakdOG5ymwiYGdI9nSaYH9cZhx7t76NLEDotIfOr89JwZWnp/w+XawRfc
z2d0EwETTLdy5+FJFsPsjlPL33e1R9WjM2WPf8wg4/8c5H03dEkXvr4KL0ecVWv7ywwnIi7S++p1
cjIHV7FFd6fOWFbJG6dx/jTxQBXikrsJnTv98liGczHiIOFzshmVZwREbMUAAXzzvm6oq5wT6vDt
B4IynpiSsO+3v3mxC/Aqg/13blhMXqTprGIx5VR7Kc17e6H0TPyqaqzI/rQrz53YgVYg9C1llcgc
gXl0GmNE0pIWb9rPzZ/S16UweIZT95Lo5kSRBZYDGTqwFWxoQZb4t1s2Sp0EpXaVNX3wmRmjTWSn
b6G43b3aRB1VtY34ay/MwTPaw0ECJ1NCuyIPhMNA52pt9j4B/H6wRr8pzs3mJwDJQjR4pitmTWNg
bgPiLG759WIJS4zzbeKEs9C5ujlFgbJNq3Kx0x+aVlQu7unwDQDg6nwTTuPLdpd/7DDtz9KZ8ckN
nxZBlDKB209Kzg++qlnjZ+u1j8Gd2o6BiOxdbms9MCOEx+n5F8WzUEwnNBmm5S5oBAHlf8qNP4gh
dd3AQqemOvOgCh5SBcgWIbf44WgWZm5s4CmjVnCToLHZG76W5CHtfsdvsU93omvCTfSJ/3fMP27M
sqr40S8qe2xmZ+QuQQvIXJGHKEK0rUlQmGVhjE3jZUkfaSGcV4+esR6K80Sc3CS51d/58vF1JvFD
FqwIbeaOw69H1/0Jw/KrM3LMKPWLPSd24Q2pap3vZd/mFJC4WI3FAyDUiEPPgGrzhp94F33qX7ho
u0ZFgocyVC4eZpdV2TS0LLhyhak4WHX+9BFkJ68/wMKMhi1YIfs0ROWPOCsQ+mew31sQ+Pk2ZZGb
UDrc+2SxNPWEWv+A7G7mDsJuDbRgSnUAn32gP8VjVq6vVivKlbwqQaC/eiGYRfur6NEKE4+4cSAJ
M9XbHcAgC37p4vJs2GbL+o56Tut82Mz8aRed7Fm/KThqI5l8SB4VjzISewEhaV/VkNRpARsh1mYi
3vMGmXXg2Gh39dnVamqQjG1nFk6T4nU1iOw7/pvNBhRDJ58QACzHSUYqMjX8NEBNQJx2QRpvOVir
Zr1i6uPFTq3TlhmFaf0xc+PbKWw5c9xBAK2tIQkG4FfpgRAz/sYYAwZuf9zsxqb9C/BQAUZyE5VB
UpHtS6AI7dCjaD98RnVXgkiTBHwpufZy+fV5rrMO/mPQxGTfozxOtJuiz8vGvK8KeCH/enWgzJNo
aNzTKGho/AMbMV/nwWnv35Qd5F0rdVTP+X3LtgQgio00VFJu7uanK39V1z1xLFz42NMS1/KMi2r4
lN9+j8vnW6aRshAw/CAar0iaNjf4IovCuUvFqjD3D8g/IEC8tSyLsuW1bKPVI6Q8oLnw57feuRr3
v+H3n2boQXEY4Oj5ufNA8++MIKl9P1o9lvtx6K5YP0Fipp/9jr0j+8+s3IdDjUOsudYBLWdd9fhx
IiiuSyxTi1AhCQ09Kaszf+5PSHLyzi1hh3uFW7yO3C1UZb09g7jCdoDG8p5RCyDXOVh6bcThIclV
saw5STmpcE8T4J9+6LrjamaUF51GgCKcwZFuVrPeruFz+3wv1KXdO8mo+8fHOfI6ixTlBuBiYEsW
cU4FOBu5ROARNa3ck2TQqvAa1O00jj932on91wCAxoIoaUxMhPGlt8EZyaO2g5s4QmpPCwikEhat
FmvKERgt6lv6QgtPB8E5DcoUT04A28BYeOIruDar3gGb60RO05qZJkZDixXSai0LmbaLeX5XoYZQ
F5oeQtDrlO+MUpsoWY3JwPZMvr1ZycJ/F2Wl3SMm1jmDTQl8YGdg75F3xrpnrHMa3a4JptkZcDMu
fipBsLFVCPjc7jlV2AXiO6bMUppHmfD6u5Ks2Q6Q8xJ6ITKyeSRYKe/xx/BJMzea9MZ7KCLDEBx9
JMcCVWi29/ji8zp5W/DPPZDolH5zf1FvmiNvrEAhTZy4nb/HDPTukPm6HgtSSMYCG4T0RbUWZCEH
Cpv5rf+loO3iVj1/TDPWjgocqk9GvC8Y4kjp3fEPcRg0e2S4KqqDO9usgqqTebMYACqcju9jXP5M
h0rhOJSySZxfcBGliLFJqntBp8fys2XOTocFyTzyMrTaRdTCf7o0vQu3rdj+na/UzXF+6HOnQyXL
XjrfTtdoxryr/Qb5S+Qe3HOkBzMC/DC+quMHQZMOyyanbPNscwv7tInxvNS0qoZS3MSGaa3JhEw4
SYN8SDTy3Hk4aFVgLseV6quxIld4o1jso1AxCBNptXsH3CFNA7qv0bWQWxpYkOvJXYVVycj0P7XN
+4iBQ7zCMQNLHfEhwW4JWCWL+hSAGyFURprlKyO7tTkB6yg3Ibo8B2eUs8I165DPFoJFYeE7+x21
SVODZ5ArL3L+PLqmDMhCz/pG/28V6Pr52T00kKDUxoPb/NwN0k9NQ6jH41NyNK1icP1saTyKJ47x
qokD+0lHBQUYIza5wUl2tzLTM82mtMLvuYV5lIb8+Cb+lmptRwD+ZrlypnMatDp2xupvUkOM5Abj
UnVV7Mr1ZqI4RIckijA+R5r2k4r9iW4TWjG+Gzvi+KJPWoKqa3188nPN7x0ntmcUjPpTi+HbcmdP
OwARQrSKCReCJW75VNRUgh+wcubsQyuHI7o8ZFUxAgcJnnmDQIMfNCKJMu6Klj9XxBufG8LP7bRj
coVuMBUxowvwoUZblETzmR4B0hdThiO9+LcmFgsC1DEamCjPUKWkqWU+63lt6XcbrWLA7Kc+yi2v
QyZ3qM8EYqWelrRTlpZETEyI4pdn+5jdLkVSp7K+QJnq4qbvCJapIOzP6RFnvlyar/c92kpQc5bB
sS5MqPNfsNN6+buAJBACsosXr3RoU+lKHATYvLY9Nd6AaqHgjHTxZvDiQ/58DgGv3nMcs//mseKw
zPozEwiQRVPe5Vy1eSAJgkx8oP0oeOOudCKI1bQl2Yp6E/p62/m0d5+EgS/0sHH6ui9jXYhQtlMg
fgV/3yOuAVPLSFXSmYMHnPtdpYj6E5M+XlTc0e9zlm0JciUOAXdbuU13mZJ9eajoNA2U1h/Vz4C4
YDmjtNlpsRmoivMM+am/o6GcNvyU6nm2DicTA4lC5MXC2MPchEta5220FKSRQgERZdvUjW/VnrSd
9jxUpLGauS9F58RAOcRNU1poYYAhbs4gUWHT3c9MtLm5BfisQSoFEzesqOro+0lR1ZVwLyD7qfet
WZAqXmw6ujESIQujfq4wpLyqOGFNLIpCQcTezhU9b2f51mfFeIQR5B3TIVgCVGuSApYPIibc5zpH
rt2DOzryZ0vSSeZ/+a5SmEIO91v6FP2pH3Db1NeAP2EsK6t7TPBXm6cVOf5tufkCaU1ksKwUCuly
NyiWpPRabsyOzx7OQnPtxacIiqciX6qcqwelZlNqpgIW0Iu2eA5Duloup3C+KjWMrfsqzBxfcQuN
1YAygeqpaWSp4fgH4EXQ8mV4jEFYa4zZdcG57lLkXKNFUWDSqCw0BFTRvqxHkkHmGkGKm8/zOI0R
ThORY77Az7M1ekw5hP/7+uehaEbIrW+vYvODjoZWkSenaUusROvaPTEDNXI+O2R9pJ/w3no5BE6I
FI5K6xq/J7amUFs/0cAie/xzP0KrM4YD45WWbxEIijhxJaTbCVUxztHsdsjRei0SHe+rgD8lhDpg
tB9UuZimc/pwwzRl+UwJ8xdpOD0ykMprGpuhRPj5d9jSzqGtOJJYN0Ymg4O9hE7KXYtIDy8zJzJp
9+Y2ObZshXMzRJ9xot51oZfU4Xz5XGBh2xREXoBje3G7OIBZcSaGoFo8j6KLJ5KYNI0lKcEWQ3SO
0VT+/IQGBn/0qDsuNrQZroV54tb+z0BjM+7JUIvy0YltRryK1Oq0sIhgUNmlcfi++XLURJF536B3
FfciEhDGa6HB9Qy77FqO+7UXjz1FRTX8eame2a5kyNDa25Y7MppvewTIa0Ph3oLqjpDXfeMYTARN
543x03I6EBXIXCBOo4oFBtB2gBXwyZgePkWGLO/rL8CehRM1ZNffKb+SsR/DoLImLydpmWIv9aBj
Sr/ZsIY6S5FXMpzFEwFWmef3VsQ1amDQ9xMEFYvEDKJXlh0JNHnvc0PgimPFHq47smBba+Qj6PUQ
Yo6LcSjhVUY1lfxKufve7zYo6Y+a2M2EqSx8UKh5CITMkYHhQe8l4Ig1xk9efJTt5OLnbhQiI0b3
iwH7LSgTnA6NLacXfQlQfnA5crMypIHzjoG8lTcNVyWqgKb9DHrpKBEj0PX2KglEFzX7l/n7hr5R
6cd3fe3KnGTCLoPAXtWiB/9TTt/Sz61z3BND3Etg+lexrHlf/66IONllGj7N85bZY+lSMQ3a8SS9
plO5jeo/RCmmVZzp3jKFSfx5y9yTJh81v6L1tU09AsayqUzQejGtuts42/mLQNA/LbG46C+LLQU7
3OVx8QIuCUir8+PZiViw2JZS4IA8lg/1+H7smKlLT1O8yTuwRw5Z+ApkAQip1S2u6+9xpX2YOd4g
rNNGtCNmkSbCm5RXAGOLmDzsH204WdaLecZzAN48DU5tGhL5ZqkKngeDqdwNv4ulQaNstdVV+xoD
RiB7zD6lIJr6bffe8QN6VZYkyMpLYBJ9q7sAQlrmVgcnEyFnjQqWxAik0igrtJ0GMJY/eK3ynTo8
mwUByhkr5c9p0ToW557EZflB1sAqjDVcdCQwP3PP/FNeLiDGTf4uwKS1r0RsetNrFkcp4SIvcHIP
xGg3am5tVeW+KCDSaxV8PM98BenPvwVXnXrJ5uiN1tpuxXUhjb+mRBJe/ipkVy7Yc9EZqdcMm38p
RjkIw76GMQQMmIWb9ZQb56j1ZDFJ4CykkKJj88G8+f3OwD9J6JtCc4l898ZMQNlv9C5ZDveoIk3s
W+ebefexk724YeVIwLbRScrbPJXb5Z74SFj8mW2vvIVpSgyAK/sPbDZWv8nHpMraUVcX1yadpgai
M5B8ZuM6p6ap7q/xeeFLm5fN3o6XHsbJm6E36z+dtk9DvqqpnV8cBp94h0cqk4JDzHOpsX6i00Al
q8ZU9sycqf2cHOK3OHY+wqjQNG5O2Ck53xm5wyFowGZIszXJDdYeRKWwDND8hdGDZ3e8PF0XBrNS
yrwXEjMHNW24cZityjdyKCOPCsLHU4JTFBqBFV1yp15tDlapk4wlmUfdVsODmCVbkt4uWsLkquYG
K8bOBpiCluMsRlOZuqoSknU8zgQLqlg+IbVHIIVIJtK5Yh5mdD3sPBk+/2KmHKYn5duVAywev0Bf
habXvFq1Pef0FJaK0Ont+Z2KbA4lTj7qyezoNbBoEY9GX1Je0SPDyOLhjnIVYtJ92ljKY06Dl1AR
jAwmnDchmYvSr3fLKc0TbW+0ml7nBjvSCR+X2oH9xic9XB9wgCZsKeoWFW371YzWFmEaJMiVMyYH
bl+YPqM9N0vPoSCi5AOOSiqKbRwjDgjvMt32FqmZXjEBpDafQS6ZnaMQBAEj6+MgQ2cU02s+1t27
iyiGCxe5KfiCjnt5NOVgcl/ZQ2jOM5XFeImnkOFOLf9WjsKtKlpDPbCezIgqddPzFeoYqREFcnvY
EUlqOznN4GuYrHQLp62kq87tH04bImWNkOw1ZFouzuuLKV3kVsZZY7MqVvovaiA1z2VxRHvS+MEW
cZPyg+RunUmixmOmvI1nhs3lBrb4XcJiE3/q3R38zZKivt3dbDH3kgk8eOOvlq+vvWNEHRERn7PA
g2HDg6jTyGqfnlw6h8lrRcF8pW1c5hlyn+gh6/uyC/yjBuEqrmVWJ1ls4zYx/FRe0lNb3qoxbJTl
2VuSAerqeyR/V6pKkj1hcGNnYydPAL8+yWOuLzARIcJtR58wVMC5K7GVx81EwpRzoIGavyzkRJPY
v+zJ6cRw93pR0y66vAtodxrDSbTi6IzrLWo2H9FZhjBK0K+aO8e1y0ytOATE8YQq+lhahDJ4VQdJ
KWfiPaldY8+ADpV6cqSzw7ZZOq2i9AF5TtyykMO1cSr5WxjI0h97iNSyHmRPS68CeKvzrlK+G0jZ
kXdyrCoiKSFnq4BCk7ybf7pt/1pwIm6wG48xyeeTTZpOIoaeSR/GVBjrKocoVLR8UZPKsRqQV6KE
TInZ5P11loCrPTqFJrfwLLdJuZgWj8DJKY8mpsgCqPhRaSsrx7G1uF4OAjLYVMB2ehYAEygVdh1K
Zoso4IWNG6bWxC+jyVhnI6pbVvKAA1xxzFb1rX+KD7ZE+veJRLDALGz2sBCvPDE12/8B0G+mnTrx
plxYGRDn6A5xeemtTD5amCM4m29YykamaROEZ73IwNxMw5CLgcc3lAy1hkZ4UxarqJAZFX1+G9E4
DKGlAy4CDBAlywJ0jJ29wnWqFZycOrGsxpXPj1UM6b4RdN9/kC0sQRC16+C3dkoQMs/lf+0iKO5N
myYm0EA9rY5t0qSxA2PYUKsg5FiQgsCHueL3l1fP7yP0fiyZ6qUqWWXeqXSbLIBXKsw/RnABCybK
z2LSNMFERPUvA6v/JJ4KxeC5VUfw41Blg2+xsXL6vYyo0+POc/IHfGnR6Pl7bEMZaDC2btjGL0np
QxWNEY/jEbC4LG9v/BehkwxwnIyCci1GXbyWrvJr0U0HPb0JFgL/7FCRgbNVuvqDfPw2YALbXM9e
VshDRB+IW9Gk+s2jYnBjI/auAN1ceja2DNTppLz/Oj+Ylok91s+bM2BjsNBwTcdbgkQ361wh8kPG
7f+cNOIJEdE2YSvU7HDhoeyOln4yEM2X/HkaukFpIaJYHq61J+GzGKf+Srvi3osj2zMC2wKN310j
lPFHJNEC2EA3jCTSVKeytWbHKjvpOjXCs/Dbs5+J7htwgkkJ3iE2zG1Sn1+S6lpx5WhCg1FRY+pO
NTAoHVDgmKLubRj7N/WU4JnM3QfZ3DlsKg3jFPmVy+QSTTjwE3M9IYRrw8jQCbgXFllHh9xBvZ/Q
dGFyFWjmDYEfxMUHlVxEd4CswjboTU/djX9Ut7QHP3ikSrSAPZdUIb6P8HEqKx+3mbmwXzVwfYZH
g5FixMZdb/sxfgm1BqTNKdoAXaU/51rpcFQt58OY2Z0UKISKGAhXTwxNxYVonJULhP+om1dNRuG+
Mkdbcuw9X66A/lFotzLVeHMuuzeVLL/zlKhiCi8y/LNq4ulcORVMRFACoiQrBs89GZJeelrRo/Cu
RW+VWmHks3pXoPvdSw3x4NjVsLTbOYv2RTT7WKn+ZmtUXZ4P1qLB92g9OPZGzXTkka39clVHe9FM
2wneQhX8GrcRZ/lqy1an75nurCB/YGDfmJGSCxOMt4Sm/EtNzkUZtsvmIJNJ6gTZH6vvUPu8EP/9
sOJIOceNPC0OXSZzi6C7NcEsWaiZwP4Df45R0SHyQ09Dd7d7UWPPqzpS94UNJQtDOEtEp+KO10D5
xIeKeUKsAtwvKvBr0vsSWzMc5tCFu6I1/tOwglleS7lMUR03OEuqMqTRQNDhI+H4PkdGT3G3zyMm
5hsLP3jHZhFkWPP0QcffSM2AWwx+JNa4+4dSIK696q/FmDcZa9KvZKVLdpt6hMfSSFYuEaDcJ7ik
GyoeVj0qYgc0aZcZewbMAIJZZHxNtINHRjODXlflhP0lrpHJG2kxEd8AyeLYWR4lp29cjhUs4fha
zahr9p4iWbAK9RB9EyKDl4cNSv0BC2KDH3+7aNAiZpVf/a5QfoujiENSd9fEnj9tZroeeSzC66Z0
j+E79DO5NJffGxiIJV7eE1yxyLi8yEwoRzpOgoPQ0/Df6tys6lOoE/hOK5M24ZwisHJlrQh0NShq
+6VU9u3nFc71lpGzFQQtGTujgF/uYhJSHjWDsYB/SSsi1UsNQF0h1P7oznFsVyS4G027wdw1sJmm
MxJxC2ZW3RbqpVFMRdFNqdvEifYX8i8KYr9i2n6QkOKKjVRShDcy5ZAeIU084hQ3+i9+mo/2Ysa2
adIRBi/fGty5oIe7C8pXXwX1i8DdDWeAeZfe3/knH07t0mM5+Itx1jjlnqFuvxs4TuEJgHv+9AVu
hJjy+IUkyTx6CoagwIVM/8OjF7wy6keR6n7xXCTGfWHI5IZHY7VEVsdcU/ZuN/V6R0gnPM4rlzZ4
4gg7hF+MoBqJs84XcDKF25Ljn4VHXlB6TOqE4yBJT84H+MChTdeXKrf6iCNylz+cCP+z2AtcKoNx
tFEYkGb+3H3/qf8G6Wr8EJksCtQSLLtWk0VgOT2V0yeOIDAMbK/Pk+fSSJ02le/Lams2+vzaYVK0
27tncEepjoBldFyX1hA8NZlJ17nmopewdKRC55j7cFKR07mBhvTDoe9ZDyPaD4hgpcFSrITrMYJY
N1LcTLmcaF+tZq/d+X0fDbnRr2kRcOl/qQjxXVn2Vp5wpdSE4cksAtvyyGCuTMrFVGYtXrtaY+41
OQ936o9E7Bum4x8eckKL8bd2tgepiPwx5KcjbKWxke+QK7I/garaDAROhvY20Wqor7hOOrUZLKTY
09Yy+iOOdDpZa2ZQzG6Ht0ggHMo5mvfkQPetERrjeARY50tZxsGENEUdT6wZqyPGBTC6gKwg6KKK
rsb5zY1z7iUcSahVsx5v8/bcChw36I78YlICA53AvLwZfhOXKwXnadWGTG9VWKAyYL1MR2sc3puj
4SGstUqQkm+F+98+8FW++HV/SSJ6LHgbvHVlSmDNA383q35TunbpjXWbDgMlwMsOYAAo2T78jG3W
i9jmpZR39Q9y2YpGnS2loj5nw5JoY4B20MCU9weXoo2in26C7pa8W66pxL9oP+eJRNQPkA/E7Ujg
b1V19iiy0Eli7zoNdQFhS+eVCJWHH3gvTyujvSrgbLZWM3ldiSnwdlMjLT6d7PNQBkUdq72NZAoO
HEj5xsemNAIIpyy/jxsZNYhNNXN21WRKN+VchO8epptsta6riqSms0lMCF2+0XwIR3xOQNZaQqd1
EXydnp9j16lwNJkm5FQTkYs4T/PdaVIaTtMOhBFyoxF5jv8BXI0hnXWe5BYdx/1J8QA2X4i2bqlq
+j2rn89fTZdTJBmBlgKrgeEtO+NenDX7/rsVS1nU/7MWzTtRxggX/JOCcAcMNlKLvgF9K6i1zn/2
4reO5vZ3suStFBlB/apUYK0PUYs/xlXhgB1WEvZawvtFGOPh0z/PBxg9nmNYRYhJ5ejeiMKypeDY
vivD2osTlCUq3rd1XQ6kAGGmnMKXa32XyvPN2+OnbZ+FvtqSG/z5ORxUsio3QAtiFEDqgEBxInpW
O91uwauQp7d9ayt/4scojT9mqpTexz0UMvL/KP2UrsYyffQ/9v52ccceHLWKlnjAS4RvBMBYbdJ5
LIU78ZrXk245zq6Bn4PKphT+rQxHE8tZAMAMQdkmHke4ViyTF4qloM1MW2wWioaTvzqA2/9hZbgS
Ejso+E4hZhU/RnAE96j95RxQG63zWy4W/CUhqJMZ0BpKhCnExFMZanPwr0ODDCTBnYwwVz1cdJi8
MLS0UDGdzmoTjcHIPr3Xqc9BMyDxNHdr86nIND9jc+FmQ7HMM8n3CnkCRnlwXgUpg439TmxtwieD
wgisgJL0myhk6Ih7qcjheps9p6diACJHSSC8bsktQQR3/f9+NMusaG2hJz9zNx89DeiVyej2506S
CZ/umsegO4S5+Hw1Jj8Py3ASLNLltcIjNvK6+QrpjoCyFci8IDlLNpmL4NDaMvp9Uy/F0SpMK+7I
4qccngyZvJCYdr+YUlryDbi9Almr/+jZhXIJlZf+poEirf7fkyM7MV51p5wNmLe05vwIh0ekRgfU
Ax0pzyyYrh5WqBrPiQN76NtC5yRTHD+7m72bRa5Kr1wCCCrjzsJSqdTzGnBhLpdxu/6JxyHBpI6c
rqsGJr324RHO0yNzaVEjqIkaA9n+lmTtIEMSdIIvVCwgjgeGzlzGZbGVFWnD7yGYDmxidxoqIuPt
xPquojYaR73Qg/ScpxnXtdiqppZLj5949/3LSzJd5+qg0N7NYuf2byMWiELXY5cR4ncfFxuRA+Iz
OUgGvVrl60sBCQd4vOcopsttQ666unmiWDkjXRw0r//xx63ttItO/AkmHYo+R6+Cfh/ODQa2i+Ay
RBTPq0ZQ1kmd3pxBEMK95N39sDpouQboT29tbabkhrOLpxa4gCogHKJYHWyC6Pmh1JlpehffwLlQ
U8ZjsnXEdUd8PGGkKAB43bENDmGOMFED48N0o+Xh2spN0l4ZYSNdwLWdJpf3tJS3YfGMm2fF4k+g
MA5GcOj6oqEN9IkP0XOMTjC48OmoR0Q/XUOdRh3cNMtmnYarWkssRoDVsBXPWwWtfnrB4NmKifW9
s+olJdF+fYhx7P/VlpdzRpqzJspCcCIVNeAZtSTKqJ4rcb6gzrUXBeiM/TdDTbdyD6ukcPGrCTNI
l4GAZqSR9cvCKPm9o45tgkuXwp60ScRucqMbtGQDqfhz3owZEFsHcPbnI9Vw7EZYcll7ExqLPs6f
k4qOOprvAnWyGlePOgGmJu+OwUeTRZloBHj72LdzHrxy5pq19yn2F771uOGEM9c/lMNHzxZU5lnl
C0WsInEN3eF0LBDbrj9B68AW9kiu/YKAOTab2pUYGkPX5ohZcgUtPII6siWrU37TMSwuZh3WCgjf
GrtfuXBWa+U0ncB1yuy2RsRgxdmSckGLveDlVqyEt1sFO2BqZ4dyprw896QvuFEI9hNtQtozc0P3
gYUuAkFoeafoxGlTaqJ1CXfTAwDqC3wIcO376G7iNRw/BnHg43sGvnG5pHPYFvZfl4JW1bIbk8tC
u2UknGTZw2EBV6fepCQ8NMjW86jXVy3QJaRcedB4IuB9wADr4QUO/0LANKQHocCvjyz1Bknw8lFc
NF/cRGvpHrc79YTKzIAhE8aQTqzVSBpmTj4mQuJCzvn/LBfxORWVNmuENhsfmLMCn3xSkCjF2h3I
s7J2T6sWDh2C/9HQGmmu+y2FgtkmCb2jKoyxF9erflptHjmjbD6/4kEjzeqh77pup0aUKGpRDpRj
N2kminy30sGQWd/MoxQZwG3eyUMl0q+aBchB4lKlGou212IOqaA9azSC6Hj6Myr9Pd7SJDBig640
/gx+9FkZ62r6IIkyKMzL0fOUq2K+3cv7C6bgqOMf6LQwXfcrd2UtIeEncVBZeBOLS2gtl2C3lAEc
4H/0GaXTR7hbt70tv/Hv6wHV0HZ0uXtAwcK1b/hVy77FM47SwtN58LrgP/A0/Y64FeBoiTvQnMr1
euvrc3yu32WD+/m6ZyxFG7gNlFbTUy/m9+56ORlUeXq6FYQ9PANl6kYQDwxnmpFptIEf5KbaSsik
Gp7mUR9hvRY/UjLvUC28ImgXpcDSm+wu5yjupXOXhb/S99sXQlH7aIXlThZ095ROA1lmFhVTyc5x
jKpJpB/JNVr8BTiyyY/PcU5eABeHEwJssXyDifIcia6BHncoO9at1x50vQ4wvR4JoNpsdUDrLZbw
3OFc+21xP7U5cGDpzekm2sPCaYrjj1VXNXh+9q5wPo8ocLu+ossaWxcR1wQQzVTIjdnTCiE1hjA/
UcIT6Ttmm+BwKBydmHOsSYuuzbpBaOPphs37KdImJBShPDDH2yK0zMKPrY7nFxx82LC163ImP9GP
ZJw4KsKQEEwMrgauzcDJMNtZ8j/vgTwaUrf2n/xdp09GPPn/3vR5g8BI/k6WYQr0BopBDYg6O9HB
3qN4lhuCOAXxFnq1ydF6pRElgz3YPzG2+K59ppmBqH/utSjS0UYhArR3x85FJSh6qB5i69lqWbsI
b/LfuRubSu2X+9l3eJZQMiRLMKjL6TYDj7L35MIOBlcIUT+4zCGJmVV4GefwvpCFyAJSAmqvgRy1
8WMkg8gGyKA8ltfEoGAAFt9VPLWtXH+vAwtwCjbEi8sTZEFFcZGuQVxj+FM5sWVsEI471bEIs61O
+n1YpedtfQenQSdnKM+vS6jBehpHkR/MfOoCsovgL24UH1dJNfG6y0NJ0x+MYO3YrZqzhL1iWn4I
sIbu8GqprApWkWZZFvwCa027U5KllVskpdgCgUGsR34x1JGgX1y6rfZYPY3uvdy3FPQtMmmjQz1F
p7yXiTMhXmO0ozBOqvTG88+D8Hb+iOGJ6KWekhnSXYFGhE1IbKhlQtGjAgzHl9fkjny2WIaj9cLR
ZmCBKgbxLxV/1Bxice9COvVfozHyKzYI8cuPNkRKEM90/yWSGttqQ9Iom7a9nXMoU7IesvLGWWH5
xdAi4wt8YgqT9sUoPZru+mj2A0WOA7TGwM6Kk+G6nHspuIzBhtS2lDxxEsBzGIT7flYc/NM+/1wk
F7JnPNAbv2Jvgs6R5sdFFsnFpEiAxiWjw3zIp8LO9w5y5XjDSike1mi4ZsIMdVLdr42c9yoyaH3x
DA2Wj2xZbraVHWLnM1bIWnrN7mWotPNCpY6e07+B0qv3nwMGqpYsxXzzASYVv/Nt/lON5L+yNc2X
5qR9FnpcvihFQ+ZdL3B7JG1qDrnlBzZp0jrx+phJoWrSvDigEVyYOhzt9Mx3x8wpJgJ/ZrK2vQvh
sslGCnARZIYspx8rpHTm6J5aQX9AAQ6r33r+Ww3WsmsNkss3goPlSsrXUTsg9hZGgUPZeT2cQXxX
W/ApeArnFg4F08Pa+SaWQTxHFEpYXjsn5VkutZ7h1lM/N8rYU0sCSTdIGBREfRBXc/FG8IL5+4pj
3Gr96KaasEWJjMMCKmKeoI/e9EXkXKCqexlCdZZfDQblnoGhi3z4UBXNxqVOfY+7/Fj21/+M//0s
O4TF7CdU2MTKrlOQFY5tFGwXJ9XiYpq/6EBIqsvNB4pzY/oSGH6UXkNDYo8Dq5GfJB2+XT8ZUeax
3PD/soyJoxHxVRxQAgiOXi/tjb9qavf54birzy00WqF0OtWSZAV4vB03j64UMCHRFmKULMhWyUUs
lc/FgKIZ7o213AUU6mIThQ6jRSH1GXJsssb/PU/L3aPpTYOgf0sGUbQPtTRgXv3qz7xaX47ECWXj
mmG/UaCeVGaxV1kBsLyRfbGNE37ccBLbZwRg/RO7Y/u+JRiWDOhH1PLxyAl9vE26vaS5hidNzmcT
kNKaDrJYySR+IORAOo4T1oq7+k/TNxaKRx5PJBY+UxI/d7kSNT/k6HjAyt9Om0+RTeqKIbZetY1w
sjkRLFy+VJlCwwpSfQOW5DxKglaRzWRPTPnXhOgPvXg8EJl2O6kZd1rRqe/38MIXvv/0jz/7VtFs
0KBsqY1EzbGDBgNBFpByjSH5UdVs+aXQvQOBTBbIYBs+LKH4pE9TDAT6ArGhNg8dHQcl5RdCassP
PMfSADyrS+FFqgBFH6h8qdzVI2BGQG/xKj5jaCZ1yeJVmUkdgo4XHzKcjW0Y/0GwtknVSJ5Niwy+
/FfAuRYv5vEHrmGYkavm83SciwAWJf8dY5X5npwB82om020cVIgJBujT9+N6Y+l+pJMHxUMfmdVW
H+IQ8gQg+g2jNvErD2hpk9n0y5qgxuMMlXCR8ANi+H573w2M9q+tGtq7Ivpn4KPPDIUkkTZ6/KFa
zu4vHoV9sYAxwYRB7ccDMGk+dlNKU43a0RnLKs3PlfCgswpqHWZEORZaFJvZcHrVUw9/lYAYjFoN
j/to0RVwQvMTzb3nwaRZAn2tSjru7LOJ8Ab0HF8nrB7ZwgFgMs5vrxkdqnAVQkioX5jbVwALsIrF
8PKOnuy0N1iXNVx7ZjAiSOKsjKlzVMagAikidqAgicdjOoYY8Y9SjxQJRbbJZLti3hLyxpdEyz0v
lIN+eomldr/CDaU6M6KwgzJGMYIkvThItouCIVr0wxATSVU3RkjSIkUkPnygj9XKAxQMBzrth/0l
5w8fJe00/CFw+wsQGGhpbNZ/0zjYmF++0zSwA/ivaai+rklRlI6cKNmr8e084go2S9+9LMP88C76
/pxMezjAbcfRQR9zQzsX8C0/ufQ/q0eVBzXXdW72/iW78BNoPVXWsGGh5fBs1Fnd62tuAEQ0fVqq
cANUB7IZoDuQ2dzqmfvE7HPmPql8iq1EMuZCOjaokAuTStHLdIijNPCF4TGg0CfZLCN+CWGV7Ae4
/D00eHMyVpeAkWw58coOC8n6442tZ0EREGKLZrijgE2wgVBs7Ly2zzc5omcqVBLUra4AdFi4OHE/
grmj1ojkTj8SpL0/9DLbzAOR9BC1XvBq4o2bAxpX6UB5xmNr0STCKQKCAgAN7oLLIOSBfg8H30Cj
cyVTC69Q6b4gxaMGmldq1go396h9piLALhS9ta+mSglOqS16ncfpY+6262uYILgoDnM1KUPUtDwJ
BW8KTMbDEUzHzN4iMF2V0o4noeMtud0Pv2CvAnBrYbF5G70N7WyKK5J5lrRvnKo3awQeK1Udkowf
fzKGtJi0dT1it5BEvFYo9L11tMILxXn9DaS0kVp17MmhKX700CFQu49taf90/wgMasZ/hX4VJSwQ
bnTXPalJRFeIGs/7yEeOVxq3xT6yPQr5ZyzNe5GAsZmqe7/8/g03E+zqdX9CQQU+syz49PsaHLhy
EGElC2Y0ZybqNsj5r5jZjtazlbuSMPnHg4kaXakBYybpYT7Ril3nNgTDm/QsIPMfheG8ZBQj/f2E
YaY3mBIreUWdHztCwVMsDTy9+NxuI7h6/VVhY40xnS7495nXqIQK2HZ5j2A0s/c9MJNYzcbDX+EG
dQIDggELhXaBGvezVC2Q4AwJDpD+9TIijDoNEJz7P12AHcVBPvrqhb00Yz94FRPbcAKrtY6uWqUW
86G49hrAFv4ncGkYCh8G0EquTgZADxSC76/jfVi9bWa3XXEN7xduxubHb2HdINEHAn1FqFnv+RXj
zA1rlqz3ME6gX2zGzt0jNdZ/BvF84DEg9CsN0SXtHirr7xVQGp7610vgbccphhdTb+TU3kPas54H
U2MPu/5cC4ts1Lii6cQ+6tPOj21ldNvapuQnmIEOELSaAYSYHZVdrY0vf87uKIbE6PBNp1az50OZ
AU1LzYNHxRmVuAuGlmUgPbYR0KrUt8aV2e4dltF4LwGayDbm9PNYbq/88OyuB7ba8c4U0o6YAr2/
cGXPQJ4rK4q0NKuwhahJSZ7sQc5YuE1AO94g/Ezj4GRJ6AD2rOWRajHbatDv4CIIAhbx5s19xCuk
t5FKqUxTsP3hR2EZskLJTcTLjj1EosXWWMwlqKK7KQVks3rD4LtQ3kmY0ONyntgr0hYKVEL6tzbj
p2LZCxpuBHRfJNlsuSXxRMe6SVRmdMOqZUoIIHaz2k7F+XpcNRjXo66YeCRJSU4PRoXP37Xq00Uk
Mx2PGQ1EnhWQHC67Z2XJ4Nd0XiX6zXwkPxuYRTnxGHZdnZvJGUEqFKgJ+OUlvslWu4ae/7szCmdT
fxhCSaVYq9bnGOd88oLwd6tJHvGoFOiEzkIHhPbZD4EVvFmbbtY6uEoIwdYTmQJZwirKsKRs7kiA
vy7qqqSUSlz+810gLN78CML2IZ2gJ7i1YryqQAsXKHgR90Lt0JywTC88osz+91Go3+N6oTRY9ItI
SzqQzOuJGUJOfszXfhkHgdtYnG3J0TcswCMick0mpWG/Y2poUBO398Rgqe9DNXaEcgj7wEO+yu9Q
bc3qAQom/yycqyHkwzA1HbxiwRJ9M54X5tVYIVMRAHlAT2QndfK4J1dchfqW3ULt3Zs4vSC4J2ES
qpfoAAdKkLy5nGLlMFTsUZqPeN2ANvjEk/wLscBmk0FuVavdt1usv/g4PRgqmpzPqfdMRwuAvKkc
gZdepQyx8p1AY7fvhPChqMl3iNn3YjDPfKGvFS/IzuzLfePYkeFrw3dduU2dkcvHAY614hZA/KNe
mAOiptDnzdKGfYdYPIYGGO6eNC2eO4/Sv5s1NNFGUCz8Qc6XshEeRTX3Koe3xruSQt7Z0P8u4JHq
4So4YzD3Vc+G8iXz9vMDrpqhm+R83P1NlJUAFRXxUXuZpH+zktTdFlRHK18tZOZLhUdVMArBxSCn
OImAjiOh2P1wac0tonFMFF44hb//+i0jyRVZWBsJC9KN1RCiF3sIX4iaBT1rzc+GlQH1h3N/z60a
YXYCizxq+BMmPEWT8Kv9vhiSVMa6qYC3XWvoKitRJZDSmCKw5u7EzIApffmubuUSlqTC8nj9swYH
rKUVjthjq4bsK8P73ip4Gch+8NVFN21gpXL/zNFF0m9CXq3ZPSJr3SkO0dUmv+cCXPi0AhB6donM
gtCMRMda8yiwsbkpT/SW09VSx2MjKtVSzLX7YySk6u7hFyYLobmnOaAT5ZXXJS81qk8hYRkEr6Fs
VhzZvzeaJLk+lAloZfQWiChVZz2HtdGCVdQmsNLOLi9XJKQpLjn0zc046NwXRmUCIeUY5Ot+MeFh
Tr9h7maC6rn1EVtYXNz4dz+RDJTPWZH3DONwforaCbWhYro7v7BPT2FLUgRfNWLMo+glEjyYsyFv
yCl50U/c6O1D0UBa37l2fbgnJl7edJI937lyfLTA+cssosO6KlY9AeGORsYUGSky5miLA5ov1gG5
q5DHEIwqUd+FfTplMGcdkuHjczl+MWsVoF1K9n2P2FMSOpLB3DGeRUriS7iPsja/hFzRaVv+6b4M
/bb182gsN4AAcuhC5sr9i4ojZ6uoFUuiRfMKIj09DNTh+otQFGqbugvBzWuwnF22kHy1uFzpWVjR
RKOQPcTGaMwDyzlEgoLldEj74CtMvzsBpxzJsERJZJ61D1PzzOiew6HPcLCz+20J3pMorAkuomXf
Zg2UftN1ecoWxT24H4eQjjSuPAo27cH3MvzYX4rrOMderEU/oSGg24yjx0s2U9KzmgEKOUXYCoeH
HiaqysPDfZ8c7ch6yuBscV7Lot2uCvtdR4JoD3maYeZP2h1nGORQVD+797h5+9WEuePafL+bS9Rx
3WFRzsdt223Ly+tgmWg/tc2iY7VMjx7wvL2TsMRMAuzFLji1rZWtrEd0QpV90q82NE5YofzZWlLd
PMasPATJ9F+y0Kq7wbeWdsqhaW8DBYtCt0tNmDRzZ0RXSPSWId6t3hemZWiZYa8IQAHtcZIhJq5o
kzX/hzQBj+XPQHSeRuSAemGi/U7qWImxnky/aqVhGSD/1z4Z/ribhr3I4cSXGbjTyDQn9//pFSaW
6saLCOr11Ndb5ZLlJKyRXzPHOudGujPxhczbqRRzWs7jrWJLZ5FaKeuWaO7H4Ajmpnvdufa5KfGS
9qZ+84IzXKZrSkEeIKZw9P96ysjUGMoNU2R8M/Jl+rOlp+ubMRWtWXA7OhDoL40m7ms60FgkoaUG
I69mx7FOIm11DHZD/MFocNRsZXzQTxGKuyOJRfic5iSayMvsIdb1K//ZcslkpbEPqCijc6cBKCoA
7pf0s4xnqePlBUTgcGXXYJH4aNXgx3wjV0P2lfdZVmCtRHx59ztYENvyZcxWQIBRbV40WUbFs51l
bz2GTxOlyu7ZhXJ37ZDBv7TgyWOvVYjDY5+VcCChC5XmwDt0sOhgJ/88Sl39hDVmMEXOBJx57TaR
S7V6qQRtBa9Lc96N5w6VAs3n9fHe9MJnCtAxZZuA1yBJU5NrAmDfNWoR0u12pBmBE/csJdPZdcQk
9W1MGy0I38hwtQnIzekSwKCeRYuE5DWycW+DBfVSj2gZD+EvztO8uyGl5sY+KCxOoKdKD9pC4kJA
TEv/incNI3azNLYSct/YSb+68TKVxmN0j30UeRMxWTlVkSEMBkzk0AWu5n1ER9I7jQBzfQpJWDfX
tBm1O9A3IRuMq0TlNKPHExnx0E5xlE70tdmk9xiBCmUNTeU0HIX0hyE5cgM0lrBCgtcQW4Z43yrV
q1TlCz1ZWWxdSEPUGNbiHm0RjMG24AGMrctGgJ+FoLcD4OMdO6FqRwnCZIJO3EAMS8cNq5iTn7O3
j2oMmFivW5FzS7YV2IKqEw37fjU8Hbvz2WlVts0yA+p/jgdeRQuPvVnLjySjvAxZASU+XwuIzPsL
JWnX/EYwYblk7TunMCbyd51DytEosJsJTrSgMGKcrvKmtGhsntirE1OIjMFSgxSrS+4NPrSAgWAB
4VyGdNZ0VMt3Yv3yxZorFPyI0htzGMwk9QoqOajV4K7i7PY/c1JeQB7PPOVb2MGXr2gPPmzUojTC
sn3RICuDmOyHGaN4mwREnsBb6am8/rvvkW4JcYXtLG2jd5d/kX77x6l4Wo6ho1QJRvGNfBTCtkIh
k5PlU0aM68x2IkJj1VP8sjALCIyBpKxaZPQmojCTOVXAOUpHm7SZIh9L8zTnsEaRtMo0M9JoDnNl
hMpr5c5/nEypHyZPsSszrwc6QFkSSu0MxpBYUcI/ZQs6LoY/k2CS4u0SBv1BNQtTIu2JAMtWFGMZ
YApL4LupHtiPvPqAjA83mc2NIk1drKTF3bgHqinM1/m7B0aVeOht8+2+xVPL0Crysi0G3xL8rUIk
9DXhrSoktVOuOAXCoXWJqKWhmh76MojYh3nTHz5l5r+ZtNRJqCTd2zwWp0SFs6l7oFXFDTtYNyf/
OvvansDiycYO6qOtvjloUNp9zPAEB8se/DCIEZt+S3PMGVkwKjvfdOuJtETOcizWcJqJ+58ta8NN
rorOd/jPLUiHEEKMgbD5m8UL9zFlIlByxReQ3obqicuOi3gsUjYJuMUvrx0srVJCm5c6/mkouQra
jaORDddFAnzat+ULRbO271l62ub0B0TwltO7Mj7kkwM2TGDzx3z0xz6GwrN+50Tia72k7L473TD3
ckF1jDPbjbgdvilY8ubtscDe2GPZr/SFZWTsbuVRksKQUlPu50TVkdh/F1Qx+X22r2c6WBRugQVE
G7iSf6voUL+dmoxs8G20tEk93J3VVGGEiKYebwklLQsor3y6Q0FzlkwA4tX6CIdqYNtPCN9co7mf
qvyZN66LgJhmBW/BbdPoKIyfVTh/Zsnkw1iC3G5+Xm9kzxuNE1Tc7OR+1uBNqfNEbgBPt4dqhaXh
uZMNAHSnKiFR3XA2x9nCtobCe3kTVN8uG+O6hFO8UbrvLImqyEzK8V+1J/ajjoyW0Iqygewfc+xH
YWTzYBp6DhOpKsDVwKDtJIPFketY/mHjIUshVDLrwvDx09hd5Mftg0CskFs6ZAjXt47QKkbmyclq
lwAUurbJ+M/Bj6Oq+FPSb6vV+KpEj+FdWTvMXWtOkzMDKvIMYCxj9bXqculcA4/IDuMvuT+YWV2R
UCx0l8hWYVK8dJnL0Qk/1FiMLTSgwKZIiEcfyccBjfTWzj7HbL8CmbtoJbOo2kp/FdQpde4CfShm
N/rg2ykn+1CBbvFNKCJBctCMwDBl3QMbb90Mfz45KgGVQWDsY8NubvXeji0IYXjgpEfEEn93YAai
YIpJawtugWz0m+u4aDftqa8fLA2+3qmNfo8srI7mAiidin2stTq39cngmOwUIHwXZcK2n1KyVM0a
r3QHetsc/hDjJ/CoHl1f2v8tK8iXEmoibkyAE5FwM5xK8cIYqPdk2HPwJKQFq6Xc+NQfqsnhe+D2
2USGm6GMocM6QBYsHiBZ3HHeSljYb5n/a/gHLZlfq3zWm/dQcoxiA6MD46FhLHAO/gJA2oIwpbRw
Lp3kdYB+rFRk7z/qUjGgrEWaF5rHAXcvgl3LJN68SAaAIW+ntllxDyHOb9YPlhmiILDBpzWuJ6LL
jaaRtdrzZJv/7uX2Zj45LTUdjHJlQflc1I3yJL2KupaRzDPWHgUL/HfY9Xesk6Zxk4qMi7jNh8Ni
A27UcI2k6NAOby9cS2e+lbbxsHPsBehn5EE+wNZ9jZDcV6SQVkJB9j5x2bw6WSukZpK0q5yS3FST
ECKaOCkmclACGHPKms8VQHiCPQIX+xm0Oex55+kNpKJnsujACZbClpS07fqqWbh0DE973Qsh1p+O
dAChF0vpb4HU/d78/uoNXM2wKy3niCmdCKm9InEGiDTpg1CbQ3PJvUQOXxgTPckln74DP+8dcCO7
KpdPrDkdUPtWRf/WcMQkSzfmN9qej/Urf8Ulxz3CsqJbQnjhtw1h5TCBZ2s5EwJqcmcUSmlQxD2f
OI5zetmAfb6fsE0jHRrJV+Z/IWxzT+qON8vYsoNGEzptT2i/bDmk3FmuEj04h9P1YUNNBCUevdkX
bFiEc50hYXRvCc/ybZ2cqkD9D2n6py1j2Mj5hbKZwf0cNEtdvZ5IkXdKVRwYoZHi+Ei22IZxTmzs
iG8AqaxL8HnWVoqk0EcflKI6lx44lwGUOO9ZO71CrgeFBgYCqFmXxZ6Byo+HWdvors6Ui7yyqGKP
TgupKaIZD/4ITLp2Iiqc61tcctlHvOV9YJI0wSXwoA/1uy/y98EC9xBLkbiIT//JP76omEqWESt+
KRAz4R7MRuddaNBQXS87+hGvO5uv06Wv8G1rxvOIOtFHUu1IMo8u7hVsKAIIA0rO54fEpXQ9ngYX
c46Tjg7e3noDI9VuTna/ZuN/dWZcntp5ZeqC+CGOoODqcn3LscM57FHGz7FhX28yv01Q1BafN2ta
LZQdxXyr1PF5C06NRJbiqRbBVEYkdoYzZKYLGuCRkLGkL3zZ/F/1mPvGj/6/UWijPmgb4vZs/kAR
pG6uuPKPnBUKEdXmny/oHAtjsLNIq7FVY7x8JRxr8bWA8/vJpkQoYvoHKUY6oqPVsR3gpgklBjqu
SvekRyTpxqJrXqhSY1uRFyuTSn8mdRPxEGhe7EVDFDPmh8Wr842d4OP7xbuQQcVzetDZOMZ61zaG
ep1gWlA+pj6ekHwLPCV2FC9u6PQpEqwtVPMndUfp+dksjO2UvuI+al1ac4lMCofsON9t7ioncbi1
0DityYjHT/EUIL320ZO1Om96CEvHVgBDjVDOeJAUMqUCgUr6b0QD8H+3VmuEN91DJ6uJolMhMpml
OVjsHrE7ksswTc+o1+Hz00pyBVlIyGkncshx9JXSGTlV97/UoTfTOZjrTHzWg9wHQDu02vImsMTq
3uq9gB1KvOmqsrxS7+GAw9BYXLmhoqBBL7H5Jdlr16L1jYztJJI6Iv0q4P7NY9zV/Q0gfJrU9jxp
kNuPbP/ZkPZfWUeXDlIO+m5PCVwlZB6p+zidviFccmtFzgZ3b3thGRMMSIEH8mZc6uVEMBT2ELj+
QNiuasapdjlXpVOOS+1kiolBSXUKcT/hQxrLldkJGhp5+/HRZfFzPE8KNr9kEIFCJmMb9K6JXDUU
X4NO+CELDkPmHSXCbl9USPKv1S/J7Pvcswjd8qbBgzyCfiocXoB8sc1HQ6vRZZ7mLi6UjQZqR8Ic
SaAiMrda1irZvxmz03AaWduRlN0EaTKrPVZGJpax3KXoTUE4wpwsVazG7CFGGxqkMEzvawKWhW1n
VuHsO9X8BRLTH+p//zIRb+CS4bWL3ykeKRmUUdvqmUoUVjmLlQu2jWGJ4K1+kdGHR87vuV3XJA2Z
9tyRNUTJphDHzQOg+X1oeq/HUGEBEOX8xkjfZZuL9FKquYFzlFKy1TVN/pJZym0COOH4eIrSBOQS
UrJp5BTxoOxYXJlqW82okU2V3/ySnye0FrVs/O6V6U3bTg7Q3Rysf8BG2EJf/hocI+KqMuCvf9/S
e6vFZmD3gzpwxLY+oiov14TnXdq5IxUYik6ifx7s/VUIxGND6ROw3UkcubJ1ty9C4R39k/VTEsOR
7P3X5dgIT4hFmggnJoCRD7yUbOcbwLK95ysOgC+Ig44nk7E40ttMb1ouI43jWSlTgluPTXj17irv
2NVkhge5TMS574ADySGIwqqN1rtM33tJjzTXWm39dSQVI6odV60p4r8eM+7jJ0gShq2gxWoboFyb
wP3yXa3nOjQ6lSvC8/Gbr7UO7IxtFqPnE1DQGTwckFOia0zeaRqfYPBeB2nSGD1onH9pgtg3qVX9
SlZLqAMTe0L7uRkwRnN5GFeuM3uI/wbFgoMwdwcbGlAtD3G16BmgfA7xRJVEEOgl973/tIyAxt1a
BnFoph0k8hLq+6memad8ICHlR07oDDuCJFsp95MBNxJREvTyKmHGoN2jYwPQFwzED+nJm0jdQghQ
rUtJZ873WIy0X+SFGDScmeBq9OXI3IHNSy0tQG8G3RFUuvVUZH0CBowUZKIy7Vdl7JP27XjnquUf
kV/4BwOEMB8ODd//C1q9X2H+PZskcpU5UlgVf2VnZYqRwI8Gr36+BEuPsA0+F3RtmTZFLDrel2lj
tMdSef9OtoTqtePGIHt6/uf8icfGuTMdtTnmg+mCLqUbXVFa4g9oQCn5Yd12nGa1rWe3SgaGUDbn
qVXK1NBpUQCbicfAR3zFdQxov3qry+uNBnVw6nOhSSkWwG/mOW3SVUWfhNr342+YMlXBY7xmnfR+
AKv0dNh+NYKyK5jvgRettbeIS7rB9PysditGRaGAv5KfaGak5d0fufVAs/W9Jb0i02yZpkHnlZTk
pUEOKe8iHR0TCFMVvLif2siW0q1ewuDRxcMeUBXWc2c27umv6n8p5X3f8yHafMs4hZ/fj3FPVTr8
wiSW+NppDdJf5yf/VQ8K/V5JBuhBEOyeIjQ0fgjN6Tuvn0g7Cev/vjsz7E2BxxDlJQQ4OjKXxLQ8
Zh6cRXfv0/OFBFSevIUjUAXhBvtFK5bmylPVglNFNZfWladAjUUtsagOcTGds7aQ0co0ZF3cD1ID
AXGruTk9shyVbEmJV2RtTc4DtW2Ik3w843dPHtPetk7N9mXFf+LJJQ1IXV7bae8kstx+NtWxsE3l
oY9raJHShLUr1d5So2JoCL7Xz3uhTbPWhr+GdKbIVxnl1L4C0v/+8487chKm+3fEk9Q+hR+PBQd+
L8yYDQPK2WIgYBeaP1RU8dW+BcykMd/YZpldLNTgoQtPcNKWhlj2x+C1of2+GDM//htuzyMe2jCp
h1OcKL8jHyjusog6IRX/i69pbVCTheelVgF7Fa8nKXAFYY8B/zMKIlSscFjkaafBHd72vtoApsHV
lsVXmXYaV7dqULWepbhEicWWGpoiEfBexODWu8OZwU3xQ6w9KKhvtjEWCdDALNUmDkqDMuBChfcX
aAv1Hve61DOWT2dr0s6qF2qjFBBcmZWoAOhgT6TtZgjzFHmqHLfQ+1FQSYpxA6Qa/DwFaXwDJSpk
d34zYhWRQVD0t14wWR0opiOv5vD7Qet2mMmUReSX8wIj3W5I6TQS76XLO6vj9FWbn06oTDw/7Reb
0R+r0IGC6LZLRzhCTbooFR0OqAp/Pnz9idssOLDTLyncBgG11jWiSVBWBi0/58EL748V10s+8v2q
A9MP/ZXrxiWk+2kWGDrxmb44LYxXtmOusl4yvmvGMeIJM2VyZYpuTZemuo7Lh3rd770cZ+UtgW60
GeUShEWrbHOnz21tIb0RggAp9D3FdjG64a5N6vYR8nNLbo1mn5YX/0l2JCSYUy7EG2P0to5hdkRz
G7RLI6PKX1pXk1ApbQ9EfnzqxjVuluaaKIz8Ljfe8D60CjYpOgx8ZGzjurY6YFILRMuPVTCKkH/b
/cWEBkAEnX7PQBtNbCv9PNDhYr2hY7BoEVKqExHa3B0OukcH3deFYCVfxEFi/GfIAJVX2baOQbV8
ilh1gMgpAEUdLyYaFvOevyU7Mq3N8r8MoRLr8WRIy1kFSVZOem+GaJjqAUtz+kQ8jEss6gvspEeh
184DEwys7FuJb3OFRTAiB5EXv9HM0aTSAFHKXqijZd7g/VGLWid8xWjzrpEqR4LuXPBttmVgyjvO
7HQOhJtCwPXFZLyhkkU2fKfOCnqC/DVWeiPeU7XIy3FxlszEsu4SJIBrFrWgV5PN51lNMAeYXGzC
uOmStTjdnPPdJBGk/9Wfal6ohh57SGGg0XU/KMdQcM+sW4RAASaDKv3L2zyYPV79N7kiO3W/+wJZ
zka+rC12+gaCoeYtk6vU5tQD8JftIigJkkPHgPS5DgPQlMn7n6w/YidRS0Eq81WpIYJeZt7IDR/u
riaQjIhxjmCim5J0amhDs0vUpU4VU/WLB5Sdm7ur85hPFqfnM9SiSHBJ6Cjbo43cRWv3MqNYEnZ9
msSriFWYi35NUKSWRYRemwQcRg09QAZOjqiMi1TMXytrzo+RtjsHo5L+/3CayiJyqbVWPQi3ucVH
G1c7Za3m12TxjjRS4ywepuj+7dvh8RzvlD3RA+xtUyslI6K8lc5/uhQWFh8XLPrFaP41CLAyB7hG
cor3fp3qSlT7Dx87u2FNEttwRTKNe9FyyS/bVMhyu+zA9HjTtUUgiCwJYKNpKVX4bFebErKyVL4f
Pq8Ln9YPyIW720Sju7fVbF2s6AX02ni3xZnI/ugMNd8PLX9wUHpCYNW5Sha/bBuvlS6PKz7TNLCN
IoCkLfW5RdySQqniaCOEYkqZY1kJ50jX2Co/u5CSGSTuiwwi29697LhJ0sroa5DDqJ2u/ZK1/1ga
TuMPUtJo2rcOoMSDNQzYEjaUDo4Dr7VT476b+5FyE58q/vVv3bOnckAO/NP8J+BWFv0E0ZoXrBQj
AJ8Rw+HxCBOVDQiAdDOmjfVZeg7s+oBiIy4DtuZJIvmnJiM8Rf4mAT/SMlqXCsHhRkjIYWWUCjUN
qatMZN0lwU1CtZNTrx4GlML1bgRq/d4yJy6imKR5VVY1nawKVnCcdAXIrEC0pFgW4tJ235i6JYPC
aRsrxJRUu8BUf+hPUETdwFUnVJVn8rP25L111D0dTNBrDVfxsjj7PCP2aniTDt1q1bloCZQpCZHj
INB/YJ5i+rzrN/qX2N6NwRnptpR6KyQFAk8wPB4Vu154CPD9Sn2LWIFYkMeur1xiC8flKYtcRrBc
oBrvkX0zShxom+McP/KvnKS3p2n9rAuRC/WLq8m2BnwsVyJxbVKLn1YNgQQktiP8XXtMT3aw+27g
la6Yt0a8pz+/8Yrr8jxIXPUtdvhjuxLgVUjwoUnVCPPyt1kSygvMDNydWeBz9LkYv2v3yS6UD9sG
rMoZzA+51eZy5iZAWzTAW+/OEDxjWEcmzqOj235hE1L8/pOeBbImCKuIN5AbDzziKHRdrUgcWhE9
cwdC9m9uvDMrCa4iiR8XIPJYNfrWtuy4S2OlRzLSNvYS/ubcsCs+L0rb4LrgUBLMiyH/xHhuCW/R
PmzADn6Uaa7diS5o1ZZBivOrZP8MYWmaO3/n65LrH6JPNRtnhVpU5IAWMJOSpt9seWXFbXsJonZJ
udHJ3x66gM9OV17Wles306MQAODb/KP5BNwMymVvXPskjUGPr4kPFGwjq7wO1XhEc9YKMCqV/Kja
gInLwpAiILm5b+3GRag1ZuhkyX/rvvpzSDAnLXN8nN1UvKD7EoUgmoonZOICmeFRvNmdopZD6a/4
2+jDxu0TDhjIL6+Jw2BSLCL6bU6NxO7J8v4ncIDlWl+zYkNFMMW+2JUWnldSahyjr/ljFcOddfJi
eMj+nkSycBRQlW8kTr8ZMUAhzwUkKmUHkN5t2v0zalSVUZ10M+E6AfiItf/M/LB6xbf0Hn4pCSTp
xkxTFiQKvYAjHQiLhfRVsCpTr27j6y1NbYqO+/WtP57Fphm+uUVo+dnMMhycuqBi0vgo7++++uCQ
IegtaYjUmH0N3CSleVk39X2bNGrZVaBNx6SmhoTlfuTJVCfDkaPTcP/FaNg5ur8wrkUZjv8GvJ7M
CmLoGO2F+hkarV1xz6W2LzY9VhG05USx6o3/IlyatcSUdjFG4zYK5X5GKwMRhycmTFqDcqvGBU54
vwxkZPfTYiXRU+1CocYW4CJEIZ5KEUoD+AjxNXsY/FU1zkqlHFjGD6aGeCBQGTog35upk5ffEpp3
6sDW7zwT3XTeLx0IIy3y0H3tpzjoG1GcudCZvDWyvZWpEmY3PxA0Mo0VPKO/wa9o0YbrNl+1nsk9
j0qtimR9fkaoPgJf6FXT3kiXWO0lSHoMuqutQwT2YW8rvYLcL0xPONbIDwAJlmrzo12SoDc2ZycX
xVpaGMEHPBI1QJRjAR3oSDq+B9GRc17fxb7hRp23/SYG7QvlG+rlNkijYrK28+GcetP+rhoKox6y
1l5KNn1+62hArOvSnbqF8t2QxbMroVJAO0/IlqqdUfco5insdDT7ho14OU2Gz+d1ArbtcE2QpMWz
EH4tujj1vXsggOE4JbhmubEktxhrIJQK50BlekGTRFRL28FD/EDIR3fyN4npCPDci1UcBxVmGche
Cjar+7tskFZ/0PhHHlg9DcqFBmwNaNgrz1ILG8i8fZSgfo/eh8WDfFlRPh81NIIjrSI8Tqkcmcar
HdbiQ6JxPdrSLrRXclStn7gJBxk3UFjIJAAXfN29Equ6QPG+YJvDBfhvXEXteUCaVjXLyQ5EgZMK
s6jdW0OiOadEEHT4wOHCFKOT6A3GeqOPyWa0Vg5bp0Q2qYd5lCzXPBGc5wfDjHl8GbwJr91TVPP1
tPocBqTPLLE+m0gZ+mxFufYhPQYOf3CbhB3hTM5Ws5x6xf6XZi455hZ2OMdJsPJk/WW20YuezcCN
cPAKHtQ9yus3v7SKnl/2R3GFW7xwMs2YRY2pp9mbYz9gxPOCr31RJHB84X8mCwpx11ulzm9RvkJs
9jzCEfcAlnT7X9WtqzPF2hiKZwcO95ULryJks0N9hbWY01yPSg+Zi+zZntEIcKll/wX+52gqVZXp
4e6JbfD4zwv61g4SQF1beR9SS6oSiT11iaSBLJdIVQcySISRAD8JhvDqSKFkK+WaNrIMBEnj9t2S
vFMp6Dj2S8I262dKICDuu6qj4F81ar6Lzm3BMNTJsv4c/NakHr3jI/Yw11UVR2iWGlO/TlVD+j6S
FagBjqEFdjKXv/3XiHa44IF6wZgnj8q78kvG/Vj62qSudq+6zaXtg/bhqA6XfuZV+grc1PVlVKvZ
kA3/H6GPHlodqfw9JQGiynFFi6SX/vBVbj2FyMaU5zgcLqzxMUlxpmvToh4QfnW9/oDp6Q3nXXhL
tIFyDqGxc+VEIgrY+YYNMvycfZAGtz2lDFuqKY7VofsVJG1PNuIJpWHR/qsG6Nf271eRigQ0CuPt
Xi7YlMMPZ5Zim/hXttPqB1irv9iBOOQCVkfu7uRbOtUmV2H9lhpeTWzmNjoR/vb0+MDCiOj30nob
hyHXrx2vVmhE9AjKFq7kOOpW9V+ly28nT5goRBoKqQ1NHZ+sz86ZA38CqrcOIwOYfES3GdcLM8dZ
/IcxaHPIDzVIVbkHAulD8jI6orkuFzGKW6Xy5fxKlQc2rtPESPAcMIbtd8KoE96xw4DXmqxxA91S
YDNmVsQtf2DxHE6angEvkyetOgDwwG65wOsFtuE6/8MHTo6zp7ZjnqHW1MSghbpe81au7bmZXgBf
feYWf0AFYSoMx6M/qsYvsDG5wf5ebbgrS8K4MuoZ75NkQ5VzjLXfYlvLOfLP9IjNwyqJw/P5T6SA
D8Ifgw0Wzi6E+iRfxDZBF56YMg7azzZndGOMio/olDub2T1OGd3dpYXA1ATJxt016g552rafJYVu
YGRTnK1uA1HF57UdONestJ0WcjuHW5A+WeYUydsZG2PPhpsuUK5VORLZXG/BIGO2qHTDE49vd0CD
h3HEKzQAiI0kCuwkutyPAMGetDz3UWKtAQQd0dUOD5fQRHnFV6/3u18ZFP7yChrPiyeGiRXbfKKo
/eOQ6u3to/a6lbCcpM2oWYEJDlRe718QxrpuWFomYk4j+Tf0cA3Hp0CyAM26ArAcBuWBQhkqn9LC
ohejgTFdMSs8+BXJcWtWRBAvue27Qitx/UYn7ln/jYHUAnmJS/AHyqBOoWd19TjvEmKbqQQULWVh
zdcFZPrHAtzpbS3/O70mV5fH9XRS6M88KT//uAd8/y1IzuaoqWLLXWfriqWUzSXRBlCbKLNhzL8Y
j8zH6vRpGy015FajYD4AQLvXGqrtY3RnkScalnK6LBcjKZySzLkfuUPPf6JfBXvc2wypcIpU3JRV
7Mp/0y2lBUmodqul30ddsPZzLeTOplOM0jQGCXH/a4aqx97B6/f3Wi1SRC2dnW4NgRB+hm+eJc3i
D5wdIfa8j3+XLXl7p9pYWQxBUdqZazQ9idwEHELpET99MuhWCl14BToNqTzKlimO9CuM/ZH2EIAz
VIwuGdaawulTsLLNXoPVLjB3UTSArVcIhrxRC/WwmBRsZboJ3Txvm55Ea7uEfDREIT0Ia3oRMV1z
+/zM8JXvdYeTwS83Twn97OeWRAljxjrIu6QM79nldcQVxIRb6Re0B3u3Mk57Af7QqVdvGzR+vD/U
qvSJEoBcgcAajkalgecbHzImXliVA4TSRqgE5Al3wQK1Lib7luyI2nGm0cKZ6Pi9pFBgIllcnPAI
VCFEwlkV3nkB/WgVVjiSlSZDXXDI83uzKH+cxgY3iJ7iDA1a4qsK+tlTi8gCF3QXaKu18Vlf/2BZ
OMMX1DqmbKVfLtA6yakgQTcI1JIa58LRPTVKQjajxfhL9iBFCbONhPpjCpiPOoYGSjyexMMW0FUi
H2iK9NcoW3uH5SXeXdVtoJnpsw+n4KK5uwezWCyCTXnaNPHsCdcE3o4ve3ik69ecIpUyuQFIl/Rf
OyfCFL0ZsuQnb+3vwyRNxi9Lx6oWFyzkPk363UNvDcc92uuO2QJVoOFEmsFgO9myOR/K9hrK2wTq
rxdhfBDavUjd3pS8cx5UEHF+oWv6GQEeKkTjtxhOgEytNqQBVzqyf3DyAQdBsNYfCC3fJt/MqI3Z
mY1VNLCynvrj9z1YX6lfFi2o8XCJEsZgj3ZLzXAZmeCTQ0LkNJYtwL2VTeMuw+su8V5Aulw+xukr
y1ZuVcCFQZDyn5n1HvLkFKH56TiGlIDP0D2Y2TFKfcCDmF60ZETJxG4FOlYCAAtzgo0c8T1wCHEl
+9APurpsTpUpeOg7k8z/n0EkmKewzN8VnDJxcdWiHltlyNgX3WlWGhydOpwtnntv2buIUfQg/jtr
uVdhqeAggNyYbkYgQ0HKUW201JiFQF6HfTTmFc4fyyo1Awq0fUxwkLuQYdhmYvpqxAQX2MJPb3oa
fu8+f37C4Cyo3RndyYHsU7TTeKbaWS0uMOC3uCIFZOtsubQv9E9orCZUBaPHUT8R2feIwV6kB1mE
Na0QiV6o5wmvfHkATUduK4Sa6Vx658lkZgxAWtHz4Zo5Ygwu4olTALb/EwLiRWy0ztnGtaZ0cQEm
qijcywakPbFgwkXchZjsByrMNHO6cTUiFHklX5hvFq+A+Lx72iJxoAd9EpYpU2FDHdR6FH7i642H
kAzsM1XJHNilMQqgYGRsHOeprS2dfwzhLNQ4NfqCB5P4xBDCUIWNXO0Bdf930qg5ETRDDs4iQr2y
VUdvlVfdQo5Xf3BOZsmcy0lGIoZsb9gUnCc4NcFpA2sn86tDNdqqaGOoaN3jvyP1gojPaDFnbJnp
wqEO7NLXgBMzpxL/j17G8R9QxXRgYBVrraCxMRMhwy65OGggPmLinhKylvfEPzi+a+p/f+cYeiim
8XW0rDdifYfY7yPSp5uC+ZnSYZSZCClthg98Hh2VINjyrYqBL3rIkQeE1SMEC+i7aPmr/u5QjkjA
zxSw8l7rmnL5UYoe/OoSOIx/VaM9Ic79cNAOUP5cr28CGf1r0UCykwNjPuw92pagWovWp5i1GhPM
SwC3ENyz4bOfXmS0Pc6zYuzQuvYgqPgJWceE0vuNf2OGzN23ze3QEGgkC3eOc40r/02e5N6XlXZo
NyM/HxfEwG2w95NjInxHTxb3wbm71UQvbdS+hjFqC41trj2eQZujZve0gJbYz37Yjk4jCSz0QQGv
cTgspdmRLnHvVpR/PBVVw3UpYuXXI8Mi6T3s83TVTjLF3Re37OJ0h6379Jfs1ZKR79iCrShT0AdK
Z6LSWuw2K5yEhTqlk3q6b3bOeZEbAcTQdTWXlQL90vScs5iWmBR+6ZfF1BZ4YWnDJSbrd5WLgGpX
dlqmGjPL2Vxb0s59CogM6eUKUAIjVOfwmAf9+ekpxz/e94i1jOwCBl9SUm3pk6KPg2e5BupQpRXd
ws9vUS28s6HyuLabgX/+RUleWNJ9hVxOryrtLLPQ9GqLuCy6OFxuQAHPpG5DUpApAGLppLrXHmNB
hpKwV27ZpKVucfAIzHdfyzPZt7q2GxoPPgWCaJ5JEwPHdsOH/jG4kc1/nUSaOPtBIA2TMiQfomJg
D4Sf/rjRrz5Tz/5iHUblt4opMaYHNabLALlZNmMfG13082cD9OUFFPgBGkezeMwc8qdPl/lGV8bx
yN6S6XEb5aJq1L0ZB/tFid/ITX/kmIu9tCpsdJeAATefspsLgSQ9OJAUqN/8O7w7godgG9rGun10
oSmHhvsL28Ply5311vQ69TK2T0NUw1aB1vOiWNQBLZ0WMMTyovhyfen2DjGuQoGkGAOpvTj4SnYQ
2iT2UVVze21VLmC9kBNw/EzqTsafQs+9GTSDkisQaedcz4OpA3ux63n9gg+DUnV6vAKCGng3PGJR
fbDT26yh4DspiEjUrJ6SQM7J01EsV5pS45dxhaCGek67crBe9+DgLUfIqAWyTZnFIkDYID/IczfG
DxsQ9XMrJqChQ4CmRslOLuvKl/tXDf04hb0Dv0QZfoQUgN8+2/L+OWRnUO5oKclwge0f0+zXiYOp
LPzo7PpKL2z8JLSZ6qSzNWpIEUkN0XKEGtX5OEU2p/u8kRHeJDkxk9HtWTGyqE/j2Ub8VOfclUCn
u5/P+DQ3GoyWXzqDG9//Wr5ptpZfvQ2VPXHB7Rfp6U42ajUvRLzt1opA/7zSirGXlaMGfesLcVLA
mQaVGJFHfBbJm4np3GJuThdXOaNkW8qEyOqXgmlVXIaLgnBOZ5AmfRSgpRa+GV8pSyN9KQn5ypjP
uIfsD57xiwnHShPX5uf682LGpXDs+uYpS3lhdtlrzlTf6uPBjlyGrx6Va171z5x9CtQ4+dBwTaIv
63f/1gFMMBOEVC+iT/+UnnvNHqXrelM9TPkIwbkfNTg1K9Xgfj5hzOuPxVN/NC2umvHz2Y8E+Fm4
spXMQUA3kIfe1FFXxC0XVW8gghy73F3RTACasSiXTd8E/NnSFgpZm+pmFOOpB3Dd84a4BN6NxF4Q
miDWTabSXzKLZNfEW/oFNuPua5M8i1JDeDubFQWNsdiPE3l++IH1biDUuf6m1KLYIxXdjFuoslGN
0FQJdyVNC+jCs1nmUX2Uii0qs8AIlzkRF20D1rBG8N2IWCz3f0KpPnLwEB2lbmOGX1veRptZvrlR
X0kk9ONcXUqbqQTr3QsUwUkMu8/H6MBHPdRO1nC+d2iqblsrH1E3aCctSiyfnvPtiF50566WazTu
dL912+5sJehEbKkYHhLzL6Y0Iq5Yep1MvFrAmr3rkSZh7Mj3oFRibAeUvoQefS/88dVL2i9ij/m2
pjb6DdUjqn6fwIyjU20IaU0IzwGQ+IHoFF/nRCsbYYpEhSzfSZSbqCKywC0XyRlFRN4Z2NUqH5vM
W5FouTdNguVw5bWTstLY4u/IcTuqnvSZQcGlH9ITDgWiyhjt43MV5LWHcUTNGZwQY+I8WLiiloAf
nF/hD/TOVUrFUPoP9zQlMhY6ykKKjgfxTxtaBv1wTyNeJHUm6N/H4/wZtyex4dxRLfGIQWt4lUtN
f5bDWM4mLqpyq0Jkk1KQxe7laHKi5pwC0QsgSqEK+gw4U77kKQ7ghNVlQJFBGba5QFavOW/P+AsG
rpxjc29iUF7/p7n3mDcryOmyOM5kR27CUtyekWIw/9VyKeVBbJPhnBj6BYUp649Z5aQ5rbDXc5MI
U3n+tc4kxcAZqQagGkDOJMXtsF0Efjc7i267ONEVlFqy8WNMWNeZEPkh1+FVXBCxoxI1WHDFNiO0
Bed1sza5KbQWY3ANMNb67PanK/4S00EhSy7V3pSaAUyGZuP7SSi4MC+mdAB3VvrdEwY7RxliuXw6
rpbFEo4j33Zlbk/farBYkwdung8fQW32+BNYqb8kDiRPbuOrP4Oy4vBH29O8NCEe947QshAD6146
QShTHkBQ6DYqOGLH3eT4x8COZVYq8ycr1RZSY1GvyQbi7cWuHO0TjtEtzk2sq1UIViZ0y9lkLKmK
RW+6EdDi6Z1abKf3qkVuDKfnLYR4Uy1O6HLt4jxnKGTZ7IkPQknLlE3KNs0xUFtmGFMhCYoo7WSO
bzItjTSeHukEHLqvnu7j2dx7IZX8FW68s2+9IdbBdalp4m7Dy5Uyqg7teRVCZwCgszKcen1+MJnj
srdXIyx5mUZZFCoF1mbkyT9vdF86G3wvd8OVQA/w/mG4LTm//dU7dGqAu4L3eev6kbLuS3OUi4cz
WyA/8Kdll7zK1qDKlAEXOgXU1+8rgpvo8WJ+lc1s8olXW02OQp+PMHds23uvEMBv/mKdgDARFPp0
ylKTkzPJiWZd3Dmz2kziqM97R2e1DnBFbktIGGm4tYvSeazrCcoL6U1FnPFLicq9xEIma+drfZsD
Py6djDz5mRdCJ7c196N/uavZnQhypkilgABEy2B1FLWDjuuBb7Q/BxUKdfRRlORfpKbrU1RWL74b
TpLEEeCsb4mylS6kEquZnOmtLuHQYI4Q0nEHY8hbxwB1d1Grp702HAB5acH4/LNIApjDC+KxlSxv
Nx1sz9LqAF1HW1wt6cVOpXa1I3F1xTV1Zlm+J+g/ZD1wO1oTGKnUZuQcjMooFJVK6Rot248iFCQD
thqj1Oq17Jx1fwxRSxpVtYOh9Ya15Sczc2CQ+F8/WnwuxO1Fd1Wzw7oQ7Fml7ML43a5EBo7BazLC
/QQJAP7igwgbrfluy2EdnGyoPVBmWu5jiUeyQDZF37wY+Fntq2UekNzufgP3YHXqXDZSG9tTukR/
96dzKS0sw62FSp5FkkYDBixH7kcJ6yTnaxGueSxtBQJCSwHwMLyymYYN2RRA7SQ6CKiyflH3DVGl
A+b7rpmsjoN4djLUXXHBBPRLgSU0qIfyNEKENIprnSANi/n7r68FDq85lkBKO/NNowg+tHNkCYVo
IgMzqFqnzSqE09tLInCtKeLl1vyiaghbiL/BupKDl1WMpVJyqyFURvvEFM8Ayit4oQdJ/0N8wFeB
Noh5ZZD+aPacGITAZ4sgly/kf+vlbY/Fwx7vKUpaHaA/ReJpgalvS3e6xAPnzXFfAE7xecf1XvhJ
qDFeqmBaQZb0dnpHkfZ9P/7g0Sz/dQhXFLPe8o0+A99AseduYhZuERNDotbSWVqCLLF91VQYtLR9
MKSfzuCActSkSGxMSpWdjbnQOzxx5xbp6Xmloz8Samfbv5J+rcpZ+Kz+VkgsXiuGxJHk9yGGIame
YTgNv6o9ZT6jX2PeGqF+KPQD0CYPjO1wGh3ReLPW075/zuz6OqWm7kMoLipDi04JGDR/z5YeQqqY
SQ7OpGn1B39dRF2kNMAWe+3f3pCyG4NPX/xT2ePiEstJxqux0geuQufOmHJ0dtbj1rbKl7au+74X
RMq6kDtPADyfenHFdo4i2B3iIXXp05lZKA0pK6i0cV7OuSHpLCKLS51El28Cr6JDAUKg1G8YbIhs
TavrkgW94Ji3Goxh8ZwySFBRBa1fFndoValIcsUuC1GVf7pwq5HzFK6RfcJRBtKAKn/lEqxV8wW+
zd8chld268PvzPM/41beCj/f2W/dlLeZWULCs+9rmoqYKbGpiKTltJ17O5G2WOlGx7d34eqLB56K
sP/RpalD0qfC3Lv7x8qwkRN8VHfm8ByEVuhYmwsxSngI7qH8fm2TvFK0lYDw51p0x6M61xII2o+w
FTsfAOJTL255NQLmjRh9j9g00IJjImGMdXrZU8DIqtSJlvMl5OPbAbdlUnf/2C1iiPjhYjk3tKT9
oGTMGQsjXbwE/Z8sY5stg9gw0gGgY8BH/aNNOSxeEhv7sqyJH/fVw3tKSe9tXNtVfPA/NyMa17f+
FdIrDNdwZ9YQbZ2v0tTGPfrhvfu62TCmvp12DW8M1HMS94CEh3lDkggg09vZ5Esdi+Q6OmQd4JHN
zgoPJJQamn6k7HVm/CL0kSFFAnF3sE4FL7CWssI5ibe8KV7wO0G/ZW45CANO9j9+Ksq05BCJJMOk
UDcPeW6JZIaf2/0B+gY2GUxjL3e82H8lz+zmbOv2fpFZ++RgmzviLdLvX4/YYrxpUkY9A7hWsJX4
HrolLF85beolmP6K01zydbCVYStmx1Skt81kpsoobOy+MZpTOJZQzBcOfizpaK6OzgSJGixgO1XD
TAuhyBILa+K/dRgL4fwkAiB4/vJNrcLNZBQFRgUzBNX0nPHQkptK5bBmwuCc1elX1IrqTbjnGa3c
/tOTc+4F2NsUYRxnIZEBHF2/cijViDOSDPwoU2OJipmi0JuDkJ15SMBo3Exm4tkUFGK7eDkYcvVZ
07yx86R8ony5XyzpvqIahCPeJzjOQzSruhpZQTcx/bsIb6aAJ23klblxAswNT3bKQIMT5nLEUiPl
s4gqls4yxIp7OrqKCbLqScOxW2Yic4bINsTr3K167KZOtykoE8iAXL/WQVry9V2qAGjiph8icdV7
xlh8xSR1boOUBNWA/cm6+CAFNW73xyYbQzhcecXZ3AiZvWIJJ460QBBIhnZtUu/KLGgEoFykfrgt
InUjL21vn55sRphleGSioh6qgIYoY+Yim/34M7BmkjdeDq0DZloCkyA0A8muIE6WZjHrQdhMSaYE
ExRIrro5gIvESEN4zroGZgMuKVme4ZTGBn1z9NprLhgZf/TFo+p2Mj1bWz6yEA8ZIIgAQS/r9nRo
YoaAMRCCRBz9z8CVp37zIrSccM9D0npBPKhr9KmGs7aOIih3CFJlItpUDs4Ibk/MHSleHMYh45dV
xZ5FOsH94UaLV3U6Xly8id0EBniHQG9FOomNdu0izlphFJHUs295UNk8YFAc7nNtwloE6GopTv40
CK+DyEni++IwL1qJnjZRSUTBm9cOJVHcJbGt4Clnirxm8vVhT/udUSM8uWL7R+YM0Asq5LVhzl6/
1UzdF43f6hcPDL+Z2NA+KVQD0Z+7xMJlZZzQ+aFunQPz+JRj2IB7oZa5t0qJoKNxH7EjinFUwZRL
wZCgILXzErV8S4yESMGGIcHzL82jtNdhH/RsP7aJHZeJzxuL77XIrncU6j7+1HaRgt7SQWRPuy56
IDd+gOgEDgAZ0TzBtuSUEwv01pLZTDwAjw+qt9z2yXHq6dtfOsaoUgHrTSjgrKGUGPVD5v1n05xY
fiN8TS3w6KBzrmUueiYbecdKikhy+KZi31UBzBko5TdBSLc0RQIStO7C/PuOZ2ebLmjemQNUOfwE
LC6eWxw4lBOyWpFFTCZF+8PY1fwcqvPg/IY5Lyq180Rb5n6qHkDbPrx53EgyLaGJ5AEw2PdIyk8M
ZxcHN/2lV4dUTJ5oMbhmVgVlHHDXWuqcK+eWUD798zyCYCmokh6kvsjfhpBS6uu6mvjtLneEwOvu
IIvqZAaO0UKWdTllfcwen0XGymeRAc05JD4wPy4a7WYbcsHvotDXIDsjBEbeJ42JCsXGUA0IBIyc
UdV7EM07WkrHzjfZl8G1BgNvj4A96tjPKwwy6RbPoTVcoKI8l2yLQz4pM3QC333EH5Jm3k4nO4Ho
1cgVK+mEtgDxN9ekfUw/lKo5N/cPTIP5wiZTRGEB2KWAwxwlM/lBA+yGAnBe4gZJ5RaVxCWcepf5
tj55IjWB4BNvjXZWVDL4tB3g8BbqoxyKIKm01Ue2GlgEuL4vcZIGZFkk+aBUKrlp0GwwU/c+MlaN
Mu8u3qaPhWk3x0LSqL2cv02YBYehhIZG91HJpYEWFfu1mY7ZD9rmt7vprRa//qs1yHRIZ2d5z+Lf
Co5rwnTFiPFa14sWpAJPlKxK8h1KHEr8I/VOWwE857nQEswfEqX0XctmRc01PgZtW108i8bRsUxX
scG4HEevy8Pk5NL0ey12XigqmkdVmBEHaO+zZ9Yg9/KsPSpvG0L8hpXPg2s8eBm34sLgTf+hnccM
nC2zPG7HA3x6rCRiRYVQaa9zwcCEXtYjSpONyTUxupDVpN/hVvgg2BnKKu4ts78JQpuPsEw0Nhye
WfQimzUv2vR+mh2MH/g1EzqwE4DLl04e49upUNbxpe9GZ9FhiZAWehWcBup6FlO9flLyv82p3Uvj
Hme8Axb/uvF1ZEch6mtPiEmaySovoODROtBcoP80cod9WS2A64Gr+fIv7rryDyjpsWb6fnBhhEpx
ssFRrOeeFsF4zfK/QQNpK+pOdfvylRnueryscgAnOuj4chKs3+BSN8fY5S4CPQXDxhMOgLlXFgeo
b4q3diIykLZjcmRplmYDUMroBzrqYLBqR28tON5tY9ZaF2tPEmo0AA74wEeZRRgimJ0bsmP/+ziT
3q6wypU/moSgKr+mO3CjEsCx7FYA5K4CEouJyfo//G7jgsqvIOkeFGdSyhrJ8E1iazJ92klJBups
iI27FH+qsRs4nNxUWIQIsFf42XH5KJItPuuACiBU+yoiG2gp1rUJlLW8b7IdbO4QOnmnb08rcJGX
i5KOarqp4mlP29Ka5dogrCQATzrDR071tsghO4dtXG4Mj7VvhoHYNcG5ymhG8ODMsruKQMObBcx0
LcnNKNYBQEnqY7oG++togs+S7y4dAnnK4WK4pp45Fxg9yfb/U/4W8+LYViTHlQ7kuoT6pl3TX5Ui
Bd9qOBHTIpveYbo36N0Q25UpLKTzVSkC2NJEgb+8uvOIUdUPDM9mBOQPaV2CPLug5znEjUl+6zca
5G67ivzayuouy6Sy4/O/HhaXu7GXruvWT/vcohpFaCHF0WzOUkpA8zBFW15AdiP5ptnQGU0vTOeP
eaZcNWdt09v31M1kuNm/oXBhYiah23or/LLu+f5ItHbctUZx5WXE5o9mqqJDEznHTixkcOs8mVzC
1kfIyZwOecoHYZnzjd+mafzh4zRdQpLOEQVc8qM9hl1SC4lDo0egYJ7Hmc4x8EyRAFoGQCuQ8gNW
PBYU+xUdu9nx6Crh7QwQOISPPhqMWAkLXRYOPgVtkWbHQmY5p/X8F4wePYoVOoSq46Orx3Hy1sb7
YDQgZ5V5Sut261TjDQd4lWPe7xVYVfmgSxb4UBmtEdrMvH8q5uvzWZ4eDxy7wag8nkoY4sYabTtQ
pyaZkXa4ChLM3vpiKu2WNvVxZmSSCsQNb8Y5dSbCYvduEqGffzn6u/w39a5iaykjmQhSTTL+AvUA
jdIp++2Sh0GdBV7Eg7e2CdbVONkZektEgkWMU8q5W4vhzvAckV/NeXci0XRggrTDbOkH5Emnx+vu
UUjyw6tqPj1YrWaKuO3NGZnzPIrujufQ9ui4xpJjmSBZE9JRKhxcKCrq2jpSsvmy/pPQ1FjlWg5Z
hDXrtNoXWIvTL7eQ2dlOoVp5P+dCLs+2WfzqvfCvV9Z7VWx7DiamuCeorcWvuFDA0jYYqIOM6Crx
+ASNOyzClHGt6+kuidQYFwGnojRP6a3i50claiXk2FkvPitJcQX3h2h1nrWgVUSgvbD9MhJnd3nA
o+JyeE0qsKlq+jyBhNXgMSC+WnHDV4gT26PxpGyeJ1+d/1/TdfmJRiqtAe9MkZy9sw0c60tJrBeQ
/DOcAPlwF3H2Y1UNoIvWsN9NVhHt1nhWqRf/ItYUFByVOhlA/L/xlltBlJwOM+l4PO73xdUgcbUm
pTyMark89USQVtLlBpmwOo1g8pUZD+nV80tiHzdcgp4iQR9CuwY3+ZfM1eB4V15oQWB8VVyPfDbb
Ad6iKuOHg/hJ8x+39LJDDwPf1hLfx3But6XYJ20GkilLRCXNoaADPWSZq/aSGymZ9/F1uWEDk9Le
9/3Mk6o5Ro8rmHzbRtj3jIIdTbLKMjo5wyxajN3V91htx1WY+FFB/Y6xPJuYX9qzKksLlG8ChD0D
/9SFbL+2mlPNaXsCwezR6INxlQ0SErCSnrXlCK7eTvIyaRIrHSpWxzSa59ZarIwsxezXLiQb6nZr
QSHxgpvsMpihwOuBaI+hPWRkdWQ2VMDBNa207L265e69huRzMUMt+4r1vnquDG11v1eEkNEjxPk0
D9tiSB2K84gxAAboiFtpYHsL2XVNSHBygOuWmUvPfGQhM9OaJJKE1VrCV+qlKB2X8hno/jA/Xoom
50nvlSc6YRvGhzvmpOlUpoPINkaFcxwMnpVQjbTObyQLM9SmbtRdJz+uLH+QV1BYz5Kxz+Z4Y3/X
PdOCoaagctKNgqxUE4giKtCZsa7r42yTDut26aOs9NwdLRGLbWBDyVQwlhBizOuYGAEeNal3XyTq
nA2lUfQY7k4lpgUR3rOwM3+Zy6kgSd5HWzGSc40oOMOEfKWzVifJiVP+8yvH4AXzzGYek5eKRRGZ
ebO1OMsNXryYpRrSyKtCRUKzXyrfGQ8SihZzfkGPCvg5XA4W89iHf+VFKwAvvcUR/YOf0wREezqr
LwVE9Eo/B1FeHxjn9IPj4FGJMI1/2U2lzrfyZgbc0D/FgF302eNIb79VqxAkGT3mf8B8cHBoy9g7
vx5RNnyewa2uOfGhro2tdGZSjB7poEs2CdOzIEu/gq45wT9wCOkZliUepSdJgVfiZzAs698LNKfz
ZJphfuP3oJ2O297SRTZhcESHvMVcQm7Qb+rCZHF/doypzrd1q9BTzgjKR9va873iAAeJ6fYkII69
oQ/02Tlfgkrr1u5eEBYsKnMQLuHW8JFtshmUwtlaX0yVhBAWa+znJ0M6WsqSIgYJgldobnnUlVII
tHvMoCTzKmqmS7s73u0oJnnIYr0fYJVF8zGWjltHk7FuHy4t9uMpupfd0SRNCx67CRVdBMPU7o8z
Ub7iTLnVOmPvbFehN/6RGHA9mNQ9JxeBsW5u9v7cnajbyT45s2EcNwTDZs4aKGMMRBwBz2SxgxVj
5t9ayCrCt/PMLi6uEMWOxINryDvgjWC2B3gW/SlraDcSVLpie1JFK/Qrd+4obJf66Wce1sb72A3G
ihgO3RZU5DmklCrWOnXF/FjwAdEnRxsFIbjVMCnxJ6WJCJIyJ7xO2KTV4R/TTjpSKQVaHkS6krAn
u/02eeIs2aF+j00bCOQxKsBFoYmD3ZxB46jOs0XETQOWs+R3h+Cut9/ymOk8o2GDVHrQ3RunP9Xs
xuHhzMH+bNxx1XbQVso8Bg07rrZxSAP9B41hO0yJGsIRsDdbN11h6VFA6G1+tRU6LupvzVPkGuRP
NU5SJRPp6fHn4ph5BBHSyopaQzjyI83HlcGD2bcsAaa4oDGPr0i6khP3SUOPdigJfHdp7du3kh8r
L3zBOp4LxxNzeueFI3Z6mwVW4yrgG5JHsLkd6yt7QENuEu59VXeicAQ75AehdKVZHk8uKnOF30l+
aDlePdFrqsela45OaGDMaq1qcftlOnZPN4mmq94vhZ0o9StBaLIUEl+oo9B5kR9K6kkiqzFoXoEB
/sPKbawcCdaKWGVa2HB22ycCfDOLn+pYWJ4dD0FzlpvNb6nI6adyfK9PttY8x3BA8apwU960Z7x4
SfSZXc1R6f2sVZhiYm+uQUzaeD/26aS5WrjJIm8z/dSC3e5Szv4eWK8hSeTfCWMz4EjUQ1bL5hqh
dlUdKpL+iYj1RHuukpn9Akiu8NeiZHGxkmYLlm+oBejsnYo40Y69dzwueNeuYUdg9QY5iy4tjhT9
/AJE0Pc54Duh4syIh1wWPnV6Zg4ELjkm/gq5qbJSx17rybMBsZOxNYrehzFZmtaVFNeM9FV2jtHC
9lNI1AlzAw9BuBhztdXOmWTT3CtWUYYrNcAojD0BVo7bs/6RYhwWYMMG0Ydn+daBoIX0ZgieeScs
9F0OHLutR7dpuido4GD+Z0+5W2Sk9N7s41sSiN1VbEX/DJgKnw7MurDnEoJiLl9eNCOLbRUm/dMY
QIDFY3TF53mzq3GgeBDfsWJzgsqK140tlcoPLWWc3x/faq+6vZbWjkMOzEPPUC5qOUV7sDqmVNl+
cqh4oii33enHZu7L1RwueL8a0BVX+gHo4BDfkNroHheAQYQYHIJnzNG+Tspl2hNapwZEss7qby/3
quiKZhglC6BbwiINZt7gpLIFBbQj0PS1VFLePwA9RXcEl9N9BndAIx24n0lL/DkThTJl6Ys5OGP7
z6CSJV+cE7LH18rPHOxd46zElrzbk0bBDEkPbwEURnuMO/sU3yoCh+qfgtMyUCoxlNAduoCmNarn
GB/MxBParq0pR3VyssaftIhA+HKDCx32zJ9iEVQ3skmKezDob9nlRm3ccZR6vJMzjdn3ZZvxr2x8
Z0Fd7ggR2cIjTPjw0b0DrrL5yPMAVMcbnUmS4yAz32qMu6VvcuYupw25tCHkJ0hH/tlz/F4bTVAY
Uuo9huC2+qOP6IvD0kNtCoBVlkKX5n7ZLg7Bkc3YKjaZKqkVleAG/3VKrptOSj5F/cWVWtjkFtTb
HNgfjhf7wxhXMN7RbXYhQVLz43poMJDZs+mWLqrt6zjtSz669m10wXhJkRxIUZ5pHC5G/SeUmKdQ
buQ4t9gAprxyDL6sIWfQDi0sbZWY3MyrWeMR+fHnPFDyQ+sH2nf36yy4qGokeXBLpWmlNxamfE9K
v6kt4UR8eDbTiZ1s2SLu3fmRkWpuoy8vQlpHs24jA+Q+s2L2TAlHIB/eje2ronoYlb9jhwmNSViX
Jssxu20bKmDlV92sO7WVrGzL29Hgly/pXU3n7xT+nlqSOzpta5jygqDLbXHOR2CqmFGvL0x9Y731
qqCOMsDkkAT92fe6l+yLHTd/qGqpiNVCjnxj7zVgvPkfxh2yAtBNEPq8DK2U3vuJrFgaTaFVKwZi
SnehE56Uc9xWzGGChB4RL6LgbOLxLBpZmaZb6QLa/jbCJX0+rIohFBSP4UVEuAPE/Ts6X21mCRlQ
mI96URV3FIpqL+ng4bILlMek8P7t7nY/wsds86Y4j3SrdN1z6bZBGagklj1vS5UICPY6xztiYV7H
pXbB1U9QPJMa0LN8ryrX/xO+3E/XnwVQQVFawUc8VFWuxEwHbPvOWnwU4Sgpp5pvdYW4LWnlxAXQ
oOFAcJJIfOPZbMTifkqVeSzmUSwyWIxZ1gJy0wBAls4RdABWPpIEeV45Q7btfpfXDahUnMHem0rh
N1MebvSUm36wmNmYU52dgBhavuSfv/LvzNt9NwUu0pplg/glHM54O68gExM+p8wtGatdogGovvYO
2br8UhXt9BEOFYWqwGrO/x64HUFUFToXaSZyviLGgysvasonM1kvQFkZV6sWjkjq6GRptyJi+0XA
3nasgfH8RweSi0zdS3eg9Fsht5STjh5WBmn4aEOWs7W0UxB+2vaQ+kAqmmxHE2XrwAg1XSJ9Y9r2
IGXUboqTjz1PbLk1cpQ+jWbMQIQ+svsVYh58rv6jwOb7QDgqUXTsbzEHCmcVDf5DDXiBurGe82wx
9GcytLa2kLhzM8zRoTIMpkCs6wakpiz9Q0q1td5sTwWhtk4Q7+Sjdn4VUU6wadgPtaKwZz8Xz7fM
Oqy50uoGCRAUC7LxorcMdbMDF6zZF8tECaboAZ75EV6yWa+CF/CHY82gEfRKw7s1Gu/OwmSPIbuB
//2B4Kmeq821b/dDNVVygJFejac3EanfCZdxu1AWUy9olq2a8f9rhyHhWve1Klo92lwe3ayr/m16
PkejIAvMw9eshTUzwpcvuBBvzlCyTCptV/uNW5emkjZc8kbgMc7HWqnCUL3OTNzRimvmEzNl76ly
edKGw2TaseGWYkqt+ZulOO4I7qUynUCPEMRQOBZZf5vxnyorTdJX88sETmh/g5Sczwr7tCImhkFY
7uLXIgo5PtEiP7fQqQazcMBPeAc+1rESKuRfWLfq2bIyWwT20elOQpYn9diPri93X/nsR5B99efO
jOZkTuisUaUQotEU0lw113Yd38oxzdMYQt48LdzB6sr4fnany+3hvJHEsdYVLwZfojjLLJNWVFnk
CxUb3MEGTGC8vgUIo+vfUHq24OHQYLEAP00armnkA+JlSV2RG37NtT0bSLvdDf/vxG/SNXNLWZXp
GElN4JvgbNaSt/Pd3noTLiNedD32rJ8VJyCoZxmL9DcLSvSsWz/FC+YYA9oHHEYqaYPut07wAppA
AmELKHs3/BeXFQ3/5F7+4oKRUpXq9/+hZAL74TYyny3Z0jmJMdFTj5X27UwfhZTeuCnXh4i6utTe
HRc15G9LPRnl0Do01tNv3gnZ9NkbRpnIuWFhY/3mcX3Nel0pfpKtpOiNfUxUokb3H2CETexCkB9r
KAEeV3jsSkiseU4oXLO9eWHnsp2hRpWoFWj1Iw0v94RMpTt60+fATNetjCSeApZFEUyCd3a1XhtH
AeDfJsQPTbc+bGu0HDVmeydMlNrIXotyJ7S0miEE6WGkdYU/w9jmBtGqFGbwtEfMCQutUGfVRTyy
JFdZNXTykktg+084I3AwSlO9P8nGaHSWg6M1xlaIflDOVeLq6SrNn7g8Sg7LX3khM4r6UumczfDw
uAaubT5uEadgLC655jupvZUvE9KsFxIKZjHxlGXh63FoLsr9wZ74f6JmQ+KJkduPPdjntX4f735k
DE7Idn9TzIVfpwI48HY5ePZbooMryJIRb7NStNWu475k/7UeKJ2JccQYAxzllOoASIcCU1x8Y9K5
DUHH9W8fcFQ23k7OybyrVY2aHbMfOo5aRKBm0WKYbshSK80FPd8uDmJvvUY56uAV+cdjTuEdnJSw
nIzyJWnQOVtE+XEClWnPgYdN5H/tICQJDp5kWSs2UnTQUmDEqcSMpJnfwCVJqHXiqm62EWIzyoY9
gHpCmJ8tCC3PZ9d0NpIZghmhzlcbb2ouwbQMsQP/wv3UXMSd01nojiOPr+fZYXV1mLLWuaSMRMB7
TbuDSmmBTTGcGD1+6/xAVXASfhMKYGUoD4QBWpvOKZtKBVA7MZK3YNsFc8GBOGZ/Dofw1jYWAh3p
0ThPX7bxwii9h4wZHj/sLMgRQmC9Og8ku4POwxNIOkLNbnGhLv/7ibiU8aanKhr9M/mOV7xlkV+T
o017WBB6dRJvG5bOGvietld4J58EJV0NuelDbItC8XzViv2UMzuuFgfi6s6y6VlJ0wUV7wyXsGM5
YWAiv4OiSh9tt9t6+4JVEKR1dvnMENz7FFSWQhn4Jw1dgilBwdaShf/uxBldWri0Jt07qr4Mb7nG
t4l/5wufGOxgHaoVCOMOJbSdWC2dHk5prR09mnzM7Sb+eZSB/XS14IuPFPYnExqZx9YIe1QEEH7u
9q6sEoA9u+cT0LYjMdx7BapYL3C0bHwN8MhfYgortouOQe4iypUM3rWlie9XsKv+iUF03FJLEnM2
eVMga7Q7MlbZYCfIslJNXWcfMJ9gqfoUT91fIwj9zLFdUWIvmYvz8RlQ74lsU5ILZXyys/HFDK4n
odhpZ9uu4SYSV16awUijaQidu9CGRVmZG1Eq1EpzvoZODSXV+fmcx68QIWtvmSySJWiZ/G2WEfBn
smC6TqRHbKyCkozz4uBw7fw6GYI19Y4jjs8Esug1fAFUj2mZ5OF0STh9Tk0UqorDGs+dmdEYwM+j
RJrIxQ9fyjJl0RMhYtY2daWRFpc4jxFyzqJX8XTmRjhsQo95r6eh0Cr2xwwGjnAUNu3QM0LtVr4h
jjocY4X9rlbBZwZhb2wxcGXZSkwHFj0TzXKELhGUjcsJw7J1JrikMWe1mUAqbJItA5Vz2IWsF2LN
XISq9JsiwzMmFgvB3QTmVXIxHu6v/GJ+lO3jNDxp6OloQYm3Hbot5FHVcF4VvUQyR1DPoqbHKbwE
9u1wEmbRzS14vylSs/nTjOGSS2tEjdfBIZ+/4lLwNH8HAuy+P43/LGR2XLm/MY4i/p1l1qpYcMvH
jFRnj73nLPrRa7terL3+14+gwa5J/oyvrnT3ahzVw4jpwFKwH2p5cMs4K50nQDv8jaQwEao03H1I
QcjVBZ7z4NUw3BEgfweXdoKYsIWYGRRiG6dyiLD2yWj/F/BLNiSAf5Yv+n4NehjwHXKa3MxF0Ori
nyFYllUGiR3V91OYxuKZsQOkS9LULuGqXfXubHylg/8tFWhKKAFl8LYBPnToK+VrnJfDiQ1mCnlU
UYnaMgwidvNhLNoNd49yZApVZOFevZT3P4J8+bZr/D00twk3GAMffBwKwya0ON/bao5SczrqscLF
Mx9xv9COW4BaIfbl5kOpyu1MTkH1gyY2DXv2uRb2NimfEuxShABDLHLiFmI2JDOXPf7OaXlyOOqc
dp3GV/5XxKsRS5sqxg/Te85G1LepELMUY7fngSwBLuZnQvJCXjn+0gi+1eamot3hriGkSg8W5QKG
j6pFsKUy2a5vbeh1p2wNVfAjPuHTIMp2F61AelpylldFMj9YYJNAqXuXkqNbwJ0hK3JOYawuEjc/
8euMSF80h1yCbnFmyfo1a7TaaCgtexm2ns1zlDi+6s9KKsDi+dX/iKslC4okfWwQ6jsdf2JEx8te
NrhLrZsRcw0R+DN7zPECdVBYehP1ebp1GpL7mJ/nAiEwOzncoeNvt3RhOYEJa3eyWkCaWDxHVu3l
nMVLw2o9SCktwlLCFS7a9j7Sp6Nf+o2sBfEUp99p4i4wl1b4I11nsrLCf8lSpI2Aol4eLvxHH9jI
SzsThRFyT4iUpIuY2BxdSISwev3i9oXzzVBfsXdUZZIvX6Kd4+HzAg6pY3bs7bTglr/BdkR45Tgs
fhykBjSxqwZ1xP+vAGUaWry8DuH3ZqWRGRiFJ6uyF36iq4vSoGPlGC84nxTay8Fh4F8zIejDPjn5
YXo5V1vm3LBP+rrC3m+GKXp+C4EKjPaeySPSkdY9Ck1auyKtcrZ0PEokBZvs/z5JXmQ9PnPIRsaw
sXJSPhZREWK3BoWakrp/NI2YodQY8DdhvSOxmO/k3qB6hb8bpWh2TJMjy1Q4FPOgd1/PLVvKLyl6
oWeG5/K6CM1jcs+u3uzjyZ3qhqoOmCC8EdfrLheI6hhoyfpZbpFJi9h/UYyY3XIHW7tR/Uciy4Vm
aE3ssb/IYocUMpLL2ZSiWt6o5vMBJnDNUEOyeTckIR0/tSjU8SgWRpXD34QjPK+Q0NKXDdSs1z9m
BX0hRSZF/g4D22fQPS+z5oHtydzLA1h0ROVkKbhz0feBbmL+bdZyFCU5rvjSa2eai4w8qxFOfq4l
bzetLS6eLX16FVl/SeKjN+yTrqBX4tconP/skOUuptiW3C31oTTYtkkwnkOJ33r1yZZTXZIvRAA0
e4plBppfc4fg8iWddD4lWyYtB+iRJoz6Xf1VbHK2aAv5MSyfnuzOjcenDPWP9Px7XrIrBnZUAaZ0
7uCH/EzRLbgHF0dwBzttwBaJHIDcNvU4l9Bt5o8rL6brgPTfQPlsTXFeBrP8l6oPCLXIUIJMMCOM
guioE6IFqzntNzv8KXlXm5uoTrBeOGK33z5O4dF7EJs+cAc+TVOq360BRuMhlN7pJO0SOqY5qv4J
tcXefco+Jeo9JRi34m0zTVdpovzz8VCuGoGAdFGyUZknCniZYF6HG0lV9m3RrrMboMq/1ugIuZki
M6t3C2rD3RCr9pKd7IDJL5YnBifClhY4XTwZGmo6bTO9WidEVBzoIqa40xuxVxFQhHVNiSRP6dee
BhW43IVo6syTkQjlwHtBzHFLjnGNNEWDUiMuGjPI4hTGE1BCULKeO3HNmsjY3xAxEbTM/7r3n2Si
uE6ornscDvPPa0xwSstCl7wDfLLJdxLAiuMC9FoumOqdNiTyhBGYiIJUmYyTRCHrfAr18M7EHjtr
poWnu9EEP1Lhb63Mh+P/hn3+fmxY7ohkXsP7qsWkf6P8syfxnaF3BWvFfgRD8k7E2hw3Em+cO8GX
Wj/q2O2Sqnq5wZMoJhp1L6NWVwpqd+fcZtJlSV/WW/CkxFn28M+QlmW5PWZ/BWDl+HhliIhOTPrx
JvNR/IDxRRoekjAbBwsfrgnGka0rYOBSEkSS4MUb6jzuqdbXXOx4IFA6lXyWWbhVhVyZLkSu2X5M
SJXBJk5mpIkqNOvWGLPedOw28aL40hmGQ+9ai0iUcyzSwbUznMUAo7qfFBB8AjfvVEZMZtfwFu8+
CbUJ+c33OhEX7EsTecGZC02kYCtFNRgD/ZPOwM7UqCx8GGhTCt570twz5G6rQF8fGKC585bgjxpJ
nV6gmkBa9IOuFA8FGQeeq5NNgz01mKsDk6t6QbWXn+WPvql/VscrRcLilMH147VkooOEQgODuan2
ylW10w7CVLTn58/zgL0dW4jKvCrblTK1kZJV+s9FBgRwbZx+gJzwORuirYnRlpC5ge6zfX964c8I
rYfnZ9BLZ1EyHoInHCQyDSKTeRxLDw+pHGyTGfnOiJzZSJmkmIHaYcpD+3qGTy2qBMEkqRYaVcvF
zghKZDu1mgYNsw0v4/Xnp4qH2EXZJMIvzn4zwU2jHFtBX4a4McF+AhWZKGwWWxbSmTvO2+RWcyMg
foUG80hK0FW4z6xuVnvFUtZb824jUQ832Zrhn/yLWB1i/LriJfg0HWX0tvQ3qvesYvnNuQN+hR52
Xc+MRSsgdANXWHG1ZjmopHsUmfpU3jrPhgxfArbL+kGfEgSKcSbqSIcZhhq3o3qmUqVYcOg5hCbS
Ljq2sMH1sdgEnRFAFRRk/T9Yf/nbsZMh+hZo+Vr/FKCLVWgcwvtWrxtDsGL356leGkmISx2avo2s
SA0OnM30fNdCHQ4CyfxoTYkFW4rIx6NspikrvzxN4gqXG2X83d72E6A8YqTv2FrTYswia7F81gUD
HkerqAefq1KXR5SRw0+57afydCSq+gin5J5bUnWrmnllh79EVDxbrOoPvM2oISrZtDGx7mA7vzcg
t+c1K0h3fcfmk+P443BV7HMYow6teHuUmWOkJTcV+wkMmNfPGvhNqGrPnVS8LA8saJuqTRF0GzV4
Zw5PfihfIpF9dll3p4QH5NRUCr5XSPonq8XeB8nRtgKeJMagg86OFMeBbMxWs+CZxsP47z1/wccv
GlYxc5apgOAcDgBjEZsP6o+l7rjHMfyyzEjsyiBIlsdkg1MmHHyGKmRvjcMuUvv4tA0eCwJhHJrD
7WcKOXnmC3T8xDJ74lyNI+nUd1jnLeCFAX0M3Scln7g+FQaE6qwzW4AW/YhMBwxqVpH3meFdG62b
ZJA6jEKPT/eH9PO63cV1zLiYRvP83FKcS1JuNVz0IVGnibSljITT09Q82wVvU2vGiWyAOHSz5hQq
ZuJOTBjrfWVTKfCAkw0kSj4jrXZbEwCmUo5YBLWFX4dMI+40mNPdUBR5KlR+KxBqBMP8xAotRaOL
bCHIzVpzAALAh1DGHOn5YJtOo6PwwdVNLSuuup5yFoK+RIaXsF4UjM/dhyEwIAtUMHq89mcOPiDV
aEGlOcQ0J9Dgqep1dOcxSpHXDYMfAMZvo+egcg4ZATqs83XvYJY1m2Zg1sNEE87D9lI6pE75W6mj
LlkO3EjQo2ikX9L0cyAvzAdl/O86gwS84Ct8k7wtBoSITSgUtTZsmWpIlUj/SOrVS0Z0gMhssAyO
me0F8rz1gUEMlPhej9gG2ng6rYhLPVAHmls/D3QQzsZsjt8y4fB+BW2Yx7vj9KnqVctdNL/HFqPT
YitPDFldZG4nz7SvvJMmxp2RluHRvVWV61j4Jbk9YhmTsuN2NL1jD14lrvWwZaM6tX3fZy7EPWEy
a8AHw/xzPMFCgdaPWWSIkJTaHIfxKBLlLida57WZa1TC95eXixO93av2DUEP6Hf2Bqg5Gwxp0R+g
o9WDX4S2fyvYJqCXO1MxUzI0pUMENfqBRGB3PtfOtti22KNwrFdIYpfvwsGE5qS4zIFm69j6/aka
67qU9Wj7dWsRAiJb5dtcea+XrZexfss+0WThZIlEb3AQHjWIILu3spDjAz8J0acpDbiH8Yjw5h3c
YcOxccjLyWAlra+84rOZFKL6YRPIKOJyD9X6u81tJ6h97A2Pb+cPPe6UtEfeLRY5vHZBBdpxYcAe
JVPtQN3GwyU/aXSUazizUy/NTRr4q4EzafVbii1pJ5uM+o0mGewr0hjzEkQzMOZTnjwC47Lq5PlW
CZqjeU2z2Swbz8pR1CZSmPjipE0yT+2KCiyyKzpvOsznaNyQrCabSsYpBxwXTCe9NBTFxDTueAh0
76BjFyn7jLcVj1zH9TeFt//fQCVjHLfEI6vDXGxEW2WpLbtsKj4jaQunaWBZmgJCgKy0TpD6HAEt
HdadTAvIYvw+eWnaxpcqVRqcAJR7oTxpQTTPV55/8NJjhYdCsxzCYqJ9zdaIUP4KCNHmVVtFQEK4
72wtwsmZfLCfHWLJINo/ETbeYrxwe59dMcaJPvca9/wZbvQQ+2/5MxiOmCHXfnuQu5i1lVZExZuV
TMEHWTTncm5zSmgqwkMdUMkSwIFbWORVIgtjzII7U7sYF+UDNTVW9Yr+e04tP40DU40VPqQSfqsC
gH5XaX3Cj4g8/++Agx3jXHFESyoN8oJHUU4r1C4CMLA1S05Vm3jt9fQERFykKE9bVexRcUySXmc1
9l7+dcSsZDXZ9W+p7DS25MliCTuLuQ3UoJRUq9witctnm2iq012pRtqTa+Gz6fDyFQZKdbxo3skm
zX6Wq/mVjkF+IXZReWRHmGGQHUhbnKB+svr65NcOv36yxY4Xq4KTX0fY14woTDviRmdiyFHjgHPr
+ImS6TBz9QTX0dJTzGL9qwhAcrgWrwapJXTpkqupcqicdhFKpHW4PCybFJTiNZ00AVrtyTggPTXE
TCa/rf3RHpGKX1il3VSGFwj2gcLIy2638FZj4yXE73VxMkGmJusTXjGOK8eQN/+RAEQw+R1KvmVB
aLm5hK/caBPXpWHaL4PmgHjgN7hUWqZXmHIeHkOBXE80kQdELq2aai0uSgOtp3rlbPp46fDeiVgE
5e2P3gCMXoy+oY4xRM116BGBMVm3RaJtJhMkexb0qKK7LsPtjZOfsuLf4RNDkfXIGOegGotag8UV
9YxS8DjRRc6RBXuVpDZcgxtghuropRgOPfh37flD5FiXzz0ebaNXDDraWFzG6zcaivhPpPSM/3lI
vE0Yy5RKkVx+l/ICbVJQjBRIYkbhRCTzfCcTcSySBQoMBkMHJ5I20q/ZujnMd/ekyboev2uKrlAn
uLedFJZmPT4jnKN7RzAq4s31s7bAM1vhpp6vw+pppN39Bw0VBKu0tFHdwkoW62CO9cNOVOCopRvc
PYncLJ2Y52fIhJyUshKd7WaSxxxfVpEBLT03QNRs/C/25QCD1WvlMwDLxrdxzotjCXbdWvrxdjfk
avRP9Jyhy/VzKHKi8uFCLEPl+F5g4flB7qwjAFoQ9z8LGlgPAYkGPqNiHdsJNWjrz3h+UIxWubUe
pgFcDY6STMh/7PgoeVFeh5pp/2XIcUKyWnLd2sIbAhZ5GwP9df1Wk8Rk3v+7zVT+eMnT8kroOWPX
Lj6WE5O+gNKbUjyO9jEStFp1pYqyaeG843PUmJ7E/mwJ0Dsb1rImADauZS9opbRQ3GSMwtZBzhC0
sUsjw73w2f7X0lfx7Jic5ztfi3l8cetvc3sBxeGoP0sssbeoNue9vTJ/uVhEr516ONVQPh3GWbWf
ul5WfV5vkZK0OrUCvoQaW11JNCt/X0YGBAcrfFphn+CVI5W+ScUHdQxTVl/DnaDfMoLLsUKgU7VY
RpFeWzTUfcAQKnO57h99+VztR3eHkrxLQF7roKtQw09IdH0PMwUkX0Bs1cjeEdhFXyFzVcC78PA9
VS9Q6hICsHwoa/FuImNSp3/LgF41HVBexQjdGdY6TSW42LH28NWZpIpDVes381aE7ZJj9GdFHlYa
hyQAb2epVpFM30kFssaIhAXxRbyWU1xrXE4fFLv+JPJPGnvB/ET8eSE3F3WoOZAoPvWKwmkNUIo8
7O9cjb31/Wxb++jxklaWLwL6fVRy2fUfRfKS40ZSFZrdz0QVK4z8/JTfSrtXWcjjfSbzNOLtHN4h
xbHdnUtfLKCQ/sfotsA+ar35pz0n67O1rvtzi6bRGHojO7MN9/DDggbJtAIJ3ztndd1A9UnM/0OY
Py4UrIalbHgD6F6V6kj4DNw81nhMGhTiloMznc2VN4mb8ahEBw5L2Eb7hM8TV8bnaz4fILcaj7W+
1p2UAjmVLVfZD/PBxif8EsUMadkqWbhrMFrYdobW+Vy+BTopFeMLTf39HefA4CowgHW/uLgp45Rd
i4VtLaVLL+iq1LpRAHNM+cSmQCq2zwIe/9wbMzMdBTwaFcb9FuPknwZvdKanqE7JS9+v6QVVfy3N
MpwRffwrtw2y/6cS+5stL/qLuQNg4xbk0J0iEnq2vGnpmZ/OLhlGOE2YVWKdkrbM3Qvyz+XXbpbG
JxvQ+dBIL3HKaPuSXkf92sx3eLe0URXqLojqFD1OSrrQWaPcYBdX7I9/SZpf5Hrstdduwu5uSI+F
ti2mayIayc4bdQYV5FnK/xIVKI7jkx9VBbDO2wqXH2gMdix8YO/ok4eVvw9QlmcwHpjs/cDce33w
KyNYEWnpIGbAFAp6D8Db9QirmtDAFvU4IQ+IOlPTElOgHalyhk+Hw6SNltPQrH8y8sqHBWb46Q4l
IFFSTwPGnIWqkORaDzPS4SvTMvmKEbfZIUDLhb/lOZAuLzqn/2n7riuDIBOKKkxucR3gHYVvbPpb
m3bamEhYSdFc/x19qlQiQ19r7xsT6fFQWSWzjmUx8e5FMTZwX86Yofu/aLkm8jXNDu3RluoRAy8M
mrBN/5Bsmgj2+iHfz/jvC/7Cz2fbO8HNqvPpX+pn5O0n6HfXLNHraBEvnvdLMX9XNy3os33kinPu
XHMDr1rBKkInxqcfuhUVnCsmXeb2N47j/66t8bOPrmwva+Ivld422SXzjMp1xZFe/9RxSV+635TE
tjphCevdnUTakadJ+ILGIv+FRMa4z1lwXmuNLfQ0TpGAPmXeKLXhI7+oIyRPJUNuo7QP3Bp15jvm
gw458xX5wCjUeGVxhXp0QDtFHKyNTlnFmUbxF2RPlX5D2M81p8Hfmvgloa/uAcfsR0m96rEsZdpI
XO0H7SjE32Idr4lhsrz6M37VeNvBUO0IGeGw6+xavtNhaO50WpWkysWKq9bzIYS37Almd+lGTifd
cbLzwkks0ji8KxMdodpbUA5mTp6ciFaRKuGSZ4GbK1LKrGzfDjQsOVxOWvWudmokndh7KftTjmdx
Bp3tedXXYJ1w+O5NRZ4Vc8z8snVmQb2S5431Cj0D/BroQNy8Yi9PvJBS1mjKjONH7MHO8t/8skKf
niquGGuF1u82f6OYNJf8rkGqoPi77kC+7FRV8ZxCMjHk7Xb+TTBhsxWNU7btI6BvBYiXuoVSpPGF
JXyNAPFVeQ7cSPFnSq9v8NYx8BPpHATwGLIW7sEBDfGAEDxWyHjdC2fGCsknACZIWhUdZADHT/mb
Rc2GXJUWIED1aU9tlXn2/sax5S3e5oy0jbjF2JX+hRBhUwNnpfcRZu6ZXG6eA66xnxcrD9v7VgdX
RrcAwYSH6+sDmcidJWEArABhCsVg1xe3Q9NfDyqkeJ67WA/e1sh6y3HOgDhmlzh8pOlPqyV2mWH3
a4+dhqoeK8S/uFEFE2JkAuxOTivUjReUrgRYvvFChKfE9p5Jq7WM9ye+HZMT+NON2PdX3Bnd9TnQ
xo6jzBGsR2fq6Z8FwEjfgE7qo941enElQKgbE7quzHLuqU3Enhsd/SC/BRrrgRKMWWS6yToLkO4h
YuQFUL7JKLaDtXhquyilTUI2epQ2ELj4DxtUAMNy4VuaFNOBql7rgbxrdzTUTR7wmMQ7E0Z8tSu8
AuKu+uQApceGiLE4T+wa5wdXgZN1R1OCfJpAUTqwz2Cc//bZNLmsPjnGWHVi8u/dk5LY9B09Eiab
DqiKNNB+r0weYwuBzO2MhMWa/bn+hvHIsw8zHg8+3x1aHytlDLIEYqH6SSYFxfoq/OkhbJPQh1kJ
O/U+foYZ+hG/yF1GBdwpNSAWWvBReZU9ldeVGDwvun1EOUy0L9NWdebIq7A5K28y+ZtzlguZBaYl
owE99H3HU6tpK/6hNngK9Zczn4V2WeLyoBA7nlbLgLGBucshnHZHtkq3KYqNEQZ6e2uwhn4WbQOF
cE7tXSFOO3nVLDjmWiFSkyTb1qWw8Y9ff8qlUUeeDrzGp7EW8RuC1FglDxkCH8T3jpu2x/K9sJ3v
uAMo2pJpQnTg0Gd1dXKfB79Mb6BOdVS++OG0X86S+ibjEqTpxYkUGopcH5PvoVGvmpr5xlhPR3+A
jWnhBV6nDwRg7/bUIEdYLXqkV66SGUW+QeAdD0v3c/MKSIRQm+ydhkB/X3EtYOWRrIk58bLWMS3C
DUgnwdftB1liOiG+UjdNhTtyEfPn2nGTtPM0xHogTU1YjREpziXIiElvNbScqHEtio8ZVTYUUb9e
GYjzkkJgx31tipflPSKm0cwBuYOGevVEKwfLpBzh0iM8cuFQd1Eiig88tnmlUL60r1RJhkG3NckL
ozMyBz9KkckEhkXudlQfDpYOABH/VZ5UiaF9IsO9mDANlCejN9wzssbzXv2SYz7fPrAgYQspwIyK
egD+sOMZA2R8ojCjUgquZf14zRpFIGFtv335nIwYoW04byY0tDBxc/isJHF+3HuXCC0znKA9yIIh
9TnjyLY8WJOJRHX81Zaxj8tLcsiDXKjsHq83td6kQPQxWg64Yb2CKraZm79PfXaa7cCo7hrRbY0z
8tmxs03MWUoX6dG7Vk0Sburu7a4Rt4EYxnPiiepTEa/e6dDuyguURNWJibiZwzH4ogFBX3cK5VkS
I0IgSaeuOuGZFfUQVR0zvWXcNZXr85vMOOnutp0dgEfgyQ5fG3PKib/J/HJKr5BlDnyix9l6z/Op
lt2lA+pPTI4qSnTGQfZDsfwCjbxREfUcAfS2fwaBzENPk5eWpZ4Q2PV5CRjJaFl7/t04ShkOH9Fh
RnaB90mWaZOl/c7r+4wYcfvfZqZxCNLaH7C7uNI0wSgry9KP2klrhB7Liyftj4GvKpWs97FtI1UJ
GuVNW5dSqScg2c7UIx99JjZMD2TpNRgf1Y7CoA7VJYO7V/PaMUMGvcKN1CtlknSloezoZ5IWJCBF
9XCZrHCGsQkpcDXToxyyducjas+IrBGVS1qeP4NrLZbjZpIerVD/LlrRt7gm3AWG1TquJIC7XaQ/
RNeGFrQPyG/Ux/tAGHVtCh0CxVlUoB3bUL/3kG8C8kQFdCDWYhVj59e33Ia/flcBTieRfAOhkXK4
bAPTrYTcam8ai0Q+/PSUVLjuSdKi0BClbqNn/sI3ja0Kt4+Sf8zidWZv8wz44AJhhae/9heJPWhy
CsyOKG8+5cZpVtAFEOvWdeOJDMWQK9RkOZyE60M0E4KlDzEL6tTsnkSGpCj5qcp9WvD7celFiGqo
ijle2/YgwIZKE75cEVv7ZmPvDeaSOnn/h+ykuCk/5ql17uIaykEa6otbaBmJwykrHk5qVj7GQ8Sz
ppZEcW1iQ5z2MbVtXSKI0YQjgnN8fIuNUWXSLqIS2kFUPtfUWIOHE/wtSYHLh0DqL2zutBVEaIPq
aJWCzNzByY5bdkQqUdhKMYm5/SLS7brOI3WXTlfuFuUlpWSjf86S/RdbTADyTZ1Wn/eNW2Qv9L6V
het0R6oq311QvLEE1oU1x/AA9xcMm9Et/FDYmKYfHMr7PfKS8rcga9tvbdoF4Dob1mtE21K3n/kl
VexTdLTfybHpDyfHJick0nArrkxtlv4nHkqbV5B25X0Ib97FLTj+83Tw2v/kldVPTP27vAKySu56
izixeK9Z0BRHOf70rfV0d7HpW+2r8ba4y8BjeAQ8sGMvKjkrgmPObMeY7j53jZzZYVb/sJB5F9Me
m+Vc1Qab1tDpUJecBI64IeSMEt6KR/VyH38prp3UBmujQiLMCUq22wH0FmNdYLk7Hsuip+5wCxha
TawdnKBq4b4YJexTZNm6Yf8mVZtF0zU1f38VM9eCSaiH1ouiXOMR4sPL2Pgo/YtJ5VbYqEa7TkxA
YVV32NcSOnEb9YyYtarv4MPft4jgJmHtGTE8pchX2q1Ks1S+TYgCVXvwo4T0Smi6h0mVqCvI/+J3
o381og3IjOdTW47lmkEYShTi8kbJpqHn3py7kp4MtQw488ejIknH7m1l5VUUPzK38J0Mi3oUused
DKrcIVF7dj7cJDLYutH6jFK/CKxz+jKtYwmn+YUadANX7npC+KgxLAnj7zIEvZom+veYXoFZ9Zv6
Dfp9ghF6sPMa+0fquMFfiiiQ2KFam8qWKTIh5hgv2SqGA5abBpQ0RMKfGZBZ0oD72e8brPljqsV0
ws7edoY93qu68cYeTaicAJzQaZ1xJy+6OJTrVPRwLNwvN9VaFH3HTIzoH7Q0AOQJRF3IRTQq5o9g
el2huiSDHd3WchTaHuvJHgz96erXoQiUIC6V6cNyWnjFzPsJZlI7FOy7lOAJcPOfDkFyErxuaEg7
V1GuL8YKByoDMNo6m7Wb+yVT/MHNF+I0heADERwGxtmhWE0HBkZA1U+em9p4kvBd6Yhn+OIJaTHu
d9UAH5ZTNrfdLLnlM07MTEeWyRZZut/dK+i2kFn4gDV5XRTBcmoPY9hYw6NXifi5sQ/t7eJl8ow3
0xyG7nBKOnQhz60KA6jayulNxewnPhTNOfFC/NK2e3EpqTVvApPSQJGkk4VWDCHQVyAmH16g8XSy
W9sSB2d9eoUVykznZLj0rjFR5xj3rME8Zo4p+ZocYEubgb4djmcCqhYj4ClKG+pVHgrDxcBPIS8K
8CcS1vsaT9fPrKa28uXsjcOSCURB3mDL/MoE5IsNzc3yqwDglm5E6FLypkMbO5QPaHD8Q8y7mXcX
PPIjaNgsdxordiSbLHssqs1bWOo5iMm/VyyvYjwAFHkeSmiZRtu0szdX1pV00Yu+/jWCajmz8r06
u3IhZFCRlrnZ6hXzvKLsumwrVrnpX99G/JSAowkF2H3Hxd4w8ET1fmtD7RFUm2DydBcmu1EhUrEx
Qn/yTTw950XWh66JOcwOzBG2omUUn9rlMxZBCNburPbH9japNuietMiksIwktzqoTvaKVKBNTIWv
F4CmDWFf6vq/GD9l8xJGrRsEmCd8QykaIQK+C6327DV2Ro8C36xw1rjzfcglunzrDQbAvktfpKHb
F+qOquKDGhBMwQYt6gWqZvkJn3kx6zd/SeShxV7w7r/Z9+YTha59x5y6SID3+++Y6srwSVLVq2if
EJtV/jiWKtBg/FemZ3QCu3MAYp0hk+WdEAaaYVj9IbggkFLQFbtL20NLusxSc10u6647WAe0ulvW
6dgKsu3Zofn6K7MGdJdQVEvMcEEEvMdKElQMGe64abDyexCjY6Yw0LqbaLh9el8A6ma5kqeNtOfV
GV5aBY2fWI3f1mBAKKAy3fC65+P6AwbQjR+DnLMfq8Nm/teZyHXSNVUMQqTen7WZYBpQT4kaocaR
gqtri8kDv9UK0Mhdzn2c2SPC9+gl5VHK7fR7I+rUkJ1NaTpi7wuUXi6cmt97o7ETcV93T2b4C13Q
+Qe1ifJ/Z8CMFCGiDntYAX9H29BnUpbijl8h2J0XMhzoAuSNY+3a/7VBR/FLdUC/Ks4E7OgcSZts
E7L0iuzAaaOBR/5lAnnqNu12i/bRmxDWh7ZFHT18Q9QpPvLdGqSIxq0tnBT9M5wMZfVt4QeatTSZ
mPIS4vxNzmTRwJHSCN2a1/tQRFtYIsPVmFB5HjBnb75CabScsFlYOHLU0LD2ty1TJdpH1Tuq8FRh
KTYD6QN09LvQ+0iRSH4HIeD6t8mrWBBRMo5pQSV4NojzNAkIizHzhacfjIQDjwcJHnprXpTfew3j
dNQlyIwXkuStgPTZ8ngNHhj0Xgy+Y5jWPZAwIA/vMZO+zp5kVyDu1ZQ3q+fEONt2qOVNtOdBdVOH
/+TA9JQxB3KFLImmpapuwBgkjU2GinuYJX3q9NU+dULQT2pDcIcJO2KmmpECIPtcBLhQ5ksjDhAq
TiSfphhI2CiDrZ7xMV4k5YICIo4Vm3Q+FzJiw6zzolFQSCf89nVhei5nhjr8DTgwLtfMIprFJ8Wl
AB0GY4sd2emnXA7ijnGx3WH0RknWVxOeCEawezBB2MawqyNPtTA4Hqqb6ts9FqPMnu14c1lFxdkN
zWhsKKD5FeeBdDlj2A3+9VTmYfiBjuvqmpK9+5FlVqqn9cwj/nzaP8lYva2/AmLUSbOwJ2XJ3aAN
pQ+R4FqcSnofjglqDmQafzsn9T4zcCVrZ6vb5r6e7fvoBW9H2/Y3nDlUure17PiieP7DfcElmIIo
SBtJL08GRwq3BmflXiDu4V7Av930G8J87TIGLgs1wImAozAAQrm2GOOYLAf9+RmAOuHz+ZJIKyDX
zv0TLv+BqSh0e8Eq/+vsGuQ+oDGLqeOrvGQRzpby8pIP4FiHRr3yAaV4N6W4mjAdATZ4sn6EawlN
xFhzXpEMnFiPgCdQMfxPTMQgjb/73R043ad3QZfV0EBnsLMDaI68pLqySHWzbd+XbTc+SvR86vlZ
Bd6O+P29cSNRs6mQKQ5jTbgU3MMG3inr7pkPk/o5HFt2MokSjQLkL7f14x0vETZoz5zSkXiuj6U0
ecHcEeYaR+P/lyz1tGbPRssY2S9OT+GLb2hTEWU/nYYz2mEVdhMSWvHg0PZ/KISXZ3JrwzAGGgPf
mUdf+kFiTLIb2f8kOntku3BjEbGiSv0N/RZHePMZXZ/pUJh1UUGDfkw52NTpnF77oluWZcvWbQ7c
pxd93OYXKZW0eW2kA2Wc7ZHsu8EDboDrQJBtf2kZms6gWcMyONFTy4NmgWuXZ9tDxXiXcVqFA7yd
BXznerSmsXzRS8oC47ZxBowmZvM9tBHNfBErm6di2mSLnarf1w9yjabJs+ottLHrQMpIEg1/tD40
zUxPZE7lL0Rd8PLvO/wHUhKwB3c8nzmk1ofwOLjpl+0pElSxwKHKT2QqaDak4phEEyqbEbhud53i
/wAFqdN28Ms6gAGSpec1VCukp9ebiWTl2EdqmuFChr/GQKDBPV289YJUl8mHeB3gRFo6lJywUjWP
dCTcqRa/5Vz4sGBbpT8AxWWU9s28taxusk7M11Q6vq76A7gcfnkG/P7Vrr0lcKpAVgvcBGwQkj/Y
QdOarLLTalWA9ZD+rOrfRHy4x0d6MdTjoRVgZ//ImSye6v/47HPzSqq4P7uPuj/YSur3dbjDWDBv
w3bjj8JzLRKohP7/SO3SoTWBZLUWyBdnEztrHwcthBmqoudgvp28043Wtb0TZifE1guTjoPraRid
iNbsR/FkiG6msVDA9UaNwWfTU15zCE7XVv1lkcysfpMT5/kZOHQob499ZZUG60dei+Rfm14Ll804
FPVLu4UJTfv+kIaznlXOJHIzyuVl6mZ9aU7tRsGBrY9VoCSCc8O+iEl+tVwuGw88Vx5c+lUHq1OG
6zvp5zB3TbG2cKgjyCQWPDz8QZg9SnxWASei9ZwtplYZlryWr74ZAy780NJe41gStvn+k6Nx16dX
2k26ybXX6DFzxGeKvLJ0V6CHJsP7drjpv2KDK16VKWTtCTXzrrk2AX/wSBWOavvsmKmYdy80Hjn8
u+vC/m8ZfbuNlUHVUMaKlmlb+o60r+fZY5jNX+QlmAR8WgBIR4vqZAwJiHUc9lfk6DKyFrp/cBV0
36SbuRYgcAGBnBjyCPizTXGeokDKuqsCbTED+T5OFW/MLVjOeNw9LWPWFQfGai+wiDtap1P3IxSa
F1QcWHrrPMTuU0OaEIv6LD516nGR15ULRPkApiQuDEIXYuK3IJEqM+iCsKCpYfpFHSToNSTJjnCL
dQQ/ZLMpIKq5wP7t9aw2uXPXP25pa9qN7a9XJkFf8i0c3LPQUWYA/m5l9mHN19MDkJm3Y9YmQ4pV
ZIDoQHnPlJrbkf1TZNK/RS0EZPmkltmo8YW5qQ3UQZO0pjdLMbFgPawOqQPkW6IxENCsc/8HCM8z
QjbJB8zEyE9fQzm6DnTwpVX3iKacwNq6Q9CTa6tXK+iEYxx59K0a05y6xsYxgmIDSbvLHFh7HrTe
wIBUmkN/zhAbJUKlVQPQzWAHh37XsJKOZWyB+ywQikPXLlxYdhtw2/0QoSW+ZzzNSgZUZXXPUgSO
6frI9MADrbDjbE7vegpnghQlSdaCpoJPBnptPRDrw+oFYq8dP1O+8jb/nbwl5hy2QR3N6o7+vudB
mZpEC6Ma0Orh4pk4hCRSwSH4aBgvAY1OMyvTN6n4ZNc3HE/nyTabItZWfZ7/zJIynKha02qpxY9r
O3cbjiECk6g8fWuR2B6/y5ErdCOx7oaVJ9XYY1ZNicc8BA+jitm2rHEYqlLQ3GYug/xMxkrH+N93
iLFR5RUXx25B9kyp41Ocea4ZMFWKrhk3yXYYQ7igyzo9D7lRNQDo8xpR4YlzUQvb9noXTKiib9pb
xwYsJlbOnex3bzshG+d+Pz67/Pjj41Q+AZQVHX8yn80j4rt3+nf2JqZB/A4yMwe1ZH46JBhgfuJS
NlNjJ/TjgtmjhAwddVXkS53qxW/NJKuU35tp1iWgrS7znrs23gqrShmUCLy6urlmmJZC0Ahvc77F
vZrJMXxtKum6x8w1eAZu8iHqy13Q51MvzNFaGdPHlEvf5c+WtDJDM5B7nX40ij6Od2SiQgK6xuF/
xHVEbp2ACTzK61GQXDLdPCUl1CbqagOX3UiGUFNxg2l15ePEzo6P323HUwtr3+JLNfyM7AmSB/0w
UhNI3T8EUm4BZT9c/xMryqqB8b8ys5iitCtqHLN/TbQpX5ye8r59u+8O/C4mS8ile+FKrcmWH3lK
YOwpzwwSVxTq26S5wBW3bpZoGajoV4rdSMSVT+cNPWfZlrSDWRXX7lWwA/e+pPMaYmjESsw2SiCe
YewInzSmJwh+jLuTa+C2XlxFxiNEvqx2yVSxvBE18G3u4ThM6P9cgRirjHBhIi4gHr7RZcshDEZl
6fyWoMSg1yDRvnyIgeYxD6U/Iqd87rnUJ1HAH8OhKSCchj/8QhDHiJdFUwMjLS/hViws+X5vuBxq
GvKDw20v55BFqKr7JckPaXKQPziuL9QdlOt2L4u1xH0hDPfONjxlJQhOvkYqVIDFoIzkKf6vpFG9
YJvo8t80KJBP0ErEjdNbWMoFshEu//cQ+scV5hhcUinQfcCvU4zMDeBAA2PDKgW+kk4OGAm1h38Z
UaaFbPjKGOUlVuefWiJkjJcFNtO4X0FpxHTG45bmENlc+quxow6d8O2Y2FDCXbgwFE2HO8+lFtRH
RNnoJ11pv/elsL5byL7TPNnRKSYA7CH5qQ1G30sN9+0ltrWethqmXxR0Gdd07wlLLa9YDqi61oou
5jzT/pVTZdCxtatewjHZnPv/nXMqIfx5q8RTvfVrA8evYJ1aBoLzydUV2BZdzcxCF6IlTy2bqFK5
x0o0V2+mIAfM0XobsWYkplP63Gx9WlGRRReUHXYJu3Cese71zeLCWRMsWPYPWaU0N68TmjnAs1wO
6y+bdRD90GqQH9JNSLQywHYUOn1os1jqeZDeh9ji+DnAflTTLXDXfz3SJWDZQv063KNe1jIlc9Vm
FJgg21+yPXR5YUpPw5yWPHj8CywuoJVbByRSK3VS4e+KZrlUIBWxkbBdUUQKSW4eGbp0m8Z/y2FU
swCBjQamevQd2Y0eB2YLLkDtIz6jjnntqlPqapci2g3av/AAUWX1DQ5ZpGyKV7lrkzNhjZpsqVKM
z7QkDWVEEQLLBHVKaenoX5HPY/jBb+dHs5W5P5EbE7eie6VjIpzc599VbxgKWIjA6hCUEfVdXSBD
eAikGt0JmRVCIgd6+/kbDDjv0g8bcoov9ip5tHskexFzZvMKX9nWDav7XOtKWWHeu5ZtbvY/C5+Z
gTYnRpdwjy148EpXZe1O9gYJNEVsIqInFJq1sF/CmgvQ8fbqFPIMFYYrdIjV9br0M4giqcWFX87X
YTdkqE3pEHuwg9z1j0CzIdhSCsGDH2yr3t/X0usr6xhAU54AYKiaIW1ACeUVcoI04w3pajKYj0zT
S9MkKU0XrzosOy4H4n7Y1xhgN/tp/wKCeTuKl3lJHK+I68WswNDwXlYTzea9PXDaN2Qh1Y+Q6SV1
8YbloHoEDZDR8S872LNWBV+oW3HkcIlmWdDu5xIyPLv2M27PUu+tZ4H11QZpCaY8BwKsjsxCktU7
jbtg0RYIu+4FA984bitWl95uueVnSzb5JUXSS9RchWNP/rRLSO6j8UbR8KYyZgcxXyRHdMx+aGfL
2qz1uyfcOrlTaASHxEireijKd6HTfx472NWrba+EEgermOt3jJnKkKy72Qe8aj7d1fAaMQ5sFn5J
07m9zxDqRKq+u8tuC4P7QvH78vY4q0CBGndESJIgdHBuEIEEiK3/FCOLRaI+/Je+ZWj13KMTNYRo
4THCrKSnZ26sDfgg68AHysUNYGWCHLDF83jC+BXlrpkLAA5ljj6NwsIkZ1Eu5xI0pUFDlonTZGZu
wdn2vDsFByo4F30+klPhxsqlSmD8/c0cTEvYP7V3AaOTnarJ7eGOWZ5NNhcJ5Cail3PKds2zl/pL
1i/SQVRclp1UlkaHUpWTYfXmTKMXeemAwD9jrzqmYDhxSgOl3APdh9ty/HnuDM0bBrw8OrGy93G6
VPydA7SJsYarRS3nsIMy8d3EMM661zFNTNuKq8kuyD/Xx41VP58QYMAfhM/o/auqop9kJlvsIQQM
Dl3gaEfpR/+/hTjyDfmW3LrOIG6oQ7hs2Il2ZLfhP6EcREIQ+wKgre1f3H/do1W1k2uiBciZwLEM
3W0b9kksEFrALhWkNpSb1klSSY1nVCPJDKJvjTk6HS+zhv4mOKhH8896Xn0sxqjSXYkI+rLTNnC3
BPYb3cJJObkKDNAxGqGL/QgCnDrMQvqFBlEB72DS/UmUS8pSy7mZ9Hh956CPpKYXx7A+pmWIHfbM
SQEX6p543CoM0IuF4HdCjKsbM6NIba9IKfJLgG8Qj/vy1GtsGY/FyaFqDkBCpRyBeTzaVXJDZ+f0
ZbPW/BSCGZN7Kb1YBpbWJrWICHBD4fUmujJUkaDXN0f3x8DorCaBJk9FaKE+iANJvuNC7W3341/C
rD1XI/N6jIG398lZqHWJgS0djb02wfbmGUgPBVOEAql/4ePJW29N5sSrRkduESofVIDLBDVQpZPR
RETPeTbf+1JjV8eGVBp3nhyi8rXdSyFOXwrp0GhHXwphUNAURXX6/X2XV8G2rfXdS47NrxuaRyeC
kV39e6elR2haUKLSl5IPznTI8s5E4Axe569MYE/nTf2PRRIICqsPzm+tYKhjgx9jnM2vLqL7fi1w
rf06vQ4weuJkNOnDYfofmCEmGS6BJVc2Ru412JPsQTxA6OYBMT961RYHYf1H7CetqLMyBHaVxfpW
KXwuyHkvsQ1/zxHilNOaBneYPqXf2VSGy5plxP3gAXNovpPTW7EIlWLutemEbTUGqFezLGkO4MLg
2YlUR7cBkjUBzUcytaTtP0S1iAfpAWl2+FeGgmit/CFYmznDj16VyADtFCOl1xZNZUAuOOqzzpGO
yyZuZLF3FyRypvMK2OrR/KsdE9JFVNtbsgO9edM3aQlF/kH8M4eLgjbgzqVYmloODJCjZ9/xTajo
rpsJUI90JN4CbmmbF+FV6ETl3iWOchzKYjxLkvoDxLGgNmYPRIuL2meFJvadkuI56mBmxT8QcvU1
oKYUpqL93h/gKGNu6KpLfOzs5UrBeoRQlDJP1bcnEjzq960Q/DRrBIRTgmK3RRoB4uoFnvZI970n
yNYL6ZnafGotkBNbQbPjxn4Fkgihy6jLBDO2cCXy7YG9Ck2Er8Na+wDkkBUAihxPEdfBpOY6t5yB
sIgQZrFSZNU5MfnRtSwKadZ01Bguo8I2b4ummdqvPBFEN00IAckQGlw6EC7SjAArpwScrm7ke620
QNFU3Bl75y5FQpwRiD5Kw6MEiHLYNFKCIxpfq7pMjru7mmEx/UvCQn2+7BdzZ2zPA9lqdwqOuPFY
hgccb86yNxEXfG4oWaFLKYkegByf+Y5dkZDh70QT0+OMFZM4ocY7bI84imVdaaVNS8ClqSlH6xi2
Q8l22SqFRxp1+8mYOusOD7RiMSZKV7imLX9eh8ocQhbmJXP7k+S6+cSpN//fG5tmuzp/hlPWDwBl
5dOP/Op3Ty7vGNPz11AAteMJV67d17F+HHP6bnqdv1Pm21IdE1Ll48o94BSdxRUpC7BtRmjqxlcW
oKzdKXqRGoiIxwS/DY78+HRHY1J7XvTekbNB048mYjTRzL/nyzqVoAw7bHomOQgNKW9rUGux2hDU
Pwy9MToEL8pY0D6WAYVPgxFmmoC21+TApRbsTt35RIstmaQV116VJw/JFarA628k+WuUz8RrclIy
cgnpLIaPzHB9BG7wa949tmd2So0I8ev/hzMZ6xXMERuXvUPH8qP5RGJVzUz71OtGYIH2as/5SXsH
PfZ2DOCc6sjRRkte4qBZnUoPhDEWwEu2HjQ4bgAAx5tNobznJYk4Obv7cS8ynF+8NIhazRScjvAK
zXzQx8j37cmkcmZS2XQgzijHyy9pfuJvhfTGxOuVJM5XM9twbcCCT21T3333AY2dWiEAy11MpK+P
Lvtd2lRPpuxmMTNqltP51iI221jkU9cboKhi/HmGqn51PoK0Jy6KSqxaim5WZLjEtcMtN61jioxk
JT3dt3dc19BIC4cvGSgBk3IgBfcsmYX5lsh8YUOm1q5PYF8LbV/G8H+/LMNrgRtY0kAFRcObGD+f
AJZdv5n6kcPsRnQ0hy5IgzvRB0jUCmvq1BACBrlQpy+bnfuaPVpe6nvgE2ilKLT4B5dQWFKmFYKg
51sZPicDAV193ggyMGhtAfezfVynssOCy7WvkRtFSLIBU5TiXrLSlgu/yITGImnNW+LoS2rUit13
xz9FvVKbvEdZEmnubrrYX628fs2LHfkPoF5BJtGyydMJtUdiETL9Y9fsuOtkzFE/Xz6G/3W+aj32
ivmo8qxgNjr/DdHHlcdzlLMwhnc1uS2RPakFnM4/GCO3vrlLUq9glEJCpSQqHvlg0oWg7jbs12fE
yjA3L38EwuDkAh5JUtF15CBGHBfE31OCNXnjx0p7l83innSc1HW8YqQ4JK+XtMvvg/cKc3sWMGKk
kW7obmlMWoZjqeV5XceVzKlN2PdWg1N3NUUC4VchYUhf+DGPCX8/vLQvZ2AS6H6jBt9q1PKTAt95
xBDXJGcL0BHZ0SCmDOSDfCEvphDALL+fuagAVpbeV9wHGhiwmkFaUwtOADJ/MJXnLd8XNNeuwFvo
p2O05jnPJszsdNsrdeTjKdYInvhdUWyPv5MLqaiUCLFpvYAKS0WLeChaOcBlxuPYc2XOklm8AUM7
oBblEF0StqKy+hQeKEx20IEsVk7nSygw9ebZNj4VIJqg4/AbOHOg2Wt6VznHRnyZY2jnbcwuxS6r
Z49VQzByu4VAUCRRFKoPQDCtxRhQX433BDjANWmHZevaMvCCe594S2aIW84I4Bh1cI4qkCmhYDzn
WItSTVvpEnNQEh4FgMxuDU3dGJbla6HjaFMgwheQR3+xa9teoXJ+fuXEaVG0NCLongW/Y5LjP5cx
IEl4sjpUNyULiiWWdOM3W5+vbZsu1MqyPjNjnOUsoqIUsgcZvSdpRuT+A0qKNqfKivWuTCUjZMuD
ZughbbihnfecY5bj/30F+QRX/acM8Il2MVu1hdJPeg/4CC3SrPcxt9WuiL5jE6KzVrwJmrgai/8V
dSHUVMMKZ7qmVcpbsuw61MsrfHRtov1JpgCYDM9LU0+5miMGf5rvo8cDiBEzm84FQYC1QzTVAH1a
b5PQe2wj5156TY7zTqhDPDFvzBqP21M7Ucxf6SPcyYK1+MqkNxH4HOv5TrqknPMZS0WI1PK3IQlJ
QXcJh8jwXBlgqn5ur642SVhEEqDQAsduLuFeUT53qhwb2ltu9kjD841fi3YYv0SsxdixspwyHpKA
0gr/gzTd8358ABhfiI1F5Z1csWhtKU7G6N7Xtngs+YyWzjlqlJqQiL3awkYq/I2VpexDEir4ewmq
Cn89ksQu4w9rciNzFVXXIjcpkqV9lXhjrHsXaMCq5Np3uGkqPAM8L7MX6AVBcUbZ8LDzuhD2+2Oa
lnonnhtMOHT46vJxDSpyx+pXOHPFSjIZbwn/2YVizUe7Wk03i+L7sr9p/KoUfnljjcm/kFEuegnA
3HbDSitBsJ58Sn+Fp3pnSp8eKCTeP7HF7gdte5RSXjiF1ut8Th6ARIkQ4uff5iYEmC/5kdFbtRrn
3bb2A1u0DMbiQd7EASozm0Clgtef3uZEvcIpNN9PcOQLBPM79WcYcETyjcHRM5bBb+GKyQULV3zq
xeb7ctrQZhkjodw++8kjiLcVWpN8GTf1XOEwl1qEFjU2PWsq+ie7KDgKLuoVHkIiiepOV1AS9jn3
RaZuLmNHvoA851UdwplwNKHriHOU6408Pf893otiELQ3lCPy82u7xnoz0RGpvxBvpUGsG5sENxmN
rx7mmnalcUKrXIVcnVL4WEQSyyfGQqj/u52DIFb6YUA8o1ttU8kHZAw2uHFzn6s69BVDVe/uFt13
4vQJRidpu2jmdv/I2aeSx5LrGn1CRu3eUKFhJZEmIWodCGjxl+3wmyPc8ara7DyO+EYllYq5NRc+
tjA0s9In5qeZimiKCroLoq8zezqcZtVYZr7j0fILqpzolivC+hUq+HhtoLcMOXfiCREt1L/ZYeQp
pSeXO0y4kZ9SVSXMsXsB8A/q/+aWkjFNMeGcHhxi4DfhFUsJX+HQ2Bl+s1vzGvdgj5/zhpAgRIGv
Fn5DV720fFj0ns4/BRiBNZkCeuogtOBNYDtUmNEUPmMZ0lW8vsAjDH7eDa+uvNnt08fcibGLTTNK
79x0hWxAKO6F5N69x2Yj9w4YHCNiwUBi7OSG//uD93Y0HnONKox82YW22BVG0hmE5K57Od/smRQG
CG18Vumm3nmjycxbvvsCcTAAy1p4Xweao3gPDRA2b5Dogn2aynuNEN33BW/XaFEDBhxPOXFS4V8V
qee0zUh5hKUcUxbaogA40a9wrPK2UVA05TBvS7FDlsEiA2gB+Pw66/q2b4+mRGFQjucnsLYRI5qm
vhV+IVh9MoGbKY6Uae0TmrsDyjYcEucVlELIXMCWSSRb8iGTZDaWyKQLEoDvjCJgKxVFEve+7036
ySFIoQdOL+OI/Z6XlZu4oHHjZEXpiwcMNlP+x1/+/Kf06fElTVdbuYhA7UAXxnvjms2j1lZHUKQP
+NcWhZ53H7P2yDgdmMJ5JHOIZpRxHaVY52kFxNKdAslanypeE53B3wVxCQU9RfI+k/bhD4IWssTc
2i+cPrI7aB0hERJuQ42zCpNPpk0F4x1P7lLjL4R4i3K/ok9NIXVZasz654gUMumi5ZFui8UYE/vp
DXCL76UGVr7N6feO47hY0wpBwV3xFvoqpWwfxWDiu+MiQU8vX/LX53WrMND8ohumZUjv477jenrn
VHrg7VaxBHyasGeZk01d9kVrD/X7pbi++g3x/rCvigOPoeyB6vqzq501olLZDIF1J5yNnf9GYBVU
XgG/nMXXLQ0c0B8M+Yu97ywjVuD4tCvmLu2fjBdGPFImI+s9twyF3oAJcEaBlLvWII54FVtsAOpP
+ZCajH2aN14sOkv7Zf/UJiGb7iD0mMtFMJZV/QVKNgKiEvPcjqK/NDztAJfwg6XBux5IcKJ2PeiZ
fsG8j3bENZgzvwEKoa8Ju3fCUGQCgy1yc8C6qEvn0PtwRu63emMifDaTkxfChALjzaCLLcJRUjAr
c4LNiccy9+ARLRi9y5jbC3LnDbQfGvSkubTKlU3lHYl17h4Sjn0rUZcax/TKCHG8mU9DwyCEHko9
bs1q33u00fI8Z8D3Hvll/lGfcRXhZzNqLdlET1B4R7mZgCbJWIPcEnCkOOc0OyUqcbRbjHc3k+9H
/LfiGGOrzf/iBYJmuAUiQ8U39wq+Y2mdtCpmGjPtibQ9C+PVbJIqCyCqUKcB+J9+sQ/ZmXb7U8Qk
1qCzxkoP/6m4r/Af1srlypgmxC8R3z8pPKLlZzs93nqpnyfDVcK55VxMnWqXEfQP2gQrX+HXNGar
EkZSOwieLWmu0zo5htTk9XBGmHhtCcUWcxzoCG4S5TRMfPMFAjvS6uYjyPd5IQ/iTQpPUNew7/Qf
pfsU8mTKe1KsdhHauRNKIXb6FK7jKjPhx96uCtRb2mVy2XPNyg5xn9NujHAMIWGzUO9Ey6+mvcp0
U7ZSNIeneJpNNWmj+d42V4MRLQuF/JIfsaJ/QNT9+3UQSvlXAmJbf4hkTCNArDYjWJzfXuYuRJzY
e6kwUnLJbP4oMwzihkHy98y2wSlnjvmRDUfuAIteARcTaM7lzbJDl41yth7Oalu5YA6oXrvPAOx0
F3drvTNx5caEUZyVOszmJKx/gRIB6rGp3eBYcacGbCdnKDmiMNguZ/Nls0MXUzjTo9EbEDya4OY1
4optVojRbRW8bkotg7VciJHNDXTL9iv1r1ViXPYkTaS+/iqWLm8rHZLudC6BRI76bV80s5LxilAI
n/4h46Q4azN+DNaq12BmfVTgEE/Omq+A8p0EdvESYLTjtaCYKrQjYR5wqxK+6IEoK4Z45uaBymBQ
3sd1hHehnLpHxfyvP73cWqKkmDsn7Uz/GQivGiOGGDw5/jqJ6AckBC/bnIV3l3MlAMkXxoZSQxdd
ALBHOmq3dUyQ3KWCHKbEqXC3XBlFfMv8clozleF+/yL90nzeYLzBtlP/7FotgURO8Ghl7pGSQ4RN
BGtlFxGi9NBRFn5+O6pgOHgysAzANEFLaNi7uIf5ewKW6U/PFLuswn+PdqZkwHd2Iw/jaxDKQSvR
Loz+PRieLBwa1gBcNi5uK72Xa+ee7alWYK007UhroDZd8rpT6gLQH1IXohCfbnP07UZNTKWTIiTp
srZG9kzu3rGnhPIBTWrISzQomzN5ilnEyN9lsWVDDFZqc5apXj0Uu/qNQzQFV9U5ZjOZPgoxgQXU
NvhHdUl4AKwjaMdc0nKt8ChVBpmYj9/S+9AOgHroeo0fOXszGWMKox7xow1k6FKkCxzuKtwlua8i
suh3yNNf+1Rd/AyvmpTMObf7cSS8Ya40oTuSDvQk3XnzMg8fw6yG+bbWWKN6OPcmZO7IehbPr2hj
RwC2fnoIN0iD3PSQ056UTw37xFOToeQQ+vK+Ew9LO9Bs9HLoeZ9vtoUOUibNfCqRq9+6mYlj0BPw
3hQEuCloopjtdpltzKj8iTN7TmtMC7bdPrV5P/8SQHMLeJUGnFvI0xWT+RfS4qvJZ84Ul5JemymL
sdfLPQVBX8A6yz6tIWbNU6bewR/rIDfKuYHonyML3cjr8BcCgqKlsZovosWmiNUzlDakwHpALdlj
VT8nxm5IfL80E0Qtk1dUTUAZHWACRn98IygWRSmWoE2Ux8K/tgNwIjjNEiPL1rsNx0PbMoOJ0rmr
rIhTzlgtCXiggv6j9UMSDiXOoxI6l4/g7pOGRrBm+y3FavIRdS20mrYUUwzuCOcYCy9gUGTe7j+o
0NuFu3sDquX/nVQQl8DsK7kAUl6RaV+XOZsnY8xCyF/RrN8qlziJct7KuyPdTyQMtZf5TWHIgFvq
hHsFx+XK2oqyxpzMYYamlwFRRil8kAlMiebMifms/Uz+7lhVM7Z7pPoIfkqsmvMrYm5dBEgMfVJd
LMVdWOYAeMeEujfQwEPYBfpzbKXE1ayZlXQlT9jAlFy/+edi1hsKyyOyDByi93XUAb/yyBwvKSo6
vyylH2dR7TlvAIFqaGq/Q0nNeZlKhhAxvwW3hd0xuY0hvVZoAeQinuqqB+j08XcK+T0BFCo6/3p9
rFer8hjjbPaNPtwY6FO6iXR7RYDy6bJZwWv4nmlQlUdLFhHWEvkSej1ymtcpL8KBqeb+LfCq4PEG
J23Xb5//6StWsYxbW85rhvBfdGFrJI/uARb2loOmkZP1n/750tyaTApXmFA//bn3sJFvYa1o1F4/
oJTFKLB/dGyCe+KV8pdWMexrdsowTHXfnphRpG3sPX4v0I9FRZXbVqn/hOMxwRSYffon2Sf7vmoH
h1r98Mhu6YROl9XoUY3nXXWhoV8HyM9OwQhofpSBd5/Fc1Qq8nSjh159Ny127mkOsDvoZJBmZIQK
wXHiQwt9+Yp9CHX4kucc2WoOiEyS8LT946mX2K8R4ZgO/U6KbHAKzKSg3xhBdk+aLPsorJ7xfXkZ
HmdrJWVAS1nC8yZt7ahue1aokGnywPC1YoqMwBXDIs7PnsFpZhFVWuhrKkXOwqb4MxtQO1dPR28T
KbS72qrF/BMYMUaZvQMHXSzxj8cXSbD6mKHkksqpgklXY3lbR1o8GICyCu78qrLss9TXmMHRhXpU
cdtCmqoJPTIPHrcyuYg3CZrsQTwDjnCwhAXkKbyOsDuPW2Kfc4Lnav8fWVPC3fRkZtB0NyTI3RXA
DO8iYdm2V6Wka5GR1RTgDJ4vKRYd5DTquDTa/WAqurmIyZY+vzpQU+giB1E4knpqDMUSp667HGKU
sYbY8sOOoE81EFA0+eZjewEUqknm/pLf38NZSfY861o4fMgTJVLw5zwk5Trf8IHBWIjeK/TXnXMr
5o4EqkVtfupk3mPwwpW7jCGQ0kgkIg3FVwemgiwMFeIw0Zv+6nWFfQlBX0wGVEGTsExgHP6vZ+zO
dUq98SXgbVhqrX3ixeZiKPNcNPeK7YOu9rPFH0Z8bumZSs0eS7dHt+dZ0w6vlGVgmcw/3TmfOAGw
2qchZ164zwplymbSVnUsry8D/kVyhiyN8J5HTExiKS/ekXK++u3ycfg67tZyuzlzWrKVnoBxswIy
io3pGH+qCsFoyZ0zE1HWPSHrXkDSFUVUpe9HblMafQdmRjM/cmbs2wtq5Tb5MH52wUbyx7Hqet6C
7PeZEN9AbPQCMPjdtsFH1bJknR/jhZFVvDey9VXOk69SBQQnTQ7Q3ogzdnxhKU7Q3pBn6iQCoKwZ
zD9Ix2Hgg95onT12ntNycA8gi303qlRcEdZPDn/FpeukWC+R35eQxhWP1EYfRCN6iRqGjl2QP1B5
bOyDoRTrK+yCG0oDb6+u1zOEmH9ptVH3MzNI9TP6AXpzzVZxH9BR8FPq6AI1NwGQuG1vwIXsKDVE
G8zxwqCwzcYYsxZeg9QZRgoK7cF8L57Bn5qDoJiEc9GJ4n6wzRJR7ycoZoAW+Mi6nAdOzGOQn3t6
p2fcNp6D20qdmYuKR2978XyE+aMQvX5/WN2zH7j3ega+T9W5AoAnCoPdNFZXLoAU8xWL+3wyX1HY
IfsASQ5bWgsw1XyPwcADclZLDPiBGOmCLZxqzEkXdrbcMWoGNSkfBuG03aqFP3Ix4cWY71xOxrAF
ATdm6hzfRglSSBqSRrR9RXE7OJHb5sa9LapPFEGdSXjIwRsX7PmAXvpi4AJMkGi8i6Ba/oAL3G2H
OSGWFF1U2KXkYRgDi5qp5yt7IBB1r99BurS+ajMzVCWoMyhKfuFlTXp6AxfCQuSZ3sD4yh9xQFZk
xcsrUR2TX3vVwfY4j0igTqSZmR6BRivehmHwzshKsl/biYaLrb3jXR3XRAuY59eKdlz+PietNXOK
xlcapk4+FClhmMJA2BFHgi+qn5x2/6LAX5Ld2TaqWG90FUjChTkOGfeu0xpouC+9JfuBR1c+u6QA
3AOQkAGHdpbEdXMKzfnILAFC2a0d/kBx+gUQ1hNStGvtpZimZkVWXw1MyZ8AjZyZy/gLYMSfGEpy
3M7pWyc4tJb4t2/fnPpR9HjLlqONty+2wMvH4pGFPrXutoldeXNXyd7ZqTgnJ3IOBDGa3EVlX8hq
KdIzDuMimTUFj3T5TyQPDI/bg5wxXx9cXcRx2bXxC4unw6PaC+4PFqLU23GRqlUvXiZ6aFpPYVIF
lq3/hmzMah3QFTFTChZ0sp/a/Nm+PxlOb/eBs//ZMI5rvTRqDoziMAT0ySNbUztuX9A/OHX9fNlr
tsdyaOfJn/+JdxvhygN0ThhZYnplppi0+X0ktv3W8refhN0Y9yVoLbpIkQ/xeNKTCJcttuwu5Oin
yB6QNjvZL9G3HjIZ04fS3SETAELCL0Rfpd6r1D0qzPASZYZjbGLBjoyjsCullZKlZa1DXa8gdEBg
pPnm3Pgyw0o+dDZETOEzsCG1GFD31oBwv9fe69XjDlRoCLKNvloWAJEvQLM5urrLsapYJqKyP9zc
dmczJt7vCC1x3JvSDlWXenQ+cJbR20HBhUljMHezhbMqmH7ZYxtNPvE2RpGHwYVkyKBp8DbWXD77
OX/KoyMRZP1DT5gt19POrIyUbWfOye5eA8AnRweTQs2zHIB+fe4b0x+L4NJ5gAffYgI07vxa5fpf
OpkTZSnx70bjX3CwKChD9j59ZfcYSHdAfcn/Jqyfao+rUPBdM1XEs9TBqN/ZgMo8GH2u1V8bKjRi
QlVIrALp74jJB5alQcV9q8Vj6A42E7CbcpeY72KG9E4CxT3NvoSnLrpiNBEnGpFT2PAl0/uZbdbb
WbsdtA7I1kttRaAIlpRDKVmTEwdKjFYB+nNTbBqDw7hmK1t6ZHgKQt78bI6WgvFe78vo4mBcG6H1
8We5LUrZkhx/DoN8dLZZo41k9oQOt77bo4jPjGq9dAhRgP3WE5ya4Ftb4l2D3VR/DuLOSTW/VD7B
sCfZyMQHYRqLcZpnbbRP8UPL/wL0weTqgGia91v+oQl+dki6fnJvx+4GvQMoj4D5aPyRMfzeVBml
lbfoPbfx2XHqKhPJ90hoh3F5D7HsnZc0Zwmp964lqkgcY5mkX2GaWPvvi0raEic4966yFREYC+i+
RTdFxWPbr1XRoDeto9JjyF4IUDcVsgYWX6jnnQzX+SOFy0J2RQPDznTz7oiAW9EEUgRLGoKMrce1
nmGJnLi7r2eKvPnMD6S3SKTEJbr2frlRTcXI0pkcFqNGd4dmy6lTn2Ef2gpAml0x4qzF9nCKN8f+
BI8OPbDGTVin0d37N+RULLMCNOwvVcdliYBYk0zlJ+8rARs8TD3+5/SpRjCktgqsrPdf3B1G+CrE
ctIr0EDPacodlfjxFmsTt8unyf8BeYuSWlCTigZ+5ZrLg3ZMKQB2Vz69za/xzp/0QgYUdtXkFvVa
Glt/mi+VQTCGLSxl3AugE2k/vfbEoRw27qiT3ugGdnl6cJQsy3QoSFTLeY++Fx3A9kt3UrJS8UXz
AkPQZxrv/ixqYrw5DA10x8N1XHgGpxl/K3GftGxWJgZrkFSmy80mIIfiXS1msMxhnqbGtSL+EHxV
UJFJTdg4G14fDTVCZOZu3iOsKUMyQ9sgqgfUVz5hJXnwz+jAKHIPkgN3D5qRFZhqXDrNjamekLCF
eZwNuDGKbYlw1SmQ8ngIwiGwwBG8oJfORH0vFC7sdnGRb1WYbbJzimWYjsAL5m9cOEkyh9Aud9Z9
JAvdhs30Vsc100qvJNt74AM3xR4wdUtgAS+jENuPw3GEJjhR+XgH51nKOKebCTm/odC+F55xVKrG
tnC6H8nwIDE4YTf/k4IyH4+sKkA2Z1zVetj89d/oc2ewmT5Xi28smwps+4JwENzuW7t/fqn56xuE
yi01Vatgq6xoWbaGgyjjdxnz9ey0TlrKVtH7SrcjyTVzTUQNsO7GN27kjvcHWXYluy6h8HGflyeT
yMrMVktXujh+kvOrTlNtxp1UmLnNZeUSqgDCKOkwZfwQgb/TK55oOOvpfYG0e9sfnEc1F4QSL4tv
sTuY/vQAFV1s3TxIgWUfOvZUwjcLpi3/TypUxlZum8ZO5nxzPixG9Sxc60TPvf5H70AMkzPdetvT
rY3+kG+bvBArjJdtd1NxHORR2mj/WcOLVLMRZInhgXz7pOqYvucTdjRpL85Zw7aqjQoir2ouVO60
pqdO61eSirkGvptPVoB2NhgCuLeL/KVtGIBR7hSJ/bTC5gUaagsa9aCR5w+wjZuVYIP+17oKBD0i
RrLOwrB+rMtmFa5U4hqxoYX//sPnrKTBFVg77y0H0rUyl494PiDley2EvrlYyNKWsBo7UfCeyzC7
csYX7o2LdXIrSO8goDAKehuotOuSEeNEuPidCJ4fGsbl/96FG1buIPwGxVQk4thTb58XQZV5k+5g
fDBg+Nb9aQejySj8C8L89HoDhKlUD7PCRWuvH1AvV3kWuSpnAbAcLvT0Z7oI8dP8TM/9mJzw8g1Q
LUz3VDhYhKyjo1vzOs541PAZP96BIvx8suS4jJJJ44fPu8ubS+VoZGOvGz0YuWupWbkGWqMEF0ej
ZHlWQAmxqtKyJp0qYZY4lsjA367O05ps89RQK1sVap+8YkHyxzYPxgY0e0YFSPZQZ1rPtJkXMuUn
vaQ/8dGqaMnXme/kZN7OdTQicje04yPed32KoMy4d85sXdsnZnA1R+1A7bHOGpMVQYZDIlrKIMhX
bYRfjwP47cN7hv7WgaiC/c/WOYNy25wHnhJGRkHRHc196s/fruECrU9SytrRXKb1KDlPbsMlELcS
9oFR4eFCrG0SZEOUOMB+BAuKfVEmyy78Uma41iSPSLZiSep49wv0wphed3GSqySQJ1UK7BqLcnXT
ZCL4eeOoNY4sqhmMgmrRZu51S03IGop9jV6BymV6S0o7CQjZt64QOvcIePGlAWi3bAzsLTUWaRll
MHot20Q4ZrY2SG7uifGdzxa6JHohdzzXkrke6b4KsUzJrHYGEQU5RrCQ7SKzaVBW99GhE1sdaoDQ
1kCpnTuYoHztfZPZ8wQKtuxZhoig5kIPqX/41k69MO3W0ITK0afcOz8I/FcpbF0DDBUvL8xUuGxJ
EGp/idXJppT1hRR+QMOV0MtAVD+lFvAUPba9gWLPvn8H+0MKGh4NQYFd+Qn86gr62sHn/f7gOysh
9tUwCw7gj/6Tskd66nj0WKnvqztmWW7ImuxBvrjcfZN68gcu74iNEHj2dWgh1j4cZuwh3YKClLJm
o5NcuYLFLCyhFMRhJLTU7c2iXBQmoR+8t8xEhqakO3OGjjSe0zCusEgnFts6SC1QUUg4ZgW0cp3l
erOvcTrr6WkkTWD2x2A4BBkZXu4Q+zoGQEw367Oo0Gfv+M7r9fJiUfcJKJcDrcTL4QR4g1K3gif9
5bo1gvvOd4uHiaNqXKrMpf9CocBnMEsklLZyzjiE5q6etmcWgvrXbFnX/cup4VIaqUIfHdWnIlCL
MAkmHXv8Y6OU95qbe0urdlTZtSQJcl2i+/s9kiiyiVW5pbPVSbqdYqGCyaDAsxICvCqwYm51CJrV
8TfVpKKnA1hOzt8S7+RndfYjeJ6qatiVUibRwV/BZFuL0b6DsTGHcopIT93B/qdaxWcwTqBcGdaD
1x0FQKQGZ/ySpSS2tGytzGSeoBL44KMt64Zabhk2XYd3tqDICgh0/sxCGl5s84dtsyzMD3dsK1qa
JQjFraR7Mj1KdBzFKGZVFOlT2CUpEmp49RinXlCStvecScA77rmBLG82ITDmIYXoqdFSiMNS/cvE
FLwXKocE3amlqIqLr1rE+0HLIFM8gEZIfdppH/7pQU9fXBkxt8ENHeffu4yx3FzXTRWNd1GhxdEJ
/JnYc79DErvz+L9jL/lgaDj3fgg4il0hrijhdmTHsSMu72jd9W0r0qk59SfZXM2oiryJjFOWz0G+
XcBRmmCYiXfw3t3hAUtgW0lhOwIeWADwczWuVr4+3clr6RjcQ0DdbSn5JMS6g5tyDyB2B7l0Jfqd
tPkALiFCW+drdGjpv07zZPa8K03vGdbIquj8VrplB+24qYyfIxb6yDayDP7Dv7w4squE/PY726dq
3bTLknOVueHVHBdMhzdQbMVB3QQP8rmgCRR+uMss2lNSD2X5YMnVcqaH6clVPlYjA2o08ijwgzMq
NC9UVBrK7u2U4yuPse6jitbq9AKWL6RRI2mCnnN0Xq+gTsU5PHujObQq53PofM98Y5IwKIzeUQp4
+5mWehfiRG4X5vYXczN8T+1IkV//loGnDZd5wQc24wtGcJWx3jQ8S3hetj24sTlI3f37UkSJxXiq
LE2+4obL3KIzIBoaZ/CSDhiNnMP3jS20wJPEz/i3FnnvAcW09PoI0aeEOPnJcUioHLVkYp0s+b1A
gAjDWySy+YQvKvrseR9HZkigpK/xDCqmBX57wpMlVNeKji8+a9RS7+7DLhDeBaRBQ+wZpZDRxwPO
i0+s2ZgTPnOoSj2X3HKHABKZSZ50KOZD/q8y14xSbl4r92UfRsCk0vcaQuNVulYFAwu5Z4hsgequ
ZPoS2YdscU7/bZFZeykb2Zi4PelxQMquH9AT0dJdhMl5ZODXfwA9OZP0pCHHeSvsPlVwHffRDgwS
HH8OZxBAnjn+J+hfcCj4OdF/MetlmvFJ+gNaCZRzTjSFEpaQmMUkaX5hlnVLav4OxGt41gzSryKk
w58cU/I53RVtNiG0GGMBzyaf30dqkTbYYU4Zg5VgtAvy7XupDjOxEl2fV+YMKrElcepAiSL+p8Gu
oLzCdHvARqL30b5rHzJuSmW4nplHYyfBsPm3GB/9vJ9Y8S6qWHTkDOt87JPqE2wFQ31JxaygRRbD
1O7vaaUQmpHw39Eh8K9W8ktC0DsSnTYy3UkKkDCddb4VUQfWtb8CqSqzAJjOmdAqr4tQPcpumD8H
VF0tkJDNruPPk8Hq493itXsoEpezCHZUKzyLSWjxUY3gJNinfO337T1nRvofRsE3/BBMHdulKY2s
y+ld3DYcMspSDNBdVIepC0g3LXQ8uaP3jmgbEBjgQCYKqN/JuXzvgM8NNWaFW7EXCH7dfTqjPGhV
iRIbNiTE+x4NtMm6GVCfR97OHkXm/wLUPNRCD9gJVnpMKcoCRRETSocFliYdzdYX+GFhddVijGzR
qT7PnNTjlKw4ieU8IwpVBhgOJx+zVLnEJWMylHcFyETyb6WR2qKOrwpSIHpauUvMqCr92Ar2A7Hu
XFcBB6HhZsNJjY2L/cig0/PXasxeTPVUyCYg73rJgP/dWqCRFzIHlSxaYTuYBlTVGfNQDvU/asD0
kuMI9trUs73KtG2NyuPssFdWuyPFqNIhQCH9Ao2fD3/1AD6uEKBFPr/PGr3ol+ZXa9FpmqgCkCAK
C8+1XFCWaK387fWa+cLnyhR+vqAle6nIa3sSbK9kYJjdLOfIpYWiSgYmLq2mDBcOztRZKg9eJgyc
EE+gCNX7VAFRzV2kTcAyDoFQlfH54d5IEnNSKq6kxgcL6kmTMBMAPPyc6VnOsfN/n23NQSgDQ16P
UkrQrmG1NtSuOkwm7B/lecr6ThVXi32UmVCqjWPk4h9/oNrTCqxv4YL1gU5tGUMVhn1QQt581L8d
NyjHkOYaU+KcCkA1lC5snRRrr23dAQPI7SDs5eQOgVu6RFiQDxCgNCAfAZDThdqJmT9aum0lYQGH
7jnOn+GjdD6SO+elcWQ4BXpFkwwHYY2H580N9lKD9BdmIsnOtZPuDc7gZ95bOCTPTRFYBGjh5Qti
ZicJcxI14CI1XVWDQUWxcVYmioj97QxX0Ob1sJMw27cuO9gDoZV46XBzpLL/NH/02ZzuloJvOLqQ
gkezBrjcyO1v+D3yZUy1LUtAOdk08DpfdAK7882OymhL8FV3uQBQ+cYxYBqJ6ZPb2zJ9ZPEAQu6g
OFqq7/gGyuoN86bnCmZ72Bd3x3R0vz7Ab8gvUVOqygTGwnoc0k4OV8v+MwRR8q9HemW1cNM6Qp71
tBPIZbZu2/5ny6daNvleV9VirUKt4y+EjM1mm15DWBul+FW4F8gpZkxLpYPiVyxjZHyNG4OYtmoT
CWiS/kr/X4dJ16dq6uYBF+U0ZeUlC7rzWPkRMS9IuAyzp0LxCMtiHCbFpySPqwrKzXxewLvOvFMt
EdNEVR2zoOYtQq0bC5QdwMaXO5seBa3RwXXjBS3v2PVRIAhOkN2Qjzvu/x4mqOUE0PV6eqwaI8FX
Evleu2tJ5oRrd7KF6sYy7YrAB/8szkX6PtwIg4BhZyD/0afN48IiBuKFnI6PoozZ0s2msF9aZSW8
CFItviHy8oucK7J/xPSMl1vAfgqQGQZqUMLgYeWUmZ7CovyvNNfAb2y9WjMVfwrcrgiaJ/3GR0/O
cROi2ovmxAWI8dMlfxCJmfC6INUSEXyNtPnd7zVlpw+dEIjwzwXu+ehmzUKQIhBMoAerSWyixca+
ZUv/XYY2RluPcHKVeumqqbrAhDSmER3B4oFLVBtgchZSpY5MQo7sIY938CE1Ydn7lJbP0JnN1aaK
ruWUHdkDktFSnjrhXs6lWjO0pf1EGmwZloxNdD5ISZKiqya9G+ixyc75HXVltMFtt5Kssmzez/QP
Tu2+03BOtMK9TyDrxAew78K3x7PXiDJAAT6Gdk2rHTH+DKurHgQJtISEdMr5HqbhOw8IOzR7XQSh
fKeEd/qs18TBP+Av8MFtE8L8JTQNowm4JmFU7QayDTXS0nRIkdfIJ2hKmo7+WDkpRXj0yv3/fuSS
1S7Qweq2rH9PNyEX/hwbjkp40FZ9SqxtCNG6xbbkwW9V7A82wOBguw7P14uroJK7z5OwtNcsCToD
QTUew2QsXQAmlbA/eSm8/bwBr0ybmj9iSs5RXvmo14DxPk2QkEtyNtmiqonjaDAXVym79m195Lag
WNM4+cJ6vKpi2b3rEG8ScjO6e8furmeZU5Yly1DmsHDIrYy7/lqOfHWj6HZB6wEat84V7DVFul6n
pS42joUlTzDdTzJ6WS7o2TeGNz7BNDzGqfUq+zD7mh+bGN7jNmdCtg4qAyqxdv9FwbtQJTOZIGSx
xJJQhIu+M7k9A+If3GPX+yJdkzMxEBvLZyttjfkZHptN80RFlqHEII/XACzP532cT/XrQcjbDM48
32W+mWyH2efrU4u2gWzYygkUMNTxqNWszGRE7JG/t6hCfIxBqsjpiXN3Qe5+WtWT1y3ABlotn1U1
Dxcxu+4sBsWbVE4U0qdQ4s4judP/wGJAB+9YNBei8sOi6R97IFZi61GhNDU6lojiiC9J92CmtBxs
yHkXKqItO/JLcZ5TTFXI4N88IEFhRHbhgXXvL/zH9aTJWPambggzgm2LzG/2BsN/gR+nfNInLOXH
0Sj5gx4lMSHBOnXIkg2NBRX+pH2bithG3H2+oBYY5tJOAEUkzse3ot3sud71UrJ9wERRjcRTZPVT
90z4fzpmfYVgIvY+J0z3nDIk8AqExxfKLPKoSjgB1Qc2xy45cUeh9TsTpN++3lY/gnex/O09DHxZ
4p0RrxasLkEyRNmWwiBIk4R2yj73RyjhcGCHyL40pjiKLEDyWgekkQhgBqmb8BZBT2U2rPsnKyKu
aWotDr/hQ5QHA0ttbBbPBtwlugrk4aKu2EhujyRMCohgf1aJTaKNgNrtLL4v4ZPWZI5ARnPjbPOS
mwEQsHHWZJol1LjFGphHyU1JJetWYpHrp/DnjZ6Qesfp5AMGhiLUppLHnzFwySeOKHCiTXBbz8I5
gRndenbcuBXGKdmwlGwQS3H+Q2rFzz3MkL3ujELjzEyRCR0Vv6jhUzlBicmCR+7U9blSP/BVvqJx
2lrbg3H0zcIkcy9nsiTGK1dS4f564a/Gm5i8lkQE8ERshQpiahEkwIsjW7NV0rQlsEnRzF97TqNC
2RMaP8t000yls1XLVfc1iMjtuNxNWooGBCElPjeLKUfXBuuBloa4CyXIDkaKt6jl/9yl6Rhgt9nR
P5kkmN3oUsASsu+Y9cxH8kTBSILPWuXaAmIBEXClrBZtjN5hXrJzeiNHy8BnRrLFU7S/2HKQbThx
3KSCQ+i1m1rpmUGQbU66iA2k+K09m29m0uLDgven8yEH522yF+ZjtnEpRueoBpK+0KhfZhfIfw6V
cvGI4w1dvGr75HHB9CQvsl9mKrnM2vbeHPz5GwQPv/j4TXYLVnuq4kB2tuae7JofZ+OA5j1kEmB2
As6GT9IabCbLywAP1Rhxg0IWxud7v+prLNOrnthjHRg01fwaYdZd1sJosvwEyYylu5bIUyBlmMC+
3XDvDxVQ5IcoRNvyoQmoxCv18z7ZJU05/sQxRnYaLXyAHw8C63u1kpMqPKsaac/iUCq7rAm2WPi2
1ZmZfZP7PnFqJNfMC2en8oqqeIGVhwPoq2apab18JnlwC3nBWPhygds/+IXgwHsaiuLQD3aJUl6e
fqTWtZUf8KG9VVapP/S+IjvyqUfVaRi6eV7RyjGh5+NqbwyIJq6zvJL8HwCa2m96nSSte0bGtXPF
x7Qi5lJzhHjG/c2pHa/Uv29DadIlZkrMdZ49Rp3Cdt5kRNKSZSGm+ZZ4LUBLUk7aqBESmtOYgGL9
9bMX97k7fwFfe4e3DW+Wmg+Awk4Se7UlFlaINLD8B0eUo9ds8R//9pOoD1zticGtmKkPzLEEVrtG
IUtIeY8yujnzIKtxPfEeS+HUOmCdhBJAzryuD7F8UwmzPygbPI7KHBqpPYXIlR6Q+a+rNvIFul+x
9aMeOnb5pGVFpxM87MjZwJr1TDJY/7M4qnQL6GOatCO4IgF/V76UK2gwiMLgOXJCNgWHCkDwslLA
uWAwVIiX191OrCUo5a3kyOTOLazHzc4a+KRdotEM/i2GGIr5pnGptJ/NgOhMeMvErs0WtL9MwXTH
0ZNdzi30hhL6A0Gx/gsw60yjVEtxg6O5OH2vAs6vMz7dCXBM8cxJeQM5IEYqrIGjSz3dR+yJvvqw
vBpOvqX4ooLhgvDj+gx9q/kZiy6dX1mxjLduaO2a1VJ1CdpBryyugdnwBviZibrGB72uDeYM2qFW
Wjap4XZ4jgDjTUWc4KXgVz2cn1c7tnwwRpgt4zNRagXOUYzMjXJ0KGwc1pwzr+FlBZaXR6I6gnTe
0LS6fYN6qIYeR7EJSzv5nboeiYwwjMcxN/uvqZd2MshPM0Yz3ibSikJShKYJO/NZbpk2mWBsXOoW
1x7+VwWgSxzWAzIjtt7DYQMHSkg3HZ/2TcYSckvS0Dz+/G2Z6XmHw9If2C+jtqxnoytiUFS5ntOq
DK+qGpD/pYhteTeZM3DloP+oZRXM1KTtLa2L9GlbX+SdlG6b08/T3IfZx1XhwN0mXrcrN8rtbY2p
pOchBNWyRYJlwtnY685b3lEHMvEEuvM+ftIEUs9UFRizsySM3dWqCbt0NLkgXb/voKwv3KEwhn6S
fMo4yq6I5ZCNJcbRtZkSSrdw+kRdgRSy2zpS8XYl8fJSgJXQ2BdS8Ql2vBMyGfTP7IPWp2ZRC5H6
knxjlueTRiVyTCQz3YlDCCLeUxD1aN6eoTf95O/gbun5YsaOoMVVMwy2yGCBS6KMqruEUMY0dIx8
N0c6s3JUtDLwSbeUgLRJMv6uA/lL6vRHBI7WD0kBU4Z7FV7aFl9b8j8lL/AfdeowGn8FRVRQLtiR
5eJqf/qSQ4eQXheRoY3HiApUp+L27OFULX3iHEpz/lOYuCwJMngLGJOKzhwAnmTohpQRomaDDEXE
GtYR05+SzwvDaacHRciPgTHIhL+3LWMdA8cYtXjUjKkQTBHW3eV6kOgtp7xP5NCdUB6uzMKzJeFT
zbJFtZQnL3Cq2zkHu8JELQVKl5SFq/zqfPOk39tetZjmcpJnBuKIHHPvjb/g8nPL5Mt0SaqJzWvD
z7Zpz+goSFl/+HEhMQeRHAsbpUVjKc1Mt/s24dMk2GW8z0xbIm58Uw4dxh5XoJFQ1IhC9ekZCvWB
jZCZqfXmu+bQ/0Q1C5YhubOgMqV/XMc/D8knl8fqWVurDr9qfwwAxi68xF6MjAU1J8I43Izwa3js
jcx3LsXRm/bxQAXGty8t+KG+rOHV/ZR/iOv+B3/DwmNuCHwLknItcracnOn27lMZR1pB+yEbpN+5
kzQn0XOZEsrPHeJUdqN1Hac2xwoPo2cmAZy0JkT4qZQX7BAMkhylBfECDmrDRlTk5NPOp76HVJh7
OBVF0LfKGdoENjnaWthUTpIqc2z6DncHAjhvB6BxfC2h5SSGdl0WZNYNv3S4sDyBPVEJf1/xw14v
3AtIx6JJ72a+99rF/Y/eUEvnKGOfbT5rBpq2qSwEnjP4Bccp2aFm8Ef82R2np67tWEUYeHvo/dja
+f0Dsd8tyzsMGCn+Zs4n7G5bbosufDXSCU5LcjTcuAdKTWevgzUVHnq5SanlfaHpIJE9Az+cpqUo
wjC4qAZOMqR+q7OjYbCJo2itNSpB2QavpJAyGr8n54cZrqR6lPEyWuOXCVfGNfJIygXRXwwS7jPX
0psKOIAUoDq/jIVOLZhZ/murlwIhwvGUcidl39d1hOLdO04bv/RFnfJdBznIUm3gBSYNfKMtI3T0
eqKjQSjsHB1LGRFf1ywUUPMREjUEbUtdjw9vsnhzI5YDgLz1FF2ve4SY1BzqDGzANdwpJQsVNVVj
Wk7vvR0zilKhrhiSOs1fgbJnRnFdjOcxiqIHlhLRMnWXXof1FSh2QiSIUBgjSOrlb8cMVBEciXEZ
5X3OzamGdxNVDc7cs2kJHC76qlwD9T7xRheBTCSyXTsys2et8l9xcFCxvtmzamBYe5+haarP6M5w
jxqYq8jKVHta8iSfqeh7A1fPkkn6tIZwcp/6U4RUnMEwT7DqOTKUGRiaKLt+KjMPGRHcxUJY7x3l
OjYgynaGg3KNo4XsQ+KRU1MzNWg+mMIvLfJvOV0iHIb6QmzSdXe2sZk+5Fbz37S/MjIGsZEPK57f
uCtL0z8kzFJlgTZXvdtlmzc5i/MDqwvGIBrulNZPW4nlQdfQ/e7rzCBEBiNSIKL9Wi/omtwa6ppb
TJKDKM/N1GM8RmwHQLajKRv4PMQNjMG6d2ulpmP9HlKvbTaaTEQZWgMR0EaNxLetAJCMox0ROaHi
nvlHAuh2Vg/0IdCK6pM65nSQgq6z0ATS0BMsDabLqSv9SDSzr+3sATePZRelb8NcMKujxN/4Ghfl
SQH1QtPW5FaAnFQ5SkjtC5QyqKcOrIcMQrC9ooemBVwF3+GZlLs64lVzop5KYCqcZz02XPBhrtCb
iclFzIEYZ3+OnUf53SVqDPTVIW2Iq6V0e1W1c4LeaqMxX4hopoNZRQmS5n5pr97X68I6+ovfgmhv
QEe7lDF+GzezdeJtQLXooeRkp/3ff3+q/kXhR82FJ4+s+5oLrFiH55F4J9gzvuLrh3CE3RF58Gxk
tYy3bBqxSstvuIX5B8OHl0qHX3MauS2ecNw+e6h8TjTNStDRJvg3/VDbuR5OEzcB4j4nc8h8JcBI
z1A8jeK/x76UbiTwTpTvfR5EyJXFpkYXP/LmwDLpSCaPG5aLqsLxc8011Cxk3DIZFERv4spBGI/g
95QG7yXK2nUf1zIQ6uCH6v7g9vDktkCpAk5uzdkMqq6/z5j7Cc/n1VeZJuP+HYRm2V1i4O0Epwcy
WJR6gkzua9WGJOOKUeMWQePpfnFRZGpvaRNz9fC5rvX8o54URSv0eU5iua3iJAkXzeflywSX02T5
9eCRHJ0oLR1llso+tgJM9mWQBBMizn9M6GOWFIQZOkIrh3BG62r2jlAhe358nO+iPAQtGUiav0M/
aIHGTCh03Tn3MuDgAujeTncqdJgkKcpscG3aCkGqgavrWnuyXD50oEMGyyGA2fpVuPKoq3hdEpU+
QDOnK57o1vhdM/MXd5+HYJBgedeiVgMxH7CU+j87K5hF79J+bQnAcxNrLmu3TLR+YkgxNey3e2aV
dmkcOb1gNjxJE03vqlnWIPmwwxwmjUKiqnWaRmc7+/7uvMc67f0IXnIanErr6TGNWqo2TxqDZoec
MfmfmoN4fYK6JDyDhKEQEZZ1yK/TbP0e91QLNBcXDKzWd90eUkQxqGr3liKlpNuQj/f4Ou106sfE
RQ6AyS6GsZp3wi2Qb+HnuXEThLkMw4zFG3zKvI8fmcQ9kq+3IkGS+KdwBvx0o7P8PVCexwwCjTn2
4p9f6HMKIeiFjOD5cSQzEBQ59+4ep5pmTetILbaFxN+TmRyVhzc3RzYRSDFegRWicDtVgWLwGkjG
34IKtpWOUSSTGEFO19bZCdBzTA2NG+/UcYgZrru2cgv+rGbSujGsV2eXPrGoH9szYWpt3x3dIhG7
/ll013TU+cB0QSz7IW8T1VYGXNtzL2TDLzrDkOnRczYfJFAbUEJHBTPJcoxFMOQKtq7dVu12zFLV
qab7E6CblICF9M2pE1YtPdKjFNHnY/pC0WkegGQfY5wYsq/Azy5zaBmTQLvy4glR/bQAjdM9nfku
nPb9pFHiDyjXnnaqBfRe3ALgHSlmLnr2zUcUsViAMovfLWInjdJZhQQnhvyinCLDCKPKg6YWuw/g
wGkUzUPzT1LEQ66zdw8ozhUZ+a+I3gx7o+uDNEhe/n9mH//6EKr+vqOOdTkAdeZ+cG+GLwauUY7i
lSX7PoKmit5E59+YKjDOm3pIUuioccl9dcNxsnnrcJk0WtJ/FoKI9C8+ZP2UMPTw/dFa2YT7rMVZ
TnoyuDShY7omh0eZQTTXMxgTcjMOlzj0WZCmQwENI0Q862tJ1mN1A/cY7GzouA9/Nd3RdSeLVQwF
ej7QutahPyP2nx5fE4Rc6B+uynEdiYTQHLAlRPrlLxfvR+1BpPbZJ0colUG18RjguECcSF/hBMNq
Kc297mWxD/UdNWaSA0qu0OcWPBbp2AbDd64X2nnHDDTSfEUhPTPE3cdQVtdjsh3QOJs3pnAWnjBS
w8+h+/qN+ZXKaijZgi9dtL2hnCoUHTqGi1S2Bsg2AD3OzZOTLXgYOvKBWTyoxu9QrEiA28uQBS1R
hliKBxkL5EGuj6MTCXOg/khoSXQcIjAnutGl2cVWKarC1+uxtZLf59Tq/4Idr/ySTYowXnnXRk0F
bxd9TXQVZ5iIfoDnCaVXVX9yAyPgzs73sq1O3Zy1AEMWVRW9tmBhUmljqDZwjFeafovXPZUCtEuZ
EOmpjwlhFeAFwrwf47Tke6Qe/MD2YCU180r9tuxYEtuxcC9p/bkVzaGJeZacIFuRQW1Z0VRLEM0I
Rz7Uu0W6AQYTDWnEBSP/ypBYdf14H1sqfj8EdbcHAJDYLmvK6Xdq3l36KsvdXSiFWDJbR4cXTd19
jhzItBT8nJClWgZo9cJ7KIVlW3RSXoblOTHx6aMAWzLg6jZXnd6osbfWmVWUBfMkuRvYVwfHVhn6
K+EBySrnD1F0hSNbdsHgJEVtFRJvFhwmbXDnWFfCfnQCCGKQWkJ8qwVpnq/acNRpTgNtLF56PEm+
mwBtK5VzsSimAOoXZr9qVkGyB+Dzi2zbCnv5emdqlp7dpIuaKgoxJZPObiRY6Ee0aCP9MapjyFD0
VaOJ2F9x1n+rQERvJtBPrYXC7EDRegd+7Z9WwQMks4MijfrfoT0gzUfR3GqOT246ig2fTsJQ93/7
sfd8lFzL0noVGSSVuV6+hbceU/Kahlqw0pHq0n6SzHsofuueJFixKXMdq6eQfqxk43Em2PTam7y5
60o0ZpC6mDHtmnaHWPt842a8/JMYKUWF4b0ScRCaum5dmBcwKAZGSWFR2Ix1zHD6GC6HGXGM95s6
Vg9zbPC0SJhzlOIFkoUiLLvlm0K/i0z2ZMmLmtE7AchKsEZQoGHJUIS+mTwktyNkMTLNRbK4d2ZO
PVjhuY1EdMJtFrtfjGEyiKelZIX+hk/n8h4aOGqHvaWI5henp5OOYfdbjBeec3fzTfP5XDlDwgA1
kU+trNudO1Ngea9vHq+Sgt5tVtad+voLmw+rt6nsqVS2y8sG5B3aU37dgfE7fykT+MQ4bX87iYfD
d3I41dOVTOkvvOilyePUhxfcwSJWEukBljaQJbxKWp299rXsu9zUJPAWlqp6LYWJipYmcg5a8e9E
BBMgM6Hg6GOPH3w5VpAlz9+lIxF+dqBqvoWEbVQPRaHMTyUgiNMcM1ZTWJu2AQ4n8+wbAtomy+ct
xMBGcB4Gb5cvhX5CKm8JnwAXnwBEP1EoTTIMkdqmpi44E9VVy5ECbXdGY9BktkwVoHQuLFF06OS+
eq41SaGDtogmzXF+CVVQ4kB9bBXIKi4mJvb85p8NGDQpwBsCDWTV00bISfCPowSkm/E+l6Gq+XHk
TU0Y419ZCWxlnfjUTDbsWf+fh0mX3k9C2FRgJsH4J8KfpqQOoRNlJML+hBR5+ZK0bsubu4GZPMJw
y8qUK6uk1c0WByqeCODkTo2YimocOAIFITfsCBAtzL8FY1wOcZN1r/38z1MA5y7ISaqlOLBPWbsr
FkbFOOwm8sTSvUoy9p5Bqtdynq1V/8Qla4Wh6AdYVEGowqb9/7E8194BBw9aQqyFrORikyMy5m3t
j6ueyqYHhEwzxQsDWDSuPm0nmMMqIzK+bmSQt9Gcx9xTFKptqQeHJ/9VZQESjVYBFF7dg2eESAB5
9TxkIA2HYTaKbxwEIFwhNSuF7o+toGuuPIuBnZdqxBMLiyxBt3ABrqEk9eWT6CNxIJ2ABd2XYcOg
FDqsXFY72P8buzFgJcaiasu03vudebyFt/AqZ+3o7KqMglJNkF3Rhadq8BQj53w5IVXo5Apiqlg9
M9ZZpPp5A0+Zxe+C76yIOQCUhdRZKmSVNtRPotMU1fBoXAaaESeQ/sspxvrDiDWelixM9kww3nIU
UgBMIpzGShh5wzf+TpLq4dN7wKZY8DaxOtLcQLUMGFh73kHbuuPtfVP71IQZA5qZZ5sahB0MhAv5
mOooDei21LM0P8CMfLWbenDzYnVso4iuXSUhi4FSi5sBK6Peq5bXVM8kdSQ1JYgI/8eFIo8TfMTN
CQfqrEaa0zDPiIJM4ACM67aVr5+ByBK9zvNbWNYsVouye9ufzZ7+A1JF+E71f0xD74cSSrFPnMNi
qRSyL8VmaUerh1uyV5mY1E4QMirTLP9Ym/4VJdZG1gOgujaAw53vweg+EgGzroeDLMbBtRv8FHAk
0GJdXQAhm91xycE+Q6G8O0r4NWPr8N/PqSr34zdwHk3iZKS6nds57d/B5J+7wbnfSfbLNYsnSbS7
w/6XTQ+kpM0Ma09ieKjSWI222iBwo90OPqmO8S4YMqYAyYQOQcY3PCJZx1s2v0GID7OGgGTnNqDT
1KFECOw0c/YMYrY+rg7lVWVch2vA0vJ+1/wj8eEQFOxNcxzj8Fg0KBP8d4qJKfc/PGX2TSfF14F5
5ErJyvdw/oL2ihOl01TJ4xI5uypl/P0A5QtuPD5c72fOhwyipxXC7m3BrnqHPbsQG5KSGctgmf0P
oGDL/FM4ANZS1XZ84E+23j4qaHFgO/xq40diNVscOb9jniehMH9Q13NbWsQZCx1Qbqk07YFuYnHX
Q9AqymP+6RUep/ePB8uO9t0iKIUncZ7qL7JjHgc6CYDFEI1Vz09EvcJD4UgNHcwpRM7/+a3LI/Xo
bbkfFS9GCbAOVww0NyAppWce2V8PviIxTDPmEbJepuFULbJODis2Ca21ggNxpC02TtTU9xhsPL7Q
+aEtVvSqtqyJoRq7RjuK118KZWZ0pC6wOnWg/99/hNo1KJ0S34W9AvO5X5ChvNu4nSTENOUHGfpv
MuhiVb9rfEtqdjvK/fmOZ85Zag18UQ1J/nWpesmkywaMGop+dVDiafgP2SS+u9vMpPF6iAxU+jUL
otHMU+SY5/HPsOU+uZXpC0C7Alu1DMmi4tXrRTC/PsT/A3u1XRVLdjoQAMS/n9MRFo8jcSOLutd2
sZHHoQ20ZMnyH6Ar3tcKGCWxqgLqHcnkTP+d/4jGorz7jhMH1ALkhWJ8A50m2JVLX+9wOYJs6GJP
FLVpt8WDYbchmplk0nmQhpl5Yp+yBpf7Qu6NaslQAAp7UwepfZzoiYsgH/5VY4zO5bT6mKmdoG0B
YW8jwNp74WhT40Do075y1rykENbYNahA4bt01J4gjT5dkl68Fzc2T67oe7LlUAltP1MWS1Y37KGp
yDQcGRLZEBZhdsT9NO1NFLWD4HrDBZnZRW9culg7ARmHRk94pVnaJFeqzUKtsWLqhWCYiu3B1hrv
az3AP28CmVT2CGX8JkpZN9UdHLX3uyJ8R+cQ/NS1e9C/7YIeA3NNU+Z+EAEzAxrVFobqmqx2xxdt
YxmoMWUvW83h92HGl0mm/PYj6n7mUlRgsgsRqMDHKhCvwm832squD3/gQ2TBn9XjC7r59ix5S5eb
9gHIfE1jIaic3pZ5lkMDjyZBdQt2QuXUU+w6sIprEmT+ICoMcc44RWeJIvHnGbTYJ9oZ21ZvMVvv
Bc4N2gc89UseoHLl0EYH8rGV6PB93+vxxTEFqTZT1AMvg3hUWP838LbkynWO0MJPF/60OyBbo/vn
SdVXOwv8+kjoFn6DoTyfiQI11iknfPbPxxKW8kREBkV6Qkcb7yV0sPeV+ZU3z5iiZk5pen0ttZXT
QCr30t8SNXt0bx77A4ZdlFkPVF4/6MMP8gXXBH7b87k7cHfQY3vKBGsfRN0gK2k4amfFGD+1MUZd
JIx5HjWk/3ZLWweMpYB/ZsYKe/mCcMIlfQT+CbWiHij2trr5XQsQqwSDODgadcWrpqRajLfO1Vzo
zwHF1X1XJB4nYs4npdmc/xNfHWfAVkKQfr7MNeHTwL6smFM0aJOLkOfCyVs+uqp5V7WouGXytMsJ
3qRYRI8bfsBc9drzwugXR/BUFDdqybhxqdIXbKH1hF8Xo0q0X2OR7cqVV7boCFKb0R24hZy7NQF+
DC9dQjPzjgkioz60/fGmVB0l9PSoRNnyDBAgTZawpAxKka0Rq1hKwFJ1kv47bxLKJNWgR+8QuJ3W
TLQM569UKLeOvAW4+VEvVkEEnvad63PpUWwzJNRwGmfeDKCS/MO/gzUy8h6xpEjZ1tlTD30fjrO/
zedvzaWWv7Qsk6ZNnKPseagFFt/ihP5lktyzKMCpANa+dPXDcs7TlHsqDDOWYFn58OjBOQPf75Jq
55qepkSiJqAjy/fvVP3Pzk0LVfus0NDLLSm2XMondPMwkQhyozROK1cm1viGBzFy2py9OdEd4EZn
tSNgdiZkS5tu8x+XA889/E+Y/mQzhNwqp5WQ226aQJ17298/lJDHITHq0fUaIkJ4zrwb2irdf1DZ
ZnBvdZmX12kwbJZ6tJPigdBvJ/Xu+Ppq5Y4AxlqCcxqXlKzu4UwTO8+IYjCI4e7C5jnn1R8pTdbg
Vcdng4Wmlf/r8fqJMKvgJL1Y5Kkmc7QlIaIDV18fqkcwABqiGkBNzdBOKEYjBUuL97CJ5xCqtusl
XTOhOAOaP05vmJ/2I+Ga/aKh7SL4VOTsRTBwqB9QwvwuZt2Ie/FyeNkfD8n9uX75HN8Hr8aswGWW
kx4t1UScIC7UzhEjMtoHLkeeqmjq+c3K1B+lwTff/xc+xyavDtIALL+FdaaDndEtN/q1XJeUmF0o
3twRnsgzhHNpCWbClAyGfwqkg8C6ERmkEjLIICEDVY+vMHS1DUIt13XLvW1HQ4QjBm+N3gaBE4Pm
znQnW+i+NI3g1pZkD3zXVYXlRmpFZ3nk2ZIw1wpY39oFA9k+9hJPYSRK2jC1ou/eGpEhxqxOVB3H
me64tDqFO0An+xVy1sGWDaTlIMryVsIPkhMLc2W3FkPJt2k2OuNr5GT34rV1zlcIfMdnl1xcnRR4
FcD/dKfC7F+AG4EfqwT5lUuRJcMhdpylpGVjoLqgXfTLwBIWAXDpFzR7aDvvlW8ZIWTsb3nn+bjj
CHGLG5N4ZTQtYVVMl4UwK2ua2BLGB8OR/eSMdmQcJb4qNzH/CbVeOf1XqY/TU4d/zkuRGYKzTHF6
pWRF4XvPcYnSxDEUjOUaUnTDXStcUE60zVKhikwcH8gkQCmp1+4OJ1E4dYnkMIIIaMevugPT+pmV
PKmpoy6dVtpSV4u4DgIu7oBnyQ4I2Uclt6XynmKJ+zwQ9Zkh3yy7LZf5McHQ0ygUYJNgRM5XdX5A
JPp1WKd1PRR/KPOhbKEmjJ4GJdNEbprk1IsUO/6K5LGkXi4OQz8qlT2S17o5nnIlguzZReyyY7V8
8P0ORcUO1EcA0Fi0z2Us9UhE4hAIuKIjT3NDKZYtIkDXhDpnpFjLlq2EKKrOUKgBkA4I7B15in4y
wreSrmPekBCQ+b9/yCz/tiaLDLCU+6BwtF8lFrgqS2mg31eYB2i7FTVI4xnosvjZly81ObDxXiy+
tXgtAWl6CUkmwh8QbbvbOq9TJ9XyZkDCAvzcBgYL41W8pdq+WwMJgkv+x8Nxgsd7PFZP6ixG9Zav
1YuiPZ3CMR4PT8NARJI26N5IcPZcwJT0Ewp8q3sbJd++n/0BqP+DgcVHVP9iKHWJnw1Km5Xy7QVl
iEe26+88dTIuxq/bcE+04azuSs8hAnYJ0umVaE7fBUhWmQ6wiATFCwTeZNF2X4UFw66X3nbC71nM
mjExU/xx34lq/1kXPOz6NPpeAShZoc7wtIUlyE+COPwbcgzLXkmO81GK4fznGhM+J3khAYz2EDrC
UwTNvK9UHGwJCov1/Cb0Y6AJx2TpmoVprwpodCGUALMa92pORjB6/aXtS6SiVhjl5pdcE9KDBE7i
/yV0TfCzuO8zdXjLv3rDoj9wmHeNHywjsBAH8YePLDAX5HsJJmD89ajNeU3R6SvrkhZdXPfxPGxM
BbBQItFcejIy9/RUfhl1mSnH7RonufbOWYPnmX4oipNDHdFgY0TpSyrooaTz53niJsbsUli/34TG
6eVn0cyz18Y1LYBAHD4haT1KJZ9xEgtEdG75rK1pJXW/LZTDvtNvxUk93OmornymVrP4q/T16JT4
KrvYYIm58v5quJiyfc6Xl7PW1xIv721T+QtffXKedrx/ClxKhNtwmWKPp+j1tgPUUOYoRBEE140E
99GS02YWf0MsKH3YDlsDFI/rZ0crE5qX2RV11Cj1wx0ppx7OODMguUp8y1bAW0s8p+Ja8BOs+7FK
B/1zWrUoqptX96mBFSctHdAtQfh8oOkIuvI8evxO/v56e2r+7v/dJrOXwmFN/J4RzgKDpcXgN7gn
s446Svf74cQU1IeGCxCD+akaO8wUTyxOc3mQu2ECdS/BWbY6PfsJ8Cb+GaQ9hFCgDcgrn+5JJt1V
CoW2YkrGmZ2zitDnC4182IU8eGCt9u0yKQWrOxKoKzDy+1+JpqQDiCzOcwFaFkaZ0bPR7VyI9Mi+
R0/R1Qv2IZeiVbuR4hBNSXpJbSWDf3D+5GyS/DXrGxwSYeiYdoJrh0cH4f9mu20HWveEm0raFao7
ntj/sPPF5xY23p91OXIHLKhugb7svAC37LRqUFBpopwXXRNWMjoMU8z9SN0QEFz4ZFevvvJm5sDr
/Tszk2tGKl7Xxneg25rWRzZ7d5tTprHtW+36G9QdNGR/0AYrUEgpob2Y/Ij7ujgw/kVg7nllg6LT
SI57Pa2NhPX1SpyIA2pVXk9FO/1kp5Gr+9Q5MfAwPqI8tDmtHn+wfMXFNRQUh1pIvbcaCnXrQ7cT
o8gsf2A15R6CY2okNOOoczSkQ5uLQKcTx8svlrOE38GBm4VOgXMUnZx/3j7om4W+L0t/PE+2XPw6
02vIpFpw0OBRnE3FPI8+1v+yTrhdBmfRPhzX8BAvH1QqZhCPmxt5BqcE0SBrdzIgUP6ObeH9aLl5
+QrkxDagAB8b4k7JzmFCZketQXVUXM4UTKaeUANWTUlJ+ua5GSsyiEL7j6+VzgvrwKYg4t9OnpsZ
MY9F5ecfZOJp3CbVTcJ6DjB55fv4JjpBxkOb/A9nNOJC7MQk3to9+RkFSwX6jBCnTD8mkQRBjipF
n8UKRjcfoa7IFzGcvikem79K5L5k96VCghgpfYyKVeI+Y5NIjVllG4UcUjAUUNBFdZzfza7QuL4V
6MSmb9/5JWOJYBE++X+Pv6f75luzL8x4tWgcvsDh+D3tvazi8SzPEI29zDvOKACgtASDtqkylIIL
ri4GLYLqY/+hLikSQeCg+uIFAw/Tp07dTc6w0oBwhU+Bs0i4PXtqBrtUU6f/wXiI/tc1u4uLtnnB
eDdwUvslws5A/kwutqXNk91cEdZYkxMuLBt0lkMAZSnjLSZHnh4sLKtknJq9MpWHMPi9GoBWWUVS
LiP1vMU5TqbMuOSDSzE5r81bCeW3xVb4ffba0FYrAMBDnEA2JBgLiM06NvCnDGXut0VCqlNXuVlz
53aPmojP/V7dpEtzfYbjWfS8NbraM62JAtBAcctCT6ert6UVG4W9tYL6/NGABMXzsv7G/13zUzoh
lxMVlyD3mIJTSGMHQ9UD7dMRzNXq/G9aDNF91q1HUR2vaPWQN2hU5HEOtqiJVwG/Ioj+agaynPeU
bW1Sd8+kxfEwW+k9xTp7W2/ZyCtekb2fADhBk1HvUjq1HBjxvZC2+iVjUfrsP47a9G1es3BJ19Sm
A35f4o3Mm5hTDpiI3kb1UuQ/Z5HrMdwLIRY29mMHH1XQzd2cjmpakDPrxzDxEyp3rSggko9RDiEf
8V0tyrC04PR2szNIihG0hyJ8USdz8O/J6A9ryEfsfaVlWxMMX4l/Vbz5IF15zsqeQYUru0pMhHsa
SSqqEgv1Frrfu9T3e1wmknocoFwZrXo721Fza2xfA3GeUzfEbNwm8eL5LmyZMiWlkNRMjIzJiO5G
sxL6+5UNo19jCo3EWvDE3y6Dm83+DECQRqggZaWD2kNEZuLKzFefC9v9koDOaGygaSIlMBjs9Ngy
xWW03NSUOroEpUHn8Ltwc3VLUo3y9GRl3z9a9ESOJi3K388eKvM+7Urt4fqqZns03LK1PlCFQwL5
PYHbMnuKhgWlKoItZbAxY7n+t96Z9twPQNAn4BFHgnGhbmgEid6kLliNF9lXpfXme7UxlGtzcIxP
c+q+m/0yr2AElVQmiQ1o1qUUmZ9Pec3vRAMjORSJqurdiFPF/X49KFbzQimjX4mk8npFiY8gwV16
lsO+9VFC4Ar/9EDBjzmRf5PdQb8A/ND0cjrcl5MvJ1rLopHrbSBQeyH/PGkBfJTAd5+b6kRGIVCa
yBnrKoN1ihDgmqLQhtjvALz40m2glk01vrrH1mvQ6JxEeLu5aLe36CD+fKJyqyyE1aOelRcWjdk5
jjXjJy7zQeAhMlAVWnjyx7HUUhh8pWfZb3iDCysCZWIgdKZqBeX6G4oVbGMZGjg3hrdWSbDTq/FQ
dU+P5B8QYQ1XyvV5hoqO7OucmP88AVZW5aYeTiRm09/qUQ6pHLbuB+c3/FCpUteMZfq9748pd2SS
jnM5H6JinWuir2WaxM5+n+Qz079405SMSSpnfe+6OAGmxXHz7oGNlHuInt+Ifxv0/LDq+aav9U+S
pednlXwshhoNHcLpjSCRJheoMMWrdUBN0I9Qn2gvybscWfH/B2hQmoDi+7QNRzYDVUbY4muPjUus
2w2YOng9dDaNlV7Lk3OYjwApAClgQ6OZt9kNy6qqPs5tSOb2qGXnz/XvaIeuLB/UvjInavpbvVHK
OpWtHHICzub9Zn4w+Ezse0ieyD7g0JyhlzroOWcrc4YdjEeq4C1uzREZS1arxwoP1pNSnTJq9BAO
WDRgTFmNcFalaKccILAbEqNWODzxNVlJMjs1OnZMdAT2cXY381VD+m4JphdNxjn/Xq5WnkE6SJQJ
koihHjHgTqxxjR4dJXE+BA9kyIVMnOT5bBVPOa6mMzmU9F5ajEJ781vDEoLcVTBtthtBKlc/eZx1
Bvd61TAEORngDLG8rfoBIzK64qQabtWuQ+4I3cRaEAIu2CI0GGe9v05pfeBjogmTjYg5dtywDK9q
G+3SKarMPvF2a26y2b89wGdrquEUmbysX/g+tFlEkBpN95nghVAAoyDLldNYW1YLpkt3kkrSiF1d
Zbc21Ux0hUtXTsdXpJEB6xz+9PgnOiR98HJB/F8j+qtq+Sy3Z1R7hBF6l/qX82rpnaQ3rEsAOyVt
FtbB3hqdvDCj6xPguiXxxoVplaMT7ZbPOTpXr8bpsxw1lY5OIP28fasJWbH1hilu3lexw7/cK0Lk
A1p7wZ3xpWfZr0rI/DCpjENMjC4Shih4zcYc8vaV8gsR3JH7t4GU0SM3xSIZpU0ydq69wQyeUxKt
H58vcmWluf7R3Pubkp9tOAJWPNV2IxLuPo0Myad6OrRyPjN7gTIzzP8ubcDxAN8owQO5dqUquXd6
70tfAuGH9CEdQ0sWvHNf2BxnMgbGAlVUcFbBDIH9oVXaVmyFAesh0wQ1EKVmtmGdTAWk+OevnYS+
qLFe8ceYG7zukCdt4FBgHJychiLBIRLqon7XKUwTmXPGP4gMFH75emS9mEMCpM8WIYogklW3TFGM
XvKLltSYql2u5j9kZ8X/Gh5bRM+Fn/c32U1ODOFIj+w8DKCWwcxNCQH0LmTFrOdQ0AJxXhFptz6m
PCXCUHaSAxtnoTUb7B/kA/b3P8ZVukH3TRxAQd03dz0MjnHVCXyJJRqaoCDj1T9miL90rscn3ilc
WXOhRmeiODhqdSi6ZX3tXpYd/E48vxogu6JbrMlAPG9FBS1UtHoIRt187x7tehjPEGUHTM45rjmu
mmGQFrEQeQ92WQdDkTFsIEVKO20HCg97/wi6pV092HPAnL6BszfvqKBmSQnXu0G9H6EOOItOJAMP
ArV99Ct4SiNwXvll5Kl/YR5cWczRJ9ztyCIl68BgV0MdNadlnN01S9Fh8iJq6Dptm1NM600a9X5L
mtzqZnUCGhhRDb13ij+ZlgKMjq/+rmZDvnasV3kG5HQqatm7ElNsX0P2er2WNV2DTEJ9nlnW1P6p
WIm8sFbB6npp2Gu0N5HweIZuVq4jHbUHvKS4BjqSqbPOjDen5X3U9snXS3o0s/WyK4Zz9QT2W6uf
J3a2q/cdUrTr+9Dmda9Du2tQiwgUlGb/kn2QQl0oE0G5fleVZvZVJu8WDqBHKLvPGlAjg8iU5MDj
/HlA7683BkDVmI4GrQLGGnq7HQVUHMOQWe6Ps6XFPcqMZ8VinOuJozez+Z6L9rHxLNxrP3c+KqMs
uqyjosyHvClhGBn2gM5q5ljF4Vd90iLnkKkaii98R+FSIZAs2pY4y7QnWFNYkqFRmtYenSTiSWde
6hqk1UGgDlOV168eb4mJKeiHfPEwH35ORjaefm2Y/6iV62QAPQYD0LndYY0NWearzCHskX4ReZO5
BBiYzvil9v8TmGXkVbO3JLsD/hFbgd0K7rmae7nHicVvpzVLLLOR6BefSLZ/qI6hM/10PmnF8lHr
Do3aE4LRtxhSZ8IOLNizo1CAVAX4Td0sarADlCMEXYp4myld3OhkvLyU+GqmGiUN1tFKIvMhPTQW
HYc2XwTjSjDhIfT4RrQ66jmXMns8rRYfYIoIJCZp55XBOFppqBHpqMkdfqhLy8oH735a2F4FP9gJ
D1O/GmKEGTk35Bx9+AHOXuDmtceQjUhhOUhxAwqqQXVh6BdrwpGvdE6Qy5Ii33l0maSCTmfONElV
gr/DLhfFpMr6UyJOur3wW7oZ3hd+Cu4RLJY/pW+/1b1c7WngsoiH9Y6OT8upiU0i4sRits6/2fw8
bgz/FkWwi5H9bUp8mhtWN5GysF343i95PbV+ht9uLBXxUZhY0hLDpptxL7GtmMJp/YzQv+6+rHGH
4dGNOyn5xzWEusZrd8ZOtu3dtQqE1f9FThCw5gsfC4goaTzO8RoLmGqke6fnu7WFJfRxno8sIGTs
sZAnP3Uv2p3GwjDQn6CkPN/9k3wlX3WnxF7aQvazm9VtsibVU9dPax7FwJvRLv9x7g8xon2wKDwv
OCcQSycyL8yi6i5G+qBLxXvP0RI5rVlXqDRWZuYN1O7L1TbZMfQyTlTAMl6SQ/bU3tYeuxhg1i5c
Y5E2fE/d+kCFI38yuNIjFmv4qdJHC/cIkBcJco1VBHpnQBs/YM/9tEsKf4uimBFeSVBLuy/ymnhD
4s+s2k+yuim6O6pSBg4ahRWmDUm4TfaAx/lz6lIF3xXLuw81PHECb3adkEMTvlDg+aWZmGtOQkEt
P8vGw+L611eRAP+f9eFzjkC4lUBuuOszN2UPy2Ic8BpmzNCOAMhpcu0QXaFtIr/at9ruCSE2tnoU
CaXFwPtfvyyBX9M3weVhvcRJL51TIlsDjkKpA6NvDUDDREAIPCC1ZkDjMhnfyxzEWmhSoo13WcUt
NvMBkgb5QInP9iSHbczNtXqIM6VNuKoGpggd6nqnngg9P0XfpBeVBfMoB5GPM8hrjIJcGB5ilJi7
OtVP4DtJ2xa3bRiXUkJueTYscuAQmhGWA9w8EIIiLoXB82OzkVU1veYrkCtIyqZGeNsHp56NEpKB
IMFK8scwX/RpgmLzwaY2dAVLNgNST3H3ZaAxy21lyDu9QtSMMoio/2xF3ugSOIVq+H3YAZpwpFnB
j87sh1I4Ik9cb4ed/3dCmUgrM6T77CeIuOfyTEpNMXTNlQE40chYFKGN81Hax/yA//Ic+9pmg8IL
XroMEDpyZErLLvq7HUtChtyzS1zBn37luXgEV4Pn/PgfFXfnD4cnvlTmlTyaVXvXUH320kZMt+va
1yGIcpfV1Vi7pBhK9Pn8s1NHtkoAKwgftX9myBgTMoxOhCmiLrU764Sjhpuqw3Y+uuCjFSvUdfnQ
myp8UESzuFQjxYXgT4bqnm2g0XjrUOmVwj87n/+au4KNoBekdQC8X97dyb6z01tMVwojfPTmJ+hH
ApJB4rNepwcIzhC96Sj74ZfejWRa0Yhvxf7EfahKfx5FXfhryVBui01P95sqKWdM5/jPkTC9AGLi
t81mi/qwoIReQM3ujJntSH4/5W4HR5dC6tAV2B6Zc9niK+ZhuJa3xyUP88V/rWoCVvdLf2YQo/Ec
t2n/NE0IQ/B9Ql5YsPS+lEsDi3SajbFwfE6QLtk3KbH2VfXtFIBjKWaPX/baCQRH8BVYScMQMmN4
0iOU7Fb7oXqLRplMrkbZAndkn+hLzs8HBiMO9ex/XteFUOm0dMPYmDWD3dvU247fJa3qv0hWQ7WV
eWrFnU9A+SKrIV6D+fM/66xMywNncmC/lGzrA7d3cW6ARR0FPyOTigkfLhV/NTXwaoQeDfglpRh8
LnrLVMPhYgtn9gDf7Bx4XsOWptkataesU4L2dR2UHCeA6y5scGy9rf7q+T7OhnVCsGODzOyaDDdZ
x6H9UNgTqHctScxuMVQ1JSRLvl8YztvLSa16o7P2tiWM6WbSHE7DyrDrneVPietkVMk2dM8U5rAP
IFrdfFStfStb7627MHnbgAR2HWSVJGDbkj5Z3x8oro7cBe7GhmexIu+T7Rif3J2VmA28XERTrTXI
s7XoAR1qkuXRJeZNx+1seW6ZRKCOBPX753RglSdtLcH436GO5PzogCCLwSOA2ZHevTwyJgCTC9tT
0ymVXVT8IZyZnj8VqIxuyHgn81/k/GzwHK5cML4xUxcUbpoCVMBMsI8gMDWmA2tokgOIpVd/9NY+
+wDrYCiWYOFndm0J6TUmI8cAFxr6HP1RVRySrftzBtdYUEJAoDNpy1Fy64eqE0S/61JaVtGwIeye
RAOnQPZnzkTebabSE9r4n/wmeRex6FrjqcuLJo1eUHljy7SHgTZIVpeguSBAUQINacXhiZJ6cPUY
dNCRhpbI3ielUs0zxSJeW87R8Ek2Lqp00ibLlxpmH+lLYUOiQxuhpAjR+tws7LN5kHquHxYTPHwF
/g3csNbwXSzv41KmyP40dRg5Ipf9cz8qrWKcoXfsZ/rGKeG+Ife00y1hLoT9Ah0n3iIPLldPp7ro
QDZx9N4rOgBydcCMehy87KKsKMksJbKfM5Vs09hMOgE7z0U57Fnufk24BBFUKEKGYkoF8ID4v2sX
zErQfHbBkUbqcPPIWnPptkVd7cSj1cjoRsY0VJdWZD5lEP3jGufHH7ClSgPPyi6OhlU6cSI0LEcB
2flVKCA77om9LIpYLjotfmKuJuICkPhywN9Vr7fypf0pikfyIc6TGeVzSWvNDeMfimnsJIgOgLRK
DX0tSD/WAjyUJTymcfE83xRfNX7CEtBYbBrsZeQyJ2ZbHCLvOz8pGM7T3wqvLHERcX9HcdzDQpt0
Vs5/7wLkYucZk4OEcNrt71rm+wYLVsMPKWGZcAtnH1YPql7dh7/PPY08VW+wnfZNBdzXi98BA5Np
aqP3DHaEiPRVD+QmANTgYjW68Jm4EKpLH4w2HkPJy+MERyUhXMgTxudNQzsrvvnGVm0yQco+BJZt
m4wRSjZVBVUY/TRZx5/HtWwGUB8nlOFAvi3boyw0l1zUp0v1AcWfdHh8j+p2L6ohvXg1qvcYV7yG
2iSQ6lXxZoO/AmTxiKuWCJVoavgq+tzLaSzIWlYqaOt+b8fHes6+UDUeABOwal82vGb8DND/M5kX
G1xUlY7jzisI65l9kvn93mHOueDIwWts5yxDOMoqu2hpSKKgFI1wq2G6pNfFFO8xwL6yJ3JPhC3N
9z/Zw5zixrZUQgtBZTMr7yQhsUE70eCufnH443UVerEU0kOlRhbc2YpQ+P3v9c/zRGhcgjEO6EvC
i9aLehIT/0K3uAWLiX2hmvIy1PWg0u6SqeQQ7FFS4WK5rbn3v6ucWzOt8VjfZX7MljjbWlIH13iO
GVGHeKrOAvIqUj3BKuNEnvJtUBnzLYAP3FnJJiI4yb7rxniw9oUT3T+LTJnEmFgs6/mbG221zDH6
MhzTE9kPUc6Ak8leO0lTovArlWNBsh1haHvnKTTZMkIqKTMc+YNPECO5hj/v55pi7/JOQtLKWeEg
G2zVfzgsMGsvzFH/QpwBrFExzPWHhOX/NaAAOU2hwvWS0r1nsB3ZXeTJT6wGJSP2ZsEEPTlCzRBx
NgJOB0EGEWVQQe0D2fyUY1ube6Z8LWPjYNLhUTNs04ARNFUMZc7I4FVQZnI4P6d4KBHOCIEZNdQ0
eHaJiqqaEHVdyrT34L8PoIbqrpBD2UY3f8I8BiQdNg4j/+s/9/iel9AYoLfVJUtrwxCFvhD5iT5x
bl4AYN53urRQ6aPQAMBbFp33JeFW1x0/XjG+V2Gx+PuqUPjDgJJ58u5mYbr5zJR0H0HI1VHToxov
YHWY3rTOi5R5wdQUtRkcccG1stwuHM4jlMs9sNiv8rislq7UJi0EgyG7R4Mp18/6tSTBxxuODzOY
wZ2xkUgVDVnw8X5XAgiYfOzArL4pjN0qb9Uie8IKJ6XIWTrsF4tm/8bq8Ff/NBbpOCXxMnhPWrLW
nTPJcLTOT75SVr6inwQBHmmPOvVe3U6WSGkj8CjOyGGwBYu+vMI+SUxppwnXoVYnlduKO9IVOAz4
KO/d0nXIabCkAZtTMtVBV+Kt/1ixebXI2zgQmFh8xqlTpDGxcNdJicW5iOKPCwOyP3Q6vwBKHF6s
nhnA0hp4CkyG1LYrxucZ1RUkZWVSz4jTFVXRbU3XeKo5dPHTenTJ8MVYFdWsg2GXlTVzm++eT1na
d7GmzaS3LOvFB76QCGq4/Euc5WAhE6h7h6fjiF+/+1/s+mdhCmDtLO1nsuO3EBgdtweAJIR4J/le
iMeHGd3Lqz5H44Ty3RL964c7nRX1qi0t3FvIYpjNat+yDYHMqDdGJ3dvTREBWRjJIvI6uVGLAtog
qV4YzlNttIJ2eROArzryb4Aa3gMD4sp38JGvcS1HWP7jyb5GKbPClCm2VXnBuRcqKwvFV2mr9UXS
XM24kj3PQ8AaMlLuItcl8jFKK3O3jWSNvKrTL13Z53hwfTmAp+dZr1GDX5cuuDvYHeWJ0pbrDCiN
5/lYxsisCZ0jdwOwQ0KqTb2vlKmyFLPszKkmfII15/IX7Jq5jt7aMQ8iwc6S1cUg8OH71fiaLvLe
2Hq8UGz/SXF0YEg3oTjctktCA21i5T0IBES3PQlwwR3BUlcAlLqsDVLcwEroL9m8wpHncIzRtOSK
e42DxhUSpH/CiACFX3a1L6CvshMW3KhRGnhwwc2P0WoIOekPRJpBvwHbVokbjCISFLlYkcSqySHs
7APBE1OjwECYzRkhzzAgCwHah9my6nAXoLcKYm+PxLEF06Y6trajOVc3MYa9/VEDcP1s7zRByliO
298Im8wYOXXMnekNARkvFS/5aygPD0v/I2RPPLHseTy97T63gO/FgNx3NQgw7q9dM/6Km71EjInN
ILzoHq0gEJI8et3C+/fvd0VtjablSMOO6W4NJnr3YuT8tKaenArExYadqiGWIWN+lwtYxwvNuvg7
1K1d9yYf1+VVr7nPt8NlVzspXKFuWCwqH0Y90zwhKGERue/CpBfYxaxyGuf543bgYX40qrcJVZPp
5yj8YQ7qWL1KetDRIhQ4pUAqOTcEu9oX/fJqHO5ifcot/YIcNs0tjqWb1jCL7idlS6XIuWH8d3Di
g3UpSD5dA/Arot+F6FIAgcclPoFzo9pkCJ0z5HnGDvMvXH70/Ldhy1X2guegS9GwTIkbLX25hoac
J6GBJ5HJ5RfVk7JIqkFTm8PJW6vLO3NQlvVwMLY2KFMV60D06fSzJx0DsVMgIpSGBHtMdajLOjE0
U7jpJ1OHN1P0k+7p52PQzZNRlGw+o7Sla3/DpwB0ZEqEoUUKtaRI89yLNTw8eDrHDNYgg7T8icp7
VMnLoOpQ9IRsGVPgRsXnzxIOv7Y48wibBaIkXuxm/xCzI3N0AwdfYOVZ8MqIGb7/Vo/jBbhcXYcC
nHDtq6nuJ2vhZI4WaFPo04S48JXOrbRXEBC7oJed98DzR6gcwNIXLtgK0tQoJ9YhQ/l8oZYZN/Mf
zTFSltos/lGeoopW59K1FiCZO+SnV2LZSxBV73kmoR2lZa2Pky1CTZ0atBAFilORDgC+YA9kNjz3
P6Aqaz408JCAKppH8gV2FqndOBrOvzSB+gPyXAft0IL7xRCFE4L7orjL+HK12u5O6+05lpDbQetV
Xx4TgUBgij5IMdFIyDcMrdg4Eej6uF/nsCoFlAu53qs2OacBirNR1RAAe8PIBvY1Y0rju1PKhx75
4tAyeR3cnBYwpkg1KcSUpxPfs8L6MMqgAynHQgVas/TnIsk4MABvFHr6qi7wg7f+eQy6ES71/7QF
nWMOpMSZRuDToausBXKnfvSib4WLyr2GjmN9x8LCaVMGG3np1z+plAJrNU3engrIMQewjMR9DAB5
nkNyvUzICSkLyahA21hVuD0WnUo+DZ4R0N8MqZn0aGxsygkDXZe5eWwVzHN7vvJe8yBGx989XE6R
skBJ/xjdnolbw5kBqzqxAmS0KlPR5lxV5hrrQnjbOMRWwSs9/bxvxHhRqVM/w8IaqSYuPDPJquil
WPFZ4MtKWP+5DNRu6TCDPxHDyVmV3CDuX15wtJTNLMl9prFqoBTbNFarliPz3UdKko10JM78f71a
MZW7rJY8UkMJkx9BKTQiQSsuEdRjHv5bTfFEldPTDuX+vSPwrpR3jrvQGP7t3B6zKe7qbk5+DL06
BYCKhD0Q6eZdt8uavFpNRTyZ6KohpwitqZOSyG6Y/XKkFLwZoLPjsMabCBcEsxo7+gDqjsZS/kh4
W6SViWKazFpzQKxQ7Ef3Puyq48zt1VHZS6s0T4s1gOXf/UAJwtJDTPxY72/ORCUbVAJdiJA8coT4
4clwhGIauX7/rUfqZsYJzi+bJbxW+FcPfu2qGjaTk+OM1K9Q7WXfoVR8cU+pWhhy5TyN8rkJt6WI
mvteYJNNDIepMtsZY8k2Oqf0JoQz7nlcs90x8lK58nxKlMXcCzeqHtsKF/QyNMw4D1jxme+BMBI1
paW01JLVd5huEBEYsdCXGxrfcfhKt1vM12FDHIthkEm32718pvsM7cvOxMRUSeaB5h3sY7uvwTQA
HBbx8LRjCaKDX7qTo9KqXc4O8jEhagbUoCmuV6EcZjkjcFmpMR7wlFCC0zFBiZ6ymmdiS44IIX8s
lpXCzxlZwu1masbZvk3QiGE5XXMfqH3xEYhrN6gdRdlwOwvmufT1x+lAOsyfE/L1M0f+9YSlSjfW
aCrhexelfWFxKyC34V9yaqzn1o8FNvEmlhEB1fgvw2Sp+881oWKlkz6fttn0tOvnntSS1RGXBZwX
MqzVXv1+M3G/rn0a61XVunPtBAw+5WiNxz8HA/ebr/OIQ7ieuha/8vqrSm4PM03TsnN35jbMUb5R
iaLH3utcttrs9xEpZ8fqUrmSD+4dnft1Ce0e8N3v5GWHeScOQd0ZpUFPS5GcVHg+knhdWalnQijw
BB0wXXd42YfScHIaNqqTcTaRnHgTShOYj+aY54IQMHXZsbOFFll/eNGjiOl4KxStIcNI3LAnEjxf
EGiNu+OMgmhfJBZjg8yKvXcj9SFB8yD76uDyKmQZ+07nyILXPsKgsatH0DVHcYNsM74Fw2CMlg7W
nDGkPrbCqvXAcRzrFAYECDDh81EkDRT39zRRFjN6xHDQZQrIQK8cXmyqoVN/pL9bqyTXTAs4y7oh
6issJ44ZQjTn5szsW6bRUhwuQqthsZKdr6LWWJW6vNUilWl1SW5Ih2NLZknmJM1OMICpEw1mXvvI
tZ82zSyxBQD6k/wHkV+K7QcSm9rIp8/UYe7ZxdEUft57Z7o6gf/FQe/Etf0CJadDF5p/QJQZvx0p
DuUW9BB5g0B1l/yPfa8nHxnOyrItz9/y58JRTjxb8Lgnful9U1T3TTPxqlV1XjnZOSQGuZyyeUSd
hJbqzJvBb6qDlX15HNvxJhqKHH1EKVMNLXsl4LNOE5dz0QzBSinokrENMWY0B6ZzbsT+3JE7zjFO
sZwB9WuBXJTo2TsVpl1cghb8n/D8Ribj6XhhoCUJYOvRex6G9VdfV1ItzFUoQhse2L92XNqFcvo/
0CE+S73HTQICfgeLh94xGt6Iaubhe5c8gMlycDpG6G3NITgTG/vPmmD71ERihZgwYs2tNcHKH7qt
r8gJaosXviwe2GKiB8Qg3Ja1wIupYIE7jhW5kwrCos1RGl5P/SmqMEtGd109UGzSSkYxpBE48cZa
peM1mYMz+mjxuDoDS/cDNctRqwjF4uexP17BJwIfZd0GJIa4fskEG1UWa8MHfTRXGyJwtj35F3l3
whWk60OZV0hJVSfwDr1qaPcFR+MTf7PjlvH3k0dtvTKQjj+ruv6Rbefmr81MOpV6EVTEAgR6cPmH
euN/unEM214z8vnKsdJt4JRbFwBSbvfr85GMU2Nszk/GcgWxTCswALKX91IhROj5RYrZo9xg+vRP
YKetJGmlyNXgdSqWWBl2BVaYTo+fgvqm/wPk3WAonl6iExxT0OnEGKLdz1TJIZxoGFTtyXJcAMkk
o7vxVI9Bq4BVuiHuzkBsB/HlxIeF1QKg7NZLiUihCJdAQERYrFVdPlLxyQmkMAjsotwDD4KXUsB0
RApKEb3iCSuSLOBgafF0ASrrAOQE8u4CCZWwDJqxhnXjq3nW2BKuPqsRHHttOLvzx3hBl8EZfwy+
0IpHR5d5yiRVvTRVXMWpyVgjUeiy6vWucxp/XxwAQicnkXqbc8/u5JBcdooSrvQmhwd5o/S53Wuj
NJ67L3mqI8v4IoSlnoFrtNbK9i7WYlLxNvOGHKWno9MeVWXVHsXM83S5eOfxccda2+gVAm2oIA2z
RdcyrQ5QtSuHzjeL9GD+SQ5ymM38lUj7k6EgXHAN94g4NQVJ5mMpeKLb7Ve+gWMWB17WGHbRaVMk
kI0FZY0EdQY5SoP8nn8frSW/XBTQsivdfGTnAuvtcnwBZU9MIbzwuD4bzdMSHZrwed3VM90MkwyD
BjhDRZ3/edOw0dk6f3ffKTQ2ecAXs/kHJuPm2zni1HLOY8+eeGHJlibn+NsKwDItPCH1Bdhow9uP
CZkT2xAJcBmfAxyza/XZMoRq3ri1MZwTmIJEV41Iel3u6wTOEYwIh8IIF9VDrawGvwmouV5cm8XM
xMRnIXZ5OBWl2QFpE0LGyGoq0Ftvge7dBz6iZ2PySc6Y2j3/C3D2/SvgzHS+a6g5k98AH7S994wQ
jHRcBVdV3X0/+6HYiJxyxHjQg+9ysBkzafGcvp/WknjI+OQ5pV/V6lAn1nv9i6nQryq17L4URvLs
4qymq3EijUVDlS6FX9wmfF1Y9WjmaSHMIrSv4xwXXAGaEUBWAUleOpgpE6LynXuOTcfOmXxOFjTx
683FOucKeomMyB4ko/GrstOy1SJ5kjzMRKdgmnVnQZsjX8KfTOcIN83kLxJ/iJdJ+HcTmX7sMjLM
IFZFv5q83lWqMbFAjFq/0177kQxLxhqqmFu1fn4jgc71dV8jD1P+LHT1d2sRJzTMcg6P9xWkEFnz
m7DnlWhL5kbuZaGlQc8WO9981xf3cNgJ+8g2MaacwOz2gnet51CUdm8127oWjYzml0Q2y7uNTVya
l5za4mF4ZlNwbmn13bXGjStQtxap9MBu8yKl+B/wJ3Q8bTww1Or/ik22kKNRNoKs4yzbskRdtawa
9K1YUYdK9kbZ0QQaaS9vbIyn3XG+axe4W5R7OTK7IoMRxNrdiq50cYEVx3LhelG2RTFeu8oAbL9i
Wj0x2rCb7ew1QvDOIIKsPpJLOJQmYqooxZsKwsKtxM/QaB0JnLg2ZeYBUMvWEnDHt2hUgKiKcp7r
YL1g0ZAZt2/AvX5hYsUEATX0A0md9o0Uf+ORqJJvul3I1paRVbtXzlq3/rLHN4zQBnZNvfcar4KY
rD5CW1UcrrHxbIJSNccUxq0jg2djwNDiOmejHYEaJ9pMjKZ0MS+cW+JcjndUnTfxqhAAu3v5vlcH
FO1uEOuEetWhdR6XhJZU5ylcMIgQVIxVNpeGKHJdNU1R54orzQeoIMgE4CSj5axRzznPhFf9SvEE
nG9Zw3t2grf15bESC38tXvEKEZhinmJffRQ9b0lSqgdS1O9meBeFVCOg5GttQAQ6HNaLW5nKzo4K
DspgtPPtGCE2OJln8hr2uhY0o+I8DEBwwP8JFnkmTuSOgWvB6c/1LHOGNWusfPtGq84BG4dOMRih
gt2BrfbUGUhhIP2uG/aCEjmFTyPdwKYL/jB8Z8wXmnJvGWDEjsKksAPTciWn60iCkZfOf1j3Gw9E
9vob7Ts8mc87v/AauKW5yXYwEw9fvMd2BdxPKfohwGtiy6Bakqbv87UGuNk12nfH1N9EI++o1mAj
9P6pHCVTKHC2Cl7jpSIltqx9ABGJqeHtbxw7ea826JXSYPn/uVAhVx9Mxvj4MLC1+quMPlyr/YdC
yK4I5qNXjCvjDHEEhm9tJLil05fsHG3wu2Ip+wkjvTr08gAaTLZuDyEGBYdnvV6CGRv+9JsvPPZY
KqswMHr/9l4NdFzrj6Hbb3yeEJwDAJmn4BJWSJTMR6XhiylwE1OX2x93is3cehbDFCr7LCMNqiMl
z1Posg4qIcKQxX3GfPVzeUGY1RMPmMlBK+xU98WFTqKaoBGoQ8IasCqdbIlqhdjMTTvh8op7rwAR
VTDGUwBpI1A5Te3xS+O8KryCM5z+xEAXwIfUJei8WTs+kVfZKYFHdurSLP2yTOqJqwI0As/rlcT3
KxNhfIIZVvDJeTtBwP7uBeLbci5IWMv9FztvVYswwzhcgqqK/+w7EKPbvRs3JEryoFBfBjxuAAHI
ZwUtyRRk4/yanQOqQb1cC/SDPNHF5LtHDRAvyWyGHrXC9Cd72fGrO156bBMQSRBaw+cNgAC3e8yH
cZL64hjLKLilNjglJOoCclEF/V0GeVKeS8n0nRSsa2tPN0edsB53ACPLQbRamZxx60RpP2pSp2e6
ahpsirI7B5kIbIQMVzcyhxcdkIZvChUFGdHkrAS3wN8rpj2cKqyE61bocCce8hkRfG3ezxaRCM81
YMSVueogy86od0M4+yZvqrBt8bkX20QI/hmJTjlPDNKplEgJu0hwZ5KG3KwgVcNYWYCFHluPw2X+
ZkN3v0nISrqGkizjtWqqmsxlKXhcIUDB/JMFnH5Xd6Xf2lXbhtOqiPxdFqc6biUTv//12TC6/nGi
nNFOdhUmI8FVQEo1/fTGRQzaVIlKiCXvGwVD4eb8oTVlros/gK4F0AflKtB7xJ8mf27Kq7SR2Fdj
I0CiMSBCWpTJQVRtGvMu/O82VkAfYA7GurhujwhIE7UevYp/PwpCPh46Hpm5POdWaxycy5PX+1+u
twOqxN1okHwjNkWlWhyIuno/fC2UkOqGbeYEhz2lJHhuI9AwEJWXpwnMdgcgKB0138lIxDI6Z7E1
FKBDdcnpvtmzZtFEKxIsfdaQi04vDKJhq5EQEf+qUiqICTgALp/uBHCnEMFH6xl12x9GSyYS+hER
bjBIAugaRIC9aEDgwdY4PAJL/OYSRRXjsG6UOywU08TkCspvZuqt642GJqEl7gLsfXcQau4TS5+X
0eNVwURZc9a7oUyAjLdgJNDPDSxmyrj4X0bHO/q6ptdFy91dpn6EtDFAqJ9OIq1lSYgw9u1OCNtF
SOGhqbEZ9p05eMKltpC/9J7W396SB4vevCg+rBaxHgyDMptM8MNlTyYz7lAOSTeg4WVLoctZ7uam
Z8yGb4caGcMIMWrgbk1NgScVKVceSkRKwNLbPACwFSaWw0YCnlCYehbfagnlVfYja/JKUtHkdPOV
EDf/4SfTxnaghoL0kAcoMnN/F+7ukcGAbwrLVN/ym3tgdhzalsKV1ey/E3LKNp7SgFPO8Zjszk8B
1gETdjiCZknzRVaTgwy9ZpSgDFtWL16SAuCqbKNy2RolWmWCBMrP7R4rb+ezMXjJQfIrwmaKX/BH
367vRDJlmLnsDfn/Sc6HbCYMYC/tbPcNGkL6bIqIguSxfk+u8W6eVEcDrmn3pmhNt4szPVph62s7
JOrszNM8yH4/yzt1EgWd0JZxkzmwUOpMLh1U9gSTiKS6oIehALgx5FTECm1yJYmldAtjC8Ub7SD0
/7P0BdsEJ//pbIEdbp4qw1h9m6rfx5OsZQzChuR1zHrgVeZ48sKb1OeR6Ws4LwmIG2QO0uuYf3NN
ai5MHR9wkuOxmGiTaMO9h+lhYtYPI2p2Ggy5G3wDwCK9Qz7mhAILWKBgNus4EJjmrXDiWDvcHT9H
8i4dyeYOcKrkAeIdbacZpPQLnlPyTNvolJnk5mdLpvo/QQgK2ZuKK+4rjNamn7tzcJ5jvzGGwg05
Pf/d/8K5jPEoPcpo22olzudiZyM4BBLBiMpr2mDNIzAILMAjQOJTT0Xk9cxTR9A5OIUfHKQimm/O
fXDuIFtmFEp4jqwhSD+X7+iRDhrj1eSkqeCnIT70znFM2rIPeQGadXA4U+ps9gqvYliJvwuahp46
SOZi71BYfgmU9kbkyAyhL4jKrdMGQ9u4IcOEHKgThSui3CnaSNzrOCHsiU2YRcujlt+8MATbaOW2
Ws/SU9kDpy8lkh4wZL3sv0rYXTziGRC809OpLj0FNPKY+HXNreWmRTIeNkBRkziNLZ9FkFiyesX0
FswVvg0p9PHdTBxGlZ4RUjH8jqLGsbZAo5gR2vDHSyF6T62oEENIbXssMAqNvmatSiQ2OT/J6g70
WnrQdXDKfeUwtKZZGi+RItPFfv0QcJl0PgsphW6RVvkCX8ETl1TAopgwWw+wR8pwMPdNdJ8F9471
nI0SKKj0sP/1mGBHLYXICkScVz5dtZU/sIdZAR5zz60IsqYTztou+mxxm6Eg83y8DFPaV0acLleh
bJDNAgcSRE5k/jKNcn3z3k+4mlVTmp56x9z6UJFDLz8xEl9/W55pxySiw6b/hNbfRqpNKHexR7rM
Howw46gc7aquw+EuwW3lq+oaJsBgsaHa7KDnrIghIaTjxOTMY4nriXFk6prO4l684Vk462ZHsZNN
XuwXb5YgIv6AwEj5AKoWObsC1VYbH3zKsliCHt4ssZaKKF18cGL5wY4ho7gUnEiLhFLqxLJxhmmi
pY5mBXv9bRvUH2n7GR23bKwRclJJv9HVxM4pvomfROuD/oZBZzjdet4oF+8U8dY2M4onU4BGRW9Z
UBm9UPo40cRpimGlrAMVXle7Qakibk5x9JReGhIOXlbX+Jx48w0AjPRZgrnRiOR0NEs0Kter3/If
wZ6k2Qz1BRuqhJ+vgyRG1oFwGu6LINs2JH5GObdIl6VjS/v5sBYewma0rvZV6hORWNZ9yOxUhGLn
P+sMKurh0TqLlHGs/R4BlRGa+KIjiCJVH+IM/qWYMJhXUZJS7KeNMJXzdTMdvs1XrTJjaILTwCgF
bUTXoCfFA6tg7JCHWkm5ImrNLPLGRW18WAmh/V2021JPM/3uCFdH4Wrj7G4G64q8g9eseE6c2Ff6
gQurZAiAMtyieQlG2cFjrf7kf8SPNZq/yNspdwHjnma8MckMIkY94IacIbeEWFq9zppneExjYelN
5dfCyPTfmYctQ+rEmJ5BihgisafuNNgCwa43/XmIQg3wYPQBAReCohkgDBURjzw4XdpxN3NuFUuK
6k3UFCd9KdoIKRWa23FU2/iUy6tmpJen9vZGrm3zBzk2udkBo6GpQk4q/Y8Lf5Yl8pznrqvQS5Cj
hGxCO1TVQTNKiToOna3inHZ7e8SEDlXXB99TRvt71AmyIie1U7AlNiWK+U+bxB7EkK4AwhsHN+8/
Kn8B7v/xytmexnhBU0i7mRfehPABZKkNydiIaE6ZigpIM8lFU0zWO/7tz1FLmytmQbU336mAlhsG
3qVH9INxzWIqG+nwHySCPne3wLDKPVCdxRzDnYi3wE8K0MWAcC1UYIxMGvEYIGUmkaTwUUKDY+eb
qobtzEPjWAfkyt+XuNZc0Bc7HghmeOLKPi3YL8fbRIzIucHZrf6ZcrNX9Qid/GAyEW/IoelL7TOX
R9d0CBMwoI9RseHS5HP9INB0233Cy8JWjxVv+zenbgxDR7hKQs6w907HJW1u5LkIWO7pTrsuKSqF
MRmi1AXchp+f5vwq9qgomCqyrJT6K6ZcweiBg/scraEaa+gQ+L5aJA3rXxwa88I4rzxAPB0n1yB0
EyQUJfnREP3iC/OPZpBsd/sXjIcjHunVFXoFN58GNn5afNB6yiLwXZ9bQZpvuN9P+Wj9LX75SsYj
D8aMSikw34Zrm8be5O+eG+6o/zYTIUij/xIXLumDKbCDAJnWH8hvVUwec9+hudASw3ZJv9aXdBwJ
K1fI6z5l3CfiMQyW1lpb98FlO1Z/9Zi7mzuz6/GOpa70bBqZtH1aLU5sIFmGK20vPPSjQ/qLw7z0
8yATxYqRHG629/KJ3mgN7k4D9Y83QW2tJNfXBecBtXXra4Vg2JRg2GuODHHxaAJNgidOTf94H0ET
Hzc8rtIfpJNrAD0bRXSIBu3d5XBN7orMEkBBbP4CeMMg69PtQ7ZeDv15dPYTz3fk/P3end2mdn/G
0aeYZJ6Cop2D9Ly4/HB39fhmd1QY2tVDc61DrEMgzE4f1x0/fYQQGwQSkE1Paa+5G+t055aRtskn
FEjJ+FTtpCMEj52pL6ZQjB18hEtYT4skpUD8JABkMBdf7lZrrsjXcPlUjGtIaHvqanPA5Dm0+IHI
LXsYCdsrXSpqkXLEVgDfphIxWvixMJol+l1HbTTG4/xVaDKM4sDaWfbLpvJZ8vmM16h6SHL88Uxx
qyE4ewqkdRxD9XZKUDee8x77Gxff5iDSUd4SNLxH4BsApstJsVeLWj8/oA4DJmINYBeF+MFD/vF+
dfzfWfYPAjR3BLaMbqbKoPW1ki3xzvrsQ5Sg0me9LVEkHTbK0g0sUqxSKAGwI3RFnpMrG7ElSfGX
LlCdJLhNcVlsd/HyuC/gS1d157MF2tXshy3XusY+NjCUtR3LkHeVtwvB8UcWg/wSDau0aNEWmQZR
4dSbrKOWHtton+wE178uEUghE+UmKzXjcAupojvf4ElHe6niKGfdsSdMQE6KgOPx5exNuSHqvZX7
9yZBaBgcDIc2GrZRyeAlSuvRa6b6Vdkkm7PGm6W892BkEbNWWMWJol4pNr1wtYwH0iXb1UPdTEpN
Z8GyBwpqb7g/aTTpraCCnr0LQnAdTQZ5a55UrPp/S6/xcbEflN5G7g/H+BE86BhdU0owCzfW95q7
VSFa7fo9Blmby8CsAXmkvda93Tp3QNw+c+R6BZoIjfsTlJbAf30QvfceZ2I87CsVE7JQ05mzgCoM
glGbM7yhrsHfSnSUOJ36Yq9KwkH933USHOc3gnQIiIyaHByN1cRIPFiDEnkcLM2BXMk+huOlBYPE
PZeYn/kQTEzCU78ZR/Qk/N25n7x1PZCK4ilFw485yo2QcuQMn3wA8Sz/K0NaQItz3g2mNN142Q3m
jzFLO/MYAjSvaJiu/QVX0cIhd8yHbNa3tbXRodibErFyZ0meTF+NxeBa2ANqQk5V32RMbcCIZBB4
+JGhE1c1RwioesgvVVRW4Uzrb9/ufB2CLJjot1iPq1R07Q8SOBUEyKkLqYSqy48FjdhXWXK2fyhX
S94uidCaHtzVSehsNbfQG/8szxfQxmZUrO/D+IsyNpdYsYcG5Li8OmP8srSGBOPn6DCoT4Ap5z/3
ThBgivEoqNbh7Q6W9a3QaXJyTUZCS6QzeMHWt3oDDwMYpal4nM1EofsfbbDjs9AllDYVBBNc5dtA
p4XA7C+/tySsbQ04KtPdP3wnzQY9sSajkTC/rLnQhMRyWS7f4fcEGGjt3U+WK+kZmMhTxkutoerf
5i4WVx/orc3I9zTzYM4lK7J8WODhY05EN06BD9ACt/XqFU9tPPEN1xBx1FIQUi2/XVkBK2XzEe1J
ZXt4rEqKw1B4QIN7EWLQO/Pr4gaAzxXLPSgYDb5OelGprCFAf5tMpSgRS3qWr46HAkL0OZq1DLhd
riKjo+V08n8WV5t1wEz5d14shngUQnaTmjtMfDIkPgmI5SerQ2MAwwO3zhiAmelDCrbx4XbcVpT1
uMhSOOqyrBoAO9jue2Rw4s8VMs/IRpqy/iQnUqL5o7CbSXL0ZjWNx6q4cn25znkYQEN19yMtPjB1
5sBQcNTjGsqRCwAo1b7QVD/GrNFrBGx2STUxhnMjE32mt7GvKefDYlYXHQqEdVUplB7+py7X0BJW
BZMkfg/ovdLzw89UDkcw3sCpFPgLGm/lReJyy6pSg/r1ocVq74LFaix1eNXzrpAU9GpWf+nhv9Wh
OZAeE8GcB0EOnby2VyHfn8XZCVxgZj7/d57TQy4To2NJPl5GwiVcf8cxAECq6XqayI/KGmjm8B/p
minBar6nInobAN6ztWuXdbPa7rBcxbgU8GJ6F+brUgp3i8EtYnkCKcjtftNy9YIO1b4YyiyZb97r
c9pDdlPjGz2FyhZ+WuDE9bcGGP3muI5aS4gV/THcTNMQmSiwcGVrC7xb7ijqYJ4mkt565oX+ryGa
wQt3E/kMbfXWgNrhF15mJetmEPPwz8GEg4iG9+6KWIhe9C5C7q3XXWCll4TtV5b0FwF8XSInH53q
cgzXAj+6fgxhM1uu7Zgaf/MSkU9OL7BICU/yVTb1TNzJuJnBquv67U2kllFabcx/9LUAuqcTueWF
npt4uq7oj0kxA4UFjiYAYypY6oc/ZU5XbjE/XEwM0mLK+UW67uKlo7faUCKwnFk0MN/XXEr0YfpW
CGEZWN9ypQnsjQtCkIAtPUm5zMEA9p/JE3QxB+PKtf1g0SmaR1FdOALRnKimIe0ioDLerCPfOcXd
ywiK2AOO6SEJDiCzsrzIxOevawWO9IsJylUudWliN1RUmOJAJkDJeec47jjVerrB9Zc5Sw7Np+8O
mjotTvlR2gpT9z7gnlRFX/Tw7kE/QOBE5D3gd3hgEixXjZhs4h5DHH6ffWp2fp2A8FsiQkpCu6bk
xVC55949SZGE0QeU9s6B++T9SObdJ5IKOD1AZQ7Bqsrj+A4VOhH6c9gnAXC1gDPJM31zHR72lV3p
2UrTrSlHB4pg7LHjNSuSh6OkzZz8tnaC4fqgIqPplwG1DzyCxV7cDLQVO4IyQZg0ELvGsOarITIE
egeby+8br0cyl5uCaS7Mr4atXbBBTMiymnkbpnR/EMWLW3iy1pM5xdQ9VhJvwetOlm3sCtmQ0cix
YCmdT1AL7OrIEZEp454mM8UysuMf10gLJoEt1AtKreWsPtd1wPFwpdbKKVyBRJIsMbt5D7x99xNL
Z3PYUZjb83Qa98KkbO07ggwSXpFX4dY2PrD2Cp6Tp1YP9e7gMMGL1Gl+l3QGbDcGq5n9+NcA0G5W
f/K+LVmh/+MeLrNp9RAWLZxa2ey/nKbUcgEJgTlXIAFDXKfHLG0EjUjb5WCR+0wTWoUBTBtASAW3
g7+ihtUid4FK3zNOOtKZ3Lx/U5fev+XEihodUJLhLMXNZA7ITAm9CwKMkRV+lsxiUEguOcfLkT3v
bVJBvx4gaFNtQmASjpHOP/ixChXV0cxGfmo1uxHKJS8FHoXjG+RAagL1CStjt4rIzU0/E8QKB2Do
kj1m2nTujhIz1caD1xDD7+Py09GhOs5b9rYeQ6jsXbuvx7rpsmpLu2XpoYnXGFXGXvVVvbn9cOD6
PWkq1CVwjcahA9Oo5pog4hFYIQt8FRy1SvvI9YjXuMizVjN92XKYXMRqxMde0OlGcCZcMpCI4hg1
FE6vZXCTu5fsX+Toqyj2+RzGVJm6/OIZ54HQIR8wlZh76atCqCYiSdT4703CObUMkWvOV6qKaVrz
cxAIJtSAST29JWBCRy2fZU1xvSG4zwQv+3wtOsRqqo54yS9Nt6DTQnauLtQa5zWfOXj/fU07VEnt
P1FehY02NIiy2FjWF5mOigNqzVr/s/+ZqhW9o342uwhH/yYuAnO8UU1W25+Arr/FR5dSUt42Bppy
k3VTvFwVs5TRRi7Tti7UMA1QWlI74HY3WQQi5UZ9QqNNZNwXJyor0Ta11Hzwsk5jY4MujI3uXHCe
NFLo96XNOcGeYCVtB6ZTtd5FXX/GGEOXdcrnjKHToQWwXGKIylqBJY7GC9gpCUTU+5JjlYbLdpNv
K8af0o28EBIGe6sgcJoXSo6pmT/URY+87GpyV4DeCZ3gMGNgP+p6xiPEyaxIPP7/l3IveDM6V7Pc
z/DLq4RQPkwn+GSqg5zhDpDlPukdnEIL+ofnk41vOVYIeR8WQrLlrVtrZVh1A9YjTYgO/0mnuqGn
XBEErTzmDxGpsfP/cdpTvmaLa6YGSqnyX6OB1T8XdXp86dEc1rEDRaa+MqVo4gPeCM/ZfPzkk0YX
vhqy2FKOkcsZ+YK8hfkMPPA82LifZwuYfMwmfGFc2COcORlwwrZV38fanBOOvtfrZ1bIx3zsu4wG
s8SWUhLO/Q7QKP3pLhehoKhr1mbARhLTG9wCic70RsHPIwQShCR9uuxDObxET5TGyras+QendDu6
qSpostXWf9U18/51qx0SuTfjVNgBg9CBGu7GAn4TrOR6LPM8Bxxs2nqoOQp+zpOceAk9owpZ2EdB
/QH20njpz0d2A5QOsgePLEMAUGklMsifFJ7qGiGugchx/FWaNOrZ6uB9zkC1hExkdflfM5f2BVEQ
bNR/PlebBnL3kFl9DVbqSR4950yyD6rWRlu77+dXOyLtHQHG899272nqTn16cDocWNf2LHUeY13u
oHrAko0YMngALv7eYBgBqvw8tx+81vq774prvQEAVg75ECkn2BJvO9R2dmnUdioeD/WQ+oTfVvdf
HQQQvxHl+17MlO9V179B7sfsU66pEGvMvuCWuIyPsBwOEGRBFER0UyRd5Vke2L7bFacglG0uW3JJ
o6jMpUcGvfM28xoPA8vJzZ2YFCPAtnqOhj1JwmOON0QYOfyO6pa1XxGuY/3uq80UPkHiuqh4wHm0
noJq9zs22k8teM9zeXF4eQ9njHWIjShgYMMOnPvz8qQcOtuIFlicHRIpWctKbQ0q0hpr0Ox8aGpp
jffsWUd5eS2eM5cex4BMTNCN5x6MblpSE9cZ/Vf13SVphy5jnDt45ZbvPMEqn4TBpDtD+AunVzCi
naU0Z3XQ+4/jsMm2C/rxQ08jY2dDN3d3TjCvCbKKdWHXTLvE8Yr1Z12LemsgWU9ntvoIecvHg0rL
nP2qI3C2ExnY0nkDfIZEMz3qgHOAXRXVF0mWeFHeHi5zZmghepbFvtFCmXRkH7bXbVAzyorcsikz
htP//xWac32Vx5EpbQADPxRknI6fRHUDQV+JjcnNZ/lp4uib3oZaBJfq/m1QCuBzWC2pOOzkyVOt
162TlAQ3blefCBMtrMkN6DUVKIsEah+ZgT7HOmJthtTd1YeaXmW3Kpnlz0K9QOSqFoVsOasdK1Nk
98P7/FhAbL4uuMr1UfW3t5w9+CrkbkweqokHfwsFQGVMip3pmWku0HS+ssQ6PMnhfXRvtUrseb5T
C6gVoJYwXfhd3vJQUSH1zDL1MtyanmGaNYU0U/gIcjD93+Brjr8mP5Jp72+Q1W0jB7A+f06Li3My
srCV7fx5nHD7DltrrKvedVr1b1jQe08eMHbcOwcWrBP8TK/mpRJOIj72bLJYBk6Yp8Pv1BR8Watl
BuVB3+Jzrf42YHXd5HUSJvTQfGsY9V+QEU7irNPpuYwNjm9OwoU55ErZzNx5YdYIIAMReRmJvwMT
cH4rI2EuyTCY9PhaR6rd89eyOpNGkYcPIoBlQdclmEjRE9ezzgBcrFtKxpsonJOi/nXmuEJ9/ELM
K88EkxwfudPqdQ3W6hmquLoLwjOT6qirx+jFM1fGuG2xq7qHxm0t7zU1fFQocDWeS6089GxqIbY6
FTL/BixMmCMlmeCXM2wXJQoowlmCSyaKUkdYgvqTkPqlHemJXwCmxBal9FyDzqdweu6MheTaRwkn
lvHAhBuCTV2ml2wDsxH3KeawF3IbzLBCwbK58ztX2UduuaCddY5Fm/CPsjaPyUaCtNglR2iHYI/o
KZ9K569mxu6rB814DMlWWg1vG8TKHK3K6IMdXo+FIIXF5nymut1XjA2dzPG5GK3tgABQ+4iHDN+O
4vlxo9wY18Xh4z8UQu2LuYTjnpM10qTp55iMDz9uRi1kkL1m2E4QzH08RPoNEo6W/3BCdfRwwXwj
MV3tIpPvcAdN/zI7wqubOn6mQCf220Jvf1tlIaJkSqg4duOfS2epNDfp5F3AFuViI4toL2atysHB
vxyS/DHd9O4i2+65g+HxbLB2XezYptBa4TksVzlCF1Vb6mUdjfuyGLEW4Q+Zurn2ngBrEdaS7h5k
VxM+NiN5JL2GmcZzcFBSR9iREnjW5tObk5WFobO8ZaxtsrCcTvDUpjKwZm/EjUdNKZK+Skz6VxqO
G8KpihrcLiCOPEhffvSA9FEw69cqtIqiqUIWVTvbyUsMYeYjorzSsEEK4xBawKmus9KWywsQBmQc
6n3WonYQNhFA1NbYlyzo4RknTkh5Q2aE+LlfvjahuMPHcCnW3/lMl7Mzoljyua8UP4d+1Ww+SlHp
MiI4ffoHtA6ji2iSEKyPQbi9SQJMacEZQYwkCgKQcQtORHk0QVSfNoU3ztw5YjC1E+MPTQTez8dS
lVRoSD7zfTzvwVcQiMn/xGkd2I2dmUFZPNfnrpQrl3F8MWL8WBsLC/M+N7wMB0leFweKBo0/3R6y
DXDmKrEBMrvacQ/WxcFqqPsC5/bD0Y18qJTlXQyzdxfJ5jK1pZaSpGC4SrZBWQ0Bd8uU9YCqTGJF
9KpJoN0in/4z874zrU4vWtba6ewSGGW8bxGT3syocHRCepfjPwwj/H292eErBdshFBB9hn14vA/Y
t3fnHMvOAuoPQekQt+BXyWWwXTVKDNhoZjCeJcBniycSIqPpBl3nUR0L9E4WxbD6xDzuFLiAj/lG
xTjLb+hpXzhipUf8asyg4dKSm66COs8ycc7x7SCmBblLgKOSGlSsezboppjA4NWRE/9gS9ULWTWi
7cxDse1EgmIA19xN4b7ATO4XScXWT0J2egQTMEGKy3COfpsJ1SmWhBrsuZnuZ9qomix4IxTB1Yh3
eEj3SryUTNx36xV2UM4OdLZmk9jTnFQnV9EgW7ObiUpr1+4bAPOZiH/F5Fm7xwHftjfa3DeQgHkJ
k1Kg/gEoiFVWxtRnapCW54FhAPy3Rwx0/PuB+zi+y0rGK1rZkzMcYN/RTXIrOldvph2a19DtXkKx
xgw+0KPc1wpN6cbQyPfcj1V2csgvxEWIMEwgZBXcL0u7VxdtOjQuyd538Icvk96umsAYtHSliBrC
K1L5s9wL4aZMDxsJYu7sm7WMQXnheHMOn8eTO7rwaDj5xh9SFMQAgAcEMRzYxgqJ3GiTHVgF/AeB
YqyxmeIIM77sAr6vZ/PfH9nB3+t5KEI+ZBrvte7rjF4Xvsny7kRx/A24i6Ez0+K/CqLp12XxsvtY
v3KW3Sw4Xl6tKU7mOfZhbidymkADakDeJ+IinIm4tRtKtJDkFpALtB6XzH1XPYM92Cee9O39zPA/
GdgGFRvyo/Da4WBpep5xelBi+MzNCIP25S4qkdyRQwr9SLgCA5NdkGokeDNrg8VcyhOmC2a150om
ONbYpywPCprtNmFJiR1wrYFEwoZrvm6QIBR3e/TV0rYb8dpuorXg1yXs+uRjk8u2w/n7IerHQv32
mwQWl+Bq+wWW1ykvCK2tuw3TN02pdXxtqGTs19YeaMAwPWVxKg7wNVIReJX8cjpTePHU9ozW4tCO
CD1PYhvAK9EYL0NXotaubOQp1ZoSJKHY9fducD9bAueoMLs9A7Gp+O5VO0mppECJm5DY6g+LH+21
FE6owUx0tlivkgK6nSaCMNFd4oUI1ONfQ+Xitaz0MnMnVdlZ3vyWFQv95dUqH5CbbBmFFho8/h8M
eQDcugYcnWXh6Tg5LLl2e8/C1fttACHbYHHlRJfX95dKnZXNj/dX0srkdq88GgU6a0yH7TI9MSt9
l8nar7d1TMotMYiICxcwFjOcHE52RTubIGJva0RnzpO0VGtnx44FrZT2El0akaodjI8ou8teV7Ol
hEkWssdp5Vmb+Rofupn5DmDDUr9YagJhAlWgNI44/VlZmI9UdDiYUSeKGPLUYPXtTAz7A7MtVXKk
wNj+/9ROHFRzdJub5USVcqeAdkHnGQOdQa9w887bGbkiGk8RW8SdXmyiwKSsNiprGgMbNhmWGFBZ
u/L6axxKk6K+cia4yx5z+yMRfQ83hMUs0SJqeEcBY4P8exEURuT3yBq8MpKch7usrYvdRtV7R3/N
tjLHqXhnXTw50TFD0fG5frJn4WZksgHtEG55/Rji946qjP40rOU/SvZTy1KCtIC1bGJBYhcy/of5
gjookaun841bKzNCY4+ycL4KNp69IwiR/H0Lx/chGbtf8VOOLDjLqtJj9gzNkPEAJCpjNNDneLr6
/EZHuumI8AgphvTkZNe647beEEelpUhPrJcgsqVviypbO6Mxao92rrA4VXT/jjcyygiCAbGg0evz
ADSfWAOltqv3iV3gAW52FlMS7u0BMRCz8NhOT0RopjkL9Bf2Bz6C2uxNtnVwxmZ41iXsdkWSaJp5
x57Uy8aTRN/tRbRLDKSmBCWQLDU1v1AdBQVVNGknuqIMG01Rzy77Ws2tenZrczp6ayL6/OoVTChh
Zm1xA6gB//9E6luM9iumO4yX0fm6RalQG5GFVBrAAooLjRPyA/CFKQPZm1po+tjjMqOQ2/nH7sd6
RBKW7vzOlcxP7DM8hAU8Nw206hfk19Gg5cq968vI0nK8VxemwXHnZsbBBSanNn0oT+06MuIJ7dHE
awsU+QYWPTbqql36s1VFPxhaMras8BmJE26jZraVZlQQe2kkGHkRSkYtZFS7qEJSfJ1OtgCU8Dvn
KatdfArRlHGRm9ImmMyFOovHSKXhh8ciYKTT8NX6BKZkaw3cqitVZGdHLRgaYHFIDvE0kfzAtIaJ
ZbkeJHs7IoxKiBUQWhEpASjQrgk5I0LYsFhKqLV0yv2L19SSEb6yf8LgWjCZfrdHNq5nkCBpzcdk
K7t+javxbuc86N5QuD+gihWZHMl2qL3HBtxEHCQRK9/LpwZ7M65eJLBo39i1Hbye9gcgTF2NOzeO
5SBfmRYFTojLDHrJ90d17WlCarU8mYEFTbD2yEJKVC7Auf3lIIIvGLxp+0feHEaSlYcN4ntrD6FM
kQ3BnNB7jnXqHdrNTmya0wFKdccRmJf6zo8EhqkPQQPkVkplaqr1C+bnwsOGhJcdjzslv24a3pHx
O3yUdgyg11O5s/hZ0lQVV6W3M3uUaLBhkpdZK25t/oHzV1yGTB+qP0ckBswY6LerF/nZcq+ZospU
iMMFRk42CIu+Vw/aXeSVaPV8RogjBSqXV5MnOMv7mJfF/lLzgVQMFHYBpGFasX1PFQBt2z+abOhD
Egt3D1JWw9nDsfBnrGx9lp/IF5srnAbrX5lBD9daYObmH6qicmWEAyzCBrgMIVtlbZUJ9P7PUbS8
TmCRGrJCF5mEVvVWhTKNwTUcLMQ+G3vZ7V7YmKmnqPywqitcwaGp9fiphKKdbGCQogbY59dXc/VP
6nx6rd3s3wfK/yZ8HbtdWFFTJ3euMaijSwjnNK57oPAsNNQ8JBJfHVj803Qs4uqgTAUgKdCpe5Zl
x4qFlxfgt65w/gD1pLPLf/ghiR2pJ8X4Zdno9BxSHszrQEaW9Ra+wA9NN9UYrZVhh0UeBKzWTvVq
2PsDPwK+MRKyyUYaZf61SDt7LXzS6d5zHxYgeC9qOyMxydKSNTxI4WCuFn9XCuJKKlH1zCedm9d0
Zc0mlC1oDn9kUhlCdVrN7K2U4VYuF0dzW5SfujIlJG1GRSm0pdgZjS7Ilp5f5O/O7qyq15wQeIfW
xm5femouiPK4bNexH7DFO9LOHhSmz4lA9Xi8oRNMkFnASsCOSU81H8jEZmUCAx4yaJJCAI1I9r0z
GgpJoqJzF6TuV4cKht6iTHPdHpUWUgrfxFvfLRCRnkQqDfIzJTbugvA6uYGQy/VONFeNgLcBUl9g
cLpgTNUf1beDO8v5IPg7HdOaLuYk8m+M4YdVJUriDqQ/FWPWj1ukAsBrBJTyY9OzdL6GmVP95wlH
g9e106WGo7jrB36tHCDljJ0g2UEPFYjzJ+NhomtHK7meT4vqRYbBGAahmcu+bfP4BT2lsmxrwg8z
3aBT6rX0zeQ6Bju7rYLcz5Xua2Xwb6a/zLwhoEnQgbJmLNitSj5pBx245ZMuNtxNIJvSP80thbhg
Dn8SE+jGGMRdn/peZpiuOJ8OH8BWmlacf6w0r3A64SFtfAdbsYxpo21/IwBlwWTwbs824qAsq3oo
cG/g8Wk7EnkY+jPg+ZbMTwIzzrHrqzo7jxormtKuoprSDbNplP9hhe701NUq/BfMI+rUGl1og3ET
y0guz3dle2/ONlZoq0pytoPzdiCqSmyk3ERZC+ouo1204fa9WAHV2JR9+HD0YnjBFYbKQr9Pvg4N
5h6QIOmQQbhmupgb3JIM54wwZmLY6dDh4bjFnW5KpGDUtPQAAR9a07jsTpmfB2LwUPxQ3AJbSkNc
CNE81jtBALjojX9nKZBWoWeJI6uyCywQCmiRB/maX6NeToBDhSwrqi4im7Zo+XqtJaVeKsX6sul9
UbiAdRRe+YzK8XNI/+XjY46VikAF2p4L2P5dnBQoXdvbwnodH23Q0oe7Z+4dO4sIuxEOXOQ3Q2E6
SBciGvhLsLcQTl5hnAsAnsLvO51D9Vbn0CRWSCMU5OCgbGt9kI8wclDTEQhTg5MZpNA9PwfHId66
GJJ75hzT4Xkk2p5/DE+dFJotvbysF4s/AjhIXrk7X3+NOwVI8dEgW4ucoSiLHv8tVXde4nY4jiOB
gAGJWdLZo+Vsb6WnD/0Ea5jJZvHU9XmWV6y+6FRB/sZEDCr/4fjO5mbeW1xriJroli3ueM5hDs0X
+RomPSJoJOtelvdcvRrRXFcFmiw1lXIYeBMUEN9dIc7FrRZjSAheDfXNQ00RzAQtLaqsqLwly5fN
7pFZfMS6/dyDUY+gCxKdY7SCFgE0uSrpwK3jkNH9bktw3hD8n0lCSFttAJqmXJNhyvYT/uvcnCvk
u07PsXksuVQ2zXYHo9/Bo9WvHGoyDC1k7UeAcP0SgT/NiyRl1IAH5NokI+4qxUTr3llq5jbOLE3X
ecdr2zeSdAuNscH7nIBOivUEzRq60kP6cCHEBasudNoJyQde6ZS3OMmA+yG5q753eQDkNWn7Iuld
awLa/OLu0sHEoeYzYwQMBIKIG0eX7IRM4Qd3Oxzn1BSkQjN7Mc70qSAxONsJkwbNXSOtHfqA4xbB
kST7CL8qURBLyN2mmZvzUg21Akk1KcRJ/k4v5+Havi/Wd9E4Np4GH2CIU871pVgh65wSyF9eMjB5
iwkvNTMWiEXKymh3fB/WnJZjqVbaETg6PzMMYXqqpIe0JJ/B5ZJyg0di9mcrMZTl7p4q6zWSRVN8
XOTPAZAsieGE7QbMlZcO28XvAXEbg4heo2K/nsGZjjwHOGG1bF4sVB1C9lwS5cBKKb/4cj1Rd80I
CvtrGKhPuLCbMccFWvtpoo56p6WOtd/OaCxx7KwqMk7xkFVtdJAnuJwdVvlNNgDcDFHEtZsyn++6
SjLew8WaGzAH1Cixoseb2+sElt4JWdlDt5oYnpB7dOe0XA0RXC7KijCSpnE37CUbs7wajYMAXCcs
paZBQ89IqJNTiwBIqQCiMV8CKIIYXysLYIkjC2hmVK2Dx22p6Zv0b1NdY5aTmhNiPZ96KWyGdpdk
J2bvpzf1islPJG7WcM9lRHdmyY/bYM+1EYTCtCbtq8NWDfJUu5Dd8H0+Yw3OEcvqpLJXSaC8gUVx
XumvkHM3yYbP7q0q6kFur76NLaZhNlFk7c/+m24wTU/9ipS9xyBsjp8Vf85+GO/bhPNNahuSDw5Q
DR9mm0dUNMhX6u94sIx2evgqOEkSQCFuu4uI/ayrZq+c+Cdq1DaHpovLDbYyRfSHCnYsMk06L0R5
zrvuOgg5Jg+UxPAGpu4wB5EP5j15c2ruj4wkg1A//MHCFYw2HuGqiMK5m8F2lDjghDZHrpHxRN0A
q3NbH0aY1WTfXP9MFfv5KC1ND0hq+kTOR/51ZQCwltBzOxJi12qdNCgvfcTUhlBnosOAGrvQsCKm
39xqQ93sTI4pVMHGbv41NqZRtkOvEfmQuTDfpEuEVpvlo41pY6dTTuAfQCu+snTcfzc9qkrJjbg+
WwJrZ/r3tywYJoXEdXQOgPd8o/8+I2i2t6JxTsnPvyTlZxUFCU2vsdtOKNYR4reGbCwl49d3OwhG
Z4d9yL30Z1BXGmCUCxjr9NmwrKBoOJsmlUhhDNbf89F3D2Z4KHcW9WnAJR6FiBOmO5GqWVK/jybC
1XzsTVOXbFfZU87ohhX6SqyYs3XVy3+qSpDir3JBK/KJidCgqXwelD1NqVKcXwhy9XS0SsvRiXQD
QKQb2urdMRrPtyWlXcB6b6NDiS9SJJiVKPRuCaLChHA8Z8EBW2PYKGwJNQQ16QauEsroZhmTPhoz
9axBawg8csLe/EuPC76+8smjUBs5DeGn/oKs9JN5ibjfDktVOHP7E2oFvlSjsH2LMIvdBnBm0XLj
faKQiTxmTFk7dGAC4JwJUkI0ZbeKs90Nf4ZrMJbjBnWBmZkvDERwXhh25Zr4A63vZv60N/jtsJEx
nAZGSuAqIsxRg/sL4t3gMDkX5DCglfFa+0v8XGrdfRP6JGaeQ5bJLoi6GKEvYFsyXu+lU0NNf2Rn
nIFrUCWBQiPofeLQ5sEpjL3QDh/8FwoZ26bsLp4bKoS33fLsKmaFurx0XrZKQoDWlwgjERn0XFZQ
C/zRGLzWnw1oCB0I6Klp4NlIegrO+IPE9mC4wxZj2A/ttswMVPf2YRl4pIkrHfPUigdQ0mboVtji
9j/qgO3ZCYxoC+T9Sgv7uvyB4nNwsqvc6Fx+gPPzqQHxNtLen3+ieRMHgYJ56etNSuyQ8QHQa8pR
WoyQ1aOrGPBOUgtPBWKG5wG96376tJQOuGEI9QNoymO4GfE1+eCiZ9EcPM1irzyMcMaMaNXVTXPq
P9wFAU+YJxmquPedtVqP12sWBYHVEKhKBtEdpexD0WiKv+vLJRZNkDEwWhc1jpkRScizBe4hlqCk
FiyPkAZ/taDTDoJIjlQ3IWaSGsCiWbHEImTjfB5Atza2lY2T0ou2StobkkChsSHYOGD1mZ3KnfdL
SvflTyzTw8yqAf3pEl/uBoCUYCbM74kg7Lf7xzSoawTSSeCUX53tSEX9OfD2OyEt4tq3FluPxDFp
BVyuXNqqMogvwVbcXEDmOtRMEKu+27RyoJ5KRm1mbyl3VA+JIm42qts2bZWxuPiP5W8ZIn4KNcE6
dngUuzfejw9cgt399L2jDCkrv5IGYZzY87PBm/qX64wylD/hiyHyl31tL1KBzmmYOo5BE3oYJxUP
hcmtxBHob6BPA11HDw4HFcTAk2o43HIVAWtjYwQ4Ts4eEsgFqbOuTsD5AJE5DrDThwuBK+CKJQQo
UWCrIHobMlpa5XNeyY0/syvhn7/ZGwwRz0cFwI7YXE93zHoPJX0kA/zSBfzhoDCiFIQCuoMuQDbw
sNedEi+fF33LOLRgNCPxnA3g9G6lAAlngIw7cC5o2CxeDBe3laJw/x4dobNLgNXbHjVDy56EGs+Q
wAgtDtKVbyp9WewT4x8TAgT2Rdxvj6k0ECk0+eCIV2HN0AKbPX0RvDpdQFp2UXgbpm9TbHWbsSh3
Si43mmQREpZsPb4nTmP+esLN1BjejhV91f0i4AQ6ljTHnEZIMlVgO9qdhOXeCxW2nyojOugi9Gn2
WgWTDUl6MJ/UAjyH7Sk9f6YNvBYJsuUErup5mNdpGtzirjtObLsfufoAOKh4gveBivHDIO8thAZN
EBTRzjQ6CC9yS2UWnpEgsqlytmptv6Px4cLzkVzmJ4lWP9NeB9ndCXUf1JgkLkv6Bd6Vy8qSYszH
DwjzMOauZ33zlBDkqJx1PJmUcJIqDNZ5+bDItdXqoWguBnM1b+SxpaEhrHczFztcKC4/z+yxpzWe
XBLlojhQsBBJ1uQLo77EXbeZGZxSsRod9B50/gRacXOUbiWV6l9YAyPDTYx0frZSr2NiVGE0SOcG
f38UGyfBfz60hWHF75pDdj7Pdz3g87FSLZ6aTicLaKG3wEgTcmN407qNrt7JV/7yTO8APfYqjRBE
7FzXzrd2NRYnf29n5/jxdw0ckcix9Z+Je/n1bnEBaQUO9b54hfaz2zPj8mZtNAVoT6wIxESsV7ki
273Yg+CfJByVwr/qsrUfwK08aJ0guGAbLiS8JYA2Y5X7jgqBz6fahtN7Gf2Fx+ydE/36jbyefWQm
v+AL7MR+nFvETLJSASPz5JO7h4u3vZEUWed+5bbhlFDw8fKtxKgzGs347s6BYmhIs3GXPADPMNf2
UCga7kYVP69UAgYSs453DJsfa+oYQF+BvEeDMJkNlVSFP70pcU9KzCGoQBZKEAxlxJiklO1Tr5Gr
Jqkl0dSuMgN+yjRxkU8CuRuTHvEsy3i7OoCJIhtPGjHh5YfqwulkbOisRiVjZcPj7VRO3EKj/eTb
DEpudyoZJzmlXY8QCli21YCEgV3nXNnsUeHw5EQVRXQyhzEKPLUhojbUhTsKqdGCwGxjt1HCb/U6
URecDg8CrermZ/QxhZBTsl9Mbeb+UxLuqFKAG/mlB+WTnLSABb6InAhYSxnv0gM1haOn4+WgrH53
FZFus5IVgsvrsKSqYI6HOkzkAzYat9YEniISXL9wKpjsxSegIl1/qP8KCfjJuVdfv0OiyFY559Lz
tlBr/npEVbvDINFrjK3dpcAsoe//puzMwGZMbCENj6/59TlyQBAeSKiJDI6AEybMMucIwKri4ak4
UFk3siuH9dn+TWxiswyUR9k/OZOpbfPqh0lGLixbg18n7t6rUQRQucGLRReAu3OVxdQSvS9o4w7J
X1RyxR70kxG4+/t/nPLRYD/8hl43g/4hkER4+SFWiDKjVs8jvgAiVavr+YBEKSfcBKx+EMsMmH/5
62ur3A2qZJsP+sVggskH56+yQjzXdGWNbUSH3e3O1eVOt0RDOZ9gegmGr7Z1qLbw687pX/f5lR+U
dvzUG+SY3+H4Is54nozh06m2p1YWdiBA/kU7urvxUmnliUkDtaFUFyZ1fiXP/PFagUZF+gi9k4Wd
Nb0bYr8NNBPPWuqHhFMsBwYySn6/RRuMydv0Bt94O1f+JOixyXSRBWT5HVQVPTSteum4ZarvrdNY
9xWXqWyvWRiR8ZHXLGnGbbuTQfG/r2H7aZXCbXo=
`pragma protect end_protected
