// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:41:01 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ko9wCFKZb5KtNbV/8n1k/ADugBRl0m3BAdE8bpLlA5SsYOL9/Z5eRn4vHy5m22qE
R8S70HkX0ZEhfAdjFHqzeG+v/zAshQFflyIz4JgqWMxldpBEz5CvwFwYQ9wmckCp
8qp34jG09DRUY9ccnQ1JKiWheIhrKTSquGs+FRihQew=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27216)
WGvx7jCT8T+QDz1RafP9VhwKLR/kwoBC4/pEVwwgSxTN0t87r9hXZThNplK2iTRk
mAW3kHnKHJGpga6K8gMXbT3tRPxQ4Fk9Ei+NQDfv3Wa1QgUQTAn8N3UIsFiG1WYj
UucgrMUdFOgx51+SZGSSUazcIDrKX+/pdINeRR4lcvY51wxUPDYCryBOxDpWLwhh
l/77HdXelE4IMU0wAzhKbz8Zh5U2zZCzrOV0/3PhV9ZxW4Gyz3Cz7Ms/dT9T3mlc
ncuMBTLg/hffmIQPKam51clPfXUfW5Wrng11cluBd2Wh3swet+IXiTWmh7KvvLEn
xHPS3DtmEPZwQeOdbnvZIvbV89UfMz2aE9KfSLNjmifG5e+/hy6j6U6iaJevjERR
TGIawlaNUOtcBc6wMoZ7FIEhuH1FWj09GaDDvuRbS/QEop/mKwTwJsLtHgQ/6VUc
ieXsBEFEWVpy3/yrh9J9kJJ/T7AKlzvEGkO8MjabTMZyCFUfCLmBxhRnSuneQN6C
b+0acRutyxTXvGTJNSJu49fGx7YPLevlXBVHVhBi89fM5K9qUWXfDukyrOMrKj1r
lslkHqnm9E+NpTXQtrIvoBIxHJManporN22tNiWn0X1EH2Mcbm96qVFj5I60ZErp
BrdrELd4K4EUP4ZRXbcbf94jJ2L/sUKn0NxuH1RhygRrfjzd3dS4Q1UlUIM3eptB
aVw6u/idbjX7HXdqqhgLDDw6EgAjVzohsHWz0IH8TTIq/+KTsWm7gEWcN5Eo7umy
MyisYYOph+knfmwVGw9oDoxtDJA84dKjZeXf/oMWgGD1d+XNExFpJkEW/yT9gglO
J2AzuS4670k3FmQIMigsCMc2TR8Ij+fS/JdYIoeg8x/mrdsssm/yUD2Kz6OcxnRQ
uApcXRWzWwtPozzXhv54RVklaCZkrXLAUEYyRDPQvaRhupLce5SMtGhjkRUxzkuO
DWW7cRt2m8cRFFWU30/PKrfe8rLFvvsWr24nNofLRplFEKGlosoEHePX+alzaUUJ
qx7a7XjHqlhMEA6bjgrgY9zFlY9Z/ZtT4e8sq4ladp3AxqUcXd6ZNH9lxOwkKtys
ozmRRyRhMp+f6HFhZhFBgNVNdMYhBI30iBMWzFCLjr6JocpYA0OLmJFNpDzr75Br
HmxHYyUbF2IePk9p1HZsaOr6lnweo4YXJqDB4eSNzRCNG7SYnw6XVUFVLM+KeCbb
n/norYKu/uPepxteLOpg4adTFdbPRYzUy8se7m+tlQ3aa8KnOEQExJ3wG9HxSWF3
H7BTdkgeHo7AUj3p5NpE3QBi2Ry0jitUx+owaoCdID6aKLL+n+7rAUDkNRA/+OFh
fXnnPUTA/G6R541IVhz4Yiw+OXihjBNOIRHT2p3c1J/br+swZM7DW1574mZhDfng
vEZ//UAXWTayWdiC1Nyf8WWhfiDcNGIuQlJpCa8Al2Jac7DaO6NZFOoS7yfXj3df
LkK7t91eThqqW1X0Qd/Uk63i/pwjktqAlGaDzo5saDc9fFzRClks3WINnHcqgA6T
CcRhFamDplP2bKqzNyZHfsBSVCIYEk00IPK0DvA0BStd0hr/tn1ypVivtIidWDst
oMZymKJMjAIPxoaSObwj48E2gLadGJTRi5vOEdM1d87sknmYTZZzj2dcOgu142n6
qii6EEaNG4dG/W9FUMJDOpuqrjDQZior3sD3vYciccIGKJ1/NtfTuUguLN33jNl5
QKcQ2D5m91+kEdlile5BIFF3CN9sjcxO5o351TEdaruuyv4WJ+IEm3R71sTP4LCG
0xxo6YmouKH4WDehZmqU8/pfm2qelUpZwW96BXCPmJiHxjDzpjY0V+sd76YgkGHj
hHU3fgJV9pJqF0MW8KHyw92gtlNKbc94EJaJ8rieTzM8wsp+k8Xuhcd1zdkW9uZK
PlB7SmyC3Z8elX52ahLMngK2DcNGYqwOsqVLpXuYEFcmQvTB7G6/Ami1W3Wrc4pt
Kzk2MEfOr0WotRBTJBrgpLpOC4xgBIUTRoVBO+8pYRpmB4cc+e5p+VlISdOOxYXe
zjbaFtvBKXMHcCJuHVPMGNH1i2YXYEnNedm7laTFRnJ7bj5ousVlJPASTvHlqZLV
ewFbWekfA7Dvo6xmWTAJl3ne3/bUplpJNl9ht3tQoPCuDSWxwjsMcVQ9VGNva6kw
5ya492Hq+KZJ41n+K8VHspKvYeHNRZrCVSLyacyDhx9ArKv5BbEK4fddhn9pVLXM
85W9ulnl/Iqc5rCIGaPSt5GnWsiUAVUUPR+cU0EZAYj/sGgxXV7PZKbkVyAigKGx
El403cHar8frSt3bRIo5EenCulPOT/QBh58b/p6V1ydmYuCoVto2TzwI+aStvLrD
ufy0hakfWKvP4nP8BdEnlcb5aJwg+2jELOrQwBc+QehElObZu2HIxwUxJKxdABx3
QLUJiDq69qI4YhCmlYyGaNUsngz1OK1w6w/wnq/bqr0Z/dRn5Xkh0P0sO9izfnv+
e7uD2/nCi2Dy57psxJ0RMrGtVGahD1BPDMONvR3gPmknqfXbIjiv7T7SeQPzp1Ws
lXDyDBKgfZiHsnTnmkVk1d5yh86Ef3VwcIRfi21TKOkUzvHrvvXs8WkIL0WTccEe
klE1X7E1LpcYdtVragYTDf29XPTngCLGkLFtbwya7T8qXB5Psdc51nrM4ZN6eTAZ
7UjbBPR+FztQC1RKU4vLrM/vprFiiTQSKYFKpJgeh5CacDbeqz/c+6NuKUUV6JJc
ZUj9Ec6hLSj9Zt+33aiM/JI9RlNs3RW6kiXlwSEGu7536XGYNO19zZE9QnB/u+Bq
It6obzroTVF1I8VIo+6kGa9qhAuhoBns4NACVcFU1Liz5bXtosl3WTkjFEQsKaPm
XfGoKfzi6v4X+cjUyd6+M+YmqvOvZQyq0SDxNws1zLW3Vaz5VOoN3SlX/xleOC6v
0vyYRLUQfpm/pyiuQK606+UuMiTm093P2O2j3R7pSC2WJDX4XD81dtsAmnotOXU2
mU5nBa8oPKzd+pCkPg5L3PGVwIZbpA9elUYlQhCNCmdXNNd7fHJBn8g31I4Uble4
F+et1sXKL8OkX+9JYt83nJgJozaQqi84IJgtrrl3NijauOavNCS2tdidWUTx+Dws
s8sEp8FpPbMsqJiaLlORYj5XDxCpeVHwxPtw4DLEkyriyS2foH/RJ2EnFkAJ+L5k
0VOCtOXnL0aWIYi3vXXGsxIZLb8sEU0AuONYk2w2drwlkoLWs21wTBKfOctabMFu
qMajFCSwwtr+aDi/oLVJ6inhfcDe9PXEhf1K4VbKr+NqlkItkORrDpecCqvKMQBH
BTY28EAVMcfS2q6nJS/3n8Un4kyCOHybJwab7xzlizsv1UTqd0SzfrCwNUuRidQe
/CQ+jV0t0VoBdVrZGTF92Ngvvoq2oCFAnKy4XUAG4rljBu6DS2w70dVlf9BBEAND
61ZJTyAX52BmyUWLEVlDnizewsQnQ44//z2DP658fri5bYTwdI0/SahD5P5TWAsH
JYNrk5eZXBnGOloHfo/tDVgMaPhrRiCP3GV9MhtO+OpMBuj80g47+bzkJ/7ZoPSh
6Om/va28pL5Wfgp59Bsy09orzRguL1ORL1FOeVXus5cltam+GhpNxq0Z36aJU44J
u7rxCJ1XWBRbofQBv7L85qMcyXFRBn4FNMyYZJp1+8k0e7WRaigIkroAozceDQZM
wPfqvKOxa8ssfvunVVhvsAohTeCHp0/1RsS8g1T9a/jyHHMefNwxQ/F9flhw5BMZ
b9gE/B5OWwx7Y7rBhyhX4Ai4GjycM3S+KHy3elF5vQfEUrKIueMuli8H+wKkACwR
1Ai9STEOYyRWPbP4Q1DnTbD4ZTWXvIMAhG8dnB7P20S1MROYXv6E7wCS4ebrbmtt
KycpOmWIsO+/rwUGhY75i9MrsWweEqexaMd+NKTNzS4RYtM/a3tg1VYt/2I13jmE
bjVs2GsXBnIt4EqL4hs81IPgaQlfbpPmvTfTumfobg9DbpJqa88FCd5S6wAA5/Bc
DKqQv7W5IComQqN0V6KB9EYBWawm9/jlyCt6GY1sOpOI6qHFxlM8j11boW+VR/Yb
rVrAPNmIf5OvQ0ZoR9G4GgwEVcxhyBfpzuEg7japxLUebEijQZcSynrqN1V7wtL9
AgavgHSln1SSih3MpntU+lNk7jPhBOr+IGUwwgFE4zX9yVRcDWw0d/Oyi6mab11G
7E7oWXrTqSiNbPnadUBF2Dm7fHenq2t42xvj7L3gdMJBZ5XKK/pz4a5o/yJQy2eS
lwGDBvttd32qUSoRhxmyHPPrL2WrNy5TFhIAAnfoIPk3ULr4QO4SKl/4mz/9qS67
cEFJ9573NwqjBt5zMfhLc1woD0BAcLfu5VD5T7133Qg+5+gcArNCdRdoipEY+fzu
uBMqvG5F2GUM++6j0VIAbDfO6mCqo3HeFj3AYde9sdf5zLo24tnGbeifEOog0YiV
1RK4qKby5zbegpdeMpVX1L8XtyYsaYH9QEbhcs0XdtxV92lGM479jiEj4KarSzzB
MxUBsejxFCP4SJFr3Gl6fllpeSK+iX81uI4GVksHSQvJIl28/z/LVznAvd6nF8Lp
YOAYCg5Dwghi2Lg6cjyUD5C5ARbJMGGO/YzGVDwcNggOokYwoFzDbvy26P19HUcL
POw3cvCglb4TtC9/mCiZ9wNAaSpduL9ne1nafirrzguRqUNIK7h65nfh3+wb7duu
DZPWkVjxgrdEj4ZA7k44kfLJYcsRRQBoFjTWRFTUzU7Kj8q2iAwGinxn3TLhCZNl
iTPujUiGw53vrQqH9cLrntQ7sHV4bMVINcdhKFZCucN9mYwLfIk0zd5PbFH40D/L
tUYOaDfbQjl4vKK5KxFMRzzTlfvSG9JtfPjlAJqgc/ahPyxZoXWcVw9Gf9MbqBCc
fU19X3cm/KmncVlcOgRPukHI1xq1hdAjU1FJYvyQ+MyDzcXLk5Hy4LC4MbgnUtkW
9gx/wDY99K4q0oHboQkTyHbGBrr8BW7qUMNdFoztj8RnhFoFrwBtVpiaCMMI7wa2
w2IVODGSuVm1+YgBCKT764SfdSzF7xBbPmwVhJsRmjgjEJcKeAI7cu3NI1tSteT8
6b9fKaEbo0KNYUpEufXcQhyupmNGdFrCmGHppWRalqDZqdY4OrlMVVQfcu/fA8eY
RGT9bhBPv4wNUQa1dD55RCAqBWr2nm1rNx0++ZnuemcHKNr+nrUWXHXjR9kQrZCi
XUwcTEW4MSqYnpS4OAOuvo2wcZSbjyg+TyloAU8hShOpj/bAYycwkGOAyT4W33ZU
oN+rrZVR7w7XP5Z1RKbUQAfMdYfIuP4Nau1vZihc3vmG0Y67RJzO5FfnxN+i3I9t
M4kbPJWEa7E3usod9MmwQ/24sacoAxPb6996OfUlyeDHoB8qpX8Wv1JP5xGVQe9a
LhIXhnK53lth4ciaWZUkukDIN3A+JkNWF9OuD4FbqC8nqeMAuu+FkPu0nIQvJ+7z
Lb11Mt0d9UDo3OBwsVE0Tl2gwXxmGWoXgo5DVdkeR4UI3wOLEI7G1R5tMxoixe73
7TJs4v+6w6f7MjjywHia7OgH2M5v2y5Lk2gWSgUT2ARUZk8EnsQbk2Z2xaRiNeKQ
r9Hz7rSFl/qrJlAuRrhp+Y3mcERR2fTSPZa+llsMUJzVW1DIskxSYn0k2WhQsMxk
MkWp7B/tV9kY4IMRqBVwPgr1L3wa0wixMeGeYKM34OOYDuSazunkrllf1n6zwQtQ
nTeHKm5MB9dm4vPbeh6uiUkR+eq6e/Q6CyHKXe6J9dAAJVPlbmEpOy2EzPEVTuaB
FDZHStyq+Cb53xbkZrialM0LqDRR3ml/xKLx4HXKy5sItkTiule5WdCW8nqgb1ah
fyiQLjugyB6wAC40/wQBWvg39ZLU7SV2ue5Ay3eNreGvK+LDhbP0RMAMKi2/Q6fy
W9P3IYxu2TpPhRentl5swzMKygnw4GADjJM3oRMeC8pLrmpxhJSOvkV1/YWydnim
SVMfhHb+o4qFMfN+N0pfaFDXVeI0t//3G5o1K23fPcTcToKAt1Sfrkops8Ahk9bQ
sdt1lSJWnvao5kGg3rRbSWrlwzJHhp3Er5ukoVSbCdWkQbcl08PKmcYIVP+88kX9
QD3xwDF6IGhFjYuTlw4wpptgeGtB52Nd1Sby2LkyBwAGcqw1/WxhPaSlimSIziV7
aJmAsuahi/FVLNPB3bcnZd24vcOfZEVTtv+5q6nMplGxwL1YnJfb8Ki6rpqm7Lvz
3kSmNnpjnYOwL428HZeULGEfVlKkj+yHppPuHRffX/1qXLE2XA4RMQg2PPJem56o
c+7zEWgLjcGC1SrEGqqg1AB87v4bCvBw6+efLqlS60x660e0A7ETiKGfbDYE/X7z
NSr/dA32aSZmvUHkLHLT3T5+PEVp56NC3FnfsmePqqpo248Sb4HBlHYqb32G8/sK
E06CHLogvPc+9G0VsEtxM+xZw6TgGBg13n05kpY1dNcd74LdUmSRrqqI1beP86Fv
rPimUwQNKErn6rZ72F3nM1XJhB6ZWR/PDcWySstUKtFpAXNxRcZO3FHfJ2ht7UcI
I92ji6Zlg9FUq1GEf7hbEEReT+sRj/4e7cvprFW96aGM0Xzdgy+szN+Uls5dt49V
9nQ7pgIs8WQ3Ptsga6a92UUrtVhkafKnnwPAFtGf5k5rCBulAlX5rww9CYjpvKqA
M4F6Fnzm8QcsumN8P6FeUb2Kt9wn1UPqw4GduXPZO0Smo0vbHmHvLuUPSza34HF0
QQKTuffK18tClWMrnHHhl64SIksBBbributWRzXi9twvXNX57hRLwlZL1ieQZXqk
sAun7OxW5dT0T5SOOA7IkTF3dkroECGhm10bcMzA0QsGfHdcPZ+6JjjkjNIF7HEq
aUoEeHKrq/WGfngfMLUQcky15PBKiIOO7E0nq2lan/Ymf9YhpNeA2HAi0Ggh933R
VAjS1BzEli3i6uhmvqbnbTij0chD1bWVHd4IWvS18jQGNhd4Z1d+XDP1OFpTK4O+
dYbNvw5aBwzUHO69NlgpH6tn3OwwcemdZQ/7Z1pdqp9aO5oH/uQhoouyFT4XQ2vS
hzOb4Eky98cIvlqRRaQNFx80SZc9vMr/B40INQmJr32nZ8UZ/9YrYYCNf1p8oWPH
vczOIoq/uUpAYEia/kXfVEM7tM7OgLVph4xR1Iq5B5il36umVnIy+DrZ/iNgRBgW
fPjOJgPYHz5O4erqfS5XCXYd8TnNuBFPLN3Q7KZFqzwm+o/wsRf1B3goZG0zTLz8
95wumzJ0MENBXTQZLr/YbphbSQidqm+bpSk1gT3L8Pyp2Yw+xkPEXqfkKn0eVHnA
tcMIpE1JqwRtz0bBry+2rXKz8HYxlfYEfRMOahY+LynFyuYyFbt5zpxnFB28WcF0
plniWPqegfa7O4VcMeTfgrm2IYR9ib0tuzI74DBEBKgaT1vMhwSsBpmvFMobfH+T
24APU3RiuBhDpYWsdoLwWQVTrSKAYRC450Joe25crutmBcTvJoMclnJUOZK9RPbY
KjEAYyOKrbajmvCT3oUJqCnZpdx/MbjRIHRSumhEvq/Sjsr9jGPp8PZmoV4qUJol
o8ypqFjbbFrDnCbYoWBfBO3P4iQ4awhIFQKZM1FYlGjJRSxfGLRRjQ5L6HI/JO8p
5AUix+nnpEg+rRNMszrAr0apFB5o2xBTrNxBl7F9gR6VmIFmGl6BIvMCq7BOM/r8
cfZAlTKD+8erJBdHnMKLQXftdZn2ernlC8eksvwT1AvqFNaTb6XLRz6HFM764G3D
5pQoEISizeetiGoXkZvZ0OWKWB3Z42pl/OUvhhUClQXxEtBuNCrjZZDb6DEHQSxf
aGRGIYa6Wk0SuEhLx9iI+1F2oJqgBSLdqyW+FMw5P0/r6PayeVf+o556STTZpy9s
UutdzSQQoyaVePFZaCHPYZW8amfb+v7NoX3vyD8kDrWJAdhiDQuGBLtfx6McH/jZ
ewqW9XLCEUxJBUatSclE6YuUDhqeHdg5pB+KEWxWz3mI8imijFV1gaZ6UIMyZvck
/X6ESqOsEu/mOFdrq18CItJarwhu6j9603cKFkS7pWysj1l1pYtCA5OSWJYTb5by
w1NPV9ugxxESdepDdlqmoAMxiKAe5LcGZT8XbziD1Gn0aUTBvFTix5ZrUBRiDDpQ
FP25BuytBFcQv9+Oyau1JgCDIkDjq9l+h+wh6l56hKHtai6+ch2vstX8KCRz61yf
RoHMVGMldckSdxGg+WMDB4di9x+sN8y8rn4RVlNwl9xsJhqraNyKjiE4sGb/KOrC
DYRv5lbhoEBkoaQe/OniNwEgudFT86El7120aEb894AM3hMRbV7waiPLznNgBD8E
ksjUIqAHaaDAYYMWskxHkNsnl7qck4kJnBZrFyePG+fZj/dZ29OnJMoL9IHxv5HK
155fyIBi5o26DUqd/IygbpWMn+8t7yhhuFtE1xI0o5yD3nxqVgZROy3SSCfl8l+G
yOUhWZvrB4xZGPjlMm6t1cwACPPmFCK0tYOjrzbSbeqYbYSFXNrcdSa1RzhXM4WL
drprok7EMJoRIBop6pfd2LH6DDrkoM3tmuIIUQUDyE2EsK47MQjZZE5hdEQwQI/u
AWeyVv0UKZ4CNc4JUU+H3tA7RhqwFMc2MNt/kMjt/o0sno7zYnc2mE78HUKu62t1
nNTPq06ChfQvjYEShlzz0aX2M0TDEOEnvPVT+STQwBxK63BcDlrqIVfjr4vptJK3
V/0XgbXxzu64y/5r98+Ia3mapmlDSNf33TAnT91vOuFzuXR+lh4fVs+/7552q9Jl
i2EXHOPTn4IlRmq6TmW6ez9cbBSz98f0mE2ZF6nMPgTmJl+jtWNlOZfjbwGrcR/d
6BcYzaeoDLQevCW+FaE9csT6yQSMbZ0Wraa5OVACn4UA1pSjlZsOHF9wVyKKUmrJ
K92ARNa97Q9Oe8uxdMEEIBDgp2cjr53sFXklDt3sLFllVUiASO8Y69U/CGNd91Yv
fbIC9u920nTRy1SQjHlikRNlU029KCCWa60dA6KXNeM/8GUStn73mRxNYnvfbUPg
YAXse2ulMNSf/jzj6RxwfXi5CQXmmTCWPvyzNLAVFb6AXp38dyMZAtm1NG9AOwri
5DHBrPOEQ0oAd8svJOsw2HKOqHZJ3jEaggjy+4fbHAMU85RPV1v3I/mYhcQw7Jjt
GXVxRvFneTLbe+GKphIf+zg1mUBUEqaBGoZWWWq27mr1GnoVrBiv2nI8Hp9Pq15R
LuqCQ+2ukAu0Gt8tzcMsDDtZ+HxKoi80lh7BKqRAlM9KcMqeRd4kiPsEthe5pcR9
/QuENSqVhOgKyvhvYuA+Il+qpXTyRUw+LOIMP9owPokpumgOYNl82ELPsqcpLn8X
9DmkMiI9CgqYSCbME8ajhlzS0uhzPlAbmLu6UWbCbS5a5SsXyOKzxnhZxa87outz
DkGICprsg8czMxsTVFg3J1e/q/nxr/89j2BK/dOrbV2UtgV0QJyXh+sWFeBoPGWe
5UGN55nqZzefJxCFU9O8bfpaCRrqAgBuahnZJWSoHehSiFQ67cdWGukGcOPIIZIm
dp9zgsZwzBdQR/+p1kSphzi6+6ZBSdc3eZ3j9jaf8mXuvKYdYnLU9MyFYs0LUeK5
bcSdHIlznrnMsLNWAyeOh+3JmbUVAy2ZOwrQcnJ+FmGVXvPTP2FLEE5RacA6Wqid
Avpje5fTu0FRlkf7S+jKUdB7GYDhBlaifXQvZ+ULbxSJdbZtygCNzldvDhaHfgJC
FFQk1NuI7mKAyvqBMqRPRwU/36Zk1LH9LXCIy426luPIC+3w1WAW8f3PQuk5ir16
vACBT/mlIS86vmp1reXlzrdgB4nEELyKIkCtI9me9HGuXXKc5wEkC9eh+HacenRm
1byBvECsNk+cJM5l8A1ZWsDzeRBvbaJXUk1kP+JP492trcRAjYcU99PeptIVOmRf
B3qUqXaCrpulcgDgpxj/Ud0IMY1u5iqPCBxsEwpuQgcjbK6BFCjVtmfBVG6q20ML
cDCvnmuvxqMgHcYZbRSpItnBTwRDeCK0potGX4gxRu41+itlSwEECg9hDbzHeQWI
7Zbr4OYDQkmYNPdXM65X5Pu7H15MkrdwuyWY/JxxIFFyjcIXglDonj7CBDmNMlFP
sxPcQxNVu/CgMFFckmrOk8VgXc+Z38Mt2/atIC+u0afvzZDcS5HKP3CoJACTyo5B
Ce3jrgAd6o6pjzz6AWCg+va5ks46w3PmEEz/yyiNthbESeYe71myiEFBBeKjH3i2
0dhzn2shm72QvyWTfhGV3mkg28WbtXnLHcJmEEEFAUfbmx1kUK9VWdXXKxaQFabt
glqxmzYX/NzT96i7RNJgY3WxhuZ621t/cjKfyjhiuNjS/ZUhMFO9kk7IsKaAUidE
IWGF2x4dwPIdRl8gzQwYCe/TT90LbSCJ+OEHBch59js5hZokm1wMPk/13Xx8J7co
IYxDCE5jgPBz/gqS8XAdbU7rZvvscEv4BCUhesCVYdEEu+sVDaNFXW0RwIqjU81Z
HA9jY4O3ABRFRx6bfjNKZZ/FHpUuMiyIeKwqn5I1nYqq3NCz95mjylQNxHhfBzj1
VUr0EWtnYhxVl7EBkWvZySZ1NVChty4TK0Q5RRJib/oa9FHGqDd8J0w5FhHo1jya
gEZpNpbC3jRWW/MD0gCH5+knGH6SaUxwScnc49LpDXwnLqhteu4cVhG6DxuryhN/
LknGfS65xFZlEsBT4sVIO7044SVN1FaLr9IzMUTneHIJ2QJxrTILC+1aOY2VRycO
n/vBbSadPUvz/K8Peqhi08xfANeV7/pb1l7OyOetpTcJ+nFFTlZJntvg/CsPNoV2
q9o8z5D8HYW6D0OCOf0tkPd+10Igc+EjHiwbBGr+qKS5ZN/HFk8fPHkcc+Xdmmvd
0tPh79glUoc/kRg1mCsWFIuNead8mpH9MQmz6u2Hk4233W9edJOUraYjvhVFJCCI
YLOG0/oi693cjbf6uj5z1xNaY9YYOgZ2a+qYqQBUZrRiKYZshwQoJJxm8prHkNk4
/z3AZFAYbg4eVoHuai4/A5fdx1EvftDc+ZJeRQnPM8n6amAjw7bLJUx5ZyCOasP5
gFkowbb5pLDRr4+mU0tJEIrVRtyfPn3e7SxUzop4w9+pLzZM4Q1B+WawVbCr0vv0
h1OFzZNiEUODsFrE7SkQ1jiGKNMyuf3GpK253r9nDXYwvyDXuQctaGoV/h+HR+d4
Nc0ComBOmX7rr+dzM19milLAtw8dwKm/MJrmkrMmNtreSDPLjugYDwLkAyAjwypo
rLzJ94uc8HtrH5RpDM6OgC0fL2q+8aESltwBa9qP0fRskK4LHnDBkJ5BEhW7977p
qk3U+5RWz/kGhjRWXqATRWUBKN3h/AF/u2qNl+98GdZ70tZJD/O+sHoL44i1ISa/
gQwIGkcBJF2nunJM8aK0YgaoBLDM8NnaA9Rw+gdgtckoJ50mXaLNTVpAWZPG7UpS
2jXjZ9sXCeZF2YVN2CaNXEphX3Gj3yXxYvPU2iHtkgOlMX8urSw5I/0twcSVFPtQ
0FBQzOh0gWEtDlAXkWNTPv9MhUGSbwfsiQECxtIepfmgjmiodzG4gFNVyfrtAFpL
bSXCpnB/DukpvimtqnQVkGmXpRcuHMWkUM+PRBMJ6wT1tujqyqHXyVrP15qEE+ll
u2PkT+8nLi60OEGD2uNP4jp/oCzYD0kSTNqW3H86iMl/0bSRU72goxP7X/V+M7DZ
wv5iWZICmdBMEQ469zva2yd0triNJGzoXzr2wi2A1PBLHb0SSmYBHBUrOIsQfLLx
KPHs2un4R4V3Lq2PxpoEm0tQ1KFoiq9m+rWpGzrpedMqKP39XUa/NBsoe5/ssUoG
EiZ+kby9Pvrjf6Hzyq/6zTEl0vireQryfgnuBYhpjqPWEDKxfMmzlaxN77jFYWiY
QoGZaOe/lhjwTzCgrkn3NUb+95GD84TD7ONoY4P1886EjZug9I4hF9WXmUavkbRL
13hdFjkZ7ZtqW+4bQpr7ngxCr36TLjiVcGUsYBEHeDRspQkcQjcY5gvsd+XD2OxW
bP4xpcbicnymSdwlpR0SphH3CmbnBEJ05+9unH6Vz/4H0EtQBDsgMY5RvaNoWcEL
sOSHRHmJLF74/h+KsttaS1nxWZ4NqskbZt6c5RB0vAsKfDjQkftxAjRpZKchyGc9
X1gT5Jgt7P0u0IbPVlQ0qfaTufZXWmgv2MmwYUOzt1wOAlDGqI+X7YZZ75lQ5LmC
wJUBkczPN2AqzMy++dz2wn7lEFus9usRpm8ppzIqgkbbEXj++GIZYJsGfD64rlhI
B1xnv3sazCEEfqhUaAWkCw5BMZTn8Ajvs+mOakEd1+rrx5Kt4QeY4khG/7blyXw8
NbmxNLJCvVlInijoDJ5nkaynYhNzWMEWZ0kIuVRNwxA2qB2QIARburSMQWuc4fy5
kTB/YvUGtLesX7Y1F+ZbPE9Oxzl+xbiNR19w0GIDGd/Z5JSY9V/n5sDIdsWp8TOZ
uVCYa9+bPxam5CGlGCQO+LjKlt/7NBfKxN1xWbKRCCV2k73QEjxv7qoocx9zlT/l
dopcLTCzeR/JdZQOoGv5vXW33bUop51c7WuaT1QZXjkphj/l3YoqqJmudA4tS7hI
sviJAe3QorRGL3tTDbNsXzga6Lwo41UtWR5ZuW9CLQfOodeeS7DQLDX7b92T9U5D
lcEH4mz+6/NSSPy9oM/uDdjeHvKPPLR1jTiBYvTX0osMd4vNBoWo8ss3ZzIWnBiN
V96+cIF9iJbIasjNX/ZwYnzDNHMlIbmQxSuebhqQ7WUfs9ixmfQD6yBSeMvPnSCg
PRdB1X8/1MJZsUiJ/wAG8ZIprAb7N4mxxgNLOSNnM89zX/8gBSGON0t7fUC9HRLi
zmIdXDMASTDkUj2ixSZZKsEGrajEIr4O7cXz7KUEQ2SmuCf8qdbSKLVxCbQ1baNp
DW2JkWQoCcsSoNTrFtRdM5MCCEv9hfeFIWUxyDx3lofH0d7zq8HgNLRDC1NDRgd4
D8RrjFXvGoSyCq7ampDPIkQw9v/5C5gFAe4YtorjexaINki/eawOP2mIM97/NQMf
IDr9iw9e2Ba+B05pTh2lIlY7BVXQO1Ft1sfi5ueP/MeBYqcp0nlbJ0I8oChsNhFP
wGV2dN66wekZFeo6lOMRs/1dSfGXi4WavdsSqkxqBm1gvhvh4FhCJTYPR3bUas2A
FCB9TNgoIYaVN+KQoqgYMkgUZtXYwNEIDQ3suTac4U/yHO6VsPsb5R6vjQTZlZ5g
IFzdWo70z68ImjU2Emmfwoi1XW11Dn7Zx+4tspbIKJYIgeivUt/5jU/CYDBXY7sV
v+0v/i12EXdKxAS2lQM+8/CphUksEdE4sSmHomDSfSifA4oKopqGg0dm4PZD9Emq
h97Lu4GT6HmU/s5jXXnbvsCI2pT6EXZi0J4f8RqtISSetUkvNyy8UcLUqfgj/6lg
e1L/9fas5pGl2bY0vcTYi1f7DDI2KXObyYCzxMDc4+tEUDTrmnFk5dA5xA0wjPay
yLS8pFgQ3ltWyewlw3GT2YfeE/1sPxOQNFaJhLkMPqavIvzRTa5PwgNWi638i38d
imJafXRduSEYvGrxGKptZU0lH8UvAlHn/T6MUNr+DyzQ7j3twg+jxbKDpRRgpJBD
D4h8iXkPITCqW+Zj2SXGzjoSjlxBiLKOhyQZbS68XgXyn1vPT+DWe3IuOtMfh+VF
RiufFzFYiP0hEmUvNZgEEccn3PbUHscklAbqA59eDW/iecyx9yXOQpqlkTDtwA42
SMUI6N3Bpj3A/6Vq1er4DNZq3WfQ32o2Ki3bKAG3wMmEFpSFA43pjDnpInuQoUaZ
OroebDAcsqnQtr+iM5ii1nRAOSabw4aLP9/j4Hbj7WDq1Bpd4JumVO0f0AG3MolJ
Oy5a6y7hdXl4XfXfDBnPMD9WEjcUIMA5hEVOdoofRtdv4/O5BnxMMz/G78iQzEBt
xFn955C3Ew9ijmITcp0zkonZZX2mMVJzxY/WXxZic0E2kg4AFZ3IGM49ZP3CIIfW
z0KlPjegf/U94pTkfX+ahBMHTciW6MCanwVK940eZNjskAEKYoSBnIo5eu5VrPwq
4AZe042XJfLqqIiN7Dv9uWtR5oOKjzfIZwguOuNnrhI6y9/nmNEj6rPG/x2pa+Hp
TkQMYdg3chOI3v4OtvdNYmARfqXBAKHHNmFjk2Ankjxk/cGj2MVV+41Qc7oT77Ax
rWN1VZJebJM+Z1m1h98bqp1O5G1etR43EHh9JD4QMjOpS6NXT8JpDbI/qLNwYLN1
RcZILa6htfHX+cYRCBkkId8AJTR1/avjGTsG4EdFGbpciYLfZX1bkzOb/D37d69D
Ita4OnzoWHvwtkUnBfGC+k5v3TgxHJt1ZUW/BSu9z90RyQPBeKMa3npvXGiD/lm4
A4q9hElLpxA6HZew3FcVic2DQUmsl23naghR4ZxeMiBXf6tUub3dxg+aAoKOiQpy
40P9MgrclDlsaqYFlog6KEvaO03TwHieesEpm/tDdpDBoOl+nO8aCdWxTWZSp3UH
Ts+F/ddTrwdshdcVIafCAUpMhzWdj/4h4AUlJ31FYnRUrrejHMZxOMJ4nC0W7rNq
wRnUhgvnR3BlzA3SGPgxBQRYqcf7v34U+5/1Ur7Mb6MDGLs0ttcRaB08vfOHQCpH
43ZsP/A3LU73jIX667yZ5JXJV2O/tcfgNH/6pu8QEswa6Z0ga0svBeQVsZ7eb5vv
OFELmcDiXah8RoC2Egab2/zJR/kYsXm7qIM1NdRTXby5UH6pgJSzdeS8h/281CBR
vvvhrjJGKJ82B/Ys4TGoeCQ+rWdcAxJNtpAlNfAsOzl/GDBYFUEC2C/bxbo9eqV7
V2oFNgJIJOueB9VSVWT/WjPwwrZp8Uz6L4WIjeA4jjI3yFQ0MtBx43IKZJNPDPoG
YnAj+vLurbtPD3/ZYzVGwuczKh0bKuLgyv4kTYEh/Du5cMeiLbs6Hx85Ig/3T5VK
Jl4u9W+F15gc0tYF/vsg5P9H7yqssBSLE2xOxsr7PJuKZni0KDPUrFsxKFfuVQjg
/IliMtmlxsnbMxMjwubmH5NgnvGuQwXmZnNj1YG0EcbWRJAcUqfL9oaVuGEpf3AS
Vd+m7FukHZyz2eKuJJ/0mINaL3dLWzZSjmZwFBsBEjTaqhAqNhSlvRfjPCXgtGNi
GVl8br5aZRD77Eg45DXhJgmJguoEIKPWZOne1ZxQnVU4IL151xEoW9O/T9yiQfFs
PJeRSK1CIEXDSyXEwDD/mRAgemnjsKyMlorzXmH3oHk0SBw3SL8EuzZR6LcBqdKQ
6MrIt00X3Su2WQSOnufZ6vA3nFvjVBw2T7b53v3o2F358taT07SihZ95wHz63S/N
IIgm9zolOJdZy1l0SWTDm0dRMzrHgD9ZhBTFnrtgCSwOiWboYFs4QrmTMzfpTubN
Gx0pLQ5A+8YMs1eqe1iHPTeiRaBvH6QLR/JZp9Bu7WnZ1e57if+5LaNIh6Hewvjp
KBGFc2A9p+rGf98zZ0e/pO/CqbOl/lVaVjID76kqzd3GuU3Dh075fb1XmMBKG0+n
joaPmxVwmWBx1mVkm4wSumJwkyFYGi/nIvZFvUPuMPUD0NsgTxYDlYPyhsujmI/c
dRiZJzM7gkOEHYIYPLE8gsy0Tv42IP/hOWFWe5+6ZVqf/ZT95bIV/xcqxAnEDPDb
ZJZxMTqzW7I/htEYBw1XVDhVSY86NuvQD3KDxjurp75TIpD7hArdZd1sJnqRnE+k
S6xH13Hg56OfVm1XU3i+5uW5Whsw+LQA7eTPn6V7/Jv5mXdrPhbmeyGfhVNcG+O+
YzSgF0CO90a33y1hBpY5Yosh6ifHjF36efJHwFfbbQxM2rN+HNyelkeN6O4WG213
jcWPT3BW0NAGw+mcBcX1vIQM0NDcB3YAVWoIXWF/KFPdZ0fkxO92Kp3dmQhaqhH4
rXUuw6ELAGU5vBHGtIpEYIEbg0MEfPNn/gnnPw2v2iHdTtQxdao7aSVpyXXHTR4+
sc5AYzoumQKQXF5e1peg+Q+FNpS2g7oOoEr7FUs5220+0bCb0Mt+BSde4R6M8k3E
9bTjvY07+hRyBZNRHq7IYcbIPy4AUbMKp1lm6H4kM4RbogHlYlg5gnjhj5CPnTem
waPE39wS4unGEiuwUiPyZz2kQzxa8L/7Jo+p4/IyXalWKZgzh7mnx2XWtjjGJ8ge
a96q84jhyP8ORLtacfjTWT4CNA5ALCAiZIlN6mQqqjt0afMKK8fP8V/Sxuqvriqw
EgktjyTCzlpSyF4PzdpXCELmjbipT18VuGXWtF5qRo57cBLZG9PtPe3nJD/PbrEV
aSEX1Cj0jL5E6EbtsqOhrCqWRdyOJFVWLdXvEWd3GTdX8it0Pfiet746F9rETX8C
JnzjVLnYyS145FGDDtyf8LD5vdG6KY7mDxSYg1M8jTF5KbC7guWjJHoG8JjuSBF/
jHfseKvCrjHt2EVaEEkOJ7kaws1vQ1f3nmdTpm2DqGtI7q4fOI//E04UXUwvfvgb
w/H6s3CX397iRvj7q8xeEwoTNSkt3pM85REmgJQrfUuN8Nr1OBhWGs4H4T+36xpO
4GcZ40YmtU/4m8XJHiwOVRwriJpUjJBFEqE+A/p8oV7aBrU4tSNgGWkirPCxfexM
aqjfcE/tz1Z4Q1L5DeFShTaNdmL1/tUtvrQDzOf0lmYs5TeOmfvhVX6nPi3cBjh4
RzGjME+QQ5EnXhLcPEx+J6BkzLdhFtBUJiJxsPxW4pAvL19sW9vZsHqJ6bvUIuvO
9MdF8Iz1hMxBolamY1HO3H1lsH561dS2jpaKAQiv4SNuGtqSiKtNzg1QnFv/BzJ0
WBpESZL5IJQ9bH7JHf1HgcIlHpmsa/Dw6wjQc8Sm2R96tUXTtUa92OJxlfIVtA54
mnLommU+Il1b6TjuSt5uSQjn8AoGhAhzQl5FqcUfIzgECDNzuXWhC3sV2s44q+IA
aimNdHhjRa9zADv0gSGTaQewNh8EMA11QT8tKuUMiqUum9RZP5t+wNnWz+CmAvIj
76XTgcy7FnUNS3wnsxL6IOliCo9FeBhWnX4Ep8rw984tFsqW/Zz2ED18LccDKqD4
kcuVNNcEoZp2t19pFP2AjNWdk6lqiNyUYxYaibffHCgkKRk546rQLs7J0bvt5Inr
+T45xgTrIuTowaZnPh9TdUL9rCBW/qlgrFihWbjCGkFGsT4PyQ8dVaCNy6navM6p
ovCLQ6lxD6SPBix2Joldbra7c0HMNowJSiwqPsbjnRE52bCLI7p4Xf04i5X7byev
pZ5lCQk63t2FBw0Ta2rlIT77/ZYHtYTzecR6iJcWXlczba4DDG2DA6sC4MDKVBza
wKLPx0pb27eWHOf2G57BtdI12Zt7STtLMz23fH5RlvEABMyuLTOEjD6PMx/rdq5J
05bzoy3S9lhVhrdQYFZ6mnke2jP/fuQNo+7fux0Ey08uUVgyQrHtoIHi2kdJow0u
J36boMEqnM/6l+ObEKD1zfz3/osGU2+sFFn7HHnkZiyhgLWTAscFLUabKDCURaUS
UOVpLNf+YpxbTHorvPDlmgYxjGeV5qYZdmO2vJhYo3lOh+6FFsaI0MEdMLV2hKVC
zLHIBXI2pTog9/5l+VSpFc86pyGpfB3h1DMhboRG4Ag13M8sKtenOwV6i4JG86sp
A1WxigceBDw9kvf9PtwPpv3FftHhaA14mXmi7F675iGNR7A5DYh1r43ecBFFknTJ
+wOpAIFAT3X1vUXvUURQ1p7Tz76KxnT/4bt8Ir/ZubrmwK3bpZqiRzlDgmCca3x+
WnZi16FEwrs2nj1DITHHq9AGAO4CostaCihUONsjNoxJl0ITpj2WdJuEPvPZnjFX
1h7QAaIY1tJAzDbdFQCr8Dd/WpmrpqWyPuGO9+w455eBwiSwuRX9a0JiYKTBSTl4
sReB8WKpWgdk91mhzSwFr/8OGu5BVh/BsOtnRCknGGVTndM0jS6qVV2c0SfhI35Z
Cm6XK0pa38DvRDASbXVCj/v31QpgC5oyw68eg6FRvF4cUk9SGXKVWTknYxdTIxlL
eHAKvw35Klw9v+wz1YMHMX7X5Qw9u5gEpo2PsM7tC3RQPvinCvAhw0I+wwF6Tahq
qEZHZ/efv89ic31NrQ9+86VVyxbXaU8UkSVmhaoNj1fpcY1ErmPkMc5uSZCnbyhR
oJVtzeWo7t4pvCR0E/bAnPJMrhOrTEfTvkGPAqS8jEcqWy7jqhWdk6Z8s674FHk5
WnySY70oNB0kUekhSvBquNtSqws5ts51LwCWfBNWh/V7tkw57q8B3SCZJZaJxwEm
nyrFQh4Ee4ZgXtJsuSVdXMeykLCBuo57GBV79elR5pIMXYqREEhJfWCKmGwCXNi+
VGvV8gEdxGgT1UG+6u05T070qGcsQV1hDiwhsZx9By5g0GssgXtkejyWpsjxJICm
C1YtbfkOz1etcyH+jz0EglKdIsvn3h3A79yCb9Kp1t4urN0yMbQscFE9A51N54Sk
wa2IEP7b9l7JApLjTon+AIuafbfElsRw4sHqKGKZRXCE3ASMG9zoeF73GKJD4huO
k1Ooro9+P9+X1NZBbaA6fXdGQqeZCVrdX1gZK3SXr2BQPlZxoBfJ3WPXFZOsq1oX
vZOm6htf+4OZMZphTmzbrHadz2WiXE2xTRQaBx/QA8O7c9z3B3ghYl4dQNjANRIH
IVKDyS6xmA0WYozdcNGMkWMEfsJ3+/KIDdUgBjxpqOX1XVzriXnzqxeHcQyK3bXE
2K3p1/7EogHdDH0IaWh8gxGb9TvDVqPuHzFxWjlebD/4qOOhGy6DVdMX0T6JIbF1
pW0i6PQrpmX8z8eVbw3OJP/FOtd4eNgUNKP+kpOvofq/u7bYn4PaRrCxxJ6D0r3Y
Dkve/4eJpHVYml2EskaXkbO+klA48M7CntTFDk3G+2l9tXb5GeJcjxeVvfgflMEs
tmT1EJ9r0N42FfM5jqWdP/byH/+nPX7EPcGYl98HPyPSskIfBF1MwtH2sCfjG0zR
QGVIpTaPyKI3/4nj+SUN5h8TV61CyGYvvJ0KdbMCavzQqkLqIOvc4l8vPVk77fpT
cU3ZW3y81wAeuMpEZlki7p44+swdTo4boBlv3DGnaim0GAiON+YFjRF2HylNNlaV
rKlYXU4YzJJbdnK772wDnmZ8VxViBH+OBsCW1Bc4xWBHnQAlJrjAmlHTUBF831VX
MJYJ09VC4/M3sbN3z7ufAlbQ+Ap/v3AdF3MnBz2xxqCNuP97uXQCT/apriQgWJqY
Uy6Qr+3RbS7fGV6ZqlQ3qDAPK1Om5NXcs60jIETQinxDiXoO0ViZfW0xYQXGCo6+
ByiWraHRvDPCuUyw0wU1GLiLDT4ZZ0pJE5RXf0qobkYsIdhSwydu7aLOtB2aXEHy
IE8cSUV93ep44qqVgs1LkNVhPr7Md+c2oJBIHHpIhaVlWrnHFeECJh/phPa3ocXW
hioym8U+BMlruywaJtgD9RajZkwAIT09e/6PCX3yRNkpXCn6mk2wM74Y0Fcp+6Ks
rFAqGRYCQ6ihr48hEF4RDNEdkeCh9Xyj2Rgtm+tqvm3NM57DJVSoDoFt3/4EPvnQ
i0JNy45gFXyebmZn6WkMUgUiX/pRFOO+ZsVhvrxlsjGZUWnPZ6qGk/SZxbvVo/bK
48zflI0Q/Lm/E/vyhUePXhDnk9r0M1rA84d9NlosRaRX+g8uHBGemIimjM7kIVtO
uGL+JGcDf75xDPyvvHqsqA7X1uALOZVk0FEzlyNQ3xGaA5oEPpqCCWAiEJr4w0kj
JS5Z7ea3UoF1vAI4QtsZEDzVV8BnXa05F38Mz2mlpBsrukS/uX2Bp3B/QhSBHA1A
dZ//7DtEWaw1hD3ecfPDSslkdV8lYa6omnMV8WT8D2/KP9ih/23wnkY9ZTZ7oc8y
jKrHXSCC1NF8BceRmG3mjYfpHs7CHIbigEShYBwocBT0Le4m1Z4wTNyyZWgemQPT
pYZUxYA0XfOilZKbHZoGnMbxEpLrdsVRr4sdV79AyyFSq/lmsvRSciaE7JXyqpt1
wM9fPbSKnU6p9QVOOsyGAV6LDsv/nA9hSfuAj55bWJtp/9+s3eJcaGwcPoRuzqNM
MCuafXiiEyb0S+Tbb1kK+96QprjwYa7FAEFJzGLWqV9Fungc9qZ0D0kuvfoiuDRD
9JT7hmq4YN/vs0b8BkdSrUPiaG386YV8rmNDFCiONBbz7NwdW490/vs3GN9ccJos
+Q156alHzaH6ktxOmBiohkHbbDzOGsecDVkeuvHmCe7MCfEcCqAdNeFB8eN2/OKn
2XxO+K0S2vEe4NmEswm9NctCEWgoAZD1NDaMtyhdvSUFq3aRPeSGOV51aqBwewHv
eeqG5sq5UpneSTKaxKmxbO6PE/f1ajg/H1z6OEb2iafe1ks19nZTQkmyglVC2AUH
Oqhvlikg+c0nG79AsB64cjSL/w8IAuLeOd+3f+COsnAp7Dj/bG5uixF23oEg8qN6
UZSVNqYpTOSIxV4xBsrCHHB32i/HUe37ra1AfT0BQpXd2yN4R2hbB/yx+5ExQieP
0ZWlj4a98tsm65yZGYg4IscW3GDd1dZgjBTH8KXZTPgq2vwAFze8s+iC5S4PnKh4
jtwwRCvP84ifQd6pSFymGgSKW1jjvO8ysuWzF0jpfEmcvwGlIlENgu9cGT+n61kI
gMEuawMrb0y4pYjySiIyU3VihsC6XoDnz2+sJvdAS04SfeS04HaND9COjxI2oLla
KQr5ox6jCQXHGrGxT3DQC4mbtKMNvh4S2VA4crZDfqyBucOAqXHuJldF77sKMw64
4CN1Pd7lQ9Y+SIutquqt8hsERzHnULUV24dl4SDeaa6ncwa3yVQohGeJ6TLsPc3X
UNjM1HYWoOjSO18Mbgj6zznpVMmY/xQhvQcHk27JW93eJx4pkHx1qdZbOAPVeU9W
4Xe1PRTnDBIZvH1bx47rKNVUek1L2deUdJyJiv9i1sFP6FmPO1Jrp8TYCb43Eu+/
hhgQPzvMZQTBUZBh/Dv9QqtARkiMI54La5ZBaYUpWGKvxd5pRrJscuTMd3hKikVW
Zo1UsHm3JHb1pShNNNWaRGusZXYqph8qjBrdjKyORotkVj6t9dHOQzLCZonRrpHm
dQmtmQ3KM4e1EV83QoSPM2avxTGA9XzN8rQfT+d1p6yUHW1wlmVWssny2wFDpTVl
MuszBV/5XI29dD9x6WcUgFVbKMTl6/rNEBWr8qvSdS1piykJGQdmbic/0gM5XEmK
E+n3Bf0di2OenS4l7krarfULSXjemDQ8qKy2CcOzCZp1GIYhONwyJQ++2BjLmqq5
q83bRpbOrUWS75Qy/pr00kMxYcAHsrupNI58yHy7jJ0Au/FL7/K83ebwthoBWRwh
8uwR1vlRJEkmFY6GOGI4WYX+hPGQ6TheRKzrQasFuuSuklI9aZsHL0HacNH+5wxw
kGXZTXNeBR1Y6jy3JaqfNQC1IB+Soif830W9CnLGnd5DozKhS9zi3PziROeXNP9i
4Uin9jDb0OFco3vOBCaGydjicauDdd+aXl/w9SK0amQ00k2++h7t+z3IXvWWb25i
vaS+ymPxjwAS+ShCLTYlGImTCgw4Zor4eulUd9IWlxqbFiHAnrqv4f4cZznxY8Ki
DvamLmqMref1hNPx2EchrY/nVV+r7cR+7J2p8YVAQ0bw1oQBadUZPNxkPhrTDVIq
Hqi05hIOgTYBcxrQWukSme1RYcprVg9x5VZ8gARHig8wS8e9dPVH6LlqLnw9NNea
plRUF17Qv58iv6vyy+nzQ4+QaBgWKwbhigBJ+tCDUjXBgyzmfSYvuZ8f/0onPZwa
cm3z0Mj2bX38sf2Bp8YXF/nMFpINGR12U6VHzhjtVJN4E6yXKSE3UdMcJcRcCDva
sBnGXSwvl6Bba9byuA5dg6rmYuwAvwPqw6Bl3QRNFPfqWsQ4t6vTvbw9FLz1aDCB
nsyBsYfX6wTDy/safFbg1tZxXAnNv75IfsgdcHZhjqNI39ip1PeyNTmHOpQytRDh
pfH2xjbLP0K0fyB3YzRZx1noQmn+GNUe71VcQIxZ9USkg8WDPxfcr9FLfq7hGssE
jXqcSF3QWj5wz+SBzsIxwRXavt3F0wCYTQw9Ht6pUz1WQDXrvL6z0rfAypCeekKC
e6vyS/oRDzKGmZMDaFd2MFC10lADnCcFVvZTl9XSJEtAIp13mbnNiSU49JQxri8H
XHQnK9oaq07H+VhzDd16wnzX1YBVRNnvEWUMp9tgJU+aCZg10TnGQXU2+nzsiveL
NfXOm5/Tt1lEf8dblG2g2yVyZbOMa8qzkrDpXZVYr7SEFzp25mYdQTP8p75MXTHe
e11wnm6ryszcUPRIPBmLz+szfMh4t/NJmMG+gtj4UU2q/f43wxYe8DJVxANwUlGx
flt+zh6wW60UZ82lcwfL6bpWFoRlmP5uPqsOPBdEX3HUYbWWndYttAzzz3slOiZR
g+mINki1RmmXqZ76IDXalwqj48GuQXms9XaUa4+UpOUjgJwNPwQZMxGA1guxljf6
cg2gBK0ElMkYD5aGNKCUd3tdK3WTE0p+ghQRgYkn1aM9kDv6aBZFEwDoCiTM+Vjr
jBJlajT9q10gEtwaJYjOiP2HbNKsoX4BgZDGhQzj2Pd/vtPdKUzihQpYHVFyyU9e
N0f3MxxT0o8TErdt8ERwqZPYdIrj2jqkjQGJRqZsh2wqokQ/zjZLah0uGU5ddfFm
F+2wFQLx4qZJNF7tsXgsODkpP2BQ9PooWdMI6OMLgct9yQD2DzTf8mYCyGFkjtv7
S0MhRNKIAowoODl4zxeUMIYw0MzqtmcQOI37ClzYXRjhGzMq5KLZdXxNfQGon+tv
Vgt83R2PNSMIMTZALUaF78tXxscZcMp4j7sAhpH51C/1WHa5qZhK8VoKBXd/HfOp
JpB3jj8fB2HDZ/wrKF+lBro48QUmc+9AQLYtRoseU//uSwjFssWWvy4zjuNLMwcF
z7VftrQha1KZoiYAjabgjRc8fAmCh38hj6K5yaC3Wo7K02zm2+KtkOBwxJr6xFU1
ZrTa1prDRFEQX8Zrp+hnqNdJHBUYN+vSeni8+Ol8G8q/LHtZDAZZ/qohN7SyAhvB
nAG4C9frZnm9TtceU8cxq+Mqu5TaWWex2Tt5LSEvapspec9LYvwOH6ea7kASfdjv
lesae6eqaaHhoox8qke3W0CtWTtGE5i0WB20hXiDumIJaw05t/DaYnMCDNdER/gz
h54IX5FDRU1JCF4xIuYThJXS5xqDbBmrEGIzKZ31uD3CqWkURGKSfSy0t528ljL/
i9xYeuPWhwcuTv+evD6Ou+XjfH0caVwO753bbix0XcKAaCJ7JR/mOM7Cc0QNVRAU
i3O9gk4Tc1Ne789qFZvr99UnKRzbx5q1mkKTog4rJd5MSOfxIinF19nbTelUa8JF
ed7Eq5XRMUdmpHGk+VGUYpwT2oaeImDD1aqDQ7CylH5QGXlL/VeCypsj6B2wPKqo
M9alw2GlHfP1k7hjWoLxQ5odQc/7oLCYBHxrabki80+P0ONRBXnIr5fW8ZB8Ji/B
TYVb602U4DiDKA03JPkrXm8tmjZHaup1h4rFfJpBP5tQvGUpZYZWwCOlVXsNCJVx
E30Hux0+v8y7pn/DYo5B5pZRH0Fii0rtGaUrzMtn0C1+5xTCpPzzWkKx9GoeZQtP
Gqdu/nMv9kNiHIcqEeuW9RB1SJikEfoTcs65RSpnqBN05ENLK4F875/sE9AxjS/Q
NjMrKNlH0tA6RyKbWG8Y2p/JMvrHSbeYOec+98WU0kwy6mME96R59vSdUQ793S26
fHMUhWfPsWxtALBxtE7LZ2oP3BNXgfdbMgxI4GBNT887GvW08ZmK49jRjK9KvOZS
g2EaDeH2URetsxZqDOI05I7lC7G36h5cRdLG347fkLtTTc8NQ+/E+zWtU/2GumuZ
HiBM8hDdlNZtY2Ayq3vgqzs/sFiGHI2jPk5mAbWfYkQfBh/dTqaSJ0PwnNcXaUto
DA+TcXL9vdCtAyP0h7xneCspR6VlvB/QYA6YEkaZzlmPJJIcpBgFZ80SOh3pHR8v
iPhStfpF36qdADqxE6CQym+v0EA4WHrb5erc9xfK1apb0A2l6c4pznLZ4x2kFBtb
asCaszKKe0+Km9kyPNb7bNpFEgtJa2IC3iWughFA7ytERQuHrgCUx3tZJk31uHtW
PyCoxe7FmDuw7a46EPClKfnhDXYFdQCywbQvAb4R+04SwFgjmdLl8bjE+tEp3nm3
9mbwim91/ILEmM/tt3ysfg4YybE7UrYuP6quey9GfsKaiFOx9OcvPTa2kYr3vfOp
hIybJC2zCGckjpOQs4kYxlpRewG5rJxVBhZVols9EmTpkfqtyyhn5qCqs9x0Iqkb
9mrPdUJgQuFiZiY9EmXC8s7L2BcM8zo5HagNsVBM78QPo28Sn/6e5pab8dSS5y/k
btO7omH3iXfZ88ALVn2IDQL3Xr2iPZxwbBj9xVUHKhCluB5ENi8bMiVxpDuWlV24
UfXTQiaJRDS4kEO1M0rCrgO126Dp/Pf/UdFvvnUBif1fNyR4vQ0FBKQYH+nF0B6b
ayjK4xs/6g/XygkLtfwjZoYTGZGXSfmHi0nhZlL7ePMPoZ2H351wdCdb9V9qIw6g
9WUgsx7/+WrOkBdaCSmWRbYAvLyAtlf4ipXqCp5h5tOIzdfZZbvAiv+narIDPgO3
HY4rF2KT2qWwx/0TldvOqSmp+Rr/HhM8pwtRgHuuW1fImEO2ce4rKl/aszM1dTrC
35ss0/eqaKhDyh+OefGANyplmjIm1wKksd+4gSLtRxWHfkH2gSzPrbSVb9KPLIyV
aeLHAoDG0YmCrm0LqrE1h53/yveIiGWdTIIhugNdyPSeh92wsFlbn0JnCLYGK3qE
mc7vmLmL5v4gUoCl7NfVAHxb5RIqnMISK0DTCl5l4RZNINvhgWk7oR8c1hG2G7Hx
kNsnkUm1XzEYy1gfDh1NSVEZuH9piQwa56QgAT0CA9GKmf+XF6j00rW/ktCvEmFR
ZM3UJcWDU0wcccPwAbxAl3LSl13DlrY4eC1fu9L50Gxd+JV2Vn/RLBki7Iks4yy7
r/SdgJZjThH56Jjc4ykWKiMeTX2eZvlkPVOadTsd8tK8VZJJMAMngXZJ7ZJsa7du
FlXzEWKmgYSYhnplFuzjt7oBrF0hSz9iBk7rcyN63w+ArO49A2fb+xabvM6fUdZd
hDk3Pr/VDTtnF9cA4D+5/1S4LPyZtKAPEoKpa0PMj1I2xWjzeBib93/c2i4sjXa3
yoB2spRMQOxjyT456VF3bxdqVfnABQ4o2B0fQqUQ8ywIvIt0cSTFD19T7qqfl3IL
D4+DqcvBgBvpDIo5u3N/jirw369z/vtUND4YQoua+I+T0Gg6HTaB9Da0DiwPVuxI
RiRzD/jjwVBbyqNtUCVyaEWS9R4GwHEllJohdkmaPhmwDrZi+NT1mZ/fzmgyxoUf
fSZAUusFdtGhlcWCn9qbGRScAzpdKxghwn68R2gzZ2GDQH1GCAIihBOTVurls6Ah
zxl7yBAE7YM+2FfVMlvBO4cRMazGNZ5aAg7BCHc2thXZeedqED5xQ8H/ks3i0uGt
Vae3t9gy2KYjdbwTJduGKZF7s+zJdOBK5V9Yy7l2AtHwnyitCUIafCsN34RSygmw
MT00AKpp5w3of4SRIKKnLvJsypuxoBwaj3YS5675VB9hzZtPohYn9SJpiMVxsTJu
7S8XiJHfZB9RaGOroFGr96NhLoz/OxLhToCuwx2Cs9WKTZp4hnMonnbUaakkRcL+
oSrTuWp7NS5utSyeTfXsVQ342qNxo6Y22HaLZp6APH/+wtOjOrt6L7o9XtGkwbbS
5MuMF8cWlRxTv326cAN6aWFk/sO6HMa0mfjzWqu4mQxuAXw6Wo7CMJqumyBlaZrz
H4X1sqDI38EH671CC7Qa5D2RiR1NhuUZuquxKDOc46KakO2QqG2qn37ky1WIVtEo
tgsI/lnSLs4ODeGhPga2LpON4+rJOJVCPzxZ5fi+ay0sRfUAoriClrsgrFgT3P03
BR2BdbjtXqNptAQJxeUQjDPIlylvUYuBNci1MY2iBnYJq9iOxs699EH7uOqQairm
IcIKSwxekrujqiPMGALTxmPzsuD1t75XSFp1u3/GRBFlcv/RurYWkinquFHyg+d9
iTskVlYs2TRK6kSNwGwU9X0ir8xRZXXVhk/o9PuuFO7HMLspmJNH/00cMRRgyzWp
G04prq6m9R28PUQ2ZyN+VVg+ui95NmTdVNNPB+j9KXsTt7HuaU7xkYSox/fEFoEL
ooTmbxO6iwANx90PLXHiDy5Kg6bYS4G2z3bMvmuSDji2W+M9y2JEKQQJYgItv2fg
S3WvQ6M5xYWPGway4Yqh6qfIhzjnmwVHB8ObA2UfiicRiYhrIiG1mtEFIt+N/AFe
grJoaqqO1BhW5w7lFwQX+kD1AxtHDhF9hhj3efQicV8KN/IsS5W04fYyaMLvBZEW
Xr/kLOEgqwi0p/Y9Aymt2WQL9MlgFsRHncZddiWvqEeyS8OSIDt7C+uw14yIvPKW
O80jXH9F9uBUGaBYrijhB49j4T3HpBHT1b/B8QG4uC5IgDKRiDSBSHLACZKB/RyH
sVnc8y0MMrAxixFj/oi8wliiB6NJtsFBMphcEBhbM1hGRgThuqNQDwLFln3r76Hc
lbpOG5NJYP8Uvar/KDqUQ2UGSvyrTVUNGIeo9/QSTFjBo14aYRYsSZcLOj+ODuzd
kgj67NP5kjmmLpENjGpIUGVJrVp2JEj266JTslbRpkwMrHCdToLXEy8IVWzNlyL4
AU4huIw1rwRlxua9cGagZNlV9h+IZ4AL5G4BJw+xVZtuICn5aa1A73wEyRZZQ5Z0
ie8sMm8BFLwKqc7HWS416Klp99QZy0XzRDJIK2+RuTt4sd/+vFoQgPmqBdNnPt6V
wzu77agL6k7jjmFhD6/ccdY6omo/5cEe00LlWai8+7evlSAje85TU+HSTJI2u/qx
9XRXmkwicPs+CHkkOAZuag/GNrJtpZSQaVEdMAqyJMZbaFdoJzKOa+tYZ2hVFzBD
/aNDoTTXOKLcmixbavKfYaUSlZDyNeY4S0eeAwUvrLVUeHYvmeqvY3Tc5LSWL6Vt
DAfXJJ5C6ECiOXyZVVNVFL1jF4DOiliQFrWXOh9C+sP4mZucBEXgbYjJdpYupsPk
S4KEMqVl8DmeFfUftTFiLIb02X5oFSsZWotwKx4KgD4tDm2g3z22pl/wglqMG/Gk
pW4W57y3hJ7mXzFKLralxNZDh76etgCheBs+abkhrca9RPz+lH/Mui8UCqqlF/hh
Uz/Z3OzcqyijlPRAjKjZXG+cL/ul8ekUjoT8Q96B4BltHYQgWOveDr64EXZ7bdEW
imt88XgM9nngZ1gzy2+VPf8IQsVJz+r54N8oQ6NsWZh9pMYTX50AoM+sucekp+LB
eHyL+ivdbcvykR5CJaOUAk0q4QOhXT6ULlNJog4gj1U4GyqL9lLRk7O+PTUd5mdu
lYOGOwlGIZBNFunul8f/gTxkpPDLVKgPu8BeV27YvyW/U4bu7KDAYwNOFp9ASTlx
zjWrUY5X+wGWzRt6SSaqfVU1mo5AfhcAcS+4x6Wn5FShboMACpRlBsLu89pJFbzl
Ahfaas6zjwLApuWgmDPFvYeOFZTZglocUeZDWFIC5/gpEGUM6xVQbEaqjcK5xPOb
E+jyoo/hp/LjsJMb2AMXXvdHQmpq8t14RIHcumIsYXoTvkbQIdyhyXdVVfBBe6mp
JJS9un42THNmdO/bJbCtKZN4X8BqBc/cJJ3T23/4w+oRy1vTQwCDp9k8HIXXvEXR
CCbYMz5Faoby2Ld9C5M0sQvUaXpKhl6PIft7kOaHpkyvbiCFqFd4Jxlhm1uCCqWV
gn05iTWm642HNaTUo9gNhw4/tDCzT7GCe3thUst6MMZ1ZeBAgDd8XS5tJ3/K3HLl
a7Br1uFEajggAPZ8k/qIJseFADQ+djY6d51mcCYML4dD+qOkVeXtggcoO0Cu7BZk
Vxy3ggUpBwMhRiFAC6pQNEid7oCQTDL4tAneXyWwJMCs0R4Y9SAp7uVA8h0Fwsld
MnpAamd0hOzoEHFpCk+oggzVnCh8uUMY9pdsOLNcWNVt1Udp8hq0QOO+EKOAvi8V
qVJvU42pyGNwp7M9Ww+JHhSoI+oqWCRfB0kB7Rd8/RMiHbMdfDU0knYApP9pWFWE
qhHGHRDzmT3U+nwQmNGjcQKjpJANbi8memubSZW+NfSa2W/BL080/wNyCSttaCD6
vQNG4ybAyF54ZuDXN32ATm73o2pUKdN4svYTZjSedi3chRdD0Ut4rFnFpjLrCowe
sGZCH8rmmovlju41fgnKNWfbK6J4O4gNZGQJ3PptpMQi9Yffku0oKaBZJIXt8MbW
IskVkdYCZ6xmmrE6iazQkekysD9MqjrqZiNVd5AlMhjzFhkVSBZECn6pzXnyBptI
XEKKY3jgKjO3F+t/hIGwzQBwz2pssTF34tkM8myvJsOJPJoQqisLlawZUj25RTbB
rEcExzfNRKapmhYgei2u5o2jBb8w3cPbtD8BCatjwwrhOozUQ5PpNGxcIu+ib7DM
PNzKUzxmeCJ2mo3b97l/+LovhvmRpa2L3/aZPxc0BlyYHfjaCPV6Qrrc/53dAc5x
i9+sA+P3xEfNX/jXGa3hS1xUJKuRRsVUUXSjpl4cXWd8QKBQ9NpvG6JTjtnRpJWZ
ROb0FJJCwXdX14PdQAU6tdTY15YxUbso8PUOBFXb58SGQLc56YR7RXtqyWNkvsJY
wqpQqMB31HXrWsKB5NPlxJsvrdJ7Zf7etXgh+d0I74xsq3BYZDoz0Wry5DDJynNo
cvSQNAr0nytY4FHVOBF2D+pd1RPEinyCy1R39T4DutZHIqKESgSLuOwpqklV7sxI
+qLgL00Z9xxPqcZE2Kp5kmQYXLk1PhwyFiEtze/O3PiUz1fZ8Pp+65dakZ4B+zVo
w35OET/C5e+uE3zUHUjj3KM8sSlEPMdY9ab8AGE4nHLH7RIU6pLFMt38xzCrd6r+
3+kVnRjmABvi1vLukKyn5v2RCRXds4TEtwzmvGmnW8f5uW5hcC1xQuMbH7HfgTGE
zKoc2Ti0iwumtyj8jnYfBYxq974TBIOg2I+3SPhLsuuyqfdUGyuYLb0+J59B6iuZ
fxxjpovIGtPlhK04+o3VT4833KJZfl/MHjpMcqC7nouts9MtWZkzeLGdwJf9AfNo
sk75exjMgwzEwMD6hsQVbdunmn69UhKyxUKDsTazvdOJY0ToQCmUG2fYrkPPFMUn
ZdPxQr33rz2jxsaV3+ucLjLaGi2SnoOSfJsOXBFp+lxiW8ACDu9hAsbuqfdXN1OL
oODcahR2qPuiZwx4EbMDJHsE3G/OF8vl4LYvS1AlNvuwo/CNl0Wyx3UHeURy0AYo
fEUo7I8TeF0TJWZs1Hgpv9zlxHc+p/a797qT+sOyI4RYkm8F0dyQeJkbGj2Sdqcj
w5Yg8Th3us2FqOL4vAQldShfJgiMxBaml3p9SDGMjKIUmvIvwSPhgdsOrRc8VfRq
asB14jCnakuWDluVECnJw99L63Kqr+pzk1LENhdiw1/0X4/7eN2AHa4hfVILx3gl
AnPEnjlZOGoWsP0OuYlEfZrfiNcvlUUaQE+ipAmx6j4pSlH5DWYH1Y4kWsjPB+GR
H/pPEyiVDkVz33FXG37hHAYVEy+W3y+/gWT+S7HchAVas/D+nKUZFxinQdNsIfA8
xtAWl8h489Dh49OWGN/jsOD5s2DeUTw84Y8bPNsQeqLH2S4wz/q0YODFYxyucbHn
Xxfi6o4BpRitkEoIBgY7FwgJS1JP3E0Veibo7lH+aW4IMiw4Feh5xQOosAbSSjAh
SM+r7xHPZgkYEBVJpBd+XoJRKMGzhfwf7upQVgnyPhVwKKWOcksediNr5lW3h4Cr
Tk/skAIW5LY0TOhOqArfg4a++xfGMiJnK17y1Rfg+DKY8NkZ5Lv6pSb3nvDgVGLF
D5CxTnsh2+r89OBIASpS2tyUkVJS2HvZiUQSl4mvZmnzFogmM5jxTzTWUTE+wc3u
1vFnDhnj89Da29+0pz85lpYys/D6YrpatEmQzl3EkP+E8xd13rX2lKGGFJ/jsZWI
M0yp58FR9NgfSY3bSZ1q8kO1JcmUyX4U9AhMgGY+p4AEg9E5ANfr+htH/EYAKv35
Nltas9U+VC0K02EbGuqmxJfPCs6e5frJ/mwzSZ8rUbi9s/pdt1wcPvvj+mcQKK4K
2vk+UELd8Csp8GHP/wygwp9ouUi8Tcg9pUsRhxydE98Ime78Nn8wXCiOjyk4vc7c
ipBVJnt9hlz//eVGnQp5cYzk+/uXMnjKh0A5BW8wLyJRa+eJWVELUXfgXKcEbvqR
YwSOBlJ+7NUGD+qIUXHHrDkMXC8YIi4pPeA7jEFqnniXKEca/T7q5Db8QmgcULi2
mIThN6FzAqnC/7teYe+0a8ZFnAKGqrJfccxX5csBKqB/W3TUVPpUM5kEpONtyvNi
1XHQrmFpNyYIYVR0KfV1XST+szKj8BhgH350sdtTP75U7MDK3yOrdMXbtzSPIuuN
fD6jC9E+bj/d1A6mA5q9i3W6WftsTP+cq/QvoROxkVBGLgoRZfCarz6Mdsju03wT
LSpWFKqUDx8VtBZPoHOFwEQYDOsZaGCBcDQJnnVZtTfgmVtYjzVr9ie5inlzuMuC
YVNZETxXzAXe5c5U6NhXtVatyGTdefI6saSOlXLkzzhiDNcGLEkvlxlFX5EmGmI5
cUbx8jHijQKQQ8SarffVwepEDes154h2wbMN6gE1ZpvBtOZg15mXOFcb3NIuth+/
6d8BRY4adu+24jaNcM/FelL7X+5P8bZjZxAYhkUI9CaCNCQKuVvOwvHS4CFA2XVK
YqlmtORFsB24zoLqLBpZeb3b8PFnw9VqTOAb/BrI2aJmXneN4iOzzI+r6ebePAVe
eF9pnT71WASUMULasPLq/1HTT7UBvtUmLKVScUPZR1vOUXwWZ/3ROs9DdmgrhLU3
Qq6zOdHaJNHJ48EcKIAAV3ey/jkTYXVjxOUysj8CdTaQJxKSSUS8IawxY1Ehmd4x
5p8E5noVI7EGBtyN4auGH4FPLlPRs/A0hhkg0cJ1Z4PCroAF3ChhJkQrMShkVdwz
s0SGAB0pWtPOKO5o3IlZQI3M5GhT4ibnfsZhXMviK450HkXn6h9eNU838flPgDJa
Pf5/lTLf/NTlUnWfqCbB5USBdRq0uOsCoJqwImArBTdukwXuaMYmX0N1M6lOIM0g
EN2dsHpcYWuQoH8s+T6LkL1z0zywkjAbXLxzzma7RC353Huh+UvMSvAwmw1gL2vj
SyeVW2HhYLvlCgAGPGVHsW60QZN01zNpyHzD4TtO5qchlYymKzywB/p4ttsJerMJ
yDj1VUBgIFhaJDGdXdjYJdy9M/HRWdVxeIUhFDMJvH1WddWI6eaWmSO3HUbGMJsc
glUSj8BHVw3xi1uQbIIatYQ6jKq4XVTpCzn48R21dzfMN3a8Xw1WD4YSGF0+P4UZ
+QMEyH2wi+rXUBLXELSa/wQRauOP175wWrYVeol6MBeQwXgdMLpIdYTLO4G+AHcv
1nk5qtv4HKuViui5uxsHledS4x14r2I+itTel1UWKet/xSvJjm/c8b26nx2sBdeU
NJ0aBRmsATyhujzATVjuEWaNN2xJST9erFHSfqyGjvKdpdtLOEafsBns956jiYAf
il57/QeO+puQ4Rn1K8EuH6TRcCE66IQzfpSqp+creP0zuOqkwaxQqPiuv7JMAzA+
RQZvN+eOuyolNQGXWxr+gNUceaY392ckJPEaKT6k+NELsvRd4IbQKEqukOD+aWZT
tjhQJbJEBlQMD4qMffSbliWKWNJ5R81DvjRafq7DyWiQTnnXk8esgCpA7DzznC8P
KlFk7V+vymrsnQdBwGggb8J2UCeNve2IJvQ5w7udqEUDFagBLvdCuCCzW4W6vh7z
8++6qLq373feUyWUNKy5UQloP52S5uQcQFN+P5btlTaZIrlb4rxhO5dDz9uj3hEa
xVH83EZq2Cw9vA6JH2d+iCSO/D/6ftYZBflz7tUwgwVAOfERGDfAm7V//DCgLr1g
y4wsJnxhFPHtP3ICSdUPa9JYum5fqHyImPss8tJ8J7d4S8mxZWkykoXBgmu65T3j
+cShqn1X0nlwmwPkteNPCvKk0+LsKLc7saXG5KM0IVky/Oqb+AS5m3nPnwkyl0k1
qoqWSTE1gVeq7DuPXtDcGoxSJniSRmcGoz/FpLuiQj7Z+yYEP0OrsaU+FCOEQ/MR
P0l3T1+kPpnv8J6yYtD0ZxBH7SXeKstJFgqgljuad5hJQ12g4iDFKCseOoR9uc5R
mA95MYRNEeIdJ4s0GedhJGZGap6hG7CMDDjm8lMJcFs6qzwP5s6TFEBbzp7wjGlV
eFmroH+2FDkvUb5QUJtw05G7diUQzVNugi0V5xcW6/Eqj0TcfGDeNb0wZV2TggkK
iFx7MHGc8NeX5PtMdwc9Wy3YLdhOLhbIq7N3neYNrA57FI4sQRnykWGoHarUfDrk
DzLsQvj6QAvkmnq8Pdue6WvuhT9L7sO4lQYNfwJtQWefNB6a4DZ3qRgJvGwfFmd/
34omVB7etznFMCvJMgGft/voU98iZjHK/gfPZLKpHUZa14+lri65XNHDGHT904nU
iPgPvF62v3Mw8SX69NIvon8QuK784hbB51BJ8/GQ9PnFh/Xi6iie/PUL4D7SPLdp
RW1xdW3wIyFgbefPNJo7Z+xMaHZGnJSjbAafCR0VO7hcrGEhCIWwwxa9ILDmaHdi
PN1t/6ig0Px2HtGLe0DFVZyIUUPpGtpPv45+lin/E4ALQA57GaCQMDJTGDx8ySTf
ZUNCYwyjd4jAGV5YuOsOWNG4Pc/VrMuci3pweYcvpT5GO7GgBQG2TOUqTRC45RDD
Yrh0ZXdfAYwtBbBa067teoYaTCxzmVMeEGv/bLXbaV7oy+HwuOsqmGu5HHpigHaT
ay8mA8T9g9VPn0Nqyc7rk462DR7zbqSWfv3XxYP0GNQzrBeEGtMEgRzCkR+3nHQL
y73z0TqBufTrTXT7nhuxqYaxBzM7oftTHr/2q9KnqBWEjsg/f2jBhVzghaYYwHMe
FodaSrfkSx+ipStRcoKlfhJpBACDbs//oOU6mqlR+3E6nJyGBJiem6banpahqgA3
I9gtf7IFCaTl+VIoTRLVI7+sF7SR6NDk+jFI7NcUYxdShwfxshVbYyvBeTPAbHFA
/j6JLsiMB5mliynOMSq9UFuW3lhY2b45aeWXmQ1to6Hrs27nlTXvdWuJh+B5/Y2U
SdCeQL7HFZAvJw4KFG2tgPnD1skQotmgBBlfG/pB90UFFMk4vppAgOrdIrGTdlik
7wOVAghUxUlGV15Ee3Wdb5ijOtSiVUbIMa0zk5V2Y9FcM41W83Yq2UeAeXfFDIa+
tfFyXsUCxm0V7aKWKDCXsRvRZNQ4XNN2aI/Uhh5j2v/w8mgFIEb42YzekuvufmbJ
opQ17gFJFxBNkJ5RdG7ky+f+X4uZjmfXqcpVBPm67/0bvn+ukGJKhRYGXUaMj9gr
KVWdNP1P7EZ7KY73LhtqOhy0MAtErkqus51BZQphSRyO+9UrrQkWLBxW71TuZnIe
+3rFKtiLumeaOvjNAgqhcR2Y7ZyWrpS7lsHULlnNT0Jm5NaoKI0RVbQYOivSfgQR
/zQoziUT8nwaQ64yUDQlNKpxrcP8jv8N9OO58djm6RBy6RINEI8Xf4mqzA0FSZ29
39bKL0dCkuMU0fbWcmMGHvU1LHgTPV82U7WXUgZrGbCsctA33VovhulESJhd1so6
Y4FBxADCwX3UXUt9bNO9mFFzX3No+Fm8lPVj79pA/XmBvsSMQXgf5sqXXV8RKWCW
bzVVntG1glIDB7MuhB7pPNUbtuSGXGnN3+tC0Cet4fTIislg+ZCp6YUNnrveS5NZ
FrY01Nr23FodJrdfyKccAJVoocWZJjs8RIoM8rEFxOd4gYLP9SJK1CfMlsWkCraZ
eC43GU9DXJw9RfYilfoyqFN6MzfaIYbXsAiPzZO499GO93PE9fr2kx4FojXsTyKM
6B7uWsAE3zJbY9la0Bt6/0sFDzoB79iVp2zyFNpgy/fv58dx9pfkUWA8IFf2Gd2h
brJNxlpf5Y5cdGZLw5YpeLz4D7QSpl0QNj2fEQtbD1tk/1XFMrfHRqMv2FQecl9L
MH9ZAmrF8pgA3KTL31YgCdOEVLdX0809v+GX07QeydKxeuBUSmWpBaTEwYCShxX4
sKGyhwVX0B+pN6aMEZ/Ecx7pg9FFq9c/nanS0soWOZyDVGSshjy8VlyRPmcZIhnM
k/MQs64hNRj4V/K8+neOy+o+GBNUetLIzlkDDVhJwC7DkuH5ViuGSxf6A559DVuF
jWkH29N1KPXvcp06gXnXUnCXy1KzruoDa33DZ3kIxbAUNaJivzx5/JDoqtIg4h53
dPsuqXrlwp+8QC47BBcemND5KcHDEI+HYMdE7bGGLbqWyPP5uhTmhYtYXHiPhZW0
f5OBi0hRNpZBGI0AQ4u92JX7QvvLBntp2MC/+wXqDiiFbCeQUmNRJqer37OApWdp
934Nl1wIiOhkbhSOTRPNgKy1uOhu2UyRT5S4zkTjQEEDWKPKZ61/gsQg7WDd5bjR
i7Ts0XczhwppZ9DAWTD/Gi09qM2jJKTKRp03Z9tPpPKe5HGKq4kRXcyK/Qvt4nv2
jBuhd1BLOzNmlcXhtMdAWMYiSgHsSV7Leurm3Uw5RvgtPbW1lbeApdDLM2SdWAks
31nHcniGOyYeYbfzkygiPPU4iycJoTLtL6gpKX2p0ZIJ047kecWwhHFK54gz2/sX
ML8NCCCKq0dK42Kwu1qMuU41Ea+y+2AKgwBkBIzT3WTsuMte11/h5lLTIAXMfhjd
VIV91QbHRfQNzk4PMLbByYTCDJk2z3cV77JxFnSa3agc9dzvK5ArWX0N0PVNans0
LK/C9dSD3JhcNrPqjzUBSHruewR2Nod4L7gzCOjHGbm50HEtWlYEFSrMfVl2DAUV
x0NyJFjH2dLGMVNW3ZMzYaDyFro6iGn0WTWmT5xWNxasQwzLErI2cuuW8CfPXfvG
iMVnwGyw3Uf0OvyJ47qg3sx8k1rxp29yiyGbjjEcpJTCSo6bbEH87x5pJjA1Sx+m
u+o82BSeWAqNoSVmJXVLZSx3pVIrpqK00ZvH2biVSWab/G+DuxnDPoXQwTb5Xmkr
NQ0YZPpkbk7AL5oGUyBIONiPB7+JOMY/3R7cBph7cQ+dMX0yPQmR0dhMOcF3P4/k
uupGQnwO9qM5z1Cp+60m680zQ0mbiqRlgMa/neIc5J1K+GiU4Me5zUcronJbCmfx
PpodPkRIcIE3Ozzc/AqEodVVsW0TQEEBZSqFIA72V9Yrs5Q/d1tEzSI5ykJ1YqUV
SI5MkTDx8QdTn+hcW61Q/iSye8pFsVsMCkcBG/QuAKIq5+WxcUkT/lBMFu0W5x+F
ANGVtekCCuDtcb7N/hK4wsu6DdzS6cKfvqXzSpdovUUyo00L19eqVYlkxJtA6smv
bwauv8F+ZKEYiNZnWyXNdkaDO+GD9OjLzUG+gTtMYyQvCyzGty6yhgoMDJ2lia4N
QowMV+c5f+r3M59HU2rBL1GNPtamQ7urLYRf+1fIMPeZIUPsbJCMcDS8TO38rxFI
EfK7UmVP2QL9xPr96Bzwuvv0PLDQ7AZosEcQxRCc3PLo+AknPznUfsTxvoY1OfOL
N7B9G84BWzQ+6HAsuXiOj8K8i4vTdzQnIRLsQGc1t0JXK04gI1fNoIiOsDrA6SMX
NdWp5adHgTsv7WdGl/xcTxIu2Q5nKkJ7W6XVA1v2yQIgdOtZLjor5Uw7XbPGMFFz
xbH0loi5T6uZWAWiLf8HGbD1UirJ6X7OMzJX2VKGUFc1ciJx9gVokRMFo5X6O/tS
yLpttV8WRwfCuwdHKf356Lupe6qM/+/8l1bmwtyr0+gIVQX0Z1KVxsbJF6kyt9ol
GuSNfEO/CCnUvLSKglsclPXWu8MI6bhxOYyK/Z2YENSHCS1SrX1HkW1GBB52clfV
cvaFjEaAz6s7rHxhjZC5okSsxZHOkwOM3/HiJlhIbJRL3lodZ71kQWc2s+tf90C4
BM6MvUoceQExYS97bG2BAqi7OPAMyueLN6bGYgSmttK6ny398b1if/Y5b9V2gGuu
`pragma protect end_protected
